

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
CvmaYyJzAT4gGJRlCkE1yXt5Lv9gJbr2gC0wBzixkhI3TupXRLTg9s4Z9WVWp43QDkUuM3VRZjAj
RVnqESt3JA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
hHyS2uxRkJ6sHR79RwG8dxYfMwySDoNzo0ZpVSoiAp/93R212I5J1LxM+7EujDw/cO/x9djlyxbz
erzC6/tIqQ2nS2hUZANmmER9YkiA1RlXlIqDOWo8pOFHNj1c4jf7Zdq7OJMDPvKF+fLgmk5Lu9Y0
15oIyfQw7L+gXpW1qEU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Cfhh7YIOGyVJiZpd5j8xa2ugbHZdDDpkNcw6vvVCCgnGCfzlen3wlGk0omzzJqyVapnfg0aPFCVf
eH/noQVGu1bQkowx0JKcNE5x1v5DKH//UNI+lq09SNF0WKlMcTAGlNSUzO8kgVv9uNbKUHDXodcD
5iGh6bHMhVPSu1QKpTfJlIMd2CMz0JfDQiVbfTaAGKvrQhaqVte7pYpnqiXM7povPwt/ntWHBH4s
XSF4J4eDVLMuQmQNy3vrqFdEUqmQFtLWgNRpG2fwo19Y2lRzT3ux5SiA0Iv55uR6x7AG21x8BZlD
JC102ufirdrREfWUzlClY8zmr+TUHpTF/SgPMw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
UWceDgHVHZAg17Yudaw03bncVn75AJ6y0RYlYeqdZU3kMG9E1W6q5REaQAI7sMZSrC2g0zavsx4w
utskoq80P2avoebtdvBfjr/nBCQqUN3AvM3GSk85froboZgk4fCQ8UtEj2Qk7ob+ox/md7d9P9dw
2YULi+eG04dUc1g45wwF0ZoZdARk7Ml+fXMnm7zxmvqVieAEsVq6ETZN/P0pwvIpAakLTayKriGC
qcrb1S28bOuV+Na/FX9rxN6hM5aK7vSdFqja5GGs32r9UVRIkX6i7uqS9pWQDR0Qa31W3z6wrRrT
+2wzEwNMDKYuWVIM1FQo/Tp0NKa1Y+kyjahSGA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tLsJPLnIUk5FSxPTGLkNhAFldHrP7oFH8h39nfqyEmnC/AmGzR3fePfCEcee3I4TYySABpWhyXIf
m1jGiCuHfIpFkF2EJqjWmBev0bD33cbw1av2xtJRFa5gaQjxChO9URfjedFvCQWWwjlxejc9nD0N
O0V2XUDQxd573YmSBuByzshlxt3bujEd6Xeeb8N8NI8c2ZsfY4693LGdb3k6gtY9ZEoo4XuYVt6n
S2tNFVJTfQjyBEXbuCPqpwGf6bPdy2SKvTE/s4rSIVTO08J6bXDaEOBUGg13XVoJJqrayiJRVuQL
LhoiPzgOqS6ude1uUaMHE/SN9X/vt/6uOsOl2w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jgk19ieS+ZYiySHKvgAHMus0OAx0HPJ59p64LMaYK8CyW0wSM8LIn++sFz9tsOBdLj2gb8IKpSVr
SOX9XXXM2pQFSME7x8q0m+EPg9m1+ghIpW4bU/w4zVq4NBjYydZCI0Hpy+X3op0a3+eENVEw5SoK
4R/zOL7aV/2nZ//wkaw=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
L/BPRr/PHH5da1O06dKRr5ST8eskM6lzR1UPuTvZQ6RCsFEjTD1HgyqjW7/ypnIq7V5TYDC553+Y
rJnEENzDc6RSpzenrYxw7NrURpUedIWlCc/PEf5Zq9gu1ESkpND7t98rc+uiAz7zsn/pHD/K50NR
q9l/gcWkOCgArmADo1Lw9usrfZ8ECIPKY2kLxeTYbh4fsrCpPQsQUk4NxX3N1Q0h3RRUCdHSFc0O
lvGip/vd24OK8zXDMaQv4fPmgToFQMUvLrJXErEUeRlkpxkcX6g6Zu4RMWwwmkNIfZHpc5K8Q3RL
MMc5rARUSXbNbpf28H3iyAMZ0y+EgI0CrKwooA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
kp+3zXmZKSIqIvl0rjsjSpE4vRXqQKS/YsQDDp8aBlfPmKi+FA8sWY8jJ4xwAjeC9OxV7C80Z1Wt
kTh+XAmO7o8b+rQsZqFT4WFgQlvrikjOraGkR9JS9gD93oKswAWicAcGe7i39UmXqUdNwjejDG1S
TBouYcsrT6NRNWPocpuSyjEGFHxQ41KPITsNapgd1oe5J0FqOEMVgKjmsvXxvjKRV1t0rKdS2rdX
hMTMFbArifxhM+RsV9faFFN3BxEdIFKgY/4kS8wr611IkUbHUrBfI7gfqg6QIR791pUWBiB7FDZE
7pk9+ash0oJzlOPWCCLhYU5erooP+s2Tr4xbSuuVz0TmPM2v1G1TdahUYsNGXLESF9zTiKI2kvK0
ux9uq4gfKtoSs2c2VMQy/gjuKXqX2pclHNtd6hSjDaG3II54nHJoWYQeqQ57o3CEDkJZ4XTJnthf
/lnjXUxgndPIYJT/KbMfgwVJNk0RKJF/xsz9B1vKXvlVUjupUOUitEn3h3bg7lRusYhtAYKlDSCE
xfoa4qdKEuNRQFQGF2OHj3Pg68llanihvL08XqxJPwCMKuVggGkWJiJS28H4g8EaVjbKE4L2goXe
X7cNkfqwQ4QXkPJ97xRO/81rTPUxj8tfulHUP1NGvkGVth/gS47sbpRM1PcKs2WL/3gBGUGEZMWi
CLXkH5vVfRAY/RtehIU3ipBomLlp35fB1T+rN8pAe3u1Ic4vSa/pBRjWq5j6uqhnlsE4CxxI1jya
4ru3MNJ+OzSF4Vn2b6aBrKoAItCNLDYcABTwdM7WBgj9e1WDCCRLOmUEIV0KKRRfnhhl5kmHQHVP
a1R+OVA7ddNgS1LDWpQd/4DZGE2QGkoGb22OmL4f5amPuKsokhWjT2bHAxX7tkHdGzBqZZocMWr/
rlp2E+FHHV5+lJ52DirD2c9IyDdQFple3OPLV9bze5oyWBbgQkZOJTA/PbF6q8aPO7P1IWs1Bm51
oiOt5o+XRaRf3wTp1ToZQk0aoNx/ABOKoSAOmYuhB99bgbdNC2bMJ26a9isek5g+TKUURJNh4l9C
NrMVzWXXgANr2GGBr6NSQBovTsyY7Lp/l8kUX1kP8n85quZxWdZzXjfxFnbK9IMDiop5VPMgqasz
RoAonIFbbAFL8IE6BIvbPxOKAOu+z3DNGH3vDpOEK2nwcnETRacACNK+4N6uuq4lxZRC1xwnvhTI
o3riHKSfhrHGe4HtYUZXgqZ8gHALs82kk9PsqKZqnkaMjD92qLs1zwtbfIKjNq66BxcosaN17UfP
uNkadtDOoRgZTbcyAqUKdzdz9Eai7PZ3JltvZotbUt1ka22IhR1WRPhascsX3ZQI5KsMHAN+NPO/
y7Xf0hVlyn64mG7dAFZwVfPZwKWhKiAjvZ4YrzHdGOCKARm6CGz9MTJK1CAsUpspbMpTDDWNJfv2
KgQGdfwZhV7ULZ59E+vbx5RvP97GFhuTB7bNsI2SpD1aBI9+rYlXbOCs4HEyCDiWuaqcKr0UpxIR
6ReOstSnHswF2TqKVQ9V/FameXt32ezKvaChZsQn+bc657L8Gl73+XCxfets/mWARSTUhcKh7nS5
rp0z4atoQzLtHwVhHlkd3BJ3Vy7Byw/hdpaMV5xMnFvg+TLkYq7QahaLsXuzZ2CF5JFZTDBmVsZ3
cJE4Ei1/RzWzdFt6+pxskDsnieWGbht2Xa3dEiIDj8D1ggqaDaPgQ9kUBYPpUkQeKJ+scNPWS28M
UAnkfONrdztyEzbcFGorIE7wdHWhCcM7tCtjgVi+gjHFZrGffPxOFuQlRXKRxUbIt3/DB6tQ0vcC
Qd3yicvg4J68wQlKpLGfYhDY0jsGRlxy3B+fMjjwX3QnE8yf6cwo4Rp8LOVYccIPdCzgmKNHUVAE
vjPax1PLs6J84YISSqGkavDKCc8emtjfLOJnmiok6uZIZ8md9tZ68P1FTJx76E7nhUqnQSpKUQt2
J7VPBAOT91rLap+Vvz4VP1jwfr0MyjT9nGJzuAaoOgzphMzBT8JG3Z6Jscbtwl8XNc9LAExB/FYc
D3YMW2JaCQqIpP0vP1BNXOl25dH1Ur0HNKSuMk4MH1tUniN6wB0ToGVP/kleoNKSW9YfbjFi1ml3
/IjwvQ9zFB05SX6ngB5NmPOUPoTQzpqUV1uERf7m9FR4IyJUmLgxfzDkRrKr4HUyD5TPPxfYVwSL
wYkxvkJw79RJvfu8ftfmuyUHJyNqoczjoHI5UiodSJgKBNWovEQk8gRCu6JWE7gRLu+8zbilJFJa
g9fkfamtqyqOeVsJOJeSwEZ1P/ypj0ggqz3NNvfEjiGLmqTroqEoos07N1NMPchYEYx/RUcgDhQP
yjic51eUcoFaI4VTdcKe+sKpNzGCc78B5xhEsZ4Wp2DrwDecRLywIPuIygI/jpAAjC/Y+FQexDPM
oyWGIGul11nW7OyuCrbMYcDxNG4XgUU9re+8fPs64dXBYZCujUirT+JHRiuu9P/kOaCFbURATzln
nu7Q/weNV/Sk9SzCZUa7dP1UR0pGC7Mw/YFb8Ye3d8pOyRnpAvBsT9AfBlArY6Y/2LGAe86OI/X8
5R9/VoC6cqi11Rt2AnhmAjQwlUjuuJIiXwT+T1Yp4LbqDffFZxs6KEUjTFYwfIGUCBjyu9gM4SeB
8jAwVIOaIsQbw9j/XWlxag8lAS0X3sXks+FJSFfJC95zFDlUl/4RNSPa8jLV/0V/zfmcTuGiEtdp
xm7c4Oh0nbQ89XHXNUziM8Y9zYcbQT5/DvTt4ffWXrM95fFOpn7YgpGa/cYPDDNn0usaIyO0vPZy
MciZa0rzaYyfWXbT7HTS+z3vsoy7HrQzt6by8geE4CYv7alXQkqC3WbLhw1ehy7ASgM3G9iVTdBk
Lww7Y5n5oR3QRC9Ui/3i0QZ23CKvEaPv02KZ6wRWstgzA6G3XoGzKCHSMo4EBUiB/sYIf72kAeOy
4vCQExMDGI/aT0cVgFLUjhfuQ1AYG8En5aMXLrtwgOX5kZeN9qVWsrlIIq0RAwjoFOJZV7/oN/v8
A2A5iqgkVCwvY5UtfgHjSHD68XWM9Hzdoms3BSKhZpAV6z5gISSWQlB7FCCJ8sac7iJYBqxcnu7s
zaIb3KrsRK38i2ShKCS0WGETFV2NuWOlJG3j636y46j9CO3d1las8akjPcxn2+S8GdnLVKM3s/93
Qdj4slGd38S5Ioa0JIcCKqG6GGlrmu0iSfPjNfK94t0tZ7NiV045qmaDzfEM+v80GIILzDN9DRPC
rwu2fD9NijtX/BgTI1dxrUVNKq/QAGxeZBbKOKJT2tv1cVKvTjKNQGA7ostefsZOI7MmAaKzo54J
WKrAMOlfgw6qTe6vVM4EF1YjEFbKbMebqYU4qOrAsWQDzJU0hjcnYMef6foQx/E6/R6633lMgrzN
D2+035aHBvCBQjBNid1PxYbm/zI6WkwBZGjASGY7bK3tNBH/0KQN69in4ggcG5Vyw19GAz9mE9Is
YOuTUe7tZD2sVQuP4QuohNmkYyxBxR647aRLgpq63zLGQCSPhsu0/sq4MuhZyPG4tcx6UPPgzp5A
9JFQcDxbUR+R6wyhMawM8K76mxz6zvXiLcCA/GX8PRLLIk2ZalVpe3Y7FYwIRJ8/6iEptwOJg/el
/RwuY+2VyUH31BTJqtpCxLCNWl7vmUEBhlGjl3OeArutuOnlTcgtMaV2HLIHYW32USTq65XKAX98
jf4sJCeFR7sNREVuCcs2oYjU1x6+MD16cHQ0n9PY+P5ovsJuDwbPaSxxtDT6CkZTGrujvE5RjDHZ
LIN1Z24N+85F5Np7eP6l61RFMXOG4lVbl//9gA0BM0CyHCpgUlcdL1QL2fjXMP8GlJ+Af8WoWkT8
+CVUFZhrRvdrRKfS0x9w79x1ad+6UsWhZlsXdNiCFApZj76AfU/2zUBTebsMLHB9NXkBCNylM2ag
UtRGyB+jYdJJN4fkovsR9EIhnR5E1Udq4C3Esy6GU0mB7JioEfTuJeOFhdiOObY8p4PKYOVlSphh
clUdcj1eYvsnA48XRVqeN+qFwxfDT9h9tZmPtf+1FQV8FYRukv0stpnandLJBIiM1Du64jsbn73Z
fPVyEyITuavZxJDkW8bX7bKftTTIFB7kEo4UE3IlpE04lGErogNvV6ImVUCGG1cg7Ak16TiizDMp
sScFVCJHHeaSTNOW9rtdsv79V4Va1jF/nkgwt4iTt4rvGvt/1U6MJihs6Wm9rLw1vU9Kb1U9zUZm
X7QDih2OI7Pefv8TYhU3L2W8Lcw5hM+gYu7xpk/+/fRd3y266ad7azcVqToN5aayiTO0WoTCFZSr
00VPRo6/0TApY+TO3dLZDcFTmWY9humpTGHgZPahtsIM7WFZGqFlKNhBOYJHb/NZVp3y1o8Av6Nd
bJSuZ40B5B+4POmUs2K3xNXxH8Zqv8NAFFaix985xPY3WKczqynSnABN9X6+NMD54QiyU2sjWOAi
YIjdEh2s2u8MOKr3HFZlIJGgIOFLbpcZhR4tF0xbw4rL4yf4i47ILeN7QMovYCyYSXrUe2euBdD+
bCDmPiTVeYbTaLeT05hSjaP6GUryO+SOAsyZNqh/gUAEfwWwPaOZaBJLrucMue3JcXnJWgg3iEeJ
S1JF3gQREu8mA/5bGJwSMkLaC+SAB0aoFh+zl3Bz9o0++aqIKj1rmDy9fT07+LXoDQyZFDaPCuQb
qhR+BRyucnvwqBWtZEJWr1vOARXkInWcVPJM5FFPBu82bCYonhClnAiLB1Fa72pS74dXWYbYMLfJ
o604WY5suOxMLjrT3J8o/ZPjoLYyt5Lv670VxSJhSnV3/zDoT6nME1lF37aESWJgum9/xiBQg/qO
yidtVNAFHJ2uFKjGnQVcABDMA9EuaMK8B2QOd3PhDoF4d5BC8UEykCVrurM3qCFoFeqCYQQn+xxo
mY3P/WnMVlPA+2sRfFFsyG7MWQtroo/p6Mlrvmo7vboJxT3lnPzb5SRN4FmGbpgVEK8zqhkp3Vir
aN3bjylxBymMR2uRAKar6v5FAHKkpqJ8mPl+HrytovQ4eadrWiO3xUgVoNODIBdkHH1qmUO5bO2+
nXEeU+amVd3a/rRmQ1VaLHvvK6aT/1gpWxFIwkvpmQUgEu1lPyaPKYbAGqIEe1BK0jYI17AWfX8Y
sogykucBIk72R8BVHPQzohDTyOTDjjxwmeDTG9DpLfEfXvzY3WDTu3BcvABiucTjLDI4SosobpJg
PHfstIR6TBQ5vp+SH2k3GGM61wU3Kqj1mztGFem2Tdd+pIRYc0zPbwGF0pdY7UsDxRzKnOEVBuhd
YFlFfXH5Hyqzv8NN24R42/mmCrmURxe8ibuKGaotxffhPMnb6Y6q1+fks59XU6epnPK/dUhh9ft/
6wYhGZW/RFALXTAJrAROVxZ8OVBEtr3e47SPIw2XI9Ahdo9honAh44lmD3qOPVbwWc3PmESga+cl
iLivA7wUb/od1PLOFF8tvBk/cxoyCy4acytse+J96DnEMBFZGLlXMAwcTcjLGm7p+2o+iB7mnXF8
hUpZzSd0Bjuc0awkq0QU6E4Pyf9fC0sdaUuSN2O5QB7FzfJOTBTv233k4SfJ0bfpFkv2z4Poky4x
lPbRPbRaz2gSoNjCkNCElIr975UNPsCYCEc3czg389QrOQH5+uMHz7DhbgtvFBZJeetaByCiEmNi
5L0LrJWzwcltb8w/8wxmGgVOFQ+6LgjxgUuq07+ljTtUYeYeKkBbDlst4/ziDLnnrL5zczPckKjT
zCSNgU+f2My2M6mW0z2XOk00kdQ234wFtnOs+SKL69p0uRzeSAcvXkhvJMRgmFks7Dw/Y7iMAbpD
ithgk/TJ/ziIIEbCYpmuQwmjzvQ97Jwuv1PeIstmG04UjA07QdFxkdvl2BNJp83fX4yKjhIGjk2S
cuVM6baRkRKp98NEuNc3Xsl2glHOR0AzqzLix9lLWuyC8gKz+feakNAWv4c0glqM8Yrz+QabC0I4
VgXOKnm43wF8o79E11HmD8nsq21lkLBfXrxoCwmpkK+9Yiy05KohrvO9XUNkgP1FqjwtC9OxzL0n
IJRSUd5Ixpe2xZUC3D5DuV7fY6l4yIGOMY1alxveAv24MvwN3HwlE7WpwisnmuP1R27YEB8nU+QW
E+mG55Ch5Rw87/SrRGdojTo3VgFdkMx92kbxhyUVbyq0ovmTB29qpecrxDfSbLr8nH9m+5JX7LxA
34fa7RO6VTV8x8RruJr+bJA938LLjUBXFROCtphwdB/2b8P+SAd+Op25sDIiqxnYsXHm20cmsy22
QKEiZQrJqEy6lZQHxw8qaanLK19lW8ui+JrjGPqaltt1on8j6tnrbSd51TTTSlkRfti/dOPkWdc5
em4if+fDrrtyYgXv1mWYQ1g6XHHlnyRcIZlAeHwHmvNRl4k9Vv1p2mhoDNevEw/ttuRoXoosKrmf
k5XZYHqrKgwsQ4ZT/Rb5HjxpF/tQyVOLezJHu3I/8UhyBrjomMj6cDw6MvwkOu4x60zFSDqTxdve
7x/i0mCGYqsE5Oy76C9Yixrh1GGDDT2PtxNUYzyxpmZFn50OBbyXNiDPQjCpJQym1shqjUhR5VUI
oDDqDQY4iLYDvQ6BF0iK1EayAVI9dahfXa1Ia2gO9x3WikO42BTfmySBPvqjyOf9LNyxTPRM0GHU
IYqxWoKFBkX+SavTb+vVXk4tJyG9etfhc7F7jOBnoadFlqM+nJ2L2ohp+gGK0oukYr9Tw0HBAQ4g
f7ss+PuI2v9b7js5B+RoDU5h5Fq91/gk7uOSUqVN1lcawAz/NyGGZL+y+2KvyLam4eEPJFxmUoFL
C1hnFtaThFgJdwbs7HjyBb22+3s3EmYaHZo7coan4DDVx2JgN+ynCmKvTy1XpwY1hgDkRMjrBIOy
Zk9hdmzo8VBiPe27Bx2IysSvI28KK4U9jpdzhzR9Pv+Q3EKS/zmVgSklxJ58JXpoIBEDiAW9jGwa
U6x8NUybKv3fiCRETKP6L8yQouOzxRNbe7uDDpmltRKwREMU9lvT0YGDVtRL97sho7VyfP+LwSAO
FjYcvRSh96VWPltLmu9f3KRH97ccUjU0HHOb2djq42aSOxvFJT3+km5goVJaGnQo0ivnF6zCrNS/
73PuYzqRBZ7r4so7qZSr9NTyWlDJmFw92ARlzT2bLl1VJikS5AMM8TeMG99P/bnRPNQEKXaOU+/9
MJHbiYx6uiXclqXmF25/3d+W7q9PcV/d5Rl7DoUZjua1oNDIK53hm1U8PbQ3d8c4/u4rB/ninKhF
Ae2XGOhJ/79je/DOfgBxyh5BctWS4tDGlSGccOgJsaqcerb2QVlq86iPhE2GTusjUBu20xpwa05D
DnQFb9MjGjdwVfv2dVm9zAsd5wDK7OiDsWx9ehdBxdsLhKP2UDpaMOre4ay+H/f68vFTMteBxloK
OFiastEei0Jjw+AsWdv8q/KjNnKL4UZaHUKcK5xn7+xT7ZG5CP5UFf7uaSqRcnoUq+pa/5OPKrEL
yrt1M3cmr3m56a34Iycz4YryqWaKPUrMbCjjUdQ28n0fnYV2b8hKioUnfqn2Q8Mwp5BwG2jReMlE
hNlILCePmUkzqgxYQh1vFuy2mtMQlcGcVRCE1a25cisAh9KTorh4yRbkLLyGakMMlCrwymFHA4cJ
hMsH4sYZVOMqZJJcAP8g9giHDS6C1VNp3uPzw4SynkMB0VSUTZNjukbiyqGdVrL4AEjm3caA05fz
ZhVTCcuT3WbRfvI+pEW6bJfHtN07szb6CpBOc86GAdeMdk2q1dMg80Y9i8sqFTNNlpDmnlYD2mNJ
IIQjX4cwxCiXTl522m5V9avcv297Hc9+YELVKza1vahLD2zEp+PjMrlx2HY8srXGH+yLxz9BvmfB
Lfo2B7O1DRYHXtimTtEhkMNKjn5GYjV0cIm9wOY3a2rhEzgd2gzwdujkRbfaxCQFiOpG146Pn/O3
lh0P0B56TCA7a3CQLqb1gOm/PwXqEATxZfcDVD8cReUrMESl4AufV2Pb4OD/54gx2q4zArYYMqrP
7zvw6FiNvkzptHwQEapLRfz5T/uvbtaEiBOmjc31Ug1Itx1RI4yFRNVrnnlWsiQoqk/2qZ4bY0kJ
SHcswCVVkxXTKmTWp5LA2MHGdoTjEbXF8dl9Dc+wqKSSCJG5D4EwzI5saZV35DgmilRv2IXBAp42
a+EJSeyblayP83L4Q+TMLcgBeWiOFui3/z5oKSHI9fHEU0rTK3r8fKVTzwZ5Pgu3fl+8Uk5x44Nl
z2IjZI8X9fOo4jKBsBhjXxDPyII+3pXCV+8607q6kQQD2Un93VibPkzs5bpSTDWXRvwpAT76OpvJ
bNLjk1UXHRu1irl0pba52L0m0fXSOUSW4t09fAzxXcBhH6typVAjQXOYThD+DBQVCGHDJ/91BDVn
sW0QRy9BqPh0TNTqHAUwjy9L6VBgimqs33NRAOAmp1TyybEuLG/fpK3r+oGhiGb5oKtTH/Hc3cZt
BlgFglLuaquZBKLFtXIf2A6JG+XpwIMNQqOV5SaZpse6K91HjMZvrgkDSaFj5iWrk0ZiN0GNL66K
IXrj/+1Rp4QEuRx2eZ5GxCztzsBsF5CVQ/5LGxfqEynlHFGj4UHQ0DOxxnQTWAyr+9T1jf5lE8UL
F48XGGtUlTRooOKigNpFkZxrdvUI4ZxlLI+ie1hZUWaMHs9mZh6RMh4GLN4+7md0DBKLLoJKxyBy
kV7meaED1Se/yCyxNnwYVgoWr6pYTX7uyN/oqf40Ml43MIMqytOs8J7T+v0RGDdpMg0JaDvTbnFI
MckTNoV1ahrkByahoHEX2iuP0EjIxoRcQiVKc7EY/clWNzRtErK8ABtaFPMpECygpVO9oGzn33d1
Tcn4IrZ3um+r5qaR6t5vIbrAzTGDWEsHIJQXUxZER5a2qVT9LzKKeRNvh7Q4N85LmYnlacK+B1+a
f8vuiG0znAtlXogjys+Ma9e9jZvygLBIE7tW/Q/Cb6VLDHNmee7juk4koYvY4DjoCrxOusPKU78b
+rCkm61/uisdmqVVt3vD2/O3q2W8KAB4mSxDo3uIQI6CNV/7skc+RpyzkAz2k1R0rWonoaLvmBgm
Nhv4vgXC65EH7ExGZQjf6+GY2TZZYjxKdRc2WEPxGAMjZRAs909hRwxlgCzCen0UOZHAx8gQgI8l
U+fmqtF9Bjftrg2rGTw3OrnuQhVHwRTNQPKSxIwOHZyjFUBtjmN79p1Z1GCnux/Y9S6Af0mHbQKU
TVAe+WCiZZKJHTQjW32RM1f6NIqIgsJW/EkbiuIGeN06snn42i6G0Q7EhDAVqnD7ODEtqcI5q9Fh
g8rfmI/WxItFJ24XHayTULcmUfx0/GJ6oyGKsX/5uOvIFBXgUcZrvyFG9oiBu3SUZrf2VRcdMoJy
mqY/Akwff5GpMbN8BXDo/CEueAgxBmc3EjW8ToEby3OjrPu/pxb1tr9vIPH1NEogn/AWgwxLD6Pz
MjnWWYEBHPedmX0Nqa8Z2xZgSR+EX05viSi/IU3YU+DhrfdEA/2AQ3MHW5+20xtxLTEFMulPzDh0
/zc8bqmx9queosw53p6fMknwsCCF9gcfoAAr6uHHC5FG/y/pvLqRvtc/AJAO0+i74kI0qgrkJ0tv
Kq9LMQw2UPz2wesi+m5FYszgduA4THnsrW993ajWIpj3rH/lSi6iSJL/l5i3tcImEg1wiYg4PpJL
/Vvr2lpe8a/WhfFKKR7LONjnK4/DZPydcR30uL2XufmSDVugzlE91GH+un+Xz3JHI2Le6BG+khho
lx6Lc2PmcNjGxm2uaaJP8VcjP/Too+aYpC+2M2Os3Zy6jmFA4pLlv+Tkn8UeVPnoNghhLoD6Hz+Y
wv383WRwAtJY7+NwK2tPaAbYQpaw9gAufCfSe8oXLTgQ90ET0ntmGw+MVfJtoA/TbZtwv6h4Jdu3
s5aVeSKIfCaEV9t/5TUGpd/bXV+PHgnjZ+EnLcZ9HBngWJqC5i/UGDL/LiQyAjqI+QwnQR7SRFh2
SNQqCxl/DLKOJ+1kYZXyIihQqkAHMGp6NwOyQ+quW5E4qkqHXjqnDAb2HtUuiOAPr7Ov1lya4/hj
2vbM0qA7Gx1W/WfgQwIRqEb6TqIEOQhpi6EIuQ75AHT5UNHBMpR30JcAMwG2uhLZXxwTZl4/WB9l
pp3vLPXs03BNujTBsvwcrmf/3QPL8VreboUV4dmvDW8PqNeHvBzMWvlYy648jxW+As8Hz269Xgio
yQ112X7lFOE36kM3qkViTBZuaKlcBD27B7mIWkS63NT90Fcp7Ci305bGcvIDZPquUiKsXETm8NW3
qf3/t4hykH5ANjB8CTSfJf16mZz9yN6rK8xFFohYjcxqy08VGMHacBvZSrWo5Sc1IQMHj+kvjgcr
BwDcqjDbvHUdL9y1NNn+BdBZJkNaQImt/6Lt23EWLUTSTLj+bAclqYptOYcbMU0dQEyiHgAnFr8r
+p5J/ckZeCrOZ0jyxgoxs8BhWIqjqt1tCpviCqNMuX2l/blEqy1vWE9xKvo+vStQq8Pn0cfN985U
nR3GUNESH/VOud/2hkr3Q+jJiTW7cfF7yrJPpybftwfPi9ifSHj+OyuNou8VNYbsUIzoUkrnMIDE
oRoT/8uEYJ8zIWs64S+Ft9C+wa6AesJPvA4VXx5k64RDhBWFUqTM7Y87xxgZxqNqpJLNYTIY05HK
R7GJcWD/CAkmvPI6cJwZz2MYU7M2PkQL60YZb+4QoF4Jsr7+llSr2lvcqHOieqG+TZ3MYWUPBpsb
34skGoWgWfxOffq0R0PIFL+zwX6ShTj241f2CHkjBSiHkg3aTJI0o5sNHPbCCLYCIMWjfZPjwxI+
UkF2yEnIOUkn4vsxUVw6nsEtqnTjYDYem/Y7j01TQx7zzwRZY8mN3vyC66euE8qu3FoYZmp0YeOt
KxZbrAWVA7Lz7vXLaa2YrUpuBLhBi5zM146u4EzDBuBa6S3ATbVWnlo1I4ULS7vRa5+Z01ublK4/
omDyXpcAfaTt3dgd+j9FBJ15PnfGfS4pu4iwA0nRjqBqxH+vY46KNn4CnHBLX9frWApbivan5iTJ
s8HvJisk//wykiPJchsm01CP4x5JgBVPjHA73kH7ER/UmArAzpuJ7EvlqnHSmiefUb3ZuJzYw0B8
2cBSd02bm66B/yL+KRK+AoR22oTTijFlpNqW+WEB2rRwt5pQYOdo6zREyjtv7ROfA66BDs4NEzcL
3RNvRDBFuUWGTm12T2fC/gvTVCOnnQYe6K/WNTg6Tq0IH90YLVUWVXAn48bZKiYNlwZKWR5DFUMy
uwZZO/8jjH08pUAYIaZk72yRJNKAlk09Dgzt6uyMLHdEMTtmbW4vaNLtFmWXcVETpVbbj8VAJ3ga
0NHh/PKWBRRYQiT8XznsP9UeYHMs5jucqfB/wNYI/cNpZK4oW7jnfSV10oDBVtQ/tcSwNbZSRFcv
9uj0zHVue33ZP7vFu+NS7KyJ/blzLsmOnHSg7FjuXN1Mlty6d27zLhLIM0xMPcofrlNMJFtYCyTA
SxR3CDiqaAFrEHGt5ZPWULe5yKwxrXxzD/6V3uaFydWhhIKYzyW83HlxXeZOPX9gEttcBKJHR41d
D5tML43xgpJMWD3zJ3YprGVrMDmlfsvwS6aE66YJgqFypfqqfUCeZJBbeoCgSSN0yzp3IlxmbfsC
2K84fgpybwYDoO+FFFf2x8bsNd8hy24Pjhv9MB9hCt7LbmKr0/lpHEJtbEqcZseNrHnOkUn5RNDB
n+5oJ9TZ7/XiHMSeUjOMZ40AGZe5+p7pUTjK5WPRPZ9dhGL8b79dFrUR4g7Dtgo3db16VV3YVggO
Ttb0c41pXtaeiTJkTeOgau8/wTlKT/yecMqfnypoxNxncYw+VlY7Cb8FP2wJI7zFRW+w9iaphkqp
BfxDzjeC3ddB/8VOBrlViBktYAgDfsTI1YJkazGgEXxjU3kstqMIaNrt0mIuWhxJ53a6IKmLUALw
2ApEzBFfINucOKPTqtyLzkP+UpDJOQa/4jGpmO8mSqGG+zUCZqGu33gKmf2RFTP8riub4Cwq/Kg7
lLJWihJXMZriC3VpKjir3XRcz4ixYAoKcXIFGyGkXattN8JEI1mt4wWmXHrW4yVuvLkQCFgv29bn
NyIYR2mMqG5c7CDCuGKjv1a9HRrIcyrK9qIvL+aEtBXexVbhIaRsC5AMzKMDDE/HA0SePPb1NUxP
XUrU9G8Y2TQbrlAcQXPWV6UvMLoRLz9IlCrsdvldQVlz8WK/zDDAB02AhL0fDsAuNQpzw+4cY4xA
Esa2t03+soH+UhvV6TeNDmJ+oj9oS+a9jWHZS+hEROZPuUC9Y9Z0Whr/FBJzuhp7/HkRiqcd2jt2
0kDwEZqsFhY1RPlCJhFJcBHcqubWYi8hLbiKnRglf9jTkUrdJ0qvojTgg315is9iCAHGBeh/WO7L
RMuj1JGCVw5h8QbnO6iG6OdW8ODItxB/cIpINNW/So3lax6L7yLoOFwvpbpolwp1HoW99+GK8/Va
8d/sXKeYyZAFgV+SSlT6RiBoqH+yAhpoHnBsz8RQL+lsUZlAWr8KH6gO4fZpeEm3D8lyGoHEB359
uG9+YT+Ktyt5IliC8UPIrWKJF3d9ydSjr98GtYFMPSXVRdUf4blx/ovnwWuLVvWKdprclcQrwc+J
UXpy3lLRTuv59zHqF33jBwnJfB9tdXfSRW+642hvEFVpjLXA8zNlm+DTIqfeql8Dn/KdUdcFa4eP
axCs50PPleKi2XJsUrnAG+mGP1BrHZFYFTgoy8LE4z9gexiu2/iMenbsYOEyayyY1z0F1w/XjPIR
Qo3aMc0J2jmWoXW/J82y1HtPlbAGMz8PDYBWWNVkOS7jhbCjzfSdy2GfPccn04E21Zx3euCKVVyv
gLhblNi8CS711gWOwr3XkZsqkgmY9YBXwKsY21Rt4EStTUp1WoJJRhTuoZwZdTXZteOLKzPWaPzf
ikug6iNuZp6V/mOybhsRWOJOBTY0JYwjeMlnaVLKja/c9sYE+xCIuJVsjYQXYLyNToy+hB9ZWTCA
VaoRuUbLJ1DhbwrA5UlYkClf3jLMBMqJEhJ7w/FROFghAhn4bPdz4pLJs7NbjBfw/eKgHvD9XAZ2
YkcSJMelhmwzGGTiXRpG37KJpHdNUBrYwGQZlAUL9oMXwXq34i8Y0sduGRD51g7BzePTE1F0rJtF
AdfVYB4MgILG7KcfoxbvjR79wmwzU9mDxB/5nhbYj3krHZ/Ssu0VWgbe6Y/buhfvTW3ts97C7hvb
394F32qOpYM2c+8eo7g1AcmV1dNyg0iVOc9fsELLjd9H5mPdzkgkXinswnYJ7YZLo6jFUClbylCH
7OWqioiF90ogtDMaoWi4p5MZ4Pvk6uof8vEBtHy1ohjvtDE5KKa9vl0UyVDro3UKmvOv+Cm0tNz6
Ns2Hkeg7saORZ2PXf3x8DYFKWJbPLPRv+hE/QJGUAjBZ+pepWUMCWx+IkUCXuOkD9M5i0HDCsOGf
J/H/5hS88utnui/lsEgdiiVGbb1sZgknzqAJ/L0tr2YbLqb4nBrXhlc9dHxCePKpS23vMfKFh6Dk
lGD/Dohhzz9Ys1e52p3tjEZmhVFq7Y4oYOUwqkh6G59qDQ+odI5UlRRWis5jVkeueBODWYub7Uj1
hNPtONnzGx6RiSn9LKPIJNxmPW2WOEqTbCvRdpktPwOLjWqpFoqnZZcVRyvMLvb+kOVimQvAUTbM
B+zrWLbKXHFjgvNIAsm3nMqYHR+lFFpKHlm+63Omlg9VYAB6VMna2w9sf1EL7MhwR+s18xPHWtj0
kDd7r4TT6PClxgtuuRqxDjtOqp/rWymgwjDPpfygWTw0HIbGulBH8Xc7zYkih5nnisEVhRyCNCif
984ns4Bbp9XskXFct/cl+vipoIQyb3fKE0xv37JBtILfQ2nN42EuIliRnH5YZiwyCEcG/J6sDAg/
sfuQ/4C6LlxEwWbectbQVnJ2iikAK10GV13BvTTVjDrr2b7DqYT7acDPYFJyovo7FEH+UhZfEq/B
ZMwcfx06kRiM/ARyU2NUGewRpVCDOhKbji6lqQZjJiCI6WRdMXPFeRObgZ8bErVJl3kNshZdPhUg
wwCXJDasWWbggHqtNfKeMlZJ242ZZLLrBh5bJhdXEqy6bZRgfmIxPoMUiOCWw+z+R80b9No9+jEH
g6M5SPhJ006zOCSqauoZnL5b65polo0TX1YNuA87FUUU6tPBObTBPFgzLbhP5y4W0VOGVey0WPRj
nfSk1Y7hY8M1x5Zza/bZcj5KIth6IVbLPNOwlQ7MhuAaw+cTsHG21ePruhBkhXbuIBXhKOmERj1Z
Jb5d6HgZOv28aPrQIiE1YsijD4na9Gm8Srg+uOtG7lfgNvpjDUBADblJnicfbZaEokjqWZCh73xO
/EASMC1tUEuqLf0A9TJl/iNyQBmWbJCd9nj8QDV3T6F/gOU0qLOWwly2rS/YrEVToTq8keclbfCz
PSfIZjLREsQ6RdifzWqXjzdj9sYb6+ouQKj0XpFljOWSY2gdF9tBJ52mcreuQVomKmPs1KSCZhvh
FLlP6eJUSzjaYRDVkGkTokBA2v3ljxaRxYxY+MTs4fSYvtaQkjJ6LnBewvmXktRpJX17zTvoNvsq
L+vEXRaFjQFRcRxvVT7wPaOOFigpyMwnZFPicdi/OFpRad8Bkl3Hsyu+0gg531wuEjFJ5sjO8g58
+HVzIzMk0AkV+6WZeKqXLX/o22bvhUXax6q7zDkw/4q3IpKqcFX6a80FcZYX59W5bDng2Zg+JPmh
vK1JHRwkJ9GKqab+Wap/OImliVCXWhLxgV5ROnDWoivxyTjyDb+TVvcqhon0rO/HbdQZOfPBNOpj
Z/lrKAswqeQRJy5ypDNpe4RYhcqL4uQMIxB1kGTplNIoKlAhzQ/eiVFcRvsErsowdWVbHDxe7ZoZ
EjKkUPF5anIHyC+KuaftqIEIdsmZTQ7l0bZyd4mgQ3dWwQ0exeE7P/+OwQAWgtq0ODxxkaG8/NTR
WCfwyujuUPNLrsA7VkmeRTv7Euzj9m4ZyCAmnUBHMqRnnPwxs6FOy5woT0zS3Fs3TGKBUGv895v9
ayffGxIPPkY/DmH/ISxnJC0qn//NQm+QmG/YlgymZ2gnL0G/2o436SL21I6ACLd4bXZQrgx6/6ly
HZtPBtTLDcbRUg7df4SwEZC1HGgt+ZkqV+rx9W5JJKh4utEmgW9LP0+PLRDlMrZkSC4bBH4JkDMQ
5koDseO2TQm8MdlogYHQZzAGrZA4o/st2MUFEgQAHjvNg1OrToxNtnD0oZ9dt+hbzhMbDimJ5xpo
jVxmM5RVXyo8EmKm65dcefcqGw/pvRjRWcrisMEuO/UwNz+KqtNI4kCR9n7ve0Z6txkN+hNqCIM/
iT85gBGV7P+Cf6WJbf4jEyGcOxwBrCF+xB5wLGvn3CWgxlrpwmefUYtN4LyG5qh2IKt2JS+/hCV3
mrMMlsfQbEafgVa8gbbOf8+mfW72du5KyrIsTtBl+yp+iNokwqud3PGF7bWpgVvVe676ilKup+3z
ESvWchZutZpGw48If9Rdv/Uch6k1Hh6fZtEice/6Eyz+6nu1yYw+yHQXYww3lqWlLJPBDjE9oq6c
7lGiAGS9YSuWRCJ8sLHaeRr9fIGqsLNFYDifmcN+KcYMhbN7RUeebDwDKSQQgUjpKMt117eJKnzE
ufJRC671jGkuQhgizHUGZSVYcqe8HxNxQXMFA8Egekh/50pJzjAi1gfR5mLv8+au3nE82Rdw/eRL
9vh14Gf+40athIIDem9ibeH2t2QI2QB5x7qEKhqoRHSqRQblbbqBOtgim2rYV40knJJPEoK3AZoY
FyG9UXmFQ5dqIBWDGKMP3MWhQI6bnWBpm071EiVAJ7g2QBEFuo1TIDb6cVwq2q1rzP6qN3+dWSGJ
tx7KmaziVVY+zZO4vXEZmaY1pNoDVa1YHsj3wXObpPUsDTHc9noxLRLc8rOE4xA01Md4trvH2Fij
ysK/gUx2IJuaWZt5RCZn+umXlnq3U/NZYbLjOWZ5EEqV1u1cLGprua04SC3GFXabYi5o7e0PqvPE
1aYYUDr5ZdQXpk6ov5JH7uCzX6fa/jsL7w891bMhWEK302/yC2j4VzON8Rao/4Dqv4OG7y2ch1/z
BvXCKqI9nKV/GcJudvuOWH6F1HnT/Li3M7rNU9HQZsLzCoN9NA8tXLgVFAeRmPf+u7oLqqsyFP2f
Q2Add0mCBB7o7x+Yyj2gh9j2ZWOqB8VEXLE4xqrbK0qKtYxzbghQVj1dwn9APQyGw0ELlQcf7v2o
iQdqFEPiZE1FzTajilDfLDObfiFChRbeDzSGtLsKEIDXfECopct8WK8UF3t1T9NJpINqISDZAfQP
DE+4SYMXMGZtVtbPk0sYYI5A5oE4xd+4V4DmhPozr7L3px9eCRit51MpWrkrTKuem15zSLXdZcqL
xelNN2tpbJ8gH0OOG0cxSNsLyDJzupfXDRw47YM6JdD6ewSQr/VcZQ12D5//N+CtIGgsP63Bxi1s
e9wjm6e2yL35HT4rFW63bZP7f58BOig963ArpbGmWMnoCsYLQNmN2ypKGEmObf2XSTaLeHlF+So4
4I9mF8H7H3EBn9k2cQLbvVSWPjyGNYemCk5nf2dOOC81N0e1/SnBMUE2//3uJ+sPZfP0BU7viVFx
Czs9dNmBq0x1bt7Htq5lWZSAJf4T2O0Lqx20waTyCPfYlc9h6QKEz+q5myrq74s3KtUwgG6XxhLo
CxEc/ra/2my8k0dml7mQdkiqYnkn4Bdf2a9lQm6mMdggRLPlkbch+ddmnXLH3yyMuxIodgfFPZjB
jnVidmQwQqXqqbvf3uIBKZS8wFe2DtFI30zoyUwMBC7GRWDGX4fqOZ4bD0HN0Ad4m1ST+/WoyygW
h/VVspAozuv+eFmQTwuIMkYKw/z/5A1r1QW3Ve5bfKNaDN8nOGQK89a/41wsN0ozp0PPgKx7abmL
SMwi7ct4iG6FfwRZ+yOm7PU1dCN5s9XkR6tqx3igZqgaoIOStrOHiH5Lbz7ja2Zp1NPJCHZ9Te8a
vjn423TORcNvSUT4BaAywUqvQVQWRaDEpgh8EnR1oDGFrP+PmnPlL75VIeGJFYmouaMx02fOLNRJ
2J3zmwufkN/CMSFgo5ItSBqz2esjC3SUNPubcxPwqJG4k9+vE5tYglXKOizgrOhHAh+nZXewmvyz
80JM16xWPYv24EZ4YksI7C2/BqkE+7wqYvDQ0sy4PmdT+1M9Li3YBYhSgeCNM6uPxo7kTaqczh9t
sQMSAEaEIo6GMhG6FnPLH0U89Jni+jWeVpWfpdgVa+yFVmntZGvqRKgU/Md3VBaeETNnuHSkkZkB
q4kKkYPpViWbHq7aLD4Mu6CKIC4RC/EIMpRaTjmzcyvUP4wYnxf0M6TGWOVmt1f2heueq26KKPuq
qLE/dGuorENBKp5973Lt/7eRye5fiAJfLJBP4YMlzipJ3Q/G5VNy8fZBSU2ZzjdFMQdOCtKP/xut
IVRBGe52XdMXDjObukcoyUDLe0EGSd5tQyBO8ii/B1bC6JTS5PIxPt8NrGBTGpDajPPzYu3WAdkR
D3q7qbke+t957bcWnbc2Z+Tt04v/1cg2RpXaO/wHiHSI9J3mfpT4EZQNqluzza8jlcx8WV6ornUo
ldorUlms7rl+VGI+vbk0Jd/F8hNIpcwDblcvRmxelJjhXONrrVr0glMXoBFLDh/K6conWx/3lTXF
4D1Z0re/BlG9+0hJYXQM3OrYxEWUCyeNHyJvF186XIpmYz2GAhkgFXdSZ8Z2E09yRdNbVg2Y21w5
AftYtL4fo3sFahUWH5EKoddlrAWvCQiTKahfZu8BI/0BgQyq+7o4ouMSYbCmDXeNND2j4toXF8NG
LmFrKRjr0KDVTrMDXRLLOiw/WwE1TnuhvVrePY7uXIUQOl5fZMlK2OYAKa31wKhjjl12Cp9+DZdq
S8odOJcYkVLy6VNFM1S36PdFQfI1Dizp6KuKrm/De83fGGHpMwhFksR+xGS52eUFq2AuHIZ8kpR5
8EA+dGCDg8iOjAUKx8l9vI6YVxo62rM9dEVyRYFwu5UTI84t2X6YUnw005dzlyc3YHicJXAdkmh4
lDaK35IQsGmS20fSZjn+m2GVeH8tERUTYjjkd35rRbM4DsBUcoKBA9zSBlH2J6kkTweBYbLGjNUw
zO3bAlHY+HrFRyu8s5BScEI/XQsiQLVCt2hdriqH1wRyZfM1ge7oAhwi29kxmV0RhkC6bE/5PbjD
H/AH4s6mrH7KfFWWoMO5GPfwV6fMgvg0juXIWZVSDZ6PKmYcH2E574J8NScFhNZPW5zArsKgX8vF
lX3uLmymmTQ2E3+i+Har2gn+vD/RBTkrB7iJA5P49jEaXgV41NxGGTOGOjSgUSWOtqIfngeuke6x
T6o4Y0/1ZztRETwAaJS/Uv7vQD7zSTt9LbhkmSWz/vfFH/Mc9OHcnE8g5Xsm00d/W+SfYcx2zOgf
eeM0ABqCNEligpLQoXnRd+65xClInq6vuVNvUZV3vfeXwm7+SmbO7OE++sFYb3494EhkoB+NP1VW
q91LEsiBDgfOFVXF9zp3zS942vnKYrnnxYlLrHU467PVLudwzBtZCnqu+4vARVZvjfc86pKR7K++
57md+lz19HEGvdTqDzZLDs6tmp1ti1h+PqWDaaHfKxG3TQpnC15JYHIePb3uqIyErzz2LAV5vffF
Pa3Ck5ZhnHqsY9jUBT0smUpBI24LBxiVjjRkO9zUUOCNPS+YJVmuLGbebhVKQ5pk036qeO0Hl4st
9WBzc242vrSUbEPm+w7sgfBwQH4j1lmrSkaZsc43MbORM/rcP3veVS4B0lnZ46ZvLVERaluk5mJf
0o7vz8334F/SofNhYzWL1+bIof2I6w1g+I2sG766e3Po0sXycS6EqOkY3lK1rbzIckoLPFhawadg
Zqc8t5JCj/YfJxZCPl6/iZc5MEY+B0z4Ozp5CJxANu+KnMxBwfmnXz2jRycokjxRfMumAz0QLdXQ
65vU9QEPRdS+b3rJmncoCdl1LA7x9MIv3tcwAFn5N25s+fByRzInjd+8lMGek56MbRXSSqxdnIaM
9YKHB2iQiJL/KWH73Bou+TpX6ltkXCJxnon6qcJUCElcPLLWq/vrX433zjevHh4d9fa1ukh28VBH
OEsWy4MzkfN+p/DWRwMJIkdpvoUecTgMJhkBoRrad5zjaQlrc8uAlOxtrgohH0vSqDxpysXocGty
IdZA6S2FOS5J2xv+f7hTrbAe06CohD0wgSk1kv6j71crOOXXWaSD/OFwRSnrhrrQIPfgUIeG/n/T
SmBxF9s/kMnAlw4ApbG04ImjRRistjM+Tt8cA3MaAQibn4ua0GToIaUUqv2zfLlbMUOjd7x8PiUQ
lH5mICahuidcdNA6UcYS2pkcfAJLz0kT7TeUVOIAbqCcNp79ciBKrk+rB5ng56HIu7pUy5IRtxuH
V4TpKKIVuq8mcmDmkG8gmR5foRVexB4Ot7F9tjldeIar5jKukvv63x7fBobkfY/jLPqpXDh4D5f+
KTHGFdjKsQ9x5CQiNfIBhHpVTW/rcg7ZQUsfsKodXSHpyEzvI2QSTffEZ1+tSO40o8idL7fkYipq
kM8Pn56X9CrwoHmcVJguDyI4OXJTWpe+tquS3wSoMGg89T9s/bXOA/LWmrELw0GOIA1nZBkPmEMr
qDL57JwwaZTuS7MmW2VKTrhVmtzP0i+ytkjieNyr9dLnBbmVHNpmEitr9Xy8RYthfr3dIQQRlZhc
ehd7u5Hrz+4/1M5FvRF+PfoDJepev3o6Zn1BT/90UQO2e2vzUPFhul75EwZm/8/3809Cwkyligjn
K7UzWpaTU/PywpAzhQqFdILxLgJryKqqQK7qoAme2MFQf04e9bR4hzozOJ9Q6/zEE83didDjX1Kj
oL5Cuwlezyo827/CqetGjzeNC7vxgYTkCveRquzD0zLCit30FtOCTlKdbKq6AtuZ7UG4jBumDV+Q
jt3hFKt+R3KaYiPkExJMZafkNTZoEUs2WED/h3fMU0Qwgdr6F3FaA/2vTcPOl2l6G0TvyyTejPXl
OQ5s7l14ArhjOZ/d3hzyO+Tkgj9qCfQtJEmq4QlS6j66j1sVBC72/06a0pVQO6fIjqXms7g6PiyA
SSw0kSyDzMpwvakIAO4Qo7nyu9aVWWxqnQHpvUOJb6DonOC2y7/BCVJiU16Y0CZnm6nmeR5lSDSQ
Z6OGjqocHvNb/cviZFUL3i3c3Y20FGDjzx7EbuRvb+N2T+yC5FY6QbNm2q6AIA0Wmq4BnGxEJT41
y3GPl8RfQQYOCfm3Aev3dAj557A7XHELqGgN2i5WfYIU/9ZAZfBKIjAGzJ3PwqOpxXgrqabINxGA
rrMcwZxMMEqJDr4tPmeM4sOgZkqecZvdcrH7CuZY7MBCaEAMRS/2eThbL0dAbwJrSzpV2A3/tcXi
SAzDpEXaqUMTNJ6M0NPxSI59mXGO2mqaWWNQXdHZ9GOMk3mlX0X3Vc3aT8cEGLvZkDtoGz05NzIQ
ct4Sgw5GcqWKVvHXAw2kWxNRtpeWb7FrY+AXuajtA6oavWwaJEDhRpBFZYGh15WAaxfzpNAd7dap
xJWNBsh9pJgpDVK7SOks++5pFKzgdP8Vi/+jYgMI4qO2W9FLFZejM4FJRrvJf/BD4Shkx/eNlK5m
SIIISrOBVxz3LnD6uKj5owVX0mVAtN6GbH2oiTTo4vyNoTttLLmoHwfUYboVdkWQFZVKLiwxXcdA
PcqVsofFLxDDb908zEwQQh9tIwfThXmbbVbgaRoQgdJ4oVWu11BM3IuKt82B3PJL6yen5QtxORS9
FntEDKoguAw26aKGRVGlmHDG3E06N3Fjm/LY49gLus5y0jbIXIUczSLB1vQVoYhPbUOud81UNyHL
2SgFbdOAQhW4zRQcmiQiXuoeB82ATtsuJRiTPh4YBOCRNSxfkzIFFNlAexGtVjmiRHBxqCSefkL+
cKuRJnpZq5sl4S1a3fkhtlrUrkwPQOLW0iaKUup05WHTnrAp23mBr4463wbv6FSdCN71EP0je/XQ
+WWGmI1o4yIBHh64qJBfuEiJkIikKT43A3ejfhYgYSUCczFcyOr7mMcPwLfs+UphHKLHXKz1i30t
5W4N11+GUUt1LZxvTAcRyO4A3mdBOTUqMa5vxkKLFqUlac6Hj8wLczohDaU1MI1R1f07zCl91nng
2ZJNpObqJVypphJ7/PxJgy/mHY/pyqsxMe2Mlvy5sJVQP2GaojpGsMxRMFiyClqz44pzMcSXSESW
gY4NFuRQFknIl3Q+LRHbbeHMChNNWsIaLDk8UeKWm0o9CmSg8QsQqu6Ytznghcw5TdEXBxp9Sh+e
zcEwOMFqbC6KsJP246Wxumhd3e2EvDFUjVOOpYDifb1f1qrL9YyrEpS5FAgS/ATEpJ+KsOY9ZAus
nfNxLWRE1xk2h/oIy1T0RMRLIbOVK0yUajCFRcbwXepD8eSoiGmYeRfKY3f3LhtmPljYgFxj/XfW
Zp1uEL+58326tAKN6tNF7ZxTsDoJYz8dp8lfu4yyULmnUZyCpOjDsrMyjcldX3Q5I+rJh5dG9PN3
9PMlNc1S3bg2CVS7bHM3m/FEsY+ZK6/iUWFWgPdr7gemZwbPAsH80cdqjWIwXcbuoFKLa2vDc1Uf
NdqGBTKICHkFD8q9SWn9JUsMed7k38aTzIyEGsS5bh6cnL6p9bbWa/pLnuEoPTrUGABZPOnkSixL
g6mBDXEBN6RPRa03ntB9qJYkE9M2q307f2vwRSb+xIaUFOA3OtlPOREGG/YOtm19IJDkr8OWEIdo
/3FVf7Wdh1DTofQkJg5R6mtWH6BCN38KGAMmBG4sx5Or7V5zmOOrnHJNj3+ZbFSbM/YUt8tbikY/
ObWfKaZPqRd17PmP8jebx4OrWd5QiGr/ayVtvtxXTcvG2yXF7qV+BvS8tb4UlkzSCQP7+J6DUgMC
KQ5VNt1CSLPjkw5rnsByOZ5u/OdvQlceu1DIBmdCrRr32Fu7tRibeZl9OavWA4+bLDKaA5ZlaFGD
fDswxr5T91u4LyS/GafmFf+JpMf6LpvlKL8QVRmkQMhGXx93Hi2xtpKK+DLXWTQD16vfTAckRXST
tc47groz2Rm1RhO13xLayPTpm+4S3aNf3d+DKMn9eP2cNOADd/KDOPteg+0lCRDxMGN/JXV82J6Q
HT6CdPVTYW8XIvCgko/dUT6Q8YIh/vEA33H6kFg99jl2WlJEWlPrW5U1VjIj5yuA2PpAMHcdOoNM
jXSz5/XXC0NdsHpjGFyJYO1WcZ/B1HPMyzoPyoiHxDI70S2KqXI2kmLP6AOMo8YAWr5NaRxCDrMH
TLmKmK5SiT95tlr5/bl1VgMl+OmWKj7muphb9qRqjh2RH/35xwIOywoLrs9YMlsIkKBD2k+vvoEl
MFuNgsE6fO+1TQz8aeBJoSWUXJrvvkwMMnAAn6aSrR1JEUtZKRZqjXWOxpPMQwjlZk3DICF/QBAB
3+oPW9U2RXZVOkxYKJbDVV2oEBGphXg+OqOhlXHXnYTYMAh18IpVaiYH4arPHn4NrdNLCZMtLQkZ
pCFEh28c4Ze3fA9304xxZKSL6SC/wgZWiOc93jFEjyXwLchl2zdHDQK90Cq+zVQ47kpcWnOtgx/G
wsBlLrN5a452YIcnjEOjVEsxyJ/dD+MVNp+c0R5+XkdVzXDOsiDhTPVwj50TglHEm/T2FGoGtdqu
wptG0IpGO9f0Jvj5rZ32HJpUW0OhOtyGoRue6d54jV8Yp1H7cRR1ybdtHGpI2CYS8hADeTDOK2Sd
Dy+NG8BhnAhrA9quwwf+WlLE1b+nXXYvmjgHnc6McLmLtUh6xYUpQqfKAmA0s7Z0EzG3F3dsSfnt
Raf+4ZuXbU3G/l6YuEAyvlLczJeezN6u3U9ccEEEPRKTJFjDjrAvaZDrwk7YWwb185ajz8s1N8Aw
lNgqSQnsqgvOxdL7PT3L5YSZUOGCBGxfxNf1imf6bLGcUf5MvGDvi+inhr5zEYynh0RP5IV1naX+
JB78boNkn/DHsENr9kkV5OZEdXdXgMWMOXvC/gjHPrSd90BetTNl6e7sN7LStzo9fwCwRY9N59dx
BKCLPANEObe1SKOjs3wgqnCxY6eT9gBExiPj95CcaaGyol0PdVK0DcEzWvdZXK6BZjONbPJ7jAPz
1/YQZWlwORRHpylK2EjSMzwkDMWNhCcmi0Ee457ukaF3AINExK9opd5p0r6maEDFiARJ306f5CVJ
RGkWqjzvzskRS7a3B7Wjq/6k8Ot2sUJ5PEBncznEcQ74Gsab8kRaeWS0TRlp7niLVrC9mZiV3nnq
+IqI1dMvcNEDS7VNGiOGPLcLQvwUSUQqqtciyU/YGffjW2cssdLEHxpSWk++OBOUgOjx4nLabiKT
cgvd0ALKQyA1zN75E6A4KYbc5rQ1EbIA8G5XjRIIm3di2cA+oe+lcACyu2m6zeG36DC+HKHabjLE
G1WMe9UWeMGuTa8WYbW5ir/wDWZVePaskuV9WyaSf8oLvNfnGT/LpzxnSkf5z/A1Vx8nOll9L1Jw
u7BQd4yIQEwtvF+kI/9/U9PtFTwK3jJLXxYtCZcjMHz+CJ6tJHBP6m/jVpUku+L3LMVn/RjQtZ5k
1SjN0sqtyA4ILLPyPQbwsHGHbU+c+MbWv2sZCJhfJPmBDLUYIX0B/dDuGvLIhw7SekNFC8sXMoNh
zDgPz8H1Sh8i9qNZ/mNO/emATG/RpGYy+JtMvj7wbKxOT6Rv5w/a9pFXOjFNz1S1/zDLWSyikfId
tp3yx8s1UF9ewUtUM7JuYm8U9Qo5EGhEbnomxEGBNTd+VlX4Ja+3+ZcCi9pCpXnQybcfDK7hxFw0
Gtq1EAOd7CrnDblVYVaiQIBZqVZ93QOPW25RoCKd5GIji3d2x30cZ8tjHttxpNvqCdRpPY5STQqP
A0ndH8Q+0s0hlowvO6v53XsWzLn+0VK0c7dwgUHz4Fs8QPYhcQepkmF5dFq2TOKKuGeC760lGkPh
ShMth/FPMMieSjD3sgUrTmvBKC36u7ZO+egGhxT7Xkj/Jz53JnsPidy1FELeCHMu5wZq1QY9xXIc
SRMHWp7y+oOjm+WqDJlQBj0zKy4YCAwqlFkGyA229/cOuZBNHKQhQm7IkGBturjNK9ECBMqwJCHw
WtOkZFHz6xELWWKIHdPkP+qlVX+rwieF/eVmThVlYlasTjBOoJjOTrcOvjyMBPSD3/xmHapsRuiu
b0Wxh4Cdj7i/J/QRgXfgQp8FkLZhavbGPbdkyRh6R3nLVo1hSqSEREQ/3JYvIUf4jOYYLS9QE4SB
rQM10sYQyXUKle52CT8SITp2Q11HC4vb4qhXWoW27EHT2nyG4iF5BT0yjo729A3eNhpPfcPG5nIF
OtTnvYixwDvSrPnbZWghy617ASRwr4WLiZVhnxr5ImLwupQClcFbQNcLPzS81cz5bYpk6UGfAh3S
2KTmXPs98zrg6ijTLlBIsylIbQyNnU6LiIiOYDvmM9ukY+FCOcOVQticvC2mRedeBr0khVlXZgHW
N26obsLHhe2JDpF3jPFDBPl8tNolaBEzJooQppfacCbZzU91nmdH5KiMV30WwzNXp+ZAqx4OZipm
T66DQxMqvGCZSFGBzQfdEGl7v9Nq7VkpcXvNwz4ro+tyLgu+MCSIazoDMc5p7cAgeUgvNbOfSapM
WFG7MnEf7/Cn4Y3OYr9N8JiI+DAXDOoTPunsAVhV+rVgdMf5d+34eXLmLvVzLCqgQNONZHYXsD44
E0Savtu0Po6S3qQxz08W4IAMMiGmww4BgUvNPpyLV5U18FNbz0yMh3r+NVSLrCuEX1K1mfc4ERb6
mcJ+RgiMAerM0Jp+7hD8bAiIH9K73SEVr0i8VufiOhoYUfOnDmjmMrbkE50tEjZObEy7d6g6MOQS
BXDU3zoNZOcRgAOK8qbb53JqI2i/d9XGbj68o3Z0Zyi/wDMbZCIxuAwTM5u8ATEEvj6mI04bz/gp
K9HAiZ6/Ejv4WUX4b9kQC0gpTLJwld0uOkQrhdEMxqE//aZoqvHbScFG2bm1AjgksewjLt8ezwpK
WstrYYhbAd8a7tToAWQl+BxXYaJN3Y7164gzIMbXLQWu6NTZGRaeAS+JywmMBW7DPGVGeUMpJZrP
XIA05xoTc9w9Qov6DkR+AKq6ssFf0zqrZk7FPFgWKauC3YN68+/OaTMZVuqZtpDpclNiGZI9ORxr
zC/O0L8YIWhZJi9QOHUv9Av60cJeeUU2QflJ8PfhpD98otl1yvLx3eGyj+pB7e52vwVe8Z4BRw9Q
KVhpdfd7MQUd8cRHnnAlthfZ3sInq0+ILnOS9XBQktvx7Mhf3E5hDccMA2iHLujxhpx4TVAmG4qW
MedAStfFaL7nh2SxojW4BVy+GH5p3RJuf0YcSBiXLooiwV/Db+HeIDgvs1tphkJkOmejATid9bM4
breRn+UDShQ4TiAvDmGRAi3k5g2JDiUTFFn7Yt6BDx9uXKFURxCvr3LCpP8mH58jz5RofiPvqgEc
LuSz82Vc9FjhJmFooPq0Civ+yrxDmcUnIiUrLkAtarGjTrVmRk1JhEL8mjbgdk9mkFPJChtQ/Yol
ZaR/WiAaCiTcaaEdVm2ZrdOWFjoCYPT780g0ZPlHdosZYqafmwwsWiKMWstg23uAztYgRrfoh3lQ
YJyvtxyYkvcZQfBpslR1KqUpylSLGxzjM4h83vc43x8mKNFlqGQY6cE2aIeZXoAQ/bfNzwCYuGHo
3CFCFz9noB9Y1DaWYQLGbnbInLmiKZ/qQFTU8hr7mtpZMJzgiXsoBPYbKBek/mKynvGWtN3yUL1u
aGE5CuZCpv1NyPl0CuP6vIJbOtD+XhvXFmxJ4WbNqNiZxtQzlqgOG4fAZwZnSnZLnqBkPuxxA+pS
o7Xz+TJHiXnjJ6cPHKz5cq83o2S5rWEU8pNh6Shh/jTheLEW+5uzGgVYKy8sryiVt1EiFfYaBfRk
InrLWKR55jfegMGNRE/8PWfqGP1YlnhR/r4fpuaDooNp8f9p182C8sSKSyTT09/UDQhE5yMRyiS/
oiw39P4jdnmmn5X+DDmhI12opXwpL9NgIA+CKriAxBUGrN47sEMpq2S8VdzS6tl9Stgh1Ncg26Bi
FEF2uTp5pY5ZM10OgG8IV+v1ZipzD1vhe4VuOLDeYNl/xH+0TgkH7Q9VsnS1LviCBAXRyi1UMyfo
k61+xmx/Vglc2AJpWIya/wbw0jUWBXCN6j4VkuzByabqLPjn1fsWV4orTfkzIIbxcBwz7yDortnW
jALr7346eeGRATDvtU38V2eop6saLFZTv93/tjziijkHS5IOCFxFzc5hMz1LSrIbhFz4hqRXC0OU
cQYpjG+z8QJmXTXItjZafCk7ALexlot5IEYVNHRne1aC9SUAAHIvFXCpS/OJTa9LNWPIfJtnghXG
XnZN/DCRC7nWG1BRtUzoUJEjiYMpXomtsg5fNSCkZ2B6ZXQwptIlxQ8ONYE6TSSjE5csU76m8Nom
gELgU2rgnBHwZDAMkUQfeSKtKBFegF+Jlkv2JVjz/rb+v+0qyUP5pseg8gu3rOsIk5Fkl+Xj+wPf
2m+1Vt6/fyOlptHgz6khMe+hV6l46Ccr0qrQTy8U//M8F1eK4dqYRRkH9F7oRHFNDzh1VNqwQOum
a25jb1Aq8ObqgQYuw0ZOz/JRN7T8ZqUe0fuRITPW9ykHZdqUlBeEEu9kK5yJ0qhKInUMLOxnRD8J
YdW8tzE0p6K1DPXBHYdalOK1g5XDh0Tk92gwQS6HsUA6z425al1DysWFy8usmVDaFqM3psWRU4Cm
er3rEi7g4H+sE15XwISfR1M0JXhdnUmUwbr5Foz+6sE0WNJRU3nGfOUrg6b7Arz2kFOzJ25OtSOb
FAKRRMXmCBzAuH+rk3ZpY9q0aALO10n/IcIpYqkebTLw7/J5kC8pMVD5uHBsGFk5xW53XZFlazPI
5YUIVLW80EbUEfMif0CPUy1bN0VtGIAeDVho/Apa6wnbkf+P9w4wAPexU9Z1vWZ7cW4+RQdFjGN+
qLG787kDYRUUIPcos+kDKqhNzYpvCkuq2N5qa56xp5MXAnMdL/xXq4ihN/19nWh5q5eLSePdvXxV
MqZI8x4LcI3z7aZniWQxUEERsh7+j8tuJH2Ou4DOox7ZrNfNRcOJX5sxxA3urqZM7fXR4gTslmun
h5/9dxCnyrQuA01FHNRcEnp4TVOwMFKu+WivNxIEzGhMxfyJp8Dz2zL2xv0z6Rv3qs+TeQq9yFwr
OgPS2+AgB3E/iCdLvKx1fv6glqTQM6jLXka08byJmRNkuXM6bHfqCbxUfy5ucU2pIYXL9E4CbdWv
R/PPRBbcopyxPGIPeB2WDt+90yNRa5rskixA8JF5QkqysLHC8sCIlSaVhh4067p8kfaM8qhvWp9h
GtJVBxcGQpkAEgYzhTDSW7vl0Pui3AjHG02ebH7FNaLMKLHh9yLA63FnyanEkf/Xm5Na9MZIG+22
OIw4XM8piM7Mr2epdTBc2+GxYooxDCGx7AQOteJv8cDXOCOIai9gNL9H34QJ/McuHcINo3vmTrcO
fNS3nTAvBH9+IxxEcmn3t0GisidbTXBvj7GA2zAbc8AFaUXSim75Qc9EzdD8MrnlHHKkzSceX385
jZBr/CpJ0704urlBMK12zlfPS7XCLmno7VI9HDr61bH7y6z2nWWpAb+azD01yO5j9Vp6avId8hT4
mCrd538uFwfFwVEiz4Dvq7n1Pruz24GTMtb8xoLq8491QC0n5MC7KycPKJHKkQx+YAtt/1XEVrSu
QBA84VUrDpEEtW5GpnGbLn1OaeDHGp1mhLFPEPuqjGNyq6ZS/NTq4XIoqb8uQmQ0uonsTX6g/03c
kGaVrPB00GeKR6vD/jQJxDBvz3i6AAX0n9TocBw8QlfGLKhUxsytEIkoArDuX7nmfIlPcKeYw6gz
wqpFyzlhvv+cE1xHLyPTxQa6GEUx2lMvmRKeEy/FlIl0TvRzK+wgYBg/mkaLWKK6bhcJ3h7Darho
frvs4QvgFBi0CY40rOlhp3yAJb4ffu4azzJHW7eehrV2EFT2Jk8C3lswApJZA77BpGMK3NmUX0Rp
67fRWPvnK8FmOcnKH2kuopsAaWdXy8Ny+6JZDn9hvY8AIBcfO5SwNCEITiKDx3xraFq0PUQ0eOHV
UBMKFuK130ZkbUmm9uf2VxoroGC/c/SegY88QrRNNXALz+tgAQ3asJZPd40gUCbLm9KKKxRV8x3j
L797E0Y7ZONzt3tAIo8UMiENG3+HfqnAJb7D+ikm2x1OHe7WLAqGXGgu/7A2v5rp3Q4Sq8Rk+IWj
NKp3ZngtoHjU8sm2LyKtIr532Wf50Iu2cq8BCzM0i/FIDHHh11p/q6KmuR0CJkLucvjy1gL7AlBs
zi1VmfbNz9qaVTEIchbxuboV++RB7UCXhJbp0rD3W3gSQQT466tVPFJQNpyzqN0XEkrfqz7XgBtR
HCFq9dvmrZEWn8ScxTRaHxecIt2U8284pihM5CG6fyKI72SZ5FRqQggUtIZHwV03MSSjA8uobBQf
auqLn4olReSy4xk+BHLk1UFYMGxjuS0YXDHBTI4/4Q+ns1gaL71VRhDfR83EFi4YJJvtHKhEpKdr
TYAg3Okw9M2WVGVxOhYMB1YLOng55rDoVrOMTYkxoE6+fjcMDh5nxvn3FKkO/zA6XsnPT8FWjGJA
2jYy1Ip6ChNZ8iyoY3wd9S1XrfJbZOHQhvSWlkPbFMLA3+5wsst4C5M6t4QvA3yjX32nIF0Mk7Px
TErRxWT97OQf+o8hij9WiI/UG8KW/W4LYs3gTvZUssMZyv2YGfawKEw2K/t0kACG9hAsKHtMbWaJ
o0fDoWLOOZfUVVbevCNjxjpCltEgKvhDLgqlZSqo8nCQ90Y6didBptW8zrtzlQbY2LfbTffE5mVI
J+P/PqDVw5YOLoJRFLN9L7mJMvhVB4YTyRWWnXINBAV9lNCjkgU/2ggOtQ7mL2Sp5yw80MQZAUiD
t/LBd60zHyVDq16Ec0Gm/jxzz6+9Dr0x+nGf1X+qukarrukHyDh+ZYdKi25Xbfh2/yeZYb7ru3IH
+SutXCjxTcyzmFmCUBAeMG146WJvs2ExYHi8IVn3vFPIRRPcEkh7UX5txUatUoLuDsaB7uYGyo4c
pniBf6p/k7aHWUThIp/gu+auJf+y8Qt4YzGsVkURbkdhsZ/k22sq3lygO/983Ri7lOYyBaXIJAHD
wJJhg43DIDweDtcNALpZCz8QoMp0R9tKh/4xDuhKtiHOu55CwNz2z//ncgIxAIttJGoiTAb5ZRvC
ifQ+OB3J65zlYXxQrePDkQZ8k944NvIF0kCCdzGgAvhSJ48Ry5iUQ84DRKDle+SwYeUJ8mCJKGk+
7lXtmZEtiNCZHpgjg7ZsktQsqYWXpQpYKt+F85mLX1stmdLHM3MMjhWS1LRIho5TnxjivppbEpAs
yzAw+Feu3ANVOXe5b39948UO1EnlNsZNkVqDz03yRz5KLG777FwIpDJc4IW5ZffQLylWpOP8tvs+
iyVNXtTTfOoZsVfbjoJ+YzQ6jGAXCXd5Ny9dgMS/fU1m8tSphwaj4cN8Y9kPvOquIeIHpL12Xyni
hL2qAHSDY7kStvLaZozcqS3/7Q3MvRSDsSicVy12pVnUAg2k+nlO80Jl5yNkFlEI4xM2ZgFWm1BV
eSfcSePDgSt2qsa0HK85fCEr8hQIqT7lczk9pVyItezAsO5ELcWWEWlEZcMOpPzIsju0yDgQ1LAE
3ESOgCAr+623r8UdFHmnbEZQyXr9vZsXA46cUtPepfB5KMY1t62GrsZuPltsBPrXhKMxyYRM9imB
iObLSwT5iDLWJcRr6tR2pToejtDNmnTHLFmT+N9LXG2658evLk2L+LQKVagYoTsKr/8vtiQzCQeb
FDP3+D5TYciIeJ0ZIT+9wfD6LPzueBr3X9HltSQouFe9umUpV4EpTnAgL5JeOmbanwMJOOomS+sS
RfOgwAnvLO4XMjcZCbK3a+0hPOxdLwW4vc6YQd0nhHSMcwNUkjtiPLQl6wq3/Hi1zPq+2V9ga2LW
6Yt+jSIm5MwgEp3rkQ7QMbbmUYWNy33hmyFyoW/4QNdzUt7OO2Qz20KOH9Stc841/1o3/0It+gtQ
uOQs9tHMiuD43MRsNO7Ee2l9rHlaBKyZqtLYaLeTDtAGe3+g3a5XPWW5yRbIRGzPC5qu96GilPXL
deJiesuxOVYkANWYYnlN0TUCmAGxc4eYzyzeE03j/joAtyqOjZjpSmYyZSdPOkePDrdpukNVx9mX
LJJKViSUzAP/FAsyDXBeFQyHe8IeZ95Pap3zjHEZpx5+LQBkK0dIAbZru2FLtY0dgcy3kOWYRapX
Sm53ySKJRzQUNhATmFkfIwSTveRx+wWRquUEMKvjNxqWfFOipCy0VKGhS1H+uFFVQXylmJJpqYHh
TuF4c4aV+olvfCYVBzsjVn2bb9A/tHk/R5pGuzQxAenR5PVOWZAi3BFDHjCNV4Pu65B7mHnIuSmz
mmWeqwk6GMK8jhDcrsxHknMRhJgG+E+5SLR+JWqpxCxPcsfgflOpKsioAyVjjsk6prVzJjVssxa9
J+1vPx8L08LJPE5kJrfmZHLG2nsNZdqGhr0mMsPWoqE2JZFzBDi2yE1B531L/Bdpm9NObVc2wXFg
gEm9TnqLjKh5xGYBfi/OgmBIU9b+3ixlpS1u9B5nTSw2ScCLfRELaWHwoOfCLLZQLAnbyrqqIdDN
k6uVNK6nXSKvAGvOqaUYVRpP6MeNj6xTgenTbkQCSOZpMaONSL06SDpkGpMKST8M2R9dk07QpKn9
1PCoLxxshtyrjsuVJqUJuaTHdpRIdHxkov7zOvm2W+GMAISoUdtOMzl9isH5ZrcRBqJK85Pw3Qqi
TsPEzDn3T2TfznJaKvwMSI0TaU8QDUPoXRSBkpMx6xrik5KUrueBzFvsMGqv+hdGb2FnzoE6ra9p
s3jv9HGCRkprfTl6EL1MnN8nf19bT/YNT/VOljSYoofkGBQ441ZAqz5PDoMIB8uuZt5H5e9tIP8Y
4RUVFSQeVCpV+j6COCKR2o4/rXjFcceh7wyt1pJcivKHdn85bD88DOQXCieFTXM4P6A6g3O/IrDP
jGupcVfpycXeyK57WFxwDauoiXhMtbGvnDs5bRjSsxCkd3zl1g+XryPDZv/nAw0mS4Cwqd2lUmGs
jXzNRR0Wb/+LDyi5sF5Srq9QRKc4YeHI8fAwYpNUHGklGBOyx8IJRE1YJlgVrd7H80XDNOAKuw3b
b1SMRdjNd8QhmqbBb8Bzdrj9GlnMLrQ3VPzZRt0+OsDuHfSy5deac5SOMxET694zGdOWCmOQ/0II
F9UtgQbvLe5qxIfWwdXlii+8txaO6VIOMhexHNouL2kqqhJHn6xbPvUd8N5JhWD/G2B7/EevmGsQ
yKuveD3u52+k6aossqwKBT8heTCcM8WK8GTpCHjNvVynEMYMhi6rw5p4sJRiFmlcyNDx5trVKWMT
pbZ63uCC0oJXgVy+hbjlRR4rCccfqE2qEV9TJ6Kz9E7TrPDGesytJXwMyDGnipzqUgHMP6K70lKn
k2HLT3x858IowsdtVcdCb1q/9peMIM0AJA3FzEvcZ2xFJzvyVU9tEnfV7k3Cizvn/gu0q/XnyI2G
gjg750HsJi1MR2ehbgKBfP7bpdzYbL/FIuwrCQO0TXvgXMD+vrYMQ2xnQTEhfM4OYj7fxFU47zYo
jGzd1KeC4s6wysHS9sZd3dtiC7ZTz8XNORJ43W7HPxfaO32PxyNxE5flAyffO0vidWWN7SR+KZjD
q8u7Rf2V9QzIydd3F+wdgjLXGV2AHr6mI967AjZVvklQ3tw0mdWmVEpdBWM+iyYL1IHPCfurknFC
hTTbeBM+XMD0hwIkIVvN8H9vWHVF0lGzONw9wdW2p1/oS4MZKQ8RkT6Cof4WdubN8kr4tMy2NQ2c
KNW+EL6VIAqp2C2Zpz7QtZOP20nm4p7XXFUaD1IpSjfq2NtG9U0sJOJh8CKvp+9uuEHGwzFG4jJk
Wyi7b8KDE95NB5Eom4pukwJB/D3njnQeQJAv0+K3XfezBMNKOqhIwYhPd69Y0QH6UY33VlVh1+xi
UY0oTbviR2aXimSEFAfJsNw3j4c8hp3qmVgWHfrLgkLQrhhLy6oOMAS3WM1WAKxBCDjcf1swsB5B
XbUxbVMX+juXZ0j2Q0bJ5T18CyLjTDRjunN+yLRYGerSf4D63QzMxmvEDQrLB/GEIcAN4rgazHV0
DrOn8Q2QOQpbPSQB2Zgi9SK6LJMClOKPFax/QfTdG75g7b0fSiNEJ4wNPNbgkRjs5Ne/T7neBuT8
/0sFfQsuzZgJeOBwGrUfHROH1pOnevWkaCiVlmiTK+jYW3HU1ldPbu2b+IQ9ixTBkn9FCzAfTC/E
fVBQMD+6PV2DZuyeJRb99glqfxroP+pxIjMWQ1AnkkL9jhQaogPuOqBvrSTZeyyVABQPWaGHRLsH
FTxXdN4fFyEXUWwFl84++1Zn/WrkHGsJcXR+aXdJ1DhbgRlPolz44/tbSWwQHZR1px3hc7zQlBfS
jqsgleg0LSwOCQj9MOnC/XfIovSQtUdPKO86+7cpVU+psEBZY89GZWZ0NPPLHfT4xsU8Ajytm74o
ko0lHTXFd4w88ywM5UjqPquUcfQg2W9LYx0o28p9pcJXhvMI5nbtra4pYY1YeOT833W1ibqyv8Wt
9MNnalV3Li8Vfd/upRkpnSm4nVHTgWjGOWW6Cjfb93MH4+w9sa0Rxj1eqZ9h5mz31DybGBD97PWY
/QeSHor+GmWZMPgdKYumg4Smj0XvExfsw7QL7MYtBut3UrqHxyBlcYjByb53G/fuZ8ooifPunEMZ
dkHhP4dLmbXpARxX/DTBxDyyPPxRcFl8gR/Su8SS8CnR13dqdvRYglCVFRMtN06WpB8W+8RbE4iJ
2GftPMu2s+UoH0RWlwZ3KtnjhL4fx9py+Kq+ZWzV/WzZ23g123tHj480oU7VTWABLTg7/9lZ0MfO
y9Sf5+29aqUL+Pq9YJFKR+V1+pMyD+ueTK9YodXc3Y9yVHZdUBxkRq4Ck2MLhsfcOaBeAh4bSA8M
y7PEzBl5Hu8PRk70JoMUE79ZeLwvJNh5DccpTG9po+yPKZRsGv90F1uz6jvgWiWTAB2aoqwl+yTW
qKQ+k35VSqlJUg1Eld/1UdfCLWPPdx67NpLAucmf41dCyU3c+1GXrmDADEm8j9ZWA8Mfg+Yopy2q
ZMCiW+UhwJ0UopnolFX2DMW8Zb/1UbsPgrwD7dFMD0wexETckiohKGtmsVZ4Eny1pvcwMOHaO3Ir
besIWehLs+jbpN9SP8Yzd/wQE92+UDGvGkqzmDeq7cTXKklAWhB344IlDRo+p15Zq//QuNOmIpfV
klgvsO/e6fiwHgs3I3z73+RxJvai0BSbXQqKvTvpFNLjbi6Zl9N1e1dYSSzVqjjDa3GRzyv/vnAy
RYqV9o4T2etkqwOH7LMrEXesOj2LO82bMywPXiccm4GoVHDfp8yabzdZu2nB+PYqfmX7aT9cu8G/
tuaAz+0XLQihgiCnM3tz2BJWuNqhq0jA0gHRgUTsKPnKKq/J0HiPdjbCSPh9DxxH2XS3U45yU04i
tzR6yMsZFCOtu58zbBGXR3XlA+nt+RwB4N/jzbRbGEGo9K2OliDMVLafbhFKAzPfBnF4uJgJzuPW
7NZHgcFtnzXb7Q7qjvieJgKaOSbAfjPRC4G/q1ALgX9qPv+MUgLTSAXj0+I3xgPbeVbXXRS4XcIs
Xkgdmzr5N/v42o5/Uq958JcCZDSQn8jIEyTOLkjjZ9g89xH9ullj6UDOXeOgfEka/JDQD2XglMf8
JMkmdZLSb3GQBJJiMvvIFWNcYFxrabvarAIG6sV9LTa8BmfqbL/subA5gx4DIWxyHKa05BwJnq0L
uPWikMMtGDDkInifOFQoskrt5Wv2SGTKbRTOmZIPUFGMlQ7VyzD2KBXVynNHtq83LN3lgEc9JQnM
w7qa1fzWGoLQe+G0cUgJJimKtv/KsKIHH6CsPe55xdVHt80I1U9ReyoHMVo1KytDt9DrYha5HJ8w
ZaS7OjwiCbdzg+Ne2wf8k5CU3OGsvWJE1TOfEuXQAzg3CgkKABRzvFdG+abUl7S12tO2i8EJM2U+
qg4R4RPmUw81m8/5b0Yd9BvpiT8LfvH9nMFLtQDb307XQSFLvYF7DJUsGZD9snWmHUsy2uoqS3dy
4t+It/VsfRrL/TOKZ9dQ2pc8/Ic3mVer8FgUeYjZ+z3VwTUp3zCiJNxJei15NG29DkSMAEJ8Enfd
Bxs2A1Nvd7MAlu4FeuOhE7WOtBZ9Jws3jtMTsy0i0X6kLhFdKnyEcMxUDSDCqRHSyHOBtROkGeFw
5TZitZ8JFNqSCQaaRcm6zTIb1AkeFHdIVTzqCQXeJ/KSrivWiT1JjOVKbshxcRs7Iq9gjAtHr6kS
o207TByjtPgxRbFb7INYv27StlNY+5QNmmR3oVQ1ZEZFR+CEjefYPd0Hzdseh5EH+A9tKFkQMXmn
kzva43rHzy2OYOO2X6S2b1dsSxbKQA7uB1tO8sr8ZqhhnlF/2A8gYginhWe+WON5Vhh8heYi3Ggc
9hhn+pm43fAlrDs+yKzE0GoZLAxVlvLiccaZq42s1ONJSCG+wxaQGAH8monk7FgnwMmMKSf7lBCX
ODuDW9ZkrbkPJkIr7by23odmZbiT+um9Yw9bPq+iONSfEV2QW9On9sismJVXvqa+YEAVjXfb0ABs
rMMggeWs5QSAXe3VlM+T2EsbuqQrjRnl1VjQVTthXWMLYv84AVJf7yVDGxC/y42tUxAKCDoB7Dd0
HvlEbdMxIRxdFakZf51ufjRIQR5ftyQmqmOX5+LNJqGkBka+02cFqc4+ZcPDTK+d5P0aMnLvmfv9
n/AMYIttEU2qVWze6ivHFyAi2t20K0qDFwPBzdqImfl0d4Pw6D07xXrx4fHuuZ6irZX3z35KoooZ
Z9w8CYxvQnBPmgbU9LhYO4V3Wz+PAm087NmQeuygAbifa8+EE4xHH13D9W1YirEQnPNOMBIuQk4M
UI6+AUjtetuerVNbKRn8/QZOQJABnB+DxvksOhongy1kSw8WdTK+S7vET+4BQnB4HaV1TGnQEyGX
jAjBLnOzWCcKRGzUqAotbOy06/+oyIfIAZYUjevbSvXnGgWeT/MxrpN2jVw9EMe6hLBBXRKwX5qL
EAaM8qWMiBvsBRjUXv7PAtRg0N94xXpAG9bC/spZ32Qiwlf536YI6XDEWB+TkBA3lECBgS0xthUI
3ky2D7RYCq6sGKxIjgY2WWIp2xDQWMgyaYg89bzTYFup4xCgj1nEujC8N/RZMtjqEXBoUtqkvpO+
fP9zPOrRxy76I/sBuLWXklW49C9U0SuRrG8+J2sy771AcbXPjS6jGgJT2argvETIKIegGeSQUPXz
gH6ZPhLBS9Oynlbxv9wTGZ8785W82DVodznyPnYL7mjPP8todiQIWZ+9Zy2yR+yEhBx8YhWZqs7y
VX/WVCMzGVzVhQ7NVcwHSe/XCIQeFVyv9/gAxhRAyMvI8Oyg6khIuZHYK4cyxWj0vjzT3phcHwLs
7tbajIYslneHNgJkkhuFESq9Z1gp0IOli872eFVB1e3y/40c8lAoGzpzBL/OLBm1ASyLgjDUQLTH
oxiHKmbR5+VWIu3my67PArWnIa1EFMUuDcFCz/gE+Cjgm05F2S8+I2QRxHiZVvaxcFDYOsXooiIT
AcQRO/jLwSNIZDJkqwYSZjA2/l3rBpzvT/Nz/h5Yv63WbXoZZRSCVpsMfIr1+lWNzHiUY3aTtdpg
NALDBeC7/87FjA9lkNuf3Ssh8/JLVk+M4vhvNAnQohJcRy9W7ffotV/vp7hHDdSpdrUKB9Kpy8GU
TRHuaMRbnsH1Ev2Z+b4vJeBnd5nqf2EwV4BFeciqYvI/Sci5u3ob972UtC/rgaNYBCsSRfQR50U9
He6gby/IDQyeaez854u0qTBxk0VxU51qo6+pSrwR0o/3Shl5PINsEssvmm/T4Nv/CNeCzhOW/dYl
ppltLKjIIQcXZpBPd7j/egLHFQ4V/2qpxYOQyIv7/bIxPu2XhrSFAZ9yoP+BLFunv8aI3cDdyJ4D
EpJ9J+4IZswUiNnkgvrVyTTQNi6Jc+kIJGtaysHFlxgYVBMxzYSVg84F7n85/xHWzQtjn48/3W1G
18VG7U32jg0XBUBKlt5NCHtcxG+1j/9+PkPhM11DCiCia+rrDTzBjuXvdWM5wPRE2Y2Aw5dLm0SC
WbzDUm4ubVlMvZy2JDrUSRkPCD6rvmN7gFQxuQPb35Mb9Xn0v66vEbgV/LDbJfnQcCkQ1IgAZD9W
zqFhGmNtBHX+J4YtbP9DmS+yu9VIljqcppvpkINDtC9QxP0HbgxhVW4fdWMDERumMs3OrgTScgsE
8U3yy7n/wWVDREL63HD4jdiXKUi7ZW+3SL9zNjSw6QSTH4l14MA6dZzNBfZ2tloz1k0CGDwKZkAy
e9kMjMEr3TDf+JZTB110JgWWPdZgaBjTEI7lYreFSlMuj6r+vEzerXtQoBCy66e1If1v8H0U8cKr
UTkGUcwabxNFVoMEiB8pRWjNNvvDjFU5wyajZEvDuaD5HHldqRnKoWtkXgR9jmt8nsS+IDJriuL2
e8Fp5ihb+zb+75g1tgf4THOAkRKb/z9/jr3TSkEsD2NqoxqkrQe+/ymFTNr8lploShWuRR/MXg5Z
+tkdtL/iJRcLxXLKFvCBe6ctdKRUdPeOZLo1Cwv6ADkgiYDX0Jz7h1Gf+C/M6f4K92LVVwSJgChG
iAAzUcR+i4IsX8c3x9PT2rrdSKGKJs+SpLH9qLZJ5ihdo1mFzw2pL6pg4RXYODGHS09br0w4AyRT
VciB6p/d5Rq6MeaHel6YAfKMfG/KCYfHnBww8Ftf66MVzug3lCqgyFU9Dqh6gm3qCYB5KsmfIKrO
gkixRgZgXWT19EaBFQwMjI6LnDq9nxoLeXzi7WI0O1CIBK7HqfqZqiH3ThhlvxCjEfb4dlGRELd7
9QUrY6u9TwsIcAj97W/8n0OVsTsdQhN9ro2x7AAnDPMvU/1G9KSoElrnJZ2MTgT6V04eq3Rswysu
hd0Vi/SOizHP8KEUxViaVfWa1cTtdYERPPJuSYCNrMqZu1Hw58Mrtg5jrj2F5NOtkLbrNst2K+HB
RkzsktLSORwBUg7flaxmi4BSOYjEC/0ofV+2uEvhGPprkniHWFkujUsdef4bdwKjG+g5rpvRqdhj
NketZNDye1Y1lcjAjQI6desOHeoI1evkqCkLIKnvtZrgsKZT768/YhhWrsX3QiqW69giBINNBVZD
KvaWBcY0InJQSzy/FNjywlojHs/p8NotZKOTjftESK/8AFY4iDG5E2E6CCxpgI1ctarDMGQcQsWz
C4Ngxr6QpjvhFgr0cPkUg+HBV7K8w9IJxAvkHdB/wQOCH6j04tS0HvYH+fWELyFrdMehtq4un29g
SIAQs3OO0lDQ2sAA7jgN35kSvv23Mq4yqKqQkOtzyqyU4GcJP45b/0Cj2WEzqidao4R5Pv2i05hY
tYY7DDguw7d4Ttt7QuSwvTAbtEZI3YWs7trVqiZ1PCf2TDpXRjD5J4BRKpE5IkZdUx7uEePGY9YA
ZaFKkccJeFJOoxFUcGKRWjB8VL1xJLZUpCgyNJ4jpt2X/7A7yIj8JVqBQY4uTnsWNR12XmnDHvRU
sc6pUK+J/OCusDOrC9ahGXGw4mubNyf4mVqT4B0EFMbgZhMNpiVXGu+aSi815F5wMB8vS6LR/ebY
tWT/fnpunX/KrKQ1z9JUJkzGNkBoKnFfwsBRjH2AAzFv8ZxTTsMMcGkphVocf6CXAzcfJrBwVix1
CfDJJKFxichFfSthCWgFWSRxbMraXfdyqcw7Wq3dhJRMLNxB1zAkidRjV1cNNyvsPxfoKFrwex5r
CdG9AVcjrsRaCYJivyIjfMzYZAkUmAoDmhFi/vD4wvs+iPAW/9lxo8ouUctayvo9VMwmphvozvQ3
CKdq1SVoNdytUoRBT6z3wd7HiyxoowdMfWb4WYp8JBMtf2SsnrJL23G4iOPlc5tfqCI9BC4dZwle
qczqzQMDiRV9RKRqYaZ40FxiK7UMwkay6TTY7aDNcCNZn35YouDb40XFq5J9ld5fblTPaI6OLIdW
3HmwUu2kLzZYsqPxi1cypvkda8rwZkn6AEii1nPJY87nj6dqLKj5KcL91SdmBGJDUZJtVo4bTlIc
v56GHuBLi2BB8sGuB+fbs7gfTLe2/MejPhSJw/3TQHCCbfJv7xHOllc2dOmqz1xJZVkQCmgFNJNO
IKyYdXvc7lqoFuH3WT21WvkSAUus95V7GgB5VW98bY6XRai40uWpHJTDECiLMlfzBvzHhAWBlKWW
X7oKH6UwfuEMIvtSpL5XxGS4UalOxFpYOMlqqKH99Z1N71wU+5MqcWGXHkersRRF4oGjmVBNoSX+
3U9Qn0Smec1dGXcsTEEuXYJ2w40VaSk2LtD/doS6jgn6tGxojnkBgq8sGJGFUDwtCZB7K3yTNO6D
EjtmQ6O/vw7/Jeur/WLrx2YgVzryqYRu7Sz5ItJAQ29MvJfXAjAoi8ROx+AIcpwaMqr6gZRqbdJd
DBUC4TTFKUfSzMs8wz+OaFg4STT/HuvZ9ZK+p8KFRoMA6TxJ1v94djgQsbF5uA8g621UGMW83ybT
cvErbFyIkKQKue1iP3m88yA2pxkP1AF+r54C2W9KvlFutAoP0L61xyd9qLfc9l3MUOKAeXyK9N9v
B8DG4QMTLJwrDB08tfOU0bu8RDnUJrWkWG02BtSDpC9Eet4I6q7hMmMnHuWdfbdTOVxJ6bWDyqpb
vKBcmLDYiBR4KwPH9Fh3VFkBmod7YloclXEuGNEsQZprPuBuEaL9zHu1MVB4RfgSPtuOmVnVueDX
muTORtsGtM79taT5v5h96u0mKsaJPyxe8xJWj6RCQvk/nHwgl965nX9RQPtDemg1dHPXHSSXJHt4
5j6z1UNvzUZjHQrGctf+9867gpBsJYWBl8mtftm7LdBy+ZQVsxR4ikBH6pMxJV2dox3u0cXXz0Vh
UNomU6TdCSrrBmi78iN9udV5BsiSv0X0OAcy1yFDWK2cMXp4W2Bsc8LMGHNO+L4SwJpMEU8bYoZI
1ovHQbYT+SDoFW6TT3RZmWEPBJFfTVhPMIwBZ99iEyVP71r/XOJeCiASm7fQFdof4PCV7rvxhjOe
7UcxF3O6XCnlzgtLK0Xomd4nIhx1LiFQWE7ujeU5WKF6sXiNT7qE5AZ7gzQLaV+ay4wRV/Y8fLcG
ZNRzR7j+Jl9uYMATMP1SmsD25z5AKTsQMSKWYqbm8yz/ClKPeWwMWUAxfqcN9cmiEOQ20XenPr+K
Ul+O4giLrmJ2EXDjmQ9O4CcK/d1lNoDXq6axR4QGQXYzPs4VDyYAMzbBAeGRBY/ZS6SNzEUKqFWj
u5n4AAjJBvhTr+d26Hvj5uHr97nSFaubDf0ZAYuSnaPD2J6P0jtPLOCOaTz44lsL8cPoJvLVq95n
Si4NA3I1mDOwL2PGqAy76WSCH3ktdyoX4STgNqdHvM1M50cxS3kjIa8eH+wDj5l60WYvW4lIXdLK
oSTRwn/ElLapCzMlw38+D3hxRAaKETD9/VYc/JjxzDHSLPIP0MBqmW+2Gvm25C+mOeW9U1Bew5Wo
oMEi/ida7e2jTopCfI95pnUv2xgkdeCjRnYCU2iWuFv/b77+cNtNl1PuOruQKBGtdeN9v5RsvPKO
aEJwkv5IEdf8z3I0/HylLmKaNEFhH2DIrHL7QK6Z4UUGxiEmlSHtpMEBrJr4Sg5QQ3lOSpfMU8+x
CXJzq6SuDk1YcHCqG5QAThY1cwLQnk/dgdzCPPG2+/uC+d9437R60/dCtXoQ2ZoUZypi2fIw2G0a
132egYRgdO6hgmx0gs4/J/d3ncwoaOhO3TeA1K9irZ5cQACtTb1HtOPHW78XVhgUZea0n3Y8ZjCn
8z6m9kQHRYBzs7py9pYG72ST37Qc1AXouFuGUOF1mYQfoTwQL953sh3DtMaBN9BQw6thCNWeW3Zz
BYw68ZbvkgHmoGwIZVPtJeMSdjaqeg+kccxpA01GxVk7vHoTY8pISHaOKqEapVw06icqystsPiUI
YReLXMaG7+HxACNellLuRO1GzDrjsy42n0SR1HyOtrNr8mVNtWgeV99K1D4bLg68CIV4qcTqDAC3
L3+OiJ4n/LYZwxPHCY/2P88sUp0NUVZv28lHBQLDLMcQHJTwXPszZ1fY5LhIzCIsnusLKbSzLoeb
PI+0g2wkGWbCcOGqO7gR4Inz2iGi+WDct/+fSrEH2zNVtmfv4jsiQPM15a96WdL0bAXCM4HUgqqy
So9FnyHz8HDevTaps9Hf7gfjxWxmAu05gQF7awd6pwRZOZ5pBzaVDyo05+PP4lHMkD57lzfWTZl0
6JmQGhets6QQnmMssSBTqueDz3yWUS7cRLIjDc2RfOteCUY30IUy56j8bApyI6FjFT3ASHeWnMYW
+WZgCTRsh5SMy/7HhbjiyY41bhnji7vBAMqyfHmoDPSpiUm+r4cWV37YW0L7FEoWgUibZluMjw8E
9JnhgYOLjJveJRSAqLqJbSvltA4rO+LIzmsuqsr2NtffBKrV5W06/jBClcT2Tef7RtMXvqRyoKJG
OYNB6KQuQECsJoZJ81t6M2Fp3WUIAYCsYVvp2d6fGf3SqT38obUHhMXI97AIMX38oSnF+l8R7TLd
e64tYP1K6MZ/iJLI41fi39eBJGwy8Wj+1nlel0RuUKAJAb5TYSMBzU95+S7INeNdSXZOipo92pf+
/j4UF4VZjTr/wMKaEV1+bX6r1nfvp9UtTqynGqgQlZYQLVHT42rjcyYPoOC6OdxfyYL19cJrQCQw
Mo/wF5BNvS7cXTbCd0AwE6+vXUZE489RxkLNsUWGal5+YxcrjtQCwY0E0+vSm5H1S7I2ocB3c/Wp
0dOKaZEFXneqFfkyl+f79bM0StcDgKUid6HRr+WvZWUgA0ixcnENUYR8eXAKo9dB2TroSiAfOBGD
wcKfSz8JToGzEPkYQp/OADOJ2F5OLJgTKtZ3f740urrQtg42CTRHw6diFQkuYekz9lQL8nG288jM
kHYZX5oDNPNxWOrb4mesfqpowqD7Cd+UqRvsc89nIYpGOtyJpiu66eoFR+JgNeXYgqYX+ZAmF7+E
YEoD9rn0QSRhoXrglixTlP7+d2eHJF6TSHoyiATFTgexm/oNUxFIwZiL9wvmhPjmszDIWlx6h+xn
xMNbS28J1NzsAqRjFp6FDORqVSzePwMQ0DeKr6RS6cqm3tkW3UlnUPR3X4NdXQcuD/bITlOOnFdh
8sazb4lnLYsKDBDg5wb3dnCdzV7I0Xcjl7CiLiXTzPrqb6co5sDyMs9y66f6x5SH6rPNDokEqhnT
1uS0fimzXuLcrWf0/Gi+/GPP6oYzKw7D3oDvMI75vlmfCfvS9eF6PUMUSHoWusNNnVGsix/NCFSc
8XkfBpwUrUZr5LWQWEBjCaQc0NLu8ejB973HIbTFeULxStxnyrlv0eq5uB9lT+XvUbLL41Db8WEE
+O+3RdT5iWGBSSYU6Pi6T23p+smo4jnmFt4IEIj4O2ofVEQGdaN6c8TA08bLc6l6fEzWxJD0oGog
iOBDsuHtqNdHuYkjnJ+kfj6rbO/rO6wRFO6oksgMSu7lt6AOf7G9p0YYI7s1EhGCpbeZ9Lx9txzZ
uotu5m5mIqy6xIiWnsfmOGmWKLWN3O7W2cnFnwagCJCZExrsX/pagAtqDrvcyXnVvstHouJo47am
mfmaRI0Q6W9QG6cpGJBdAq1VreVR152XSAYSJJcOJ53e2jrNESKcR/Kgq97lXAWfbzuwr/PIImts
gYy088otowZRUZaNs38dZLsFjDUnBZGSfiFyNCKER2sEZ9B2JrHry7lrG4MW167TA83Qo7ES7VRV
ebP+Vx1ZiQ7TRtqH2qhwbx1Uv82k3iguZ/Rg5DgSMcEvHdlo96TrpkO8Z9Cwqz3vUIptrkLEaee5
uRyJZNc8jV0iqNHj63dyXTgyE0sbg2UNPUwi5FIY+BmPmMTBtA8eTT7lQ9Davx6g6tmyR+aZAOAn
AUJPEubFiW+OBhRIIuQB7kA1NJjiiXRaEYvb9LLCYFQ0q4M0bZY8xw1csItPOc9G6CzuCnNSV2yx
ABdUTpQc5PIx9ANfX3prNUbnIE114jtZHAkr7RLh0bcAER3xnSrtJsY+7pG2s1vAdDA8Umj3aFOr
+Pakn+x9Q8G2bxPKOJTPYCJZ0zQ5rQuSX/hvXNA+vXbW22Ev0XbJfH42Fdoa7JDqOuHkapchXaOW
rV5f027taFzZtHhraUSWSdQRouuhpobpntH/m7PgQqxNMTp6GOVNMTHjl7Z/dzmHZluXps9BJ1vr
YRPuHHNwMepGUAYWPkl5Av01jxOF6xXEOH9kXacDTgeppFpKceukEfy/tzuVCU0cG/68eHsClv3r
p+zJ0ZL06APsGdDcm2/hjtbgO4V30d3kz9w2RR9/v0lX8W91AI/RqqHIzW+T3SuKGrs2KIlCDCxe
aepMfW9+/kkb9CPzv33PglZKPwL06EpEJJXtZC7/V7wgxvTMPPo4K1zcR3MbC9HPH7VSI5LyfkaH
0yAGhQeeR//R9MNoMQ9A6j31a0qRqtGEg/oeFLf4wq1lgfuYadT8Mdu0sgWIx2fJssFE07LIcoZO
M6kKchK9AjAxrPxmPR0pfYrmyzOhsVGzbegDIZj3zIhzoH2ZD0U+LL7OgAFMG9MqnHYxgU+v1BLI
OCQg1x9HAh5I+samMwTnF/l7FYjdnCp3fwCXKOeQsbB0Zo/7YaZTz3/aKoK6kX265rYDGAOsz9Hk
AbSY86pXS8E+VLHC3lCtlexZTC3UHA803YTH1oqT0HZMI1ZhVOvomQh9WPn9Lfyn/kJaHi6YZqbG
muQ0sr4xmpgZu41Dn5QhrK5ezyDNeDALAJZ/AazrXr7FaBwQohcac1/U35uSG4ksBx5cM29EyRgN
frGulcYQE5XqvLCpO3s8F5tXsXNySj51vxOsOiomYwi9d0CbrWSCXGh52hllElzygqDLJV+YXCMK
vg/XXF3hsQ08BoewdBiz3TcmvYSWniv4ijHuk+Mr/MyLRtNar82lh30Iu2b5aVAxwzOkNyIfXPXi
ChRoVnli3VF+q8IeiQdY6O70HknuW4/IghMRJ86huCyaAu19H3fm6WBOnftI8+oP5D/BK4o3o3j4
8rj2c2wmjmfHecZpkZ5PTRNIsJa55CqXg5Y5CROmCit7aBtlW3DLJ1pAkFuDQOhujLL2O+eDq6MN
uqJ1iuJ18w3IPRS2ZykPI0AqE+YICjjbf+DQom1vm1sHReOd/C62/yzZqJL66KfLZFY8EpV7ZW6u
HoR/zHvVS8MJIdaFLZTSLbkK3fR/Iedr5DPGidk28GquLCUfqRSxR4rSx0sRQpwvKw/gxD+u5+xc
s+XogcgHw9JuCKZdNA9I6jDpZiTjES19CPiXTOTVG+FKUeYHcgmg7yvdXpThnOe2Z4vNSFkD8JnV
mfS+n2OTzhwET9B/mPZWr6Mr9peo5sEG/VwGuAHyNxeeKrp/I0NSv5WN6IbtDOAEHezxA7wK0aIN
WrM8JFHXgb0pGIg3UewGgTahGgmv/y0I20nOuLG/YxB6sXqDrvYbP4x8IE/ghEW1UWy7gudpyzg1
qd+ZGVdvjCnuTSh7iv/rzOG+v1Hujd/ww4uMlC9CdXXH0lqO1ilv9wOM64zKS3Of4LFHCyM0H7pA
BEU9bufMLHaJ0YepDn+16l+S6Z5bEGCFZYks61UCZgkA9uqU/7h2Jf9UmunpfufL9sFMP8toG2fx
O6Hff6T2sa13RL7YLi882zy8AhhsICYFXqUQLK18wfIjDp67WH6ai1V0498Zys9aveWIbufDLAay
+hq0ssWIzsdtgg/Ge2HXUDpenr2w5SOP59PAzLqYJF1g8NTsTLBtwtq67gd62RjMLG243CbDT0RO
QAX1cMM5fzKoCbWXUdf/jtYyoeasW/UG1aSoDVG2p0uu7pRDIKDwsj1JxT2xcXauvCu4W8wczhGK
Bdd/+JUySbhsbJSNRQcyHbpoKqmWh7TCMcl8tcbPB2j/7e09ebgXFyo8DPMCuJ5Sm87Nwurk6L0P
sGYdeQqnMoaZgSC662rydvksA/C8gszoHsq5ZbvyFdvpbPSnuPAD/6lWA6VQ5sV42yKei0SxoY8d
jS4BVZiStMBOhUgPNSAYXUTqvMOyUf4vWZOMxl2rF/ysG4jijGXmCIhTeS1l7oH9XDqtms7pJg/b
meWc4YUcNsTqOMAkB/bAK1XnIr5FzT8DBwNEKPxmqrYTuYH4dpJQzZ+Z4ARRfA9sOmDPStRUdnxP
lWEYMw1R0LRz8WSb/fz3D44s1huk8hxIfNBScqSgMcLKgl0uLVVjir+qOuYmybLL0tTu5bWo7YQc
mhnH1XJ1YOFOyTj0W6V5zojXU95xZujoH/sgu1TR+9AWLK5dfl8o7n7AmYfaZXi1sMAGgwmlzhQw
+yMC9aBoK3v41AY5sl5FG8FIzrsVu6OYi2CLoQanSE+q5uOcXwfL4PoOfcMhERCVNX694PQO9rbr
LVFs5wq8XwKjh3Wya5QHsAbNsZOTdl4ps0hlHG3ovN6CJzk30z5+08xRkwNjvGKKkROGTY4PBFDj
LbX+hKD8VtYmA7LJj4Rn+vzg2r7jQk16sMRceDNzNwQWFseNbtPxoiHTeFxgeMqPQF8Xg9i16YWi
FNPJZF8SkiBBzrhxlhHA/UcGydW1G+j34lP1KlbrKu42cmJjtw7Zw4A7qVz5ICv6kB/g5Ea62Cg9
uUKsKNjMXSNtuEZR2N0qh+P+SauVek2QGmNexvlNdhhc0OHtkd3dJHDPTeCHTuM+pCLdV5/IOHX1
Y47yTDjm0UYLHZ7GbPlxVPiBRMhrkYjIvM5bkitjO8+hHIdVsT451ayXVW3C42Ys5gYHJU1OA1nC
BHSrP6uLN2O2dVl3J+mXb/DBDIMqPH4Dyv/n8mYUs21QSy9n790gUhPRS9eO2/JOOhl4IMnjp7SU
blOyorv/6Wv+v3hW3XjQCKhKg0b2Q6ysu4+3g5L9JmnY2/mLqfzeqmWG06/R84/LXAEmG2sTs5AQ
Fvx+W/+GwUQ0PtSdriFsb89IxDoSTXmnHn2OIqB5CiNu4l6z/AW1g4u07F92esoViY2rNEQAjw3C
ZgZ0Dod2gVUCMRfk7cKykmrOb3MG2tfSBrq6gfYcbMzhp1jXGd1iHwOuZEoEnKzV6xkJFg5LoDtR
I08kVuaZ76wTGyhBt9Fu8X9tanESLO6oTGgb80i9yo5X07FyeBfLNlxXSi0nOyHSbHAMBf1N5rz7
rac66gJd7YzANsOvsth2G2LB0ynQDEA/pUFrpPfisrB+JRznRox9fdiRpoukCOL7ZjKQh5eqbljk
kmQjnF8GyG9J7hBYfLkss2r50UTk6w04GpOLT5htrXBlsTI5UYs1RsnDrlC9O+l/O+eCczUshBsW
1AHTNxNhY4UeCS/+hksxgAVR8/pGzohcj2q+fdUVNA2eerdR2azCY4CVq/LSARRmoEMh1ZNgUpym
KRWq5jpdGHd+KN+KOP+dql170Ld4++ERSYOOpJPtkl2LWl+B4Gmpdf3HXxJkXPYyZeKic11GPVDp
5wBSC2B3qPK4maUsKKU5EcUJb5gUFcyjyMtTMExnnEIPpcpEL22C5TlL0PW9trZ7RwRqjRFw4TRw
YySeTXlq+31lqSwD9+HisLkq6qWA/iCOovLmu89SSrfSlihK48iwCPK4DmPsk7SeD5084SB4EyrO
rLzOsZBAqP/3CBjGTVRfka33TdWFmdmW8pkiknMZBQEtVdws8JshNskoc2duYIQEYo5BfFCmr2iW
zbTeR8aEiX5lgsEH3UcJ/5skpemgXGt16Rz32I1RT49hPowioXvigRLrOIz/DpwwYB9YsG0MpHgB
Re6IhuwhBnWy1t+YL53oVbEjKCG7+3i4eOF4rlzYp1qvzU4NYOxcIIo5aw+X6SuOs8j6JGhmK9J1
QmhKFsOARWDW4FyQp6nEkHV1vgVWH0DCnNuIoaEgYuqXOq+GSxMkzeCAiDBvEiDlsDK1ZLU2q8bT
GKBSrsUEj+S8wZbhQ1jGr5N+/VREYuT6e78vwwOcsq7gFpKBhzJmfkxZXIkV95rPo+/m4cyJWt7f
GIFmNK+Rpiy7zzOEl5/zdkaRDUoTjn7YpahpITjkgVttURXbYMMO/x7AJvsSrczsmfKCGx9/fiCs
MSxJFvE2IyomEOnJrV1pzNMKs81xQzaUgniuxDz+3dLouR4FlZvIJKnqQXhPcpXgk4GARFaUDvf8
MfrO0YbvblaujqkTV4cDXsB3anQBrnWazOf/JHMznYN5Dycjx0AhfFI/9xdW4OxpvQXBG2oCTiqw
JxnJ/O7KD7X+rT+rdcXV3P13vXCghO8BQN2F6eUL60S7EIwD/VQhc1cODprP747DzKjpAC+scRSB
vF4jupmclQW+o0iWkSIjD8nKERJOO5PaonhzsIH8BKtB6AiE4YR0XQfwMaf6wDwF0DEEakqiYfhF
Ry+aPepLimwAOByFWu4g1nSYWJvocCL1alqdBzHhtjsmQ67pUStSikwiaOZ4B+WIZN3GnQ+e4nB9
qUAl/9h2S0zUWHv/RYHzRvjXNjcmpS8mgjRLW7Vb33ee0KmxQpJQUk2SmtSR+Jp2wpWaLykkzJfG
5lJtb/RyapftMzwa8CNrE5HeuLm4H4X+vyQxqPYau+Zy9bttQW4oD+u1OxQGG3J9edDeScY4uvu6
FDoWvNF2Gd6MZKeG/yOK0cYT2aBrk6Fa1G9+7w/W3hl82dTJaVmuWe4Fhy0crfqa+b4mI2KRruqq
4kVwedvrd12xyD7MvPuAZJv33tQ+2LiWmUQXGLJOObENpxSJcIGfISsxpIyOaeWCnvwa8c6KJnh2
Vy6/4olPmwIOvUMjIHeI5Ta6+37feyxgrhVS2bBoKKUjz5NHPE2A8G1yV2gA6k0Xx5Bj5++7ycnm
5qXsmMwdpIcYFVNl3eT707f2VvJRDYdjvA8RuEhZ+R6aEqLGQ/W4/WnECRLlRlSeENnMQkCFhu0c
H5Ic8FI4G2sBaQtjyBp6s0YaH04g9sVlvwdFUOof4LQDQsAQoPWA3Fxii41cA+hvu63r4JqlqElQ
vWhGRxseAwpQBR26zNgjZAj0dLGV757/G7BekPmL9yUAvJCuy1KjvRcjCrMSUINP2tAmDjhugbke
ftWbfpglHW8/9m4cTeC7pTITxSSQwkJ3YUmdUyunZqz7ovRAzYbTcpyvd0QkjakPkqzGWtr2klir
3puzS4ojnbmrTzrHpxxzRjBk85JfiLerV1Z2wxQDYeeC6IdRrgiE2CPQ9ADTzfAknshb70uunJyP
2CsPZBRnUG6vtZ0cX1YhEXdc8Nrx8ypa98vsWC2xQj3Qob+Bz7YfXSZ8b4VJmOmjP0PVmA1Owx/+
kgBKO2eWrWvksL+8SsTZb0fgGIz9AoIQOeLgCT0YHpPaC0ey246Hxl6+ydtsg/R1xGWrTlHBQtmT
h128XWUjDhRroKjWyh8Br3tJX4aNU5CAtnISnuyk3Fk/J8r9GwDpAqlyzr5H59zjzEZGYbHJZzRA
XQVcN1IVIHpARqMoz7ZciHG3hXAa3mDlnrb9FuGDrKr81Jev/TdBkll7gidE5tEyBr/uJD7JpwsK
24Hn5g6aH2ye4RWL9Uvmw4zJxDeMmGZBvlKo9LOr7Y5b/j9aEiKKo5RmzonwQTEm691u9UEgPU4O
ZaD0QSvNaFCNY1Jc4mI8ne5+68McEjtAMTiTCLIcIeX5YKeVrw2voYzZqS+jecZ+mksMerFNqxwv
Uv4+n1X0GUYhyPylKHsuRMlozBIWbMDnP/+MtMHXE2gR2dAikLtV/UcVPD6tER80HHEZICghjAa+
JMSLdr9d5Fwgrwo5Ijj6A+LFJXNkoEM4xjoBXhOsAqY2nTE85y7RGNtjNiCFRncBb+tY+D33jD65
TE03rqECbjoIpAqCDlaEZ76krgZ8PBGjdc//aCCRE2fV5WIQ1RA+XOwIRZXZrRmhyqElrp4OXPf5
fzyMe9vrzzAkFML0wO4ahQ5hjEO3DJ0yXQdvFBYRNv1do26nHxifJJERtK+uEIV6xD9SIRz0uqWk
UdsVgRB553UISyoehUo+SParKSxrp6wXI2W2ts6a/s41G7Z/+KsCbgZP4QvxaNFzmixiigG7RMmf
YNo0wWNYRJeNH45xW3plBp/XGwY7aRmteY0ISoNUatVhI+b35IHCCZreA1oklIehAXP7ANNIysTC
2Z0ysBjQdCU+bNKzJk/bnEIWtqdM/2gtYZlp14juypulB8bmURhbHVDw0lZOS6/7JqKNiiI90yEU
IIj3W63eLGbM/8Wd/hBEpq8OdYB2rhlstz4f29PyAZs3Zq+nZLYvK+nwRzJZfBxV92BO+C8I1DoP
Zd0aymrBToDEeXv8w48fMk1KoLDHp9lGtTJ881xeEOTXzfsF1O6nUVX3G8ff4XLzQy9FbHa5m6OL
coB74WGE99wQ/4HB0qeoHINqlsV7psnLvfVGNlqv4Ke0rcl41gSQ5tPsa3TYFhWJOmkCoMboKHdW
wOX8+RKeC5wS8ItoP1N4dY7grl6WqK/5yrMgprRbzql09f6WA0v81xaQ/0PvgRgNBVuPkFu04NUQ
S8O5IMIUwica0dam0EYiw9++nfYYyNJdD52wREdYLitbLXObaYVK6WtmihNSNBo497mF/NlrYxT+
yehyyZ0prIqkEVcR9nF++tmBbp3OvmgouZI7V0hXJ9Z1GwTpJTBTiAWzPp/Ukdp+7GEQuoxGECbu
4rZVysk0VD2h4LwB5OPNN9udFCT8NcylhgJKXw+D+Ng0JuEzcpdofC2TA9A40eQy9LqzteVDYemn
9RRrp6fyowI39FUEbMwwdnwBac5ZpPKCx9fGSbJ+QVHKg93wHem+bHRzhVCHljf0/aSlXxQrOvsW
WkUYwpVYC7ubYOyvKI3HySV/kUaLhvL5igba29dR56AVZIh1rlZ7a/tTa8LIXwUN4b3y7Kzm2Qby
3zvJjVobXh27YsHH4NX7nEBwTCNLyCbmFnC/8FFECfHNrszh887SLA+1rpExxAJwLntpjzQNi9ie
DmH6Uo8nupzksot0CLFQS4wNThxt1I3CfyMMmwgsJb/wOSpAA5mQ9hvA5QcGk+BGPQe4i4EhrPed
lmdXkcp15POmwBucJAPPDcHLoXtpBfIbrapxkO3xDv2520S1PMDaryBiXgNvNxLGLLFBnVF3XGzx
Wp+KdDPGQVEvq7OwFyLVpU6cZu5JrW0LIq361Dy1UoyRTEZ9ndptR2m2y7SDxvgW83kVuAxAuKXU
TeeRnHjlQiEFo+sKdg5AsIqnJ9bEDXpkg6g8f7v0MR9pRH+7O5oN1++F+VdX+/SyzJzsQZohZZee
wfrr0gkmJuNUmU4MlCxzW2zr5WnrXSLu0ztBk0HQQedrSuVb+kKuLLRgqywsu/fLDnzcbrummVmO
LBSnS4gaPT+uFMZbx279XR8I6YufW/aCXEhCZhqGAPM8PiHomFRgdpzfOQkgAU0sM2gO59lQ/Eg0
EXnSun6r1TneuXi76P8Co1z8Cb+Ka3I5ySOaIVxpEn3xXl88eQeE+4YwKEph/SbvDphLiB8lfCh5
XfpfDMN4b682YUlnWYTHSv1CXviDh8kkscEqrYHYU03OlU3WvB8ES2L3WsG5ODzzwqfvlYCEoMre
Gmog/SF0J2iYunL+ufMpC0y5t3+5C68MiZyyCas89sNd3bnn5mYjbG6oRcOH/Ci8r0vtLqmr0VeC
JhBPkpFhC+cMecinAJuu7RlQhH+w5Hh/PWG0tlAtYcVTGMZbQ4xATAYef4rk6Mg8DGO5yLSSRixV
W6RTMh+hmM0tLVKOFSxLspxaNgcdtkc0lWOslNHZWvfXkRB2ncivi3I7ZUL4Upat3V7QgWEnVp1B
Pn10ybk78vhmyTcPEcclEEm/8ipGBeddGmMVsT3pj7ThWUT2/zzO5MsXqqu2mwQDzHDRBOZ2KUoN
7xvAqa1lZ/iV4jvArvDbZmLLKjZys7gmAygbqimiBAfYoQ4oEPCyMqjoKnfOE/RLxAhAeAbBlXan
P0a8+U5g6mAY7RIivRGfi9IPhW/LV4Wx4WTySa2OPC01DSla466NBzMn73V2YiJfeYenrb+npvJM
WKB1ylmjiePv3SSrDWk9jW0Ri7nDO1vyuOYJUVed+hjwmEW2UCQKaz+H0XRgPNd0lE5IXjwm+rrt
hlDt5nvkewFQBsIlGuvyjcv5+8vY1Ad1sNcz3URweBn4UbCEXOQ5wPu+nc0GFZPC9GIpCWAs7Jzr
YfH5wUOTqZusJ53cruEGO6DqYsZ4zVhFDNDytztcnhjjC8sU8j5VQ1Ajzk1RiUO49lUNb0Lje11w
y3JxQ4d3ScMmI6v0di8Sjkvs2fnof0m8uDsl0/cMAA5A0BxxY7wiH35B7kn1KSqg2/6TyRitvc5Y
pHaRH50xMbIzZhuQdRnympe/uwVFsG6dDCbpwpgeblcKnnWzS0YTzeX8uePaPvzkvhJvoTmFoEdA
+I7LQZZ/8R7GHZ7n+z8iGuT2nRmowaWU9VeWJeshNl99C8ji+yvJDcgsNnm+w2vVGhXihUD+5ZM0
VdnqeOlZe3cz/pPkk/7UEcXHC+KOAmoWPess2IclGBglwDo4CNgwh4ioNf4yf5TkfCEUP4TMV8sq
GXuLgVSn9ZmtMGQj8PV5j+jsorxfoFwTxeLt+o28DyHplkPHdImRbxXsmzDYnU8GU/Tbe+KphKg6
LWoxF26G8VDtQVuMpokGNHE45mJju7VPEZIjBl/+FteAsDu9v1E/POCHr5HWwJzpZkN/l/KE7PiV
ggltCxV8IbRDhpGtvOnpzxEEKUfsJq/OH5Lq2ZsUASd7bZVVQQeTeC2+GKxU4cLB6IgTC7c2ABf+
Ml915l7M/IyupNxevLJ6N9ZiQ6s8WWTV0krpw/Tn2m3QCxOQriqf99bkSvhzlYwfsaTATwYBYqLs
stTbCdsaWlthvw6jgv6GhBcDcwfuKOMskTq8XX2U8YBTqIKKjzh7RquqrZvpG9Rt+O0LPZjb9PRd
URVMnvSr5aCaYursba92LevdAEF1kz/EPdSSYsZ4TUC3VO8pqPWnHsdaui2DKQmo9l2BV1kUfgOm
oY7CPbMEftIk1fjzDA4a1mnJA4RXpQLWRPatJ44NxnKzUV+MQ+GNCIPk7w21YbamncAQPKFMSEqo
HOUDKVqqtjBHI1gxWNCzZTEtSLRLwu6UlW2rsTKcJiQB+1SXVsl26zcdpS3yqCrqnym9LDhgbPeG
7sM+7tnQ5L5lepqa/ZnnL4EcnyZA4iWoJ+Hj1+xDQtQHVvjNyDsr9kW3gG+YtN8GMMBYye1pTuhg
K1es4kCTBGUDSQ52Bpw08k0qdTUuAi2fYFzpJusvlev24SsUcq5S2+yAl3e2jOO6jocYJ9v150dg
89b6V5OWacEKuoELpcy/rv9A4MaGN2okZxfDG+AFduVV9aT2Qyo3twx/2UUDJuP9uv6mNq1d/HhT
SUBjygswkBYKlEByJW0ZnkyS9q1mOCjCgrRLeqLnrapO7XM1JBRo5ESROp8b/3Vi9v+IVPQlfLDf
wdO0veZzD9I35+LW2kGW+dNej2WDT4L46APHeCY32sOGmHR+9Vmkwbu+H7LyXPBz76z7neS5ztpN
eB+AUgPBhPDSJtPinCbkT5fn/LYGTp1nXtIA31raZBp68Sb+Sgfx4HHpZ7CZgGmIKi3DeA0g9jGy
C7YDs9fcPJAszkaOpFJIi1QIvtjVq7gIFWcQ6eqlm+peq76qFiz9QKwFZWXv1cpxsK1IX6KkrdNq
wOOC3mB1Cx19zG3SO5qVxkKT//tlx7cWq/EiSwx1VRG6wb/D/vzVB6phktJjtlNGnbuUt9HVkh/g
vOy+qtmNdv9O2sGe2FJn3xPIkZHEj7VYjqb/m2DhMFDSe97NkBLcbB2iYMR0p6X55hP90yox06M9
cO2Y5raDgeztcYaz1xjAyEVqFC9baHrNz2dOvccZly9us8z/o0s2Fv3GSvBUbFRWcohPSR8UhlO3
ooDNK1iWQZPsi3rRVd8R6iDZyHjNxpBSx8u+12ABDmJ/FG2jURVTJ4q2HlOMQWUNxXxsEFaA1UsP
f4CY5vmuAQMBoNqQJAi4n0KO2rDUz1l9IL3U3hd2MaSaGsHR8UjohsQnRnSJIWfPiRS/+UFdtRel
kWeVhWbHw9dijXu55fWhwMYTkxvrJX9lXGt9sBFN7goQzbGOckwpWHGDBl88+eXO5Ju4zChD3nBK
jG82b3+Of3PtVm6seIdsPPbPN3Cf2kstAo9TEA6FcZCKFVJcjOOkVcMRL57fbFKc6dqQKdqpDN63
1L1/XEW7qt+ycFDRHc8r6urU8JWdfbD/ITUAOEUKqMelOJxhVEmcauyJAPF9eoGubeYBXQGrWiUy
81YDy4sOWtcc6ab/iQUYKnzZm0Nnbx53SSTbXmKKX5d0uiNqz+dgas5eMg5PffztCDuVnU1m5Z93
qJPgoqvLgGjDHLsYfy1JT9DFf9U6VFro6i5kiJrh1zT8tDLu6eDzDKzTnDxWuQAmVpioffpIhGIp
H3bGXBSoESLFHhDKUEhunnpHoPo0GwzZPLOQgSDGNdPoBLLtEuZNMsOnTdSpBMTH0fPr+w0bu47u
l1tHADpNSLL0aVBXWQnd7bJsEcg/6xbe9Py3hU+K7QHjMk/4OQWck3wynqiLif+7WHQRaKXsjyDC
sDMH6zNzQuc8cutag0an8Uy1NDrtTspt2/3MvNSOEjtJ0wx01T3mEIvSpQOwdAGm/uWzalY3zhQ3
AGFEnVOZdS0zzBbUwdD9n0UdcAE0gZ16PKtb6/jTJl48KA0DSb+T7yKca5grYthkmup77NoZCx9V
mJAUcMX/JOqJ55xhS+Udgq7uWpKQCSXFDbKwEF5Z2G43GSDrgbGUcO8xWVCpapA+A50Il52XgEEy
deVUcjRzPVubzmzj3L3wxa+LRjAGgSURLsqVQFn7ENJX+0gALzivHGqGbLiYCFWyOBRj0Q1DXJel
E2ZCKKA2s65I+dnXEVrMmkoB/IBT1q1UP12bJr8OhIjfUzzakTycsZJrGEMctyVUUOkmDpCd47dL
gCI6DU/ivjkPJPr1elTWP31CfkIvNZzL54TCdcX07g6HFNU+j9P6xHwAN7jNTkhfee24AgCEWUAD
YB3JjRhI2cM62GPgtf6A97YYkxFk4fDw+zHJEAC/ek8uF1JBFTu2gzznU3zrVeI3dGgftjcB3kMI
sa0r8Dwz3aQcLJwYyJoVL3AU4S381WQvaWILLP2h9TMxH7MW4JxSSk2wNMVz7F7fWOvX8rJ34XTt
64y/XZaUc6pUMFM+qQr480RUuALq82pyEhN70qn7MI5426C7awvMwohsL8Jz1d/MqdifS4PiUSrS
LIhS4RrLwuW/xGEPa2PtxKJaAovRHI9qGIgfo2gtSQAxkXH2QZHbXrgYdTZArXHlwCc3Vbcr8t64
59LLtNwdj00ugYZg353lNT0BY1dt5S7dQhcI/ELeFdP8ZyW4REKpBzD7B+JAXlGXSp7dGNfVXqDM
hdmxTvZLoqsT0PtHgv5e7JrSLz5jh/MFmDvq/1lrI8NU7tdrm22H1fC+4sW8j9Pkdcwlk69s70V1
s7az8OVPtlVyur3nRle8Bjd2k0lsKIBBIyEuYsm7OEWQdsCm7az7LsO80HGHfr9I4/C1e1snL1Ed
56qE6SaxIbDjgF+fRgq1CqWxFLhZeHju6iKT0K2f7B1cFn+viQS83yG8wFa9WvvFSpwlKSxap2bw
3x3XTMdRDru4T+R80VUFGf6CJBwdrjyIic9inQcviWbYdgCQIWKyUPU3IJzq6y8CtdD8QU7fWbSq
tNWi3w2qIy8+HHKR7MSwB6Gb5kgjUTUFUHA2vbTmBTYirRnG5SSA7dmWRXlvGCBgseYeK1T6XETQ
RaCkJ0sFK/OTm2QHEMcFB1sTuQLoTLpgs2emxN0/Y4BjmLb+K8YLRnePOYzKKhrsRt3nbns/LUEC
bwd5cwelPSowi1XB76/8y3sneRXrV7ipMk+UIAv03IaSBbkuKMi0mKj+1JftiDvbi2orFCa1YAkO
Q/OqJpdogUcdkDUE5clQmTHJ4Ik1Ty4Lk5FnRhnFYMWwuhIxNvAOdI1KxhKle86a5fKW8qiIPAAj
shRSPv0uFl+/Fg/WU+tQP39pxGjAd50s6fl1SLGRn1FrXG9SZVHuUIaSgrNqLdk2fgIlf1MkafzN
W0EPVTXrEVGELItwlG0fcvfT10pyiXHO2+7lg0mPvfOdle6Xsli5Af0rUqWeLbcs6s8n21l15c4n
0r1xF6AC66Y0M/4oykYSJ6E5bYSgHpNSsKt81B1C5VOYtn6qWfkBeDzwNtXnmShH6GIB9RGE6lrd
RC8k206bCR7xHXa4+D6vYooBveMy1q0MDQpftCxRbNORu01XOowrQmySLYvQuZjRLWjwOcXFLqPd
ddPnKHTmL70kVWucEl50wGjRI0PDByypFHVKbiXfYClNqa+vEfyXoS0Q9axcPtx02FBWMFiDXzH1
Jz8tJy7/puOv/qDQ3lT/X27YheHzo4aolrpjV+kZ3DneIjtyPZIiNhWHIycct9bIZoAKlryK7Zc7
rllKN/WeELM5Z8JRqjkl8COI/Bzq104tUSthEdsp1BNHQUVOW5QYn6OsFFIvcz6Ty/7MfXKSGeHo
1vFcC+1JDwBiMSoKmGPlnnvJ1R89aiRI5xXTm0pgrOWrJFJaF6BGhc/cWabYOcPr10eznL7o8Ty/
9eJO0T5sVw0PkkW5Y9juyqKufc3e2hBbMu7odUrh5IG7s7nGbycRsIAUih9KBZ+ln7xiiscW7uIV
z2BnuETdGhhzNvifwmjGE8FhcJmaIdVeC55N2v+8BtbSmBJBAqyb8f9Je0rS6o4LPbyKGxjyoH7B
bbbVNwDPggRUrr9MekRCel3iHtsfdodAAB/YVd6mCjZcoPgJ1QQh0jFTQ0K1N12De4Gu7q2XYB8a
H6bZmK4xIQ+awjgkd2uWM/l6LrOVRd/4tcDiA358XYi4SMZA1Z7IO4ggzw0QtjXO6KnsqyQAvi5W
aDVtQaFeji6UfMZ742xNElTXHJOEAy4FDVrna++bstPXC/rXxN6NT+FzYGo1C7aT9WJib1E5W3lf
KyUwEERhj1goBD9kHpxMPcIJYLgQbvhcn+LJZ/u/yltmqPNTNNtPcgHK9hDdrW9dJNlAn4yiUFK1
lsawguMy2XMD/6GkaBG/Ig0mezKcne6Vsc1YENDmH3Cs1uob1qJZxjTj62yfTZ3TlIhmCA+3/dB3
GHsLajLfZ9LpBzTCc41X7M5BWmSgA1RjUyj47akXV0tFMijNv2++U6dBZ1oaRRdBtngAgChxdV9F
lAyzrKNH9s7XOOnQhShGXUAE1Q64sXH8qeNbdooRlS/DvEgMr8BErCw4ZhcEdyP5lYceCwMNGETZ
iHJQHUF61soGRwkRS13lFo58MhGmoeY+iPoD5qPaA2v21cjOHup7pZKwZ11WB4RhDcdQndr5pRe6
vhBx8DK+Bo530JNjn0N7iFrUP6kQOr4844idjQSqKhJxctd1PmewZJmoXY87mN2Jxn3vuxLfBq1r
abOc91PBq+cj0pPx7ah06TcQOkZSg1DCskIw5CNObdMasHEYu3KD7lrO6kUzhuQ5c49sN31BTgYA
oakXJpv5gHKFJi1/mmYU7u9/MmliXRk2Ep+a+q43CWrFJ8RJpiFlufgdBwGvq6xYtOzRLC3a4gdL
tEK5Uod4JYXVMZ3WC51ecRKv7tazbg/e2kR3FovknrT8vSg0Nm5tce2P9Tk4TkA8EJNa4IkGbtK+
jPIvWJChbbsh7X03TNpEqR2ouyDDocmEP20coZRW2kT6kfjOWzJlSf5NiHNbul80fLt8G+089/6+
g5OBrK6UYiFnjxrMDWUTuJc8xKsupangcWs3OZKw210RSXgsiXd2LMB0GbzCT1CYkX+WJHQUDD4k
St1r/y+AXWP7zIiqZsZtNJXbXfOkz+bGrUJcJbIsd/aoj40ho7T2C9u4/S64stNtH/rs5tfmWMNG
zlsvj2r40UbzFipp7T/WVmQpR7Om8OlAQu+BH/PTKwmN23tPIfoX3+ZGkYCJItMz0iNnmBhthkIx
8eJQoTdTpZtlGDZSINdmYFiRB2ZRD8eOBEIGUU7JnXjeUxQz6CIkSaf1NNhmB5wQyK1yRxg/r+UA
dlf0oYrn3ldaK/Ubxcz2Ni/RnTQOsQDRu/+9tEtJJ+gx9w43ghHHh5NlCB4EVTNW6Hjc7nRjwjON
rs1u8oiylfbuR6Y4CVd8M+fNnmFBfxokhXj59VzGWiK7VCd1hyfBZLkYiY5CZynauf1KB7Bfh3Qf
yyrLBlpjqX1Z2bBn//+ZHefTkCH3atwaQfEN21IGCfqs5m2/Y2EYf5oYKc+uVFkAanpk+FnLCOIQ
w8QuL/w3OcAofC011EvhmXigGitJFxapM9dpR8+lfmv/TSHJ0g7XZzXtP8P4JvL8T9RnK4VHDHIV
C6U11CefcKKgfUGuINkzWOHKFSaOojzJOgsgrbirUozudZb3hjPl8eTmgYqr0UCYERss+B1XzJqm
t3IkF5LdC1EiLMWQXj31ewlw8ATKHN6eBD+fIXUdYd0sblCgWP1aiiOnpwp/9nCp/mUj1X0j0zh2
70goG1S5fAeSl4KSDJa0MBJWnCwS5gl8zTp9B6pJfcZ5qTDpTP3e6HZHKO8SdfwEEjOtH36JsRed
zk0zqZMotHO695tsr3DK5pu0abOQ3y9VyrWNrO4wJaVYW/zwWjz7ACm1H8IYBE8F/jCKZySl+hvB
KoKamSwK2m/IDRyCmeAIxZ/loyJxxoieEHQCC444WEkpv7HY8KRCBGNHXjwV3WAvD9b7k+wi/Xkf
Vc2gkD74EhPCWW/cp3iJiu0V6JsHVJKTn1p1kYgpLIzj3GSe1h1uUmYJOdQhGWHd5G9J9dL7v75Z
sEp6zrCu5xoa7kS2RYm3Ig6sG+6E2x28iunc4LEXQSfs36FIhmp/0jyuBdNUUVleMriXRazddbZo
h+RhqHomHRhyq/rekAfBCt/TQTGS6QNOYL6KTLKjmreD064Yh+XqWvd8AUiHV3Up1PCmlGeCy6x7
PFnCBkAMQTiRp87TjqOxkdeBIJ8c+Gpa3Ec1D4sd5pcHjum51A73j8qZDIobjr2V1kuvBeCWCBWD
5AHwHVPJyQAP8X/SDaZGwA1ylIJS/77KE5InxLKxRA63OmoZ4lzisuhJ9To6248hGxqwW7dbBqLo
G99WwDxgYzBtnqpCHp+n++wU/mRlncV7zzpHC/mkO2GfNr22IzI5hPsBPwPKuGVPVBI9W8EIM1L3
cRP1UirYDeVXTbOSkV9l4GSr9raEoZSC4gC7zoLL8N0lg9njntjlD2wePI+FaCBgQgb9CjopBNEr
61eY9AHd1ljz/s4AjZst7BN/d+uT9icesnZkBpomiGTmXpIjhFP5uDC73ApSC9x5ocMpbxPou+I8
fQ6N3POZRl1wU5Pu+E8u3yk0pU8nBt4v5d8xEy6DA0bu5Lft01+Mr+5kUooUs8S8aN07DleVuUSS
Ckhpw7oMJMVCVSSFrtm3QYCRsMOF3jdSwQso1LwoIxEspyJcrZXZFREWI6t+8/CV0UhQUoXBDlnL
PtmrsvjI0yiDpqRjEcgNaBT2ehgexcxNU3xWaLuB4l7jOfrY1pliF5qblF8EdLU/YT0js9PgzxSK
h+BRu+fGYKMMlaRAcNDFMtIfu6MC31gcmyOVF32m3M4bi2KK4hkrUj33xTCNYmBDsrdYaDI7pKIi
9a8CVkaPWnjey5SvQFIb/fLkllXeAZhWLnk6cCSkS12VvNIDaAM+ZLgR3z6GjJFmq7MZ41B917i/
RsNs2Sd61D6Pz5eDrEX8oWNGh0sxQSyNyfJcAYg0WWHAsSzTnjR2PYGFeob9xfzyEuj9dP1N2jdu
Tn2h+KDRNBOwQb1rFWsBMPYTWImNsdqQU/sHnc28FEq64KHpPd01hpnin3nuxIuCtcNrNrUvdHjs
XRgeEx4TPpH6/iUOZXRiwryc6tOJ+Jr9T8K+z/lbB1Nh65CtQwvDA2Ld14+4Dm1NG4h5P5zg+gFO
Pt9yUdnR6XHC7amTCZ/ZIcucABVaJN9yaqwdJEE2IKX54uTIiudycIcUDPU6e954qcl59GZP4+t3
QB/iDPx9NbibGwwju4P6R7iuLR1t9bwER8EAs8AASbH9lz2ox6VF7oZ7HjC+vwkJu9h/eAM5gYyf
D0Xcxs7S1K8rvyncIDNs25/jeWM+zC4PfeEkxF/DcIbbYXkFDXn94TAduA10vHmjzAd8UXugmVMQ
szbqKA+nZlNwd1OTPJC3M2LdPGJLodZaKeZICZQUqASLWX8IsbjuwDJCPZt9etE2aYSnEhUcxgUh
gxDfjbCQz1I9/lamOspB8wXNWwjqYWUfY9BmOPXWXiqUztgh+vdla9nbXTbwQuQldL1LYxQnvNhx
ujroAT50M4THoTNqbuewHQhu3bE2mu+FyvHxG0r7VpQK4EJe+STutXOqb4G0nEpRZvOc9cPSPolS
/meRBr66bqmNo3XJc+zB77EWI0FgrCQSQjj6nQDikNwCWgxdJEDrddgkEvydYlWhYyM4RTQOjX1F
/ktorffNz2YV5JmoVIOmipjnXHrWO9ZQ6pOgkql/66C3Mj8Mf9tIO+7QajnDhT1Qe+ok0DkTCTp4
9GdMERJ5w+cfvOPy+yIz1b+fv2BnIEiQiRSyi7a8FyfJ5Md4cTPJ39bXa8KMiQ9mU+MJQPFZEcFR
qkWQ8/rHr/W5CQgWMg7NyOZkbFvaGKzTKYXEokKuJgy+Xkxd4G3auxzoQy7viOIE+vN+UMu57d2S
2Pr5oj1+1ASiCNIoO7g3YFOEVUf5jE9OZOM2Q9bhr/XdsnUo7F9h3oojSoQQBtWd7S4jN7E7BUjo
ZymNPMb5+rZllUL+SkEooVRBi4WtPETyox6xOHHCx6LOelSo/OZ7ZD80PpjjjZRgqNTgGh5FOyzV
cuP5un/rz/9JP2w3yCq4Wi2WvsaBf6FWY2R+1CkD2QJd85VjjEeP0W6ZVm8JVNmJIMNc9g5SHSLx
hW4XdHc3DYE+jdyhXKbqE+EZytA5mOLYFrxmnnwUOrJ3ok7G+WpamFipW5GxgSj/ebiJZPHlBXVc
pKk23i6m0I+UkBPvNxUaaiWna6CebE9FBRp68vifIPmiO2rTWv3bCvz4xVEi1KD+2mgnFJO2yeYt
Xz9khJmEftM5A+5ZNTDn7qb0WZ+mqSUld5bQXVjuj2zUhOL5YpO7iHzsgXiT6+pNHUAbXP1PjvF3
T3HQa9tklFNTVCa35/YXt/h1apSuOicP70IzGa5GL01JeZZRjOFgsJorR5l2pKJORFzn0oLUVuMz
Ka6zOMA987RTwb7QtvT054pKgdYJWVRKSsfxdzBxp/50tKx2N+nbl5bmZqF6Y5o2gdEc/Ae6ft7Y
LpAeOdvWIFtkXN8lB1p+WPIXLAeqvW4XvfvAK6ZYgmgaLfDmumhOsPDxqBNUhC6QS0MM1qE6yjwu
3wyVmak1oNCf3s2XhzENwfU8XDUPCY+slUy1txUGUsnP6x1ENWOxiih/jpRKpq3z9+P4PUJkeKEG
VOPyD+aOW7ytexQFOkn1rX+Ww3Qgy37KFXkrp1F1+CCTtX+5tUQrrdYNPlUoZxL20n7arTXCLGFq
g5fQBEZpQx5xkjPAt5ZSlR19dG+T0i3CmYSjnvy7AMHrUrV4L9EFpYtsjQvgRWcwPyM1uun7DI8H
KJRzdUmLjfB1/BWudqRe4y4/Vi5KOVSarrIU2cy2tAf/YFgP2HuH7OvsyFWHnJ4b9DPD0SkVfUiE
3Lxlp3CtYZ9PeCIbPHHnvYsj6HwSt1oIfMx41tlwMRjOpdHulsqrX3fTU64aN2RYgv7Wjwxl1cDP
Bgqfv4hoLowAD0Bmmkv1RWt6LfeKBBtPQRyplJRcdYLgajHnApSR0XCvU2CVHune0sST4ggQqHjh
tm14MruaS7AKaNiBVYTYeVhxW1nPNJBpxRIsKIGOKVsaiLyGMVnc1aiBu5PFTGLVM4lWkmvOiuK+
BCGX2Qqtg8tMBy62DJ0sDu3ksw6mWMMgNtgkVv2Dim07akJmTlzEjokHzytWFvCC2LzKtNJ7sYt3
tWwhiRERDcjcw9syzL+XK6hHZE0rTYMWHpHAbAHwgLhdoj44ciUyC/dJVw9vkcldoA5PH/GIRwCX
fo8ujw1k+cdTDa1ALSitHZFbUz+6XaZZmWt4Kmq9TkpvxKAy0cPW8MRkC4zCZ0dQdbm3mq61Hz2Q
2t+kGuxbQSIpCnu0VuG0NUiTFpFnoL05b2mRWDLbnhMxUEiwBfIzvxN631uAkSzuwXw1lzcjQ56+
86bu9TW3iBmXXSA8akQ/W+YVvOPjjKwi8Vo7yQfpQZfArBrACwe4Uq04VsQ4qfiMR61FxhFv/6j0
64fyjSKR2/c9qYiwvg188bQccxG5PH57LI4gdpihuZblr/7bbsDJUWR0QbDrCJmQ0Cqm2mHDt4tE
6SsNHuTqVDsyBOYPVMVGoo7ovLtIvR5M5aCMqycovW6p4//wiOpxgtq0udmH1V6cfGczxOqicRNr
VQFjDf8vDXoUsD2uAaC+7dVWsA6LGS3AVJImZPpSccj/RJoEjQDw3eBlVkh3QgB9zdBhn6s4nMPU
yJHEMtAU98k8SYPLgTYCo3OZ/Ea/bbSy0i8LAHkc/BNTNOGM5LZGy9m5e+NbAKmIuYs/keyJKsgq
w2NYSvwPmcAFMu+Ud9x8K8IoXZcPj6BXVshDzPUG1zSywNeLEheMLtp+KF2kAwHiyyjRfca+1fhz
ahfqflySS5q2covBams9YSGjYvuYnv3R2SAq4svZEZm30JFmnWsxv1VcA8hdbPXxvQUE9cOJR2tC
Yg+L9fTXpwyatrqd7WW/xkCXIo5lvAym7fFCe1F3BIhL5p1Rnh07p134pX0j3j/oljNPQA11nY3x
aD2MaIan6II8Q/6x+QDsa3NopEgchxI+iFPBCN6lL8NFtVKHqBJafXTMUHQXl3sGLF7zOwsO6wQX
FC9FRHWFW4vr6Jed7XEKQcwnBPwLKj8kOEEsqhR/1J5K+cOmKd97NkEcbjZ6uKyDcOz8LPqrBt6E
hzF29P4Gk3kVOCAN2I0jOWw9DGleqkTm5ZzghD2QFUY0VQPAmwS80gVr7X5X+nQpoYfNh1YthxFv
K0eWlpTmuaDmhbpHMEPx1+yO3AguHEHiUKB5sQoItB80MsEviz8JJt7cqEXlOqaEsRQXRyHLV1g1
uXTEo3h1HK2AVufEfQ/2d/8Dtah41eiGWmqz+qtx6KvmrkuOPy6RvNYN0FPD8CKQUvvKX3hHSI8n
Ea1VIDz5GCVgBWz0IqXKRUZS/hlLZDJaUrrI6YorQwGngAoDqual4B+rnQmTnCQGseVkYDDb6TbC
ymYFHl/pEa6lpktFjc0/FuteyxoEUubvlgYuh+KvwP/qmaPhRIn05J5Ye1aYvJyCg2tx2Zp55XCP
2WjAtDaw4dSICLU65UlRRjFCJzrQjyTmw6JMS3SiSsnmAiSSKoe8Dqtep05/mJmzTo9ydUaehvu9
OKyV3/huqMOzE6Ztq8Z4OLU/VUjdUQ0wuNPdCLg1jgwt1dHpVSHBQo18PFUj7F7NuGZzG2/aSEdI
dXSCLOFn9ymL7HAFqafrF6Bs1uLG1AqoJIxpIq2OKzHJhv0ifBkW/f56oVlYMyBHbW7QVPRm2iWv
4kyXK3kG+6AbRkaoynbKUKAkzMoezhI2kg0kLuerspgtt48cVEnUSrA+2AyGVi6K/6w2S4lt2bbt
hOjk91VF/egH83l/Cbx80E3GzQe7kD7kcibgrVaebfylMm1ZV7Bh4TUnMsFEGhn0+CCBUVomsUKP
i/mC2If4ANHbtAXKQzoanM9SDDy6VT1Nx8Ur12qG7jwtKV9meNL1OXNWmrh4MnYpPIEXDgW9ZA1a
hsQSer8T1NmckdljiMajiumsNFpXQTUL72NM/uVcS94hWwj4PzkB7l9sj6AChQ8YmGyKFOUgHSkb
2hjJl+X3ueJJ3CgJWPUFwhShAcGVM9UBsQ7jSwlG1F6MgLofReGpw3OEnNkxWf8OB7uLOrKtSp5H
rLehUCDlXB0WO38CmgNRopw0XvEr5L6+/bcZq0Zra7nolmNS91Kz2rngGT8Q2KZ4+2vyOM/xey5x
3GY/TYNh135rxa1HkVzSNiU9pcmzZ5D2Tls5N5tJmyxXLss/eAJWJ2QWimeqQ4Za6J0yO7uVvm2T
NSiA8kgWnY1/tfhljk1FLDOP1e3WlVqRo6WWVfkDbwsff5IHjC3ooIQCcUrRF78En9IboXrFA/p6
O5THvuUTgnZUheC0lsCFc08bfSPP11Kdjho2qJgIqIOiUrV0xbS2wFG3h168HfFvRoN7icpI8ykr
cneGiSxiGjThD8zBQD/O6w4mL0OfxdQhb0pGJ9s+gemeia2hWZJAmRfzwWAxvDL9mdGRoggzUFs7
M5y7EclfuScq8hyRcfLPDI/WDrLY3cewe1xX//UO9G2ReYs8L2QVq4Gss0O/GLgFPMESeDLKL09z
kHkJRNxLiYsdbS1qCr800yaJaTuI/39ciVLvkV0X7JAEelURw2NuAxef3ooj05+T33yLogpZJePs
WAL3hRU5qjoDDdVSMy10bm1FXdHxHUZOHpFHjShaTxssFXiTTTGufyo3/dK+pNbLCMgHre06VG/X
pyB5B265J2GOy/GC0gZYPh7W9qHaSJg1Dh1qgClR7clHlta15p1wXvpUXyDDm9oKkOXYM+DiJM71
Usai2EeMp2oaN9Vip3j4bfQGECQeuxlJ7NQ/RXu6HwOLg4vqOLKCt0/URjLK7Oyf16pvwRL+QzUY
Cy07/Nx6sbSefAOuib0kVkehNWUrkdLFLUSLnCBBkLplf4irWPqQHWEauX/sDNSPjiVqO5BnySC4
1nqb37YcpgLa+XQTQ2QqEyYI8H8Q1YqxfwAGLDTB+szz5CkkOZNf6a8qcKSkzMWEAkoYtQY+INWg
zmMrgEavWgJt/a4SMcAJM5mp+p8RK594ep9sR34FHQFUiwxU31HEXXWV7Y06ytN5TvZLP5A9YUF3
XDlp35zwZLeFi/weTH6Tn4uPbejta9CepGJTs/1QPZuVj9cOdTKC6y2YsnKZaIhaw7SieR5sJNTf
v+qcyDblAvT4h6KDISNdcog+9px7BLUvWTNy0Dqk1i2HxMywdzEnYMgo3nIuP/2BejEMBBbd5/9Y
yUgvhSmY4xgpOVPfEQ7NExSLuXu/2iIbw2cdtzt6H46si+2YktWSbaCy5vLT0ZfC/XdFMQScQyEM
laiTiQLR4751UT5MvyYCI2jJL9vhcoAs1OLconicxCrkkHt8c5EqBdM8QFMTklt98OeG9+DK8nsz
gulOnFG61JqAOMl8hiSZCaQIEVQuP1QZGT4wNWzQjZ7rD5Zsn4Xqsk7HMuQUz/jB6rxfISF2xoBT
+qfVR6SSZ1FTyq08Ho/t70oeVu4cYUIUvCOhITt5pm/G6G5Li8HBWtfNCCIt9fJp9fjpoYfC0qJ0
RZ4My8ginkmKBWt0mEdyPKK0/nT2QjQWqyHrWoq6fJiRktnWCke83JQhRbvqOrL4Y8DLr40AIEhv
MSSYSOweIAQigcawccamio6kDHGFpH5MISIyMtCVb4ZexhwBNdQGAYY9/PKXAA/322Kom21kqHgN
+2pYutVPMF3q4EGoK+12uTuWf0ZYRjRCulsbWpRF1FiT+MiClQ/8GLJr7d4tSXHZy6JaFYPFsVmU
YFwnbAxCVRY5yGr1lwbx7zwUzlNLFHFjtO3YYHgjMZqInXRA4XD6kQVjavcU6o7pXUi9FMDqYqnI
q3r86GwF2APFN63Shvsv8muhZdCs5T1zaXpA2Df7PNO/c+iqp+16iPHSgTI9qED6H4laMkS18LBj
dRg4n8QGdcEtvuRPUOway1ZDV+KudGeu8+PPMgARXLbBKK3jUmYzLMTV+j7pwGy0DovOBMVhFsae
vI7oHIBnAYUKodMytHVoHi3JVw0CwDTvCGeYpx8mnHiBdgJSytwNF0aJF+JvTta39yjWmWP6S96y
3IV/aGmUO2dP/TOL6lTGiDgA3aFRMwvqimAX6AxOpypLQROLiIHWBFnkNDPO0mi/QADGgJzUGICm
8Pv6ZlxUrC9pxa5DjPg0vnr3TPhBSqMKduZ27OPpNEo+7YNygPOUqG37/v9gwJkh/VCn5xqmS34P
9dgRRWT9ytXY81Cka3c3ehLZzPk6URztfUYIQkjpsEjoKLPh6kuYTj8yPYgQKZUBQNs1RBP8bVKB
SoC6ZkIBPzywiAs53IFGnZVBJJd5rAhATysl4s0Z8ragpAsv0GPzGC3VE1slhHtu+guUlOsucGsf
5FWd+xFdZ2+XyzBmbsVpsbeqPesCtXPEOBxpmGa5yvyMXi+ObtZh8tkqAWHMAUoWsIoz6m9+gPPW
h463uyliwdaz576EsUoiMPPJt9KKu9/B5a6CC/75BhZC2sCMsCQUMz0e5zhyTVYjDujYuVqa5Q6R
DolWEXQ10sHv5DeFiR2jdHfmugSdviJpC29o1aQGBIgU9j7fuSxH8ZmCcIEhYcRCoATdBb61xIcd
PEP17HNVd9/ANQHb3PrCS7POeng6yg3gUaUQcmXKxO05zLQ9dmNLy5jyvc/yyzmo1Xm7smc6DcA8
zPBNWi51au+itkJv7tHM0V9k7xDtp6uRr6CcEwBqPT6KSyh4hMxXkmUJgr2IXiSnrF+nr7Til9ye
/Urc99u815kwUALn4u8edhdau/IsvW9btmcsA1CNx6SHdYfersYLSPq2153f0YLFASyztW1Xq/ww
O1SeybVj5OBBquM81oDoYO8yNa7byFQxlFl++w73GGZjHmD3LgmPwaBlfWBXy/GPtqCVXL9vq+pk
TuomF7godbRezf9jjSYHhSF79oUplhKbtW+OTbnFLRnlwzCoqbdnk37u1/pVxHd2wasvKDhVsA6D
XHJN6StHwo+i7pOK8U4Lx90ntdaZJ8cadq9OvwbYd3W+jEsPVX2MYwdu7sVyxpfW+4+d/h86dt1n
W0U2HD3hs7TPi4KACIBog4WfOkdFL0/qOlkT4hRfuS8Yk9y9oqqSJXiqPFhafRWLt8JqyZCXrTo6
NgS7oBmtu/tEgmwStgUICvGKU5lmeLjHcU+8o7oeMLvYOwQeApBzcstKfKT/N5GrbiSy09Pn4A/Q
hqCx0hW506cXSAC+W/VWigdFKcBgLf6rmo0+TNxlhXeIzmeNmr+0ZKISLCTo99NvGdWCwwM+kcsb
oRFSGTPfb14wnVab3hysNvwSijcBwIwOvWam2Vo3vQP23UlXwhMBGE/f7iJILkn3MMKuT3kKG/NP
tO2/B/VTCxTMH9cGsWsMGVSLeSXhyIXUgeL6/7ezasPSymb4UJcY8s3KOLFtt6AiOJA4fYjlt5ix
0hcAXxgZB2UmYa61jpK8Fn3rxPR79kw70y4UgkOjXB7aY66UEDpqWUNooNJAFPhQg23FpDpLhcwA
xT9C9OLBbjZVMcWmpWeB94HeeTZyQ+K4AhZchpLl54nRbD0QcLtdP6g+76nGSdIWvCDwhGF4lW+t
s/uCHMGxVdWtY9xvcjKdUnTlTTV3cscPXFpzuE4TqQMLpTdjFHWWso7VuiUXIVNiXncRMTfg0DSc
ERm3VJuSnAH8Z2iog4v6eNl8ZqrAHNmJVBiUMVKE8dYMi1dOHEK1Ct/QXop8NCHwJu+Vxznoyw/U
cZvH1df30G00vRzvaUZ25FTlkL36LPYTnIZ5gAxY3ZoWpOISAGYBtK1w70fbmcoSQ/jHQLLeoNBx
E9TJYSXIAnvUBux5CaAGOrV412PS1cxvyElknfSqh6YD4SjN/z65FkfySqeygWvptfh3pnGR/DOX
kqHsfDP1JPgxiOHYCAvx9XjFye0RIpQOqDABkUQJCh0sSPk5+ntFlo4JXmMy8vZwr6f7TSHfk0Ew
ZCUwG9fxbPXypz3g4pvMHQuc5j02xkbrY/lIzvY/YzVXmtP9M7qv0uF/Zm0eqSu3huw+uTvf/9ey
qiv6vw1qdYO3zcMMLS+LERVsLr+HoT7Lxkwn912T73d/vALMdU5itJ+wKpUCpA3niNAOiTdFrQtC
rFkZ7/PZ/dpDttaEWMptUpHxN/0t92wP49MG4MN+XmmtJvrW921R7um5v9BsnAoa0wwW6gP3CXl+
uKOnwEcDZ2IvTmYOK8FZ50gkNQPh/h2A08vxTdiDx4uefEcmqh8mqTe6pcOc/58lnK3rrzpCKMfb
ij/balFFkqZQuvQWWUA6jJR2BYezj6CynFBetIqmTBFG8iqxRByhJIBDUF5K/EcYjNhWj+9YbqWm
SA+LDUsY9TphIdXg5u3h/3ySZNPvteu2jTXtdPtEpp1llPTk+twMvcLRFrhAHPRpS6+QVG+Y/Tk/
EUUBhGERpNb9oEfaUL8BOMbQDRLtMjOkagdJ1wx98JGWyF1+R0VVHxHzW0sD+0/XB7ZmpAyU81w3
DjRt2XmiP4TPyHOnxW0QNmHXJOT+D2BRkrEXlPqsJhxgYluJJbXNxsgkxLZBxCYraCU8rPk1Zhkd
dGhTFow+A39YPr/7cn5TA0TrJxVD+HEPOKTRq7BgrWpbAcW7lrcYUC0ccdubhuIkUmgpN1Rm0hVE
QcndsKoYrA2BB7/Qo7v02fipBoC3qof3FAB5S/H7Uoe1eh/zfWA928yUpBAzlaVbk31zI0RwltaC
N04RhkOhWHqBJyOf8iB90MB9uSoH+iAd38tkuBY1tjmvgHJizLt7XQ01zwYImcKtaKnJE/WcOMrD
dDwzsN8uYhibHuIJCs0v4RUBXJdMk8a0Sfz6XqZYjbL+ENEijF9JO1oSb9GWDbdlDT4EKDZoAyzu
I5KVs15XR0gHZVNTajFbgRmkURKrwO0Rb7g+/JqDr23AEui08hsw6R1EKFZ1KiTRe9Nzr3uyNEk/
3kDTaYIz9nVhahLlM2O0fjH51rqMoGRAf5g2vakL6buwrvSNcLIG6YQdnfqH03q9cxV1NyOoRMon
8GyhQzM5+vBvAZccEK5/4xqk3zCDaRtU1C0+E00hoVVpAMCvaJ/53MERawuWwYMkHxAFNjatMw/S
bT8oYJlvtgQk1Yr8paWN1mx0o/rSJTgaVuUeXfnDfUcfAPwhWYJvHvGYnVPRa3GJmz0JKmvSVD32
OUm6dP7oqm2W50Bu3sxd2PeTyGtyavMhnbXHkXteQy1O/VetUgijZM4BPkJYwDNGM/CvgFm3W1l2
LPIxeV/VEHuqOPJ6M7JlKWLTqrUFbRFiKMjvHZhtw/6TXa+Ogy4rwbLt2hFq5LKAYdiaHwN0BZ+n
yg2WxEfdPyGR+Gt6le/ZDfSEkHnlccbLVQGGmA53niWJ9BxLJskRgNfa9oLPt+5sLGZ4e5iGbJfN
AaS9XMqODG6PsBA/F22TfTb8iSSx9mzfNZTtnNw1VhzTuCWkV7+w+JMHtsAnF3vzBXFHgNZjBt7P
/ypLna/MmQxUVYouCSBxpFZcryDFep2PCoJJRQ/olejmstYg4IpsbJzbTuG1nBEtiOS6RhbgT1YV
Aoka/x74h3CCEtXujia+fmk7ty0suKrOcDbQ/WvfQotPprhWY4aELUCIYG3uYkERH9SWtvxFWRWF
Fr3Gw+q/yQebx5NLyGudqjOdzjFMMuf8XsxdyLg/DYmXCsCmYQb9HvgW4Upsm0LiRps4dh7bviFa
kCIN5eWLV/ymEOE2bMkLY7m+GGIk8X3dogG4EUTzBNp289eQPN6Fs8184ZLPtVlnDj+dh5L1545G
skxVUBeTYuiGgvgnFbc0Zaj610tUK671EhlEdlqdNxODSQoRNzN7mh2UyEiqfz+BC8WqCPSkNtCP
8UbPf4Q+po1IyCrQOWfyg/EggMmN0ognwU6tBQgLWRwk+D2XSIfWd8zHKdoKZOuCes12RulPz+d4
d9FogIBuxhvyXyorMqHW4rKEib2rUk//FjalUZ0GudZ6ZjiCIpOqYQGsqNjJUyFmz3jpng8GhZjj
uYNo5PAtYL+kGRav68FiIxQEN0SlxgQ0TBsVE9FgnwMRRGQNvYBJah9tLCUi/tBFA85akm0VOEE5
QBuSMOdWh8BmkhXeBR4520C/wUrOSiLCAm6hQV9YsxinGwZhtPcVLHElsls+98FJSy8wb2jiCj/L
ry4rVT7HLhbWkDZjCf0ltz7VqDY7qExEsDNVv6EX/MC+LMI00j0xQw6oPnOdvCUuFGML+uabzgJC
jeRnuy6WikOanq4OfODUAiCZGtpGndkInXmFY6lSNexUClbxYMDwoVqba7xJuurlDLvSByG2sQgR
7F3TNAmOpVaSeQX2VYR/LstMrijr80+L9SDu42iRkrgVtjzeGithzFynNRepqwVdunJwMn/Nrl5P
YJKKXERzoaKIoKf1Vj3KPmrOjI8AoqQ442aD+M8YtaZtqe8DTZqLOpHUGFGWRqYImP0lAYHabpnf
zyGs2NrB153Onpj3Q94TSsYHUsWAYXvqsomM9CDYtHUetwBip5zFkbLvfTxKmtV4kprKqwGojo3o
IrKzorBf4pKBImRrEcIpuYUOSryx/NNvfYYRVmkOgLMPZgX2veh0eDl+CJ3TiPLOkzGpCmMZIcOf
XKab5OEHeJveb0e/9G9aaGhIhJ2dRSxs/YmfCjDTYw88FpepzBV4WT1kUS8OWRqmCS97JcFPf4vt
MboxhgD5p1+ZbAP6OR/aDxnlxAtIa9JhH4dIjDHiIAqNrxTArTPpbzpMrLwJr4bH+jL5WGbjMbQE
tL97JPH2kiiaCH8Vio9Tz27jS6VooTQeXSHVl1eSsKAwVBr1qu+3ziBFBiwORJvcOWeKXShpB64r
4kzyc0DHGKnP5aHX9gf5yYJ8Hw3EUVeVbZsz5PZR7BaRRRJjL20L4tidDdXF3XKxAR51HiP09Pob
l4qT6/V5j2g8n2mCGBDFusU9+OrjbahY1Wqmd9nwDfsUnBFSdncl3bPSw26F5p8USqBbdExbRIFN
wM3JT2LoZlmBvJZ5QRQo6rMKcS7Nv5SjWhnT7VzV+Drqvs8XXYRcQCukO+Jw2w5c5NlzHRJc7aJS
x/3HmSZef4h73Kog2UcJpVIDU1xBygNSIi3lisvjvjHLSFHOSwHugFVFVMZHu5iygoUXO5ncs4d/
IRWMeludmCGIDgsoCgI7WUEZ92Qsw2UIGWiMNJQ4dcEocjrBLOIefRnch2jWOFsYQ7WsdnT7IqTY
YJ30NE8dXNeT0R9hJG9pie5di1I6Oj60ya4mdSZoET6bVF4F0tiioc7bACl1W7Wcg+Mz0gp0GLkj
USyxye0uMbnaJGIziXl+4Ix4MEiryLl20FRvIrz0PnJO8FptA5a/k2GR3bxx9JV0DlM6z3lDtaOn
UFS+8mnuRqkffT1w9+tLYNgbAw5c3J10hwxzNEjv+KC+LXQJdXj7CulF+IQIwEaekd6Zuh6o/b9y
yLcpUYfTBIOhpWu9rgm3KfueJKdim3VDVawssbBkdDp0VjySnGWJ510B8+f8EeXHqB94o5Gxgi0X
PVCdT1ODFLC4mCyn7+aMB5tBYkldBDg7C0bH/sbbkN8RYBjEIcBF9UMips0SSssY/lV+ExMhoIZN
JgWbodtMXyYWexCQq8wMH1LAPHYZCtQBmk99WAHAl5Iqo2E4gcvRHQOcl22aQsR21oGKVq7YYBat
KG7q9YuvCGotObfUQnURhzgF5IXYKJ/f1b8XkzsSct6QmnPvtVPledYZ1hkkI3J4ddBw0mOfKxCu
d+XNfMk5rICSrbaHR6MLirX1IXiwFOJ1pyjSHOWJ/ecMVW2EXmy0Gi1o/mLI+W3LhKgNfW6lFJpr
YjxrrXsQbAO5/uhQYSmNtclVFVNubJqKU9QGuNPRTrLT3tWTMUI5rP+IjCEZuV1DqKcLrM5ezKcr
VIP/hez+Nwhnc23Q/hdiVbgXb2Y6O29H5Ik0SOJPFGwDszMDpeJKCO3mXxoBcrkeEWTPaZb7Xclg
9m+61C6ZqTT1jIDLUsWBrFgolIIf6z2Q5WTJ6bnjtYQTrZbf4ED65GrK1dwes6GxkAoeRfLalW1t
IRj/ctLSDrK/AWe2lC8wLX0c6B8FUC2uVcp/ZHmi2DWY3TQ8JfL3qc9t0a3jd2cfQdqk0/5JD1OX
Wei5yCIjZ8KKOHiaoJZcRVoLVN9yB/+PbVm9jkb1QFaqmi+wM2KRg3ZVIYNH88oIVKOsbhm5VdRB
p74Bx0iNMOX6e5kKUpaFZ4gCvePjUX+sbkOKfXgZcI97P6dq92JVHRhuigEvhHY3BHBU22PbEvPl
Tz0r5uBkJD4ELRZkO14hf9fMdGi1IWPcDF6G8gFhmfufBUSRqNAGqPOrWM5xlIDWPq5kMeiBN/Kx
q37ZiM0iQ7vGHbhTdroemTmZWXSDtFWSFbrsPOVTu6tNDnx+9dJUup85k43Sfui4dmWrMYHU6bOA
Uf5ZNQ8eclQeoiTPh1VUgnXPCo+JK+9kfw7txxIAxniEc0WtH4ZHGSuPKGI4r2d0a2NlHYnRKzud
rLlOqZwSt9HuRFM5K8USHdMwOWqRwJzMpNvWPl12m4sYUyLUo98Qe3nl8Ee8S8RM83OmiNJCNYPs
QDSejk3bKa4Xsebsx4bpBYD8LKucPo/0lYnMUxlVk92quW1ad0UgJAQ2HdJ02Ya/1/v6dQ11btUw
imOfo0WrsC1rZG3VCuD9G7QDSxJKNTrJaFDkeqiRK7uTZyKeU8MI9BBiZVHq9Vx91k63KCDYgC4d
yw20JQHAyTrID6QnXCRchef0BSLhPQcyYDuQ3WVgtMMSKzGIcGhnF6SiOJeqbIOqqylmgCT9gflk
+76jwweHR8ZTIwJ0yRd2ytVYayvqcftDY97xWy3N7IKR5CtnQXajsqlMyPZBoqqaQrgPD1XGQbIh
9x1A9EuY8J9s5Ccpd3U9uATfrQBcgjf1ZuUfpMT1sYSPNDinrsE8jIBH+AIEOsx6ufpGonK/GUGG
eICbmkyTp75jUlpUAGqxf7K+kwgXyJ/QRZmtYaGMdTZAvQLG2plCfQSrr7/qVu0l55KwN+T2txaU
n0stzpuuGT3KSCU7z3ChUMWlpeEt7NmALqRy6lta02HNsK3otKLb4d1BN1sRelpZa44eqdlSASFz
ZolGwdTVgRk+2h7U2SD8iHqmfNp2LL0+HmjUelG/RwDdz9sroVblDnxTXvJT5GSyemlCeHH5SEy0
ux0Zit7WTvLvCs818iiHUHMTylKQqg18LqIPuCw5Dl2jpERWv6UXdX0BzMFCp10ZbjkRO7Q3oJ1c
cXG2FViszUBRlpqoYlOBqb6Po11zRFT9CiqMB27lFm3MTyVyJZbHv2CpI6khaKUI9CAaU198Srgw
KmVALsJRROmy/p6VNHDNk6RzcK1A9Jq+3X1utCy+dEDsahwfvcl0MndWDQgdQ+F4XW6mLXdLLpll
0VY4PofGooOwODbhqS7YmLobokZ2YYVUqwFSK9aofv+rMN5MyK66cILTvnEVwpqGHRUqGNyEOu74
Sd9zJHzvRfH/fkp0N8DBY1UScbSltV1TizR6MbVilEFcx01eGutBEKEL9GK9kvq5GPvbx1Bk8JCG
ZrGifNpGRAds7+8O1McAfuMQOy3GsPjQyaQ8Ba9xXkWFjkVpPXzZsp9TFxtCJBpg484gpCca7Lq7
VzcLGjdxCtxRVnAbI0J+OyT4nWBB8sKh8rtBlgnqUeMht4oNHthPTzZXBHTBQUXBVpXPPYhBRrks
tD/QE2RL0LX6KbhGbUPewx53y7o2pGsZ1tW8hau6We3NuOPZw5R3mpTufK35VL4Aqe2rw55HL2Mk
o4eW+U6GpPhMxdaJIos4IDEzDC8Sj0pq9Id3wMuht4BxxEWfTyVp/4oYhf89iLCdXqQQ5i+M0PYy
sdNiACgbs0R+9c9ZgCgoLFGWVXY2WMoo0tt66eeteZYZf0T2GhTDmsqX0331B+UiQbOGgSNqsKPP
pRpFzvfKmG6ClMhXHkk3fqA8DLJnQtQW1fu0A2zQxeTxK+E0lC+jECelTPKjksuHEtnSIB7WepQW
zDmjHq4vt+mUfaTGcFr8euaBjnjB0VTcs3UxNWccLiSq7VW7tdmXoBRlaW5xhU02is9VFw8ZG3vi
74KoywnXKnMaK15r6XicLZbzXruY0G/JUHfId7zPUoA6hgU8yWmwnXqqJ7pBfktAPFVxpRwduyeq
lSn3i7j7BNTgCbQn3AZDdG2n9pvVNkRpIAx0deJPmq5KjxCqYqWRWEz1S+WEpCxEpUDgwTMztkeW
wRUQaBPHoVpnVnEAAiY+8zHKk21KUfKM/5VoV3IGi1Brc/xsZnXycGKZkmRIl6NMvlC8Si59uRPi
uwK/4DGdKYgzzO28sXpbEeGgNP64vzwjqZ/JxDW+rJgJchHsMswGMtca511Rj5mNhZytanNL/juq
KTth1oYNMCYQDJgE00zToYRzplhoAEgu45io4kIdj9cHkaGTaikxDxyKALW83wFK2oepkTcEE0lf
jshDLe9r7uUlE3TG6C49kC+wVvxG6ognyB2r9J/PvxsLf4RfdyOhFjDjBuwey4e0Po67v6tpsqsZ
/UJU/vSXNpXtNujzX7C39+H+i3BI6lkEugR2rF6i2u5TA5eZHS5JGnV1xiJtWt9Lhs2zP4UaRANA
L5ZUp3FBuyktDj9U/Lk+2bGWXUcMoGLpDBMNuct19lXJENdpjYny0CAJzr3+25Un/kI4TQ1IulJa
DwElyxHjSfg3lRRyp3epiXq5yBAma3ouaomcTITQhcvnrUbfoAaviGeEHBlJFoHkPNE06xKhwo5i
FZPEBf3UONCgNUS+DSmTRvjseyYOh20zaiAt1ZLo2U+l0qnSm8+oRGg2O/ZgRtdcA9txzXhysQWt
MoI/lYyR26hTg+Tpc8wpak6c5lH/smhNzFAQ/rGV1OUAP2D3ul4OL2gIwzl7Qrew0+GsugH0ckOC
64tBTmjeEs1i6CA0urLcUVzPrEoD1EjX/BLOlVzKNDOQ85lA2vAnon65acgh4goqkpM+LGPp5pQH
gLeYLPBQo0lXesFtO6LylMh4lHYEciRefFHTQoASeSfEQixVyiA/9EHpk/2S8FFVBzzGLHaJVAew
EWRaxp/P8aumTGqqt+/vFrAtdImYbK22DJOzvhaW4EMNY9aQ6uraNBgyM8ZfCzzP9L6CZp/h1mo6
mWKmDlemsq7MMs5QePkHp937ZmFvkez4z98lHakKmAKZ54gdMiIov8k+xbyPBi5oOJUgBcKY4DHy
9u3ZUJZsz6ZjHF5PGDZMarWUWX2ySr6JuVB/ZEDCDNM8Eryr2NVAtE+2UNrtuufehIeV7fN6bLkq
7chjrxwtmKHr4PesGJb/4Mi0yb4w+V+rOr7ft6nvlLJqPDpYtpq4RbshUsV3uu/NC/Hxu1mcs+K4
8UlmB1X9oKjWxDXvPJKXS8xSOw5AR4zbjZyPe3zp6q+RwEthYlOM4zkT3OC8Hbj0bREgrz3A5lng
u/lCGuAKH8Gq6nqjqGUpWeMriREjqAXKgqmKzh6eg0siygb6YUxdtXp9okGUjVaPA7tcY1vjeuDb
fq9mA14lXOXPkjf1WY5PDD0WFgyjpFbBbRKKS4jEiGBloz3wgXlUDlz4piVSxXMPMOAzLFWEpCJt
mwZw0Wnd/zQqVVft1Yc2u2ntpDaMZ0R1JmCpeQMitFxgI0udGGuV82PWLXJOID12CcdHZs4RwibT
Sk4LOHSmC9v1pXJxc+dK+lpaOLtD9NzUmrGPeDiKzodGF52Ybph5RUoBcWtnlTsJNbvtieViYMnc
76vNfWZSF2N9/rEcfjg03zB+N1/4VLhnF/JTTLPfBjZ3yFlERotv5IULKKXKCHXgIdqVcal/SE8a
Yk1O5NWdi8VeStuxE4HxFyOmc13aPOVcgtWQcnRyCqs8cDYNE0e0TdY6ZPXh0Qo6MUzcBIEjRnR7
kqoakcrssN5jrLvw6c8MrCEbt4wm+xYVKfgpZCtMLsotsCU3YgEchC5O/8GycEH/k0FF6+SJYWh4
5wBkQE9rXaSL+tg3y4g8OulYjKtFcOAfFP3bCCazX47hu8wnNH65Gj0GechZk9MTToM/LNvwWwcc
DkzFmtEWH6AizPYpFZX2IQJk3Oj10X0ENkTSDErauXePdv+1W7aCGB+rB9HmOsq0XR2Ue6hPMdsv
OO9u9IsGjMeaOdDtZXLrqCa++EoV03BbSkNvcXl3cjTePUj+UkshuhceZxiJQVrVBcpQBp8pQXCk
LBa7eHnznsaM4dY3QbZRmbXYxlDuypDKmy6L2sgDpjSIDeNQkOJ7CIwDOVkavLzqGQhwpI1Agkl6
kDSBnwUMWDtzbLMef+iP8vJRQdSL/4FwSM4v4Rd70jCjn+xPp0DApHJ4Yv3irGiZhDCaeMozsqMU
IAzKeJlVgbFnBSO85i0p7O8LjiEakBkUhl7drJ4bAzgcxPS1Ak4MbgquqkMviCKfRCbfzB526d8t
uSn7Z8BEbgmTqBs61bWvvuMuvmVNWMHAE5cKtR8tV/6CIboI2zpfgbDmt68aUGX0nTTP8d5ZJe9s
oJj8EvzgQSND6MGylxvCX9g7FixTaLE5pbJPjajmoDixy5YycYvry8kGzjx0VMHqYRKhBqnwBRzg
xU8KDaL/KEj6cBD+rBYJcZ5AjtM6DChIl4C18U7Cp74wNNn+d2D6eAtuGxQjrckMXGg0fczawa1G
7T7UswP4o58qZdclM0hgwOx1jkGGFKlJETEKZozjrnpgc3GKn9I66TkRfGkjhPk2Gs5EAwEhf+/X
VIBrhcnLSMYg3SsH32ExBFLS6tqlrJou/157sdqaA2rrzKoCx2N1NBNDdr37kbENmyOMkKECjsXD
dRKGwLGUf6zV15cMMOGN9aYjxaL6yNMRQopkGjpGP7ERBbnMP3nFndZoLFE101I6kBiq2hiAGcom
fODf6SqLGqernDbBNQ5MGe+IFwukV15jXin9TlW5mgPyqxCa1RtIgxQ+PCh8uMcrPA+uS+BEYSMC
nxW0TLCp4rFjSKr7qUH3FUCGBY485M8riHuhgXAfoNXEhscxjji0V76tbiCdFKXMX+77YHLHkz0a
VBxLBA9/9fACtnQXa9gULtE85MraE1IMNtYRa8BvX76QPeZcQ6f2kxtcuX2cL3f5rr/30R2xa0Cw
w860nbUqWStu7W51xIWR9lUgeGYVpD3DxAjXqNVzEI4AKn1UJqogzyWJK3tw5315GGyZXx2ewrOf
WRd5PtpNPxBEqsp9XDzNRlhQ4eJYtBrfx6HMMgSwb9KVmN+52ap/3tisx7kZqIGqjuN15odfZEyV
/OghYdCXV5AVgTZp+CwgN6kdEZJk2Nv4BQ9eJLePJFvPdaGJxh/6kdDbz4wEnY4OxqVvAtX2OTyy
R0EVazgquh9i/luenupdLxhkvJjVwPrLrhsovJl5bbHY5tzppv3J2LTfg6py58VAIL/5zAhm5cow
bonN4mpHHb0tgzQ9bBu+D4jaPqunXji4A5i7JgzKgunh5uiV6cr33btPIgI38Th7ySu2SdRsXQWa
6+PkbeAQCDGHZ/8Vl6HwfJI9sSzfsiQR7W99MO/KdTXKD5CgKrQPdIB3XyRAYqV/wvo0/CfWGgn7
w+TIcjNU4CPCQ/Pd7hxkcPrbmjLGk35cc0rNpYH0gUH14MJRpjvrzz8rruEjs2eM2Fw+GSlc0DCD
W6SW0mRUGiM5liBeQOfdUpeusR0SejeDqfmRVM90w9Wh0g2Y21RhHkJKQH8lyR3sIiHmBYNKxA3C
BwDgK+Is+1N4rWD48oeKmCoku6hWyTdl4F78xMVV99v0w4D1NYXzILqxe+yBxOOrOT1Qer/6MTb1
5zPyDZbxZ+JwkXnN+qYUhHaj7fHCDUmjfQEvZGfuomkS3FLA99pHCl1KRoYXpQcWy0MeAD/ofphI
niM7wP2yjElSZZRXzlxcKMwp9ucru1XFyUHP6zxAe+aYHifr4XL9z9teC9y5Ro8XVGBkKeK2I0f7
1uqAcEPlPkWNTJI+R/iGgw50LFhuZq9VoIW7pgscLzjIB2/cAYQ6sydgvgpWLaV1B500HT5G1rZq
Hxa9jLRiVQ+fXMbM0CFHkz+hhZZaFuDK3TOSvP05btKRy0923dtwLDRSIbDSUGCf35JWer8ibAUp
uUJPemVeS3Lqo+eCpiCqex2CyS9H7dSjb9pIEt+X4wANR2hrDYWpE2gOYyhGwXceQwxA5fkJHiiO
hal8nP6tepIEl5xCug4i5xOL3A3CQy0qs21t6/dgcFehiG7Z0wDdAyIe79xOEEqCY1K5LQrHLHGk
wiFMXFOE5ewLJ8I6gf29DDjJx5/DKrfXKsiheaOphQ2SKnIKuLxBIjHwwZJcjtlhXw343jTEAF/S
b7vjeF+qMYSWls+bvzGb/xoJ5/aMM7C/i1eZwBXnL/IaosCmgh9o71cpnfyeLlClvkWqQj7jNRIL
p1TkPAtEr5p1mNCeIhPPFKQFL4HJIjaTdUsOp0bzedytzm4bVX2gRrxmOX0OZwM0YyopWkTTVFln
+uE2hc4AP80SuMIXgG9oDrmjR1sAUSfiaiwkmBhSYZl1Zc/c5JZuqChu8E13RgncJ429KOPsvV2S
pfjtJ9jWyHzjy6mGyogu24EV7IcFklWe0hXECIBhtrCibZ6OZQglGx0OlX7oHf+b1qlF/3JbtkYH
O3DfJ839CgxCEms7CqbVG8Ak7a2GTOHspi1lW1/P2cxvm/bsb00kHuEKDArOR0hNlVhL/zk/RZIX
yLbjC6ErnD/gO2GDEK/VYZN/t9mMEl67LileZcf1yurVpvzuPpYBM1X1mXK5oZIDVAfd78c5UR1H
3YTguu44kTJ5KqHOdz6zKPrU3Ty5LFdcAv8VSXUl+JwEbERQ57CJlroZhUJ6/pBvEfe9Wyz3ubmp
KHviy3/Mi3dXb7708q66oPp4pJXPZx8O6ozEjBYGGSDTSZFSZYnHOlJfCO/MKRq4XY9Vh355w6Ga
w4DsN1c9HmbVqXhqel3MYfj8Dtk1JX/iKU92wqPvRZCWlfSLybPi0aWhBhx/JNQopNcMtMSGYRfE
jb9MZbbdh7S573WmBLcqM/o6PRzjbsmOgDwiLaG8+oHea7Fl7x8PqdZVbWYNk+TzEgw+HLVR5rP3
MAxSApfXhFjvS9S9RT68x5/HgQiAbLYDpqpUP1WZAZvL73zGvdWIZEiefTEw7L77dkcZG8JU2nKq
JlP2rz9DX8RusczePAT5AIsz0/9Gs4eLbMpsTYtOe7iysfjrHXt2c8zLse+tzogJT4fL2Tnhj7Pr
GREOyPDy7MDIiaMzRBHBY6x8mXLHZI1COvdbbxi7VD5cYhm8ZIo3PDYgrrl/5YTEQKkiMoZscBB7
yoVsiBQqXUqSGqsbMCesJTgGLKGgIJbQkW4Hgz4EplnDBFE2GwKkzrNQYagNAJVwwMvBwJtgB2pt
jDmhS3iIv8K2/e4mJdyrXJUuEr3SuFalT44KBoXOclvBPk42stQ7qInA97lFL96kjQ6e8un8A6MD
9fmRVwMN33TXsnlaUFdtOnnoj5XcBBmO5iHSrnCmn7m/usxDCnoqBmmetrBf7QvasKQL913H0oGL
oUY1N9CVhYrqx/Z0bl0Qetmo2OuGBxzUrDmkAj4Sro3GGUX0gMXV2h5LAEdAPZdN6uzIPysmtijM
kbRND4aNWdTH7J0+/79ZB1xQAl58w0jzV1jkKrsAUalpwgFwrBTExo05B9sNRrc77ebgEpYuottz
T/WwQTw70C1UknddUwTEvHZwduSeloaQopUgpIgo83BP0UcPZ1pjhiV5EJtutXh5Uws6MgVLLVrU
zDkiVgn9WdanSLVFtWYI8x6Bh5KQG6akj2r6QX56g4lKpaRMAKXbxMoOshOV+FjtJNutr0RI9rvN
6lotS6Kk5rSyoTQ14RGgEOB5NgiXitOROyXcUFA1/ldeVsZsYLPEGqMuqeoKzhyQQRiPw85YFVBu
j7EMFOYWqELR+F/C2cuElCPZhXadA7ZzudDxtXAv4qPYC4cy0UeGEvB0dtX1jEx3Wke05ctcero4
fmAMyIqZ62ITn5CSZ4vGJQ67A5rgfE+bYV0QfkO3ToJQYrT85kE/AaWaMFgPFvflUUQ5ggm9jvdU
kIVsuHzQ/kBm+5fB9c5ibYiE1iqVZshVWYoWnejI9qCGSNHFprRRNSycKX6XdE7AMapQ8UB/TT26
5tRFOc+VXx8VMwpbUJEyptJjzdM28hwfeQr7E2hf+2cqIeR4kwAPtTpxK6m9Pj7665EQTlnGs8co
6Va1hKyC154zo2NslCTskqn+iCamKj1gveDEoNbqbDBhG0kA3rRERz65JcvQHwKpVr9DcpHpvq6h
1KlTT/127bJx1DqAzp+VOwOMuoVbUGiiy4Tqg7nldicuuG1vM3ox8XcnOeA5QsB8zjWDIuVQN4sL
XYhVVfqVEKMELvY2dsbJ1c8ekkloAjH/OzxE6w39IL2XQi6NAPwTaXqnsl6l7mkkX8uO3oyOVq7v
KlOe/8wZCKDcCUeBOO1DjB2fnOTAJ/mxKG4Sm4oD6x4sIFY2h7qOydGfF7xHy3h8Jf79OOAqZwI1
ZlNi47aUVFSFmj8ZQ7PtsmRsY62N4QOZj0irjXPbgpJT0FHavmIYjUH3JLPtXDf2I/FhJXHgvlB7
p1oSd2VK2yVm+y5In/yFHfb8dIMoMWad7W+wh8QzY+1m7IvEI3O2VNPQGkaPgWnm3TnO3VZDNPdA
guphPjCMz5aJ7LazfPLa0RItiSjrFv5JOKEf/5g3PiR/vt0dEYqq8nCcoNdnCj2aj/mZgos4Ipi4
KRICJ0BVsXr96XQ+O5aGo2e9qTHHvQ4QrNGmVZqPWc4y5H7fF291qxfhS45SkpEgb00DQLAYJ8nw
v1iJdhYuHJSfiDheHy5oyHLu19nhrFNLiH5BcjG24D1bxTzVD08EjZiqdbntpWK/okLG0YL6h2et
1dELD5VLyIGYPbfRDGXijfo5x+p9mqHiTTrSUs1eOPjyHKaBjNN1aQxD4dK1WZCTxXYdQBemE11F
3Jn9Z/YKSyssAlw4AvNy6XKL2r0o5Wui58ENtCwW7P5eJlbcXyUXMygcwoMDiu7cMjel2pkUiZ80
DBjmNqgE7WxEdinRRfl6tD5Zlw83izulBPkc04s0fkxkuqVpSJHfVtsLLqfRUG17FWgvSVwJe8HG
XYBLyGm/zAHDOyXBIo2xpbMy0WbNxLFouWhS+gNX8Dbno90caWgHJzKHvcIFTsdMgpy/rSqefyAZ
RWdkvwcLjvV/upVeZafOoAVPxa9DGh0F1/Gw2I5mVPdMBomz3N6HVhCV5KQ5+Y+5Zf64A/gqR1zJ
UoV1zlWRDCpHoSLpTVG6IxFgTZ/o2IUdD3N7ODFMX2uZLh60R+F29kyqQp1RdAI79XUurPGRdWYC
WbiDtx2wS1yr+PlrPEta8WJNpcTmpGJsjFMayQhjLiv+uSCOTWm3jjm1dsOeob/VtZGnY8jn2F3C
S1AeGrh6WVUsAv5u/VhqCB0Zu7mLo3OH2yKsqvK3VX/S2PfOcTw94sCTIqCrPWJBg2ONrbxDlk1C
YlRV8VJ/+J+GzMqmZqf0H+mArO0LnDzsVoUDZ2c77J8D3yjNFh6eWx4RlBErW/27J1uErDWI9Jmb
qD26/JGZsbLQFscHXOLc5DC9Q8beUWkJQzznF35+yIqi9xaRsJxg4s9Etd2cfhR/mm6L71jTz3LB
o1hfetvMSG+tpiANXjNBs62eychObsnIEIs7DMk0nyCVvyzD0d6DTUxJZ4x4kH7LgwB5mHGkB9Nb
M5HBW2qrZRnwoONXnY8MP7eQqjCApDfUaiTBfde/ix6/FRgSnO/KEbDELrYAKdBsGlk1jJnBqTKR
/5YbN1+D+a8WZigFqtKtWdgVXZwbhSseee//3GAWCbqQ3c4HOEIkzYurTp1T7Oux9Y2cD4ZI8laX
fUrm4paiEo9dkCTQuo/tXn7ifNtpFwDv2CIvBeeHQ7wU+7x2SbxG4zCi1JdTx1d2xHyvPtKqXJ0z
O0qvByc4NrO1aqarCZF31Lp96VSpNQeMGIG5ODYQ2JD7nUwtL1JmskyyT4sJfI/ft3I/ENAJl5X2
MYOKTiD2gajPEov16f3EO84bJNc730M48W4ZKQCi81sTWpzGMF8EDH1cyyWm5r174tOvjtTGbvjF
zH4J7EK0WrKXxh5Uvp343EJdou0APQD7868YSHYdods0b/S+tu3o2VmiU6b9YOZ/MojOAsED9o0k
jpw9JGGglCarDgX8M+vR+yCv6g66r6H7sXDpDSq+vw2NnNKWMndz20edGhjk3K3BylTHWyFE/LUb
roe/C4eE6YjFCmpZm6WuuId8da3aX9AfK1SHJTeFkZqSWeqEz3BO6SRnaEhCj4/hD02Vvq/ZyxEk
ON0kViJALluGJWMx1aAwTTE2tRA+7fUUn+IPH2jdug8vd0SqOh2yfSQxSpJVjjbgvriK4/zO/TUq
nvSXZR83N9eKoiGl+eur+J9LPq5BiMONZjRaO6v/VJr/mduqmG72Zpsu+OdWJJERL96em2hNoIhU
V7k/05Zj1PqtyPVCPlfx6f9e7UVlGGlyoTLRvJzkuLJS5kyqMhrggw0BUefGmH0Qcr8mFHjFiKIR
urH6CXLRpaTjsc3CdsbMRZHELFJ80cWQ0mJ0IOCKGUTsT0tpprPamRar0cRUDSQY/eUFxDZKc57u
h7IXeGUyya5DohkSUSejfd/B4fsqE6DEs6UN+qo9NOUTByTg/7cmDae9kyWPQL8YIBddEAZszn1f
UF9RvkujvF4JHUdqM5sd/fZ3WhSFxDFyjP60XkzMtZCzUqW0IT4e5Rbi3ghbGMs/JIMcLOCMtJYp
l9+yiuL/64rsZJO2J2FllsjTfN5pHqJ51xjnLAYEW7XiUMKz52b+khWguHe9p7lJ9fW++oowlGqj
1FcwloXfrDuvGQFSmc5m6vcIv806M0ONmH/s9JD/MyFUnh6/p4+cuDWUaLDHIn+b5ptJdW2x/EAJ
LIrc4B5OCWoCZjmeu8Y3biTcfCr3f/Gnx2pir6XmY0JjOvawcZZOik3nA2ATHgZmt7+A3wkp12YV
h8FFP6M/08EVrTUvRFALXiR+BiblhE2e7fCaDdtMKGE5v6nOhc29q94KOT0SBPjRQ1OjwVBvyzu8
LWXNKpF1gJZfX/7oI0I+m6zpPynJTzkizOJSXWRtKJRKgMclMM8ICXVqykQ7aERSE/R7OkEs/VdJ
lWsctLuCg6suRj/nC4cDzzegrHQMU3mGao0kMftQK+vXtvZE+j95AjlGWiSHQzHRQZAVs8b5T81T
bl2BFvync44N0AkMJfsYfkXUT+ZONXlZlrH/H9xVnGaj9FvVvDUHBbtKlVuNHJGs44/iwfgoQj/0
tgHe/XAL3JUoZy80eIy5V4i4UhofUWD4ChsmZREh5Jh89UdSz5bXzxWN1oLU7P60RYlqQVBk65W5
/dOQtoZh/vs6fYS4i+kxiP925dzxfCXqhhNu0IreSOHLZBkI1GEijFTRx3JTtOVX9r9ijuGGnJw5
AhJE2hP6WA+vyDbZKGzqWWbk/4Be/suXAepPZso7K2+IPT2yNKJzPrHYKva02EIBiaEGiehtUa2l
XJ1Ldo8eHIYde/CanKkujfcierdt/CWIlx47PlpKPN1Fl4F2uz1aNwLjDPzCFer8Y2KYl45FHl80
BTO1zBxPugSnhrY3ZzQKA58WLotIL5thjaFf0O3tkKn2hjrnbSaG13Bc60jekgjpIDIQjokVmZx0
FW6+xz6GAcdlIZmmwJdZ5PVDM3h/Utrz3Esx3skA4dYP0weEpGFgh3+l+wFs/5DVCeXCO+fI5X8r
cptn0tAHuEqEytn/5d8QNc/v0kwFg3+J+DGRFq2i4rT94E9hQIHxDLx0Mn3Y3GnP5aOzCqhf3Cr+
HoB1KS3V6OiagxeW3iR+ZewnOSRGOwVR05C4v3Z4s2HQf/A/w7/r3wYiafOkdLKebxWSygSDiufw
/WsyoxDVhg1BETcKKFnDDngpGghPb5hvr8UCBMI4NjOsOdqGU4jFq4zZADiAqeMjVwNwxDrqdPP1
HIK00NzwjcBZuwZv3yCQwjqiaE+EMhb2ckN9Vpdp3oQ80tZ/7YrD09EPibOfTWcVSjKcBLomvl3L
XqsyyxMUkv7hKQ8wQTjYkcQMX3tvwTZxecSPLOFfvXtLkrd8T0bXRIcviRf0ryuFVyZMfNMjiWFl
RgId4pmEwyFSA8VTJBjtdoJrCj4B4RFmz6OvvSKgnoZIg7fJEDGKB0rOmfOIPV1veo5jGmIVeS9f
Mw9OhCB0ixVw9Bjcw8yya2fH/mhBiPXvuKP1oInI93dmVwGJf29ZRAoq0U4cAIL8EfKl766b7gfr
cLrhCqCcHkF87eWa/mGREFq43aYRHwZpo/D1Wl/0ju1Jnt3od/IsCGYdU+JpIVQkwn8HJn9bINuJ
F2sqnD7YsVSSK9js0AxbFy+h6joVXDgRZUNtGP8duYkN2jFMWdGYtgimdPMqlGZ9yd7TX2kUUdkG
gFYk5c8QHMXR9idcMphwcn9EsJjJc8EwE3Iqk/OXK95fKVJEs/caIXlsHrmnoPRc1glHuEHcMgId
BPd4dXKnsQfg8eFiO3se+RxZexBUQvlf+9MAD+GqQTXzUbR1Pi+ksBvhYDAjub93XSMQS8eBNG6R
mQTtdoRRVXigV42+mkaVZDhwMenLJKcmBngcGGWSnis1kAmsTq9UioRKTsAfplXlfonAmvI71MB4
4JgUadBbBfxLd8zZlYOoC5h1ovz/hkd4kxkqgi4nfGSnKtIPEy9/yLQYHCT5sOV3oW1NBDeuwjfn
0zzDHOF/wF00KMy6/kzlNzE1dznc/brg5Hs5+0UU9GJJZ7FuMsVqpL86ZBWr+u6ZonBbw6jbSkr/
Fd212FSQluzKaWNS0jOJc5C4G88kc1wkNdu7GuQFCyJbTtSI7TP6cMTPRufzhQWOs/+eEvQ4Drjc
mfO3cN/AXjg1wmWKCkuvULNLigM7pvHA9sgbc5LjtHfDFnliY9fswORrx13AhZVJUDwuogWjV14K
FdFCXvxIeKdcyr4o3Qk6q0PlnPudfLUoWyUnAkK/qV6+cMAAwGDfNDzjbbz/hs0TXq34E+/u5i1A
8DuIGVqycR8DNATT0wYsA5q6qBp/ml779yHjZJKrkAtU9StJxjIalOxEVlquN/mr9QPXBkHBEJw5
r71Mh5VbJPMyNCfClmjprRTrM1lQTjYKzH3HY0spMgG1/dO1uWzxCgNm4YiwaPxbmGfQvBENuPe2
je2gFVdPUv3EymiwdtZEEtWKb4Kiz69uJdvwUVsOUrKCPTe4At0W0p9pnpgstLc9GaXE55OC8/Ny
8Gb07c9kjndxAOhqpyWspcI1dbQcakRxR2RmSjFl8HzdN3vVZmzODdpbDygXhAYLEuLJlXcVcjkn
+64BGeCpA/9a2AM/ziOFMbL+LsP9SCrmsrIPPiBFc6/t4JzFXstlFc+EyyT+uY0UKEYdkbIcTnDy
heQRLBbypPJ+zEN4InlmPYWook6grI3RMWmj8Y/6gZRA0PYbFflswRDupUjykz2Bx2WmpNh59dzp
lIjk3H/M/2PEepgPVgGbo+tTuAeI5mSOMX+3RvUAXWR1pJKh+nVxDl4b1q/rOgWwOQjOGVnrtP2r
Q6sVSLXVeiGpO7y6f+02qolsy8q6qdtKshx6BIz8PJ8GmXhiUK3rihSrYHbZHBYTweyuHhsyDQy2
W6EL8+tAX3xJS8zK/3cujz128He/lejcUa60fepSlOKhXAx2k+BYKuf738+0VEcs8fSuxy+xEHSU
Den6QyadrjSDBqxif0dknvIjPFgSFyFRu+ZyisiaUuUyy79xaKDI5zlgbY0VYiSWW0wrzwuDvhag
B20cB+t3nCeSg1GaI2NRlJYJZVl35jxW1iwaZdJ9b/Mr+lT09ALmLZLOMTuwYaFq3GoQwNHGmfI/
444wJDrhLBt/i0wDpNX66OCgwfB43YYbORyYDMcnJ0rZYqkmsNo2qBYOWUaujlKtW8jz/eUKjnTw
Nn5GZu4yhltYBA28+Ig8JS3wCPePuMtBN96TTqrVZubHUJE7Mprt89WLB3/K0qq02N1bpmKMTanZ
VzHCW9nPW6HRY+odFTyD8QFQvZnc4XakmY+YeNSrleTR8pEFgdzTX5YtDD17l9AYEQvS8c/hFNhe
IXF9SnCb7rXymUfXQRQKYYSqANUBpKeAqFPp8iXTJKgH5K91GVFd9GQ6tXkOgLPN0EiJ5F6xyEIF
vREk315KqNdJrPG/ybRGzVkLpqP4rytZzLceohG1HyrmC/pvw5ATpXr+2QM2H2RJmJfqf+H3ag56
fXo1wkyst6d+fL9Ze4av4tbxHRTnMXb2jmStWZeD4T7dMJo8OvdFO1g13O98Jaf3ml9WNHZU0P6Y
HaH5FU9g+a0V4dGfoDdH1fLfCuciCV59+tUfoax95SC9M/z6ad0KLgagqBzZjEuTHDVx6vlaqktr
hXyQ05wtKFshSU3szxUHcfJm2WuGFoG3ckDbSa225yRHsmtjiJCvDywgCke83AZrSv2nR2+rURNS
598nxVaDzOeU4MhFuHeNjYplYbI1gkW2HKBkwbG9PE5LW+eGsab2HwHh2ECS6F5gPr2IO5V3QLcx
3tTRlrPJEREXBFtK3v+VtatsnnlDiz+4xy3eoQpGe24qfqqEY8B5l4QGAb4c+99wkqz6IhjYj+pa
WsSO+7PdJqPRaQ+Y5jz09TuJU1lPi2OVvqZXXYqd6B4e9oStsogdQffyaRzIlujyG3WIh0l2gZl3
O1DG2hI37LIO17YDORIHEEIAj/kB1tvHO7V3DG1cdjv3mvmTmvd4j5ALK0HSB2DBGf0Mi6oP9FYr
zs4FF0/2W1m60xtOh55qjLzzNxt8MRXqbhowIMh6s7u6+eiV371G1J4UB0OvmKpr/t3xHVH6OMTd
5p5jrmPko3/ferJiexYCYD5KzvYbMxOc6fBQTONHMZ0axQxYYo7PjumpHj7uTK9BZGwxi1TTMA59
jt/QDnDnZ48rHZE8wL1t7J+Rcip2lzK2vV8e6RLfeWdgXGgcv5QMBedTSesbl/9nB/9m21iWRSA+
K06hlgz16UGLhxkHO4ReVUxy2YJyXgH8v4KdllkzJTnMK0cQia5pGyrCDz+TU6erQNRgr1UCJRcs
9hJV1+8pbQm0NuYUZWnE3iVB9eUtFXlIoo5Wlj9++BqG6PV2Ugw/pBRtPi/YoAFnLuOFJ1QGpPGv
IRKb0tTHvi5XiFJaoLHEEFULri0Gzkgko9CxUkcUEzfHEM7Y3yUNw8RT98FMefUc9WW4Fy9datEr
mWfamI4mCO+TQzRJHozBKdgLv0HDaKBU8GQuCNFMm3ryc+o3blQq83qB+G+Jb3BegttE/jSIa6VM
DR7ojFNph/fyO7EoFSASbO2QUQKOSNRXVkkocXjyNYpHYmFoH1XK/Wagc4kLoJP/RisoXeIo507g
0xEqS/gr70fVSqqS4JG/IOVdYIk0z11dXZ63tdX8T2N8jfQM0UQ3eiHGheWg9xJmzglS7SNWy6d5
yODHXFbap+3Xodogn00WFDwKXrhLlpIZiioNBoCZ6l/LueUd19yNEx1upAD91Tqc9k/KZn2ImthW
vHlMXtwk6CGdEgZfD9lZcMkQLqfCGCZGnUq7J9Yu5Z78rEI3VIeI2QcbXYvSO8zJeoLknAiinZ7k
YlQj1prif4C4ZbNtijhORbgMU9+AOnchvDVxyU6jpyKUanJmBYYvnjDNyozqduc4nTDQU6FgnHvy
ehSIkJ/yi6hpCcln9u/sF0zHVEkwoQ4I9NnyTS4ohs+CXRkYQPjgvA9ZZWBFcAZbxBY582hOlq0f
GU5VkRxdqv717KNXFB1TeBmowg6VyvZgTd83d1LtoOzlapPGhrJzzbYH4FlM0CDCUP/w29uIQ6dM
+aGQeEiV+0eoO8qPNe1zcayUajccMKoByKyI4icBrLy+uZXy0tMSRDk7Kche8I1PRXBg2tJ0dJFh
xx9nwX14Gpy22NYWEYDt5YyFXR14EwG1uqPPT23nUBKnpKbvM4LfaR+VfogeaOwb9tgEdfQUwhgD
9SukbThB9MmxIl6QIGaPUY6ekY2yiFIhRAL9SdVthqzEdKgrwpzMYXmMjpDonHSPMZYIpldDbFbu
Zq4vqekLcXN16Vo4UJ6/j/UHAUovIO663N4jU38cB3rXeYOoAKVcwU4kILKVRmm7qZSCWy1HmtGc
VJ2DcnEY8903zhemZVeAcc1BhnNSyOIXrMGIi2EjISQNVk95CjX+3v05aypJjfz2gL2n79saKelQ
fHjoloXvDFQXBeUxHGDRggyVBBrcZcz8Zjxw0RPhopulE0m4qJDGlMQCBPFS7g2BG6kRDrfgvjws
p0h+vylW/z7rLH2gWItIAqtzUeitQkRZMD830EOU+fbYa5lq6QWhWmzqx8dCbZcIf7PbdYkg8yv2
miBs3duI4bYcRLQR0X5lGdAeOc6IiiTFS6Q9FkfL3s7yTKmYMIe86QQBJaBN39WijoeB2k7cjiXz
HZM8Qk2VJdXEatvwoa9voqd03QDgYWuDnaRJ+fh8hXwl+FQLnhH0oiaTKWMBomPK3mzEGVOt9+Xb
XCrSmjv0qDh9ILpfndQn+loDrEwTTH0EHa+fEcj6jJjXR5s0TSurCR9cPa7w6cBFWIlEwZQWhMQO
VEpmVXqSWo6HZM3hazCOfcBIQM65lJHjw/QR6lW4NL32dc0dT3Duhw0Ki/RnS718KRXtDTaVn0Hf
orhIMAuHclCpoteZojbxlfzui9UFDo4l3JZYDEUMb0A03a3WFpGDbnambv0zAWra4ZVon21mSIgY
UEPgiw5bsiU2A3aGsYkBuWfnB2RnYzbgYBJEnC82yd9ctvrvNQXEP6R7r487r3VeSDMUBHrdGXhd
vqQjHfDwUVYT7fg9yxHwllIitTLFZ6+9cJB38fsyZm+VBHxfzVQdv65+qVcOvtI5S10CWpfhlH2x
ps9J7QsEtCXaq6HMCk/Z68OAy1XvcIXw+oOzNiVUkIlz/b6wpSpT1l1UsZunl2jN27oEk5tWkUuH
iz6tSqounktfw23gYcGzDcL1wP+il4YlaImxVG3E+kUu/VZt2Z5PZY4rvqXmzaakAbana9bRGAT4
mYgOzzLgy5HGC5v1UaFxjpR+z646Usi6iJxzAEZEh8KkPud3fntEwH+CldWl10qtur02L/PC6QeQ
4BCZI9Bm3SwKXCUeUlAinhrD1Hv0Pdy9OVCt40owkymb0JS/Sy+mCfyhIsCnQ6NGBGzG21fFYvHC
3FiU1AT93SdabIICKMl15fs3IE7dpinTEj5MxicihrFEMXClZpEKwIlI1+4jm19RBYCwn306Jpos
nNr7beNw6OPWNTaXzLilbYYcj9yNckhFXPGL5vGbi8nMWb21uYFqrZuZncLT7icNsWdQBUD6UStY
YYJuXSTIqrwPawnejIVVNc/diKBbAlOkAubnbqX5Xy0CSs93p1cQ0XTjksRdmrbiEUlc3CSLz12w
VQs5MwaLG1AyWjvV6ASelozNsi3L4kpbgx7w6evtZPcMdf5XwI9hiRp4vTxWhv9aMQi1VDz83W2t
zZ3YUo8FO0vhyJV9uTr9SEAUfQi8+mCbHrxCKn1SM5HZecN1BnbRhYRl1POIsHHeM9WE1Z5FvxTn
wzBEkRNQiRcT/I8gdSwvvAjtQeC17k28oj9aPuJfwLRxlZIagiPctp24GQjydw3j+QMciqYQbhUC
8sHX7YkBYJjO8Ocj07njB6nKq5nDyg5VvmUzJb9RAzN5GYF8QOp1TpYF+kTBcRk3w73EJ7aq2UfV
J4zRHfY1Lp9XtMDq28rZhoU9lR8oPTDtI/miMPxPcJu6LiWgZz+htLTSfGLsljifMLH5xj8szkvx
bTDWe7ly4oGdtlY3OAcpKWGrzy8atxrgZnn3QoxtdPqErCHQEW44dxije9o1oBud9NQEgNDa4mTu
24qplX46uWNcxBYGD8U6YeVx1bKhuEJnSqtYsGFvceVZTnkL6pVvr9cQyl33Y2vDtR7myVMTkvtM
rHlF4Huvy2d1A3sKk3+uSF1Y4yn2f2DH1p6D8DnhXhNgqGAhrqvLd3cLn6JR3El1eYoDy+7X+aIl
FxLQeHOPCRSH6kK87tWWoei2MN1pQIBSWYJ/RBoKmYwiX0imHE2+Z3g+2uqMGOCxjcemq2mHGLhS
1oM0iPLIqUHeKNgKJgHCaRGvlq+OSmNu2feqA+L8RpnuzIicVL9HdEYW3MWoruWe412BCd/XBUHk
LH1gKDa7xfFgIWcmS4dqvgi/LwBkKOP+mx1B9XSSSULWg/g3M9sJCSyTYA9LMzmpLKiR1Z1XrDf9
95rrhW1hTKyF8lOtjOLagdYApbWx8jvpVdJK57KyMcoU/VRMJhs3wfep3medFng474jtBv13lId3
bj21A/7a2CtdSqagAgxrpNEXxg0v3OccD8Foh17dhEhWgx2ICqrJwHTeJ2bhN0uwVmqZXxZeJuz0
xBRTLaeuqMLBcHl//dVKXRyUZ1DC8pkXxHlJ15/JgbKBq1rc1I/KBKWG9pojQgE5sTU3EWJDZMjN
IzkC7nsB8ecJKqnXcGSVb5nf8wvAlJ8Ub2Lm7FRFNoftyWSCm1QGc6Pp1X5Iyb/Y1E2GoDDxKEKc
4N40oTKiuB27gTqMKm5Mzc050Cf9lKVr/hkHp/g+jCwmhwzX8P4iOkZLQzOZB1aM0Vcf/grnuvKH
hoB9OD08qLsUPXJq7z7XXMhnv1l+Z1GhBi/JjvmYsMuD4myxES/zoB3hFM8g9zUCvfbEIHp32K5i
R44UwruT1qmcTqUzWHxqmENhxIbG3QB1urQ6SZbg1rcD+t3HWo7xSE4O2X0jpEgp35h9PngNfRuN
7PIs/zYnvC5zPgNGsvEX3hV5WwvrZ+TBSO2rJriWnB12PVE8BokEOVj1KsQ86+bvtUcTrDENiaKA
oJUerWsaeiIUIg7aCzejMc0BJccdjIkQmNWQv98oZE6mxVYweZVty0EV9NuNkCVVy9zis70+DDJ1
3mGESXjqn3sYjivUeuw7ofjBHFH+R5LMoIp/MH7u7NumCe9eDN/GOVm/1O4RLWGwg/uNUdnaZ/68
r/IqDCKK7RCk0xO2BdMSY/JEaHHaVlPgHV5XmjV8pF5q7ldlMIMWXerhjteWCbNMmkCbxezkf+Qs
RwFO2wKQGUcIReLHESkoKodmobQf0wofB70xLrJQpgbwnjboiss68zm+vts1ldLRBvJu07Ti9/3j
x3MBDfssIlM5S5dB7jPwMeIM5HgxpaqoTtVcUJNy7tyy9CKgzDeu6tzgTZvkbze7Mn1HNi+222qI
xTWrEDMtRB3+6CtxM/iaUdtA0WhU92p9VVu+ozyQsSl8KSbJmTwMI+MyIZEktNny7GCgpP+Fxr3J
rf4qhvkoJui9FaxPYHRmtMXP3Sch5wtNDTKYqduNC8gW5ztblLybmv2K2AkdPnG1gXBy7Qto28l1
1zA+mRZeeqFNf96i9K9ftAwgutOSPHS+FbOIi3uQPJ0+Amm7SJ14KU0XpsJDCvRUq1owLuuD7SET
mIiNKp7B8P/eeSkrD+OzRlbQNJF/Pq2ruCNlVl2ScN36Vdvuqb3HJ5JaKiGFAx9vSaZkGMkK58cc
UQyMPzovwdllApGQFBwfRcRRWf7zwJCLRAVu+R51BrsIMjjSyB8O6WFM6CUAHlnbcfinUysirTKP
TQEM9rPZGW5S5chvDxsVH+kNtAfcoTdkM+3VG6sFGn65/wA2EIAY+0qqukh/I65llLCtA5QTPzM4
DDpTyk30eiwlZVrZwvIm31y8twZS2EcC/QihRaKmRTVfJgN9arFkG6VTvOyQWfiBLH2yHt51oht9
+I5g/Oz3zp6WQBM1yfc330IM+5kSWYeCu/CleSXzRegVh1krn0pqkkezfvmYrIcdLOSGzDOZyvgx
XkAmLbuIxNBqrrTggpTGg6XSLgIzRZdfKkcNngAW4wcD9ZjWkj3fQgf4g5YdBACrrYXIkZv4WBYU
IuCh7uLitZzYmr35rsi362IWEoZoIDBQ2EwuSTRaLDPRrDVziU8CdWCl53PFBzE8PcN4W+a/mt6w
KTfSIt+6LOLu7vH/UygRTe7j+9yXDduk2CP3aCH4wCzf6w6T57I0Cidsx+ghSnM133NpBu7Ews1/
wk7NCTf0t05jGmSG00mbX3W+j4FDCfw4n55INaiTYeyu60NlXUu5+M99aa45wsOp2pT3TChDmUkw
9XQWQ/0nYdxVAPhkW8yoiiGfSE+uebTSV/vLl6iXtvUv7nBYAOz4FDR6o7I9TUVYoY/pJIEUvvtQ
B2JhRNzYOpgURPn8im0o6cx8QFSoYwXzQHORimNssHADPpKO/qwlvmWQt9jZS1FvcLeIi6Qx8tcq
xem9FZT2UrCFjm7W6wkeImhqJDxz6VAdWH06ENhoOt6las59JpnoYdWKNYBvTFCyi1Epa92xSJJB
LQhYi+IYyo1sHjaLIR3ziB8OzE2cp0VrB3SVAQQyjLCDqDBNefg+hmVbl0OGG5cfCsUKP7ntYvtB
8C7HX3uY8U9C463zmogqw2LYeMkXWNaFpaM5wvr8tebNrlfmFnhyMBj8co4k6NM9nEM+WDKhjNxA
Fn0W0YqbTKn64wVAiEieZMcDN43hazwggcrinBd5a+8l+4+774OQ5P+ewbL2A7SVwXvy8RanBpiS
6V/jL8SjxJGf7hujgZhnCly4KcVWbTVI5t6TxN1rBtCcAMlvCIlT639YHsyv5FnbqOvOsJEcLzk8
/LcPHvd4uvdSg0dzBdzOZ7p8wJ+TFJxcQwE5POZoYttpYQPHV9FaTJu9uobrtu5Erbmr4h1p4WRQ
P4Zpxjli6hJZcCpfiCFUHe6NwNh9KUWK4myVvIZhBFlamYHeJ5Q0epsULsIIxA4RrITybIxYFVTh
VBaSubVE6sclzyZkwaxmp/bVOh8yEdUiOROGIbGRcmfIEnLMn+a3+Td7g/lIYbx+OI5NaDHBmvK9
snqEwf5+s5uTouuuto/uxIg/riqs27MYAjbkJph1RRjhs03U0qAIu4Z7t/2KDG4nGWmfrWWBPDCR
EGKuirmMru2mVtm7BxJ/TaAjgIfOyupfk3yOsSN+QNeP4qVFHJONsK+ueF8Q7OZ8F0V+74zl2VsG
65Q7tTFlZJZGZx2OIWm6MF84Z38ssSxxF9n+C0XuH4YTGBv+LrSa3WdnFnaja3d9SqYH7mYSsiQ3
xLCK0F4YEpnYVBCVPIjON4fRD7o4exnIxzy4v8QwZGQpnFn0fhAUZ7rQ6uVuDb/e1NwZovISaQ5r
KEJz8Fbdtq1b3Ce4OcFIYNsVTTLS0vczpDzjL2P7LLuQRIKT+9Sl0DORuJWnR+yo9u5BCazJUC97
7dlcmTj3LAOBqxufCY6bpOLsDBXeX87PAseTCGqMF594CPRAV3gEw1VcYIawr3uP6OwXChiRJkfY
Ls3NZe7zrJRE7SskjX6aTpz45JQbr0E6icRGUiH2qeDTCCMKAkfXj9n7YYghC5EW/CYXOJBfhE+L
K419qz0zA1nv0jOK2JQreSzoApSsE5ay6WSN+9vKUL1P6TVJYPdnug2sXILjwTVEcMrEHIoD89H7
T8mzGGYugJF/p8wBfDDTXZ64QIhK/6vD9+XOE4WncMMSmaWgLcQ/944PcyDmBNk69n21wq3LavKK
q45fUFeGUHlz920tph+O25stvxdVe8wKjCN5SIX0qxf0vcZUSfHsuCvdt95BSr5RHf4QkHd9YYnM
ieT6nklK3PTcROC+PNm/sk8rcdOjF6nTlRy57dXzwMfE6TugmWNuZZgM+obzorHoIFGAuZz/Esa7
J2yRAzWsQjZ7dx62AA3YtvhlPXJFRlgFZ0meTlD0GDp2iPjXrIGTLA1r+fUnZtscGr+smh6nZsNL
JK92yPEhs1+YAhASrUYDKfGtCFsGSHawfe/O4dge69f7EELufqNY8a+svobF4557QvpyjCl7KDDT
mIRZS8/yvuahjBvwiykFlm51PMnhL1B7ai+Q3w5rB7/mLJPAbFrp/GGHubhrbd4D8l6B+RYl/m/L
ALCVFGC02JSSRbDXCUuIaZ+9L3zNIGp4chUgGYWOamYVXXxjrm6k4xIqHzve3xnea9eR4F0uvKCy
+GjpwtWHGib1loHdB683Fd43B2/z73G+nr8NQ4m88MPBCaRNgO/jIRSMwWqEy4h7N31KaKJkCe4X
4tlOqYonayfpnfiTsDAJlTGcwC5S/BvuC7liwQSfYxfTOkLzDkEJOdYeM0h44bn1TAm+eKvz03JF
2lknGy+ras6dPNkb09MSjau2GgAwu1v0u4+RRODB11Efws8a4BQzrLYFyhXLDP/OjyH8SLVfcR8d
hotihDRA+lnsnmgJ5iur2m3qV9XQZpk45xZ7rPlbOqVRfHdWHw/kmekYt9IKJf586ftkI3LlP4xB
a9PaixNtaIy+KaPCu5nBIh6EXGy+/6m86/5rnOypEM0GWWOgfRrNqvn5qyVoWHyiSzvPTLSSvyVl
Jss7ANIVe2TYp7gU+tLWAnZ74YgZBPC6hEn9GdFuidA5zqdO3HFtd1et+APPonl+QpVDEi33QlaG
GwBD2lWyRzG+TCDKP4Ik6X0S5G3ua2zFGa7WTTmzpbQhvEaAu2Vg+b+NOdzus4j0s3vgggbNdDlM
3QKCR3yE9JI6sHUfYYUrKPemyVmtPM9WhtuYeFvCt//sVnsJdzxIvNGxlcQ5RDLGTFqnB3xMNZlI
Rvf28LSmBMzrarswUFuDeUViD4NgQ2nRPp0mHnRUCUJAwWbc+UCKS9UQ45sc83N7LlYbT9z2kMK+
SwkzIflG/9/1ummiVia7tsrmcfLBi0zYvquSxWqrYG5JtU0DzhhLIm3wTKVxNk/1HHgNbzdVZPb5
sOr0V21PrRl7T28pYSxG+LEkBTVmM33HGQW/lFFXsJPd+z6rGBrFIpM4MyO+51Ijv3CoO9wg9d/y
e6BLg0QYf9PTT6BCnTwZIRFCgIU5PZlMNT3ofDTDjBS+NCLc0RIE9kHg6UoISNRXIA2Iv+9Bq7tk
Sed4lP6Mmst8/VvwsQdToqIJJOKCgkOqfMIwNh6uXnGZyjxmHIIj1ow+OmLw9hTMmdAUejFDaXzJ
bpQ2O/P9DflH8LhDKum/B+ySSAYAeHD8hXdm7HTJkzGGPkzAlojcQaSl4/oLAWwbf8jMWsaDJi0g
rCj/bc90e1R/7pDwaZmT5DJxCQHzB10gn8KWTitIF3kClHfDD3r49o842sx6ZuAIurWPfGPwcS6q
rant88ej4316GHuFU3sOXVGpelZdRAl+Js5YWWFfN8xdvoIcf7dJIij3aqisy6v2itZp4IP46zqs
MHsaJlxARCL3NrJDY5cQyjo21wufg++tMTNv8ik1pHbNG6lXD0gI2L1zwrlvfAM3y+QHLp4okqgo
VeFWGkQ8QFeyShUqeiQcsB8yPWa5L9CYQWtXc+wGR+hzarMpLUGrjS8hkbiBOD77VV9y33wnaCbw
Dk3aoveZNTcq6moJeieul2IoU0yQlw1um+1CNOJW5OOVtnpArf0mXyY0p5vXesTiaCzufVguaRn8
AcgW0/Rn8JZY/ccrWaLeUCco6QteXPNfkgkrMwZX3emfJXXdcmkEz2fuugCdc6tC82z+e0OUIlVl
uhFpj4WsY44o/sBKe3e6f1qYLyppr2LD7nwihXkWA/AeUaTI16WBHauy0GPgPLhO2zc8QxmWumDL
AETKMNQJd9O468t5HFlBMKoYrbsHrGoYClHhoPDfR6LRxjsh7W9pnCN+Lw4O/LbViJjDvvQfOqsu
OU2UBAWDq+5B/AOqTm75fZYdeze8Ne82hw9Jj4f7mMoa4knjE1OGB/jtFs0d8rEg4ulQRCjtYQla
G0w2lEP5Q49yHsMqCKpLZPCgu5Ns9NNBg/BpsK9kVPQiAWZ9ThVcKB90DP2l9w5Tdpqr+TdM6Ghq
dB+Xo9SlOW+J/DVLJBV0zNI8tIJlvVbLEngAIDHDD9ziCmmzj1hOTker/KtLt/IRzDzE8Q9YeL5P
FrVzFfLOhqEsEPiAzlIhqJIpDKFtmM+m7rPNjoyQkhBRi0EvdAOyW7wWXherOk9fa03ETPsHyGtm
i6zh2CAAct3P8QftPqW9hKpMkb9GgLA2weJNXql94WAtDro6iPLXGyM1DJDIMTn4oveMQhBBq6SU
Yw+HGeIzkbzILxzcIcRIrNZEHvz+7MV19S2VoumLcPyWgh57qEOzgAgjtZPgAScbjDIvFiKdU0g6
/1tbS/RAwTjEfkMgddSJek8PjYGwYPuhkRRu6iDL6gJhSs5m35NcVd7mwl10qaWahft8Pi4CEmwu
d0AIfyX8P2FuR3a+252PCfPqRJi23YJkeiGAsG4XnIchGzSRHwK8CXAgmb/UT7d88shrEQ/Syk43
M3d74JKG1F4FMF3PN2L/KRQqLr/S9A8ijq4jXJxsxuPkw1OUxkpWUkhoSwcisjxzVPdFuR+RcGVI
ejs1kkmeVEcbcXF5PN07wmi+F/wP1bOu6OQvNGFws6V990geqWtn3/terftWHTJaS3rVzd4nW5Zt
fa2l7U1PiXc3f2egP0CK7x7VcABojAzSMtCRZtmQ1OjuX5KxMrCaj/M/ATQuS4mRE2CPf1fLhOjE
m58fdngnfYjxXM1abrQXSbPBKzDFvaLJbx1xHsbzg1MfuWpddCJ5r6FSiewkWAjxH+VWfuD6mROv
gXp19kHXTsYtJt2Ka2S0e+Oe2aSZ6+B9kCmtFB2O4ggRMvP3cM1VUnuaU9x9c1T3gJQsxK72iKQn
5cXLQltLD+2D6WLpfD+gkShLC0pZxkWV4oxV93KUlhkzeShaVVjFox9InZy2XY69ZDLtFe7WJrVo
8ar2bvUdFjtMzE5o+ORbx34o6IQp1cHyrjD9LSrM/ZzsxFj4Hu2O3ybfnMDO1KERqeB0De14cmvg
QQTejqUXc7lDohQD1AWYdOKDBMwMjruem6EB+SuGZ2PohK8147lPH+PAwxNcxfC/vJByfwB1BQGY
gddkcyWxjf/nZY2Yu6yQaESIN5HKSsPVMc70io8VuFRq+NAvbFJJ83z3VcAyttvb96eqe7mtcJK5
XvBv3cVc2AYmDpkD5g1Y3J+eiYyNHr6nCCuwZBZKaLIdk9wRgXq/lXdv9ZZFAbZBLNVScPRA1EaK
etOOe1kXjrU18kcUQ8aKKBM0EtL4+FiXBzOd9N7wnizGXRlTE3dHLvtH5SRuSSG7zT5XJYe3kwRp
M3LCZUbMsWCarrhPsW7Lx8dhn9JgGTevb3XfO2crYE0PcBr4SQYLCAjKZTwW6YwRqG182Sk6QQdT
G6Nr3nl1q4zs4655Ymqeya0L1uzooL3aGzGBeilAotd2gqAzYgTgPftnwbQwTpzQXzpNjYzCMaPb
aFJPEdqokDgjC8TOttK52XvAtKG4ISDzj2Vl2Vyca2M0CCZemyw57yVZxuqbktbQRHaJXQdV/7zA
/HrIV3tvpWHKYh9cKC7QL/5/nAE3UwekqdCbfs9rDvsCEFvzuOPTv6jx3+H9iwt6W631yTdA6B8W
KG18ICG/wcszUsT5ww9V5Ni1F/XoO7mOz9cyyIb4qf2IH/5N2lxzfu2AGhS5Y8blHCw57IsD75Tu
oBG1d5Tb/i2aiDMA1yGXWhH7iFz3qv2cJXBtvwzO3XTZpzZEPTpEt2Dq4REaNSQKl6LSEgONGYTi
5cRYwrwkdKzHRb8MfitdhtmeP/P+VLrH3mCAkzaPpvHu9c/gXqU/cDu6wIcH2gZibdK1YTzjFlXD
YP99X+MpvjaibVIwRL4dvp1Lxpvve+6OOChBnrLFN7FN3ELwgh9wBjWM/Gg+IBo3c+EN4fdnuBoN
eXH1a4W0CkZE+OAwRr8o4lxDq4rUWyaIa3opuUKOnxPBR+/rjLPoAKdVlmRjI3YNMJh1LsLjkncL
KxAIa9NR8kTOUOzvtl6OaEYfzZjvXNGlpjZxDwXYVaNgwin8C6J3yjdjvF0KJBJBxciF2VQzsf4j
iheDkDaK4Ja6tt0w3Ny+xaowNUXz1b/6MIXc0uXO2DYECw96lU5Yb4OhMlizrlUcDjkrEGPXjuAQ
TswChZzJprPA45m2+9pu59RAzSghUn+tXsveq3NYanm4IPGmWA30MjDFnThaU2X0CwiaXvYWXDtk
AKIUAusd+BA5ksJdwY/QC7m09Y9OxJdCf2sefsiFi7KhM1o2IW7xLr8d0c5hrALzRBEjng/L+tER
F1jkgqo8TGUFQh/dAA+5LCDHpULVCMJo+mu39bW25eEhFa4fme6Mlu2u4BxGeAUeAoBDXwr2iZww
nSQ7VjqMR6Pljh6Sz/iqWtZ23tdmP9p05WjxNUSk1dBfAh52og5X6Hhsq/51Xtwb57OYgJ2XPXvH
Ca84SY0vm0bX+Ec6BeV4FPR0k+l2WljY56RGDw0lEnsq6Gqm71hICrTgyxLLAksh/Sqb3AuaE8aK
5AmW9DSs3FNElJ50h+y2Q+u0ZA5jJuIk9wO/0gG8HAgA3k9vTmoO8976UHLLyjRQaCP9yxQJEvFk
y+IrtbxEsfvQECyNeSm6aSLurVdEQ2RvZ+7D6v19LTq1+Gs6kv6uBgHStXpgYFl1aEJwXokvhbQi
U7lLf8NWvSTVi9Pulqf+1I1spPXMK7FbRGM0pXs2zgN7Qaec8PKo/XmDGARYZwHicY+X6fz0oABM
iZagocg8GckvEOE/m0x5JPz++AxlSNlmrxy39Kl9A/2St5OJ++YGzcLW9BNxmCE+VoNVSb+FPq/z
7reib5409oxgE3b6/e2TcUyl7AzGqSqOaI5FE5WcDtVZbcDComIkTr4rDuWdUJhYTm3I1OEZIawa
O+ZdDO8ETxO6HAk0dURtBkRRwN0ENAc0cuDcXUDw8a34qQVQkvvkV4F4Za+RIxzYR3uEzTqrOtx0
t7Bg5XIdKFlUkH2T7FfjVU6kPKpEYfMXXoENfDgmpUPpxioOphm80gOwXA96P+9CSlLmiJC0QnTz
Lyo6hWSyxznUGuPF+W4xCPLLPvZmv1z0Q0EaFed+kwryDG7tOmtCaimGkHW9G0zBvOuwqpbyTCFM
eS7dYkpcjQ8fJBcQPHUH1r6lRbkLCIFpB0zxGJDsfByhegB/e2JyT1MDpTEDIVmp6bawMyIwp+gG
ueMr0pdTAXS9RVzNFv9r2EQCPMahriSqRVFiYwsABO1xQMrrkSDX6JU8M/bfthRPjjnYJknCqqLk
FA6ghLfVBPNOpTkMyL19jtYFmGP2BMGJGrcZsIk48boZ+PDkxFBtS2ekBn0xqgMsRPrfd5TsTbPe
BMwKBKY0V73AEJ+4rN4I9UGNPCmQrhRoIg2RQfZ+0YU+O85ZsRvnjlzvSPSL5GubiYPoONBqE0ss
g4jlBXQ2V2xZzYPkoOAfRIiKo6NDcNw9aMiY1xSYVAkMSfZrRvPzDvMk5NF2lOnq4Se9FOwV7IrR
yXLgXeFtDArC20Uab4ngOuHMrZMfcNdcwXdhYesXynP4oz3NsN2cWa+GEqHVv3SB4CSffR/RhNoh
FdM3Ytq9Rb402WhivMLJgeOy5imS7Xbp62N50yrRM2Zk27MHwPO2Nna059GB8PbGhxfpw0vQLohx
0dJjfYoZ+yoR5yqiMuZjJhMnxr7QWs+nGIKux3La+xvedCNEmmL5aoAjUPtieDoxOaBg7DjXvie/
ZC8ItWTa0yX3JDPG67bzdu4I+Qga7rUYtI9po70fUJtVsMopkW3A9XJ6Wnnv/cf05Cus/l7E/vvb
ykjeb2vq0OVTvAqs5BoIrHzSKBnJC+YVp2eKXAT2w7OUgPhkEr1dNogKBuD7PLMLjbW4HGSSTwux
auGRzERIun97jwlK/ouRaIqNuzb5dYAoXWS4LqQmy/bUElPmiyCw0U7q37zO+d2IuZ7xMrNsuBVx
6m8dA7Sp4wz35mrs9/J9SBemgbONmEW0CMBFgpY89IJf1GBpeJrTrKhNw1kdNsrnk8qNGlMaw7+j
ME/i2lFyO6/85QYHGXpbJFtywvL3CkIAddPr1//JRofPHcCK9NMpKIs8PVMBmDdyHVj5vijampOh
6c8MAJPtou0e7Hvbb4YdDpEaksrdvJBbBJ/npoy/9E0ZS0IzOPK+3jnwVo6Hkozaly83h+qp6qmX
4JQ7Vv3YEOUhzytYn22l1sq0eAo8LSVrLeKnu3DwqmMFK22V1UouxCsgIAjKtsc0wIUeh7yH/dqJ
4NZPraSD6IPt7aM3ZRazJd2C3hypFUjEAGRRVSlQSnbpH78GrBcC8TlTskMM0Z1C8IsXS+7LH3uj
QKeNiyGA6X1seIKf18p1MiuLbiwGfy3X5kelq+lYr1GvGXnuV0kJvTVtnbv1koyhovQOqe36Hee5
Xf9MebbPlEsi/UvD/j8Asg6Er/+00GM4f9h0O5A51vBggh/94b7bg89sbTAQDFpOCtXR7w0FxVjq
cbAWhtAGtlAlMjws/F98FKTk6iOCPiU+YSbUSbMJWN6yxSW+7rdjC6RxrdFnDL870k1TRGAEaZOh
9DrnB91HFhxKLKbunOiaVDx04YpHyDa0vGK17bz0v/OFBdEXlP99Mq2o2RV9nxr2P1ywu/ZBBIwR
0sV9i8tP/UAkHxjNKxkRvLtPWCpFclrc9f/be8iG0WY7o2dnp0edWP1h3GJWyRHwpI+DBgCxHmTG
KRT65XATk/UYhA4h+j0Yy12PBpFkrYpuLXBAUx2lcFZ0d++ir+dNPc4Kn3VfMGHSIM1hKVxE+9TW
KHhdGTx9WJZb2pIfaAuDiw8goUDZtk0vdV7HC693ejRI6Zvbvn9+s8rPF8rTdXUulfSWgpqnWs7t
xhbOV8PUoFr26UiqlaNCUxtSe07P+ME9tuN8QRX5gfkFS/4bR0H70uf74L418TKgtnbjOmg55RKV
eRJAY6Gr8KMqq95ggTFgOTW2rtLcYtAgkk8WFMppjHmWbHjYYVfzRDPTPMqUVw3oaZNPnLkYggob
ANTf3RH1ORcQa6PGJArIxYhMTSE15sebRX58sEZes51laCjlrOl6JVHUa40fa+/teBlkosQFyue8
8eXsSgLc7NHJUS1UgQ/n4LIVJkrKl27DuBOOjhE9nmPCVA/6GVY1E/D8nAV5n5T0Fl4fHUPN/ktL
zy+LTjzyvwLgC7jPOKWEDpyZoMV1aVh0Nbz7PMX6hlL2lJxTT9v2gCZeETLE4gL+9dsqCcjld4le
KkmiG+KhFcZwB7eNVwlD6O/EwdmUHcId5ncCvE1wgo2pirpJBpLc70h6vDEpqDqCs80/AqFI+Xgq
5ULPd/z8MHz3XbLXXMwemwjhPD2BnsoqUjvaYerCdsGwCjNqQTCMBeW3fUhaGlK8Ea06wD8zSNo3
PUKaBDMF4pmEC0F6d4U6RDuyZt+aSKjhx8Ew/lhB2ZGEMUDJcABUU/+BzPUp2il+lfN0oGbFTCtK
DjdT/kZVt+OFY7lpQDCAdJpycSyTeSCTcbfqsHMef51JGe2nL60glvftfm3EiftigQUiUfX/7FfN
Ov23/nfCchjZRTS4SaooGGNTukS6pBeYnURE8C5yUVyo6QqrkBbkfO1F3vrb4SucHsmaRziH2ToF
QbZZjp6BEaQTRG7G5bUw+dPvw5zhfeAdsx7yKRIqh6JJrAa5ea2YDrgB9Wm1OhmbpBIoW4iYmZTG
7KDjx/LERXA2d973HSmVQiugosLwKTH5ycxQLqift/DtXoihdLOcNzLx+j/7arx117iGS6Tzx/Uz
/vixWYktYYxNkNmkGkVf330sYA2jGjcCOfR8xzANldqWCnm/6fp1Dxy4/JO20A07Z/DwT+ooIjy2
0p2oA0+R5hLIipjsQ1lt1wM4oDBLFJxzDsmcEWLdyw2fpoXu4PqXS+n7kGMFujgbDZpzS09hLx9y
yLYU9Cfo7wlZrFDAtq6+k+E9snl5jd2IEDALMuVkEmlrZWWxe65XKJ3v8nhKusUsVeMUoznaBBMz
oXfKSxqi77FZeD3wrpQARUIhthkcjorsy2QZIdE2ZnkE+NhF1nivOLCpuXLDaG6rmggwkxmtwlYv
giatQg41YudIHyJV+cP85NQAtnmg786Oozbs3KC+VhDuDO+Sxcj/tF1zpRSuoNM7X7PcwW0Uy+UY
qAhFf6DJuh5CNQNgfup2mWEijbyGF+Ff3kLhzgrKBeEZ8D6W3LMhSFhnsCXLzY55SgYYr9L4Bsmp
5IP15MNxYxFao74D44R49LB5skvvAKDnSER2iyReC7mhF/4MHU05CNT5sAEBPy6DTrjapMkChDhO
1WYgwDy1hKrejh3O5YzGpJ/3QCxE9XnFfQaui7c/lv1eIeWlRKUwWWHouMwC/s5BH/Z5CfPvMsX/
QknGTIIK459KE3wJfL9PNrPki2ugCeKeb/t/byny8dQ20zr3+UYwaLTiVN4ot3amY6O6CVq2slUC
0jIHu25yptIv1POnyrmwrTujXM8lvH86R9iStm+l7bKWwzt5wVOdz4//L9MsdyTbwrU5onCmaM5z
mIW4anAF+wRcQ/Cl8aU05uswDQ4Pn9WaBtB7RH6YoktRbb0+GgEML5o5yuVrZOvGZM03TOmBn4lH
DOKoaS8Po0zfqJVCXCJ16KmXN15WFYsaExSvzPdwByI9OQ/KQis0SuT6kC4y1KGrq3gq/3JNqTqS
C2dX6xIWL0CDr1umXVyFEkppgX416ZkXB/s0CsFp4wwj+Z1SL+vPDv9SeC4EDaRAjKB3iP5dwAwd
jPWaTDlO7v36i6qH+0aVWVlo/0XZioeF39tF2dGAoYfIkNCwzCRDvlza287Umc84ZDeyv6kc8pi4
jGx975P//kiDUUm8G3bWawK2BQ4U/HDnFd/mHsp14++/Ms8i1HEWPIwueSdnzZRz7Xqm7h54wTAO
K+LvHUJ+c6two6zScBnA9UivDEtbWrv3y7UmLXxBKS9/l6aR7EyYBjEjmoAkfzVv3jEt2f4seeOG
zyLBedaS+SmUn6S/fe4SEJDNS3h3lO5G/A3X2RfJTfNoGK6SMWMVJtdalo0iA/u9Yzu0f4xcW4tW
PLEjGsT6/GtfQdaZjMfOGRsqb5D2Lc+BWQHdnMYFkP+VyzjvQhExtfDH0RrlEccaRkoQSxt7q+mf
6SOE1QjjZpWqN2grvL9cogu3iE207JkHUJlGWbA9VES7vplT9/6Zl0zmHNRUxC94azjf3siyTNjG
yy8bFE1blJXkMCHvx7ajO24z0D0L4iaoOksfNiHsRECRnKPZf08GJCGbAU5mEoglnW6cloLjXKxT
IELIciZTyFVKOBp3gaw25TzecZCPgeS64ejuaYXo74pAheXVgvT3TIaRKn4iXEQ/vp3gjjjU16DQ
NV4ykqgmqnhBKmzq+Jh7F9nnYw6cM7IUAiBUFWpIL3tRR+cijdkuAGht7BvpRvTUNF1oKt9+J0q6
PeR40OF5NpqYwNvCY7pRY/HoGBAFxeEu+6KvJnx+IXZQNvNg2WokRzakZxr05Z+LUSg5+dy+z19C
MYaFyC9XN3xyGZaKUVQOAiCdSkU+fChLYKcc2YA29QvDeShwIyYaLM1rBPFT2AL7lCLGhlStWfvo
GmNuzR3Mw07XaLLxb4oIROQ94SEyUInCymV7xajDb7mJGtcyR2aWi+FeAT7o3YuCqqn9DyVtEvai
b2iJKSp4rJBdCTPD6k1GxsCgQW8XsRuRnmdPFupKWAE9EmmljRwcfuSClPjsJCI5Ch09MqBeC4DZ
xzmmEf+mBN+mJ986xoOpvmH2YDh1xyUQOvRsINWCCUVzFw9P3r0fkiZdGg96uxTf2lRlpNsXXJHZ
yy1EmT/DZSqDxBB+Kv9Kdg1DHmAb9sdGrrzOIesonsBGj8GSb6+VVnll5auewOsFVDhm4mZ6c+UN
IrzgQhLJE8IWaI1keHcmBgeABGoxwnheYsAeVbQxGvp/GDq0IXmkytHMW/7RSYFm0byhBY7yBMey
yR0gRNMOtCA5ddAq+5W/Zb6Z74VlaWaKJkSRnnEwvExI6aiTAT3lmrnssewgM7gLO5WNseSBRlqU
NQF3RbyUKkZMFqrQYf9b+viEx4FKehdkeUIp2JJwlD+7ruuk908UbzlRmpVQ50u9EI5BIMrZFlsi
pGEM4X6cnbMdBv2JeXQC4TdRx/B0JZoLdG8RwS7rCVA5p9GQG2HnjDuA3+S5qAxD57Sg5qK2rfJh
L79ywp/e14SFBtTpvqtoPmVfRn9sWBKAZeWQQG4HdKmzj/PdDqjdC+NqQo1t8DibyXZuK88xFveu
Flhsf5FVCVPZzKUZCbOpqYHQ69BksCRbaJILIar7QWzDIk0IGXd7k/k0UIcsmoQSpEBRudWPtdbH
AGUMdR4XdHO8hGKxLSGbDOu8QRs1vxIrHBzG8fltTEaqLiwvu8P23vcEc2kiqMFCbZBgfkXL8C1E
MbKZ5Dzb+RtqE4YB7FzS+5OZCFA7rStRG5se/h0DgHqUS++FiOreMWGGrfJh8VphRkiZ/ZLamVkn
z32ZOqo7UPZHad3KndigUPG1ppy6OB5libGsVFagbGhhrmlC+lsUT0Z2YMOPOQMWqBBp/aDaXI1n
XVPNMzcunxoSjJQm1HWLD9ip26VJaUTudsHuImvJYDVzzqdFT02TMlVBIqeXgbkqLzQDFD6VJ68x
9E0dqHhH35G8SdHWJWnt97gEd2OaqPRjRIiabG2EbbdbYftNu2vjZjP+OwUW9QOAo3xVW3WVv0/l
60UCJW+NQRO/6poiAb/xEso9Eu7ccVafiZx/UJrZQKiq3vtpToEQsR5U9Gl4Vav1l8ItiEtZOlyE
CwuLM5Qp7jFakSKmr+7wlc8bU9TwXUhNlywA2c/+lwSrfp86jp2CPnQ024HAJbFbg91hbr5zNxEM
Dz1JzGmH/X8e4UqhIaDhweWGsV+e2EzdoEyQ0LoZqbrYBOCKM0Z2MeySceHatbbXkTh6hUq5ciMj
xcRwMMm6v5wBw+0Vm3e+uyO2pyLJLS1tXfN/MQAOh40YxIvwLWTuYLuy2zS4vqG5GyqZGW9/QySd
Z8VSz8KjbQrU3INfK02sjb6QSWmOHh5FSy8YOn3MBsS3bvt0KXaGWcz4GIja99FwItGt1f3szDMC
9WAEAtg57szg3NGxEXSCeZHjAdHaByJRwhuXUQspEJ99KeE9UNF6f3hVfkNIb9JQpuogPs29oiOw
vUBArmpkh46tX6c2v/wDfSesxM94z3o1vHzV/jFTuf05oTYK6EsmnVTzmzeCiIDXX14p1w6sLUCY
uYR7lQ2mMtfVHX2w5P/y0xAIUkItRYvltbGza64ArtPeab/Cu3ZsM/2jTVMM9dFFKDCtpvvp4aYl
j0lyjyRXzV8BGf484aGmeGh9xLjbCmwV28I5havw8qh2tKJidYvJEO9ZJC4zlyxRz7vffgDW4vSf
0Boau3CVZwIENbIoj3govfMV9Tp19idK6CJmq+S5OromlEjuxho3EaAtSGsTl6Lo02LzIJ9QV10m
oo0Qpw2fCBa3StrNz56AN6xyS/Hlmcgz0fvixb+h+IYGuvWPUFlRJjPNmvYpu57OocQMyHopN+dv
v0kyiu6uteyS1mu5TwcUXH/zJZh7QTqxniazvc5Y524UiX1azvkKbCquk9SrFKGucwLlPLS/0PF1
wpJ6FGqaBwg9YOU+onQMLb44dKNRoRqkKLPjZRw85TrceRqSSiJ+StvDem+I30lf+YSJnVs09pNm
JSjw3UD9X32UIMHgVzptiFGCZGwFhA+Wr6+JqgjHFze36bDyz978BYTk10VMX5gDv96ngIrtKxRN
2mSBt3Kh2NcHzsdNgxZJKi8SWa+17Oa6dXuVazGQWajKK+rp4mvLdQtu96GWS9D14imxA2S4Ngvl
OtwaLnjKSxl2dxlC0R6Df23/qtGyWm5B/sC75EP0+GYpkbVmlffU81XZw7t/jviFgRydv1bs4hOM
8/6mrrZ/f+PDvpZUMeIWAjxxfWHoLsFtRmJHJ2J3KHF3rZex4Z0j7D2syr8PdmJVA1ZjWkrjnbM2
6mhJLoyqcd4J6yiT3FhLlbFqMKfaV4vNLHM8pX/WqsFy/QRJJcod7JXceBa89oV9mC/M3Uo8t7VI
FyZ2GPU7mcSe8W225QqKVPf5Fq0Knz4VEXIPvgsAAimi/ErK/ydHDW2lIjES09oQ5nPHN/4DWOLy
HYyVC7Cl4WNtMYla1WTLYXuwoEJJ3jxDKdQF/VMIndVfcTM6K60Ep9CkTK3i6QXTdaOeCRLESei+
rwOqTJowslN+LL/ASypObEPVmDbpE9m8e6vmVeSFVrIffGmiO7ESST4QgSDneE/O2+bkKQ+kKa0S
OjB3OPabUB0IIupqnyhLE/ynzU++10vUYx8uDR3/d6ftsg+OBI9mlLDi4KctuPTdxu2kRVi+9BS9
FkTjRZ38G3T+IJEkuOsiGRr8tJ/npyjymaefVwrLBVnqF1Tf+GVbO3IlHvCUci+B14/HQTc+Kcsk
+2L+nSp9NZj8VMKihLHpN9/SkxNsOGgNCkTSDjMCPzZVYcmwYDJyYRbsqadLcokJnzLbFhSX4qfz
NMIh6gxPLzmNwYr6eOex0HcFiY7shYRgZbFvbe+QuGlKdhlxtymlKwr6hPIxrJruOn2gJU+7sQBR
PnmxajL9fMS/Nv42qS+HrSiYiEGZx8FfUAN/jqEKYGu+OM9vBvV6kygB3s0eKVSbw9CehlIPYIUN
O3G2Su2bzXrKVCO5PdHGoVAddNK6PGTET1KddCH99MJG/KaL4oITYeN3gBtLb8ET0e6QgGVBJQBj
7u2THRdv/0yHoaDLqnj5zltsboBY9V+rCNu9CW07o+EkyA2BxckFV3sEx59qEWhDAtSfQlqaUEbo
v0eJEyta/Qle7nM4BJnf5HUHlykE79G3olrrSoLtM7NQBZHdlA+TWNXOTX44wWtugL02X2gdrXc4
sDtnNjaW4DlcwfKNo8IrUyPo2Tv1V9FiLXhFdhuNxLxkOzppLO7stHexZ95e8soJz6gFNCMwsyVp
pdK3M8SMyf2mBAoHotC1bIokskhmcZ97DKN0ol7vpzQhraS7S3Md79/KraiIHo7/Y392bYrK6/nm
YMiopDsyrDM4CAL+JIaU+RpMl/rD9g0E3JnY+2i2ptiZUpvfYJgoL7jvt28SWyUTY8E1M27wGDlg
W4msaay+n5IygSR5cJCz+n/xxk+3Uhsxmc6V9Kz9C1IXmZ5oWL51XApdTYEVraQw2tKXwVCU3HnM
RH/Wd2+3G/vhLCazt1oCJ/citjUMeZKyD+2g4t49tTOWq1bCeg2spZFrwTZ7mVSuWhpF0ffuXuL9
sIaR8Z5f+taGFium4XrH+XV1Q/43Vet+yd5sMM7QvyGSFt/moI8KIv6ugrkdh0fIvQjg9m5VHnWS
voTGMua6rYHe5fbBA/cEfw2/fAp8fTEoT5mVJb02O1fa/4FNiW3HkY1q8BFdg++b9x5ghxeBjFda
XTVL4LYcHKGXNDjEMj4PO12ebk+fYXXY9X7DYWGugrZDeoLHiE9djzVDRseBwy/Q9rNZ0XXXChG0
Cs1Vuo5/6Bt0eqqaqjwRFHl4NlFS4R/9rIUvDyZxYGWE+Ov1sLRop9JZYGnxdvOK+sE+uOha1uVc
TF5wJ7hITSjglkU94EzStwwAtWQGPiZUuunArPk2bIgBHCevo+pJvHlUxfGa2E59kZJNiY9pKM9E
4FTX67AISzRAe36ibWWvhi3r6qci/5oNEv5+olM/kgIBbZ0S/r77vdi7gu0Uh1Y0u5b8YR2F3MrO
XsJ0ax++t2FRKDKRsM0blBwFtiF3IsbvbxE/XyMNMBbNrPgB9S9zdYl+yahN0MiwBZ2px3+vazjA
KR+lvRBIi0+FLOqiTCxCw7UYmbVYKKFfqxOzwhnptqJYRvdSVdvg2CAtiFP8Ipf/+ZAn9Cur67Dp
elBPB6Nknv7F62ICehN0+zALk0pV5JC7SlLkRHJih7yXpXsN+fsLW2Lxxp7fVJiCwBnoMeqN+fBw
QEOn4G/LSOMnEYFJMpIsyxYZrom2TojwkeUklbj1YICqNfqvbZaDkeL3lWvFibYbpu1oCHxnRWKx
0IwqPjOa17FYVqBMB4qYBkxJaMx/YQOhOSeYYOsJ+MBuDJMdVnCZRg5m0obFw5a6jKvxpCD7eopG
c5981x1sHmIqb8enFVEUrSJjt1CoBCwLQFaNPTaN1TB3WHiwtcV1CUfeDAmwZ3Zgt/iReOwkYt8N
25B2yQOSqGjbFbAOP4VNqYXuLA3/3XUSHZ3ky/HPIsyF//orpomXc/LJhmknOt1OQEOCRvlFljT0
5Bqnbhdz7c+K6rAE7U+vXmB32r2F0CVRK9WCl8z+bv5J2PbgdTeI7c7J01ka6YMmhR69mJRFOTeD
8pYTY9sS7t6NfPb859VnqroiJ7/cz0PbUzq4NRpYC9VOtmBO+Wt/NZ08DxKyUR3pGW9VsovI7r0k
eeovocjDLfTgbEBwcycxDnoUvVTlOKVIo4qkD41kkQPaa1qWnjDU5nfqzkR2FtNKRLPmlU+0Jtva
7bPFdvUQarkQSr2Z4Zv0gXtfPCodt1KBFt83l/sLbOQUX3Eg5e0tKDZ0bBcueKpmgXqXENePl+J/
aLFsYDtKxvmxDy1GCIA5X1uFNopKkgfc+oXXfqeNlWvjRFh17SOlIt0YTmMRGiT4o7fcL4K+4geb
sO8h3iqpaU+L7yJf+lWkYlzaihuFYmAnPO2al6KRpub4KSSxvrCRz7WcL966W8b1abEh77Cz1tq/
AD1oLXKTqy6UnQUyAWuWJCPfBaJ6gXc/mmocqW6SSJYHM4lIOwGz873dZI3xfVJltbnPy2ta1fci
dBIUaUGFDEIEqmFPDWNmwxX2NvR10OlO4EC9K9JIosW0l/hQEgn+JHMoDh4TqlIz2MJg3YwHEtOE
6gfDs9O/EQ7yjPJW2B+831G8xI1h7oS0hoTiajHj3/5omihm4TIhFwxzrHMSlf1ldh3S23MMHFAg
eIzH7hsNLUX6zTTNeiz2NcIG8HaeLHGDMt6UlD5/qyKkpSL5ebZ7BmTp/TolxRDee61898CKq7OV
ahlZpNHzmjH0K145FrjwGZSHLlGM2rvDXQ9Z1qIobrHQDjIa/quKdZ0LKo8xNcufOYUeknnqKN6O
nfoduNI9EDZnPPPi6Ixa46KtT/mDB8xpq1CgaRnE52z2rMICbG3VUw5+x8YyI6EethXq93/qKn1m
xaofzW3EYjzdBlve6p9ZVZ4K1noZ01fDbd37OgTvUQLW70AkIIGLBbD+npr693kODhLTJ5LWJSWJ
yWFC1s3WhutSQjgS3nYYtjbfkRT7laolkyBFdT9/x7YNm2dPv9zXfnQnObfT7WajKnFQNkJefB7V
4ut4KiAEY126Lq7ISuamhcp8YETsMpK3+9rbyYBwL2uFZELx7esh+MO8O7OO33RHujdtw47825xb
HQBmVXqy1pISfMjf5OQApChEIkQMw96Yh3DyvzW8AV4J8KBrZ6AjbLxeq+PmXA076VoYHwHHCqPS
VC47SLAI0KOwH6Odn3SDsM+q8QPXjYNDUBq8fnjNQLnskv2tcm+VfbEJwVrwWQ3YAlfMncHwHTAz
AZK67hIN2Jqp5IAcJybrehbDhNz0mnEURYVmPPL7ELjXLD7Si8LFija4j4/SgarJ+G1JchlCYb+F
tagczMMhtOY7d3IeFwTQLlbgbOKBuRLEmjmk1Ck3vTmbuqwIQiRvVPN2tUH84psdOYR9HI8AjTPw
I6iOAIp5V2NvwVlX2eFKCSFVv9LGZzvwP4wOlv0AftMjJVRL01CEgq7teKISW5jxjiGxEKfcFPsB
yo72MOqjj5wSdYYZb2M7IaEbVylX7qpoCfCgkS67maFYl5LcnYvmnt0Ajv3DRmOr8GMXfvxPtWpD
f70fvUkNWC8H9xe6dMLBVDKnuhEO/vUBaiRM/Wil7CoKFotN/U4x1VX0u6h67hkPbrPYhYBpN4QN
zNAFKKHGHJMSQZcG8xP9Vu0PID4O0BYHpFER50sYfHnUiY2VHKysIhJexe3qbEymj8BZylC2dtco
guNFncx6f5q1v6Fo9rTPUoMqmomA68HLVlOscc0oE4qXW7JyVMopYRUoQBIt1AAWwjOnFOs5BMnz
byLDVs3876LBGeVe7Ztdbl1wEdZ0Uf9FCmLhLe08i75ge79v5PsG3l62aQtcWVQ96aloSltPPnbt
VMgTMri2mDaVBmtTZvaAtED8xO9jpmXk7WU2k/cEFOinJxhmH0AkLlmWR5gqaPI1J1U7JfM6r5QF
SVUrl7Io84/u0OQRtILWyo56pAK6Ehj6JAWcWCqRqOBri0LE+U9YNCbjJ61QTnTkhEZuWVUiLXFv
VTkrSw9vm91CWSpA8/uI5QUanv9lKKSzYICuRCNi3zhVpWAT+oiC/qQKNV7A3QYew8GInWdxRVe6
zPEq/Mmo/XWN4aDWhMHNEn/c+3ZcVXB/1UvabIzVP8R4sG+PGv8zMrpJ0G/6Jgk94woHHsCx2rjJ
eql4oocZPEVz22FDqAcETXyAhYTUxnm4h8DxbIihYrbuj9lU4+0Ta9Dvg2RpIznJT+qNHdCQMmCp
CQFvfoTkzhGDLAtgvi1jtKgIufg6XU9VRZVTshm9PZTqwkN3LpWOsOmWNEgB3BHnpSfbXc+xyJG4
ArEk9O3ITVIsFdYvnvfAY4jAD5CnC/ZwcLDhPtfBANuWe4Rqa1RpkZunzjukahsAiNsd1uQO5JCZ
c6GbaKUBQNikQeOcgTslb9v9X8s7It356CzkbQ9pVuivjYjpx0T9kdL7AsE2mOvEV21OCROTo1wz
lnZQ/Nrg68288dfi1APPGJcdDKQM+yWB0EkVclmWQOaHt8ZZyAr8S80M0mqD4SlPjRqi3mkd0gN/
/J3FlCbOuLMc6kFC6+DhEQj6NN2HShH94W3AZ5xqxWhvLJr76fIafya2O0o/lJlFEUwKcePO2/Bk
qsHSRQoSXQRfp4fRdBQXquVevWO+vc+Ewhw+hnP0PDwyK7swXNGOcLwO9G58MaMSk2BXUW39GOvU
xUrN2hkLjwebK2XsiSI7N/pBvV3SXaSp0UMlPnq89+VRS2NJXOPE0iai87rv+E5pJk3H3L1LLRcp
GtHB38RCF3YG61sTCGd9T3+P98WNYl60wns5GSEzNQI2he5mDtuyW7B+YIa9aF/4nc2dA4HU0aby
JxtaGhAZ7GBUoSv3n8jN82wjElqmPVRehZMea2TvWgfY4PE9mJBrISCTx3xf43rYaau5tvHI3qXG
T5BuhXeVGHv4HKE0boaQEILLC1Snun2Qa/fbO3jG70RyC+jj0QEVQ6iUQC9SPf9lvZZ135jyUfUW
vYFiSNcWjFlX9T/VfiN2tIbT0P5azhmgFOOwHEVxYU62Y1HrAhk4y6VDT4mYoIfE9jLyDnXZ2LSz
L+V/B0Jrx/wxHzs7h0MV7FZBf/jY0j8ZFLMYyAR8hcAZngdKAU5GOBRNORiU4PeYKLeX9xvxg+rC
3KNXzkzmz8JKZw1PF304sfubQhP+pItkbmhV+iQeozzgJPJ4aWgO+doWp8jRCiSn0FU3XPy4dh/m
orftVzEbPyyyo+Bdi9a58dKNjQ/ROClTn+Nhb1UwIHjAmNmdt/0FFcqEXb1Pq1PqNE/aMyxoGcWe
Qxz1mW8CThubhVhFbueIOB0KQ5iqk6VEqNcPfMV+mN/wWX/gtWygLOIhS1m0yVRKoSBc6vqXk22M
W0EoPYoV2Eqe+ltkcXAIPgZliCxCyFN9wsA5gWPSViu9UP3orQKwaRBNWO63GeJ2zFfX+fiuVK/a
aKw13Z3k4aoFLtWtXb2l2SdgfLwKqoPqZoLNut2yPn+nHJPWXn4tSDJfN7am/uF5S35ylOhFUzV1
/volyGoGilVGq6IjCWQM4eqm0LZIdV5w2JxMfCCd+w4+v0Fj9oE4/AvSeetMNZKtDmzX4b5aKK2l
PSh3003Zmm0Bq+rXqzjkIg1JHZCFfVNBjtMWvkkuudYgtlMrPB0+8XzCTFBoFhRnOiKOCYI/BEex
3rfBSD56l/dUcitx4afjHVlmqeqrbY8BsnpV8jMoSEBFhX6R68au4kgU3Pigvx4pWtkS9BcLF2Ix
bGzPFsgkOn3GqKjwXQv0CiXwVKGRbK+wg45Bqlqicvd+ek9o2HXMV6Wt9C7kaq3UFZwI0kNqnUZn
T3w0RRH1D8Qawkzmp5HVfBuS+GK9i73oiGLNrUrxzBSRstQwqnn02uMb4CyRdblDRHYnMcAHMTI1
UeZvrD33sSABPxmJYyrDn3ZqyVCD2QYZlrCkRsPeCU1PWNSiOsydUB3UYHqa6qqYO4ItGTs78ipA
G8dy91slcrl8a6L9hlPeHORUGdw8qUCAi7FJXA7CfPIIFwKhYr6h2HnIaOWGL7Nq+T06GJ24rvBM
b8pLZGvdrKEB7L+eM+91sjcyKu2GwohPFbQM+cwcap0+NfT2NKyVAm9Lq6suXpaG8hZ6vFyt6Ql6
/bHX0dFUIgIjWVd9wR2MZbae8ppT9n2Wy3CU/QC14BbbdC1DfmDbWSlm+F5softoKm/0b2CW1yDw
TiGHsA67ZOc4UuJ5JnBGOKdvHIAGdoTV5DGMbL2dzM/SghFh2SdrB67gtEh42PDtJBIyuLpreC0s
Vz3dRDIqdD//n7BOuSh7Dw8tZd7SuBzkHg3bd85mWxrMRPlOsEsXJeu03fpGN2Qy/Gd3VLFKdCjI
XlPuU1veId486im1Rp0M3Mc5KFLbpLrLAaRewKBDiP/EiaQsI/ZxZ3fm33VH3qqQwoQTqwyhd0oo
8C2tPCa0dEdrIshy/vACjfRTnQI/70jyXCQ7Vofl2GXmlCZ4xUbPSaEX/7/LXIdGHd1VydcPrYXT
+ukHV97mk2z3f4nuny9mC57EjfUZWw1MWvyJB5mVp7cC7MDu9/FlBXDbbPFDJi+Dp/mR4LJDscm/
tlO//5y8t7lU/EVudrz8/xmmc+jTBPvSEMB0WlXUVd14q0Tig+9VMvvofZmNLiPOwvZ8QESUFtvh
1NjBJvTqp1vK+OLX+2PDIJhe1eO9uRKb9cwIFfnXSFChWja8/ZgcK7GiRJmB6vb5OqtIMGibV4GA
m1L2bDfnDD4t74jzZ3W5U6Wy+PNZmF0DOGxrQvXyd6OBwC+6c5NvEo6+rtNC/h4E1HuKKIJNP8/e
L+BEdXI3VmWnxo5a51SZuR7oIY0fBBTCT9FPCWLP27+OequyhEdhv7uHsiUQDTJHB4bWsvfW5tSV
d2tBqRfd8Dea3FlQFZu0j+o7XGj6TSvoha0Vp3TJseVQRJ6WcCxU7VU+rlybnCtPt3jGScLHzfRX
Adh1hzwkRG2Ybg4IntdZ6khMIZW+aLHj8gVYwTxmTPgEPD+HhuEtsmJdfNzy6vACsgFcIRj5K1QQ
vE9PJ2HdMG7eGEy3i/e+gtQREfbr7ozn4a4eEv/gGMIge9bps4NbIk7XOqZgSJk0aQszo43+1nXu
rmVhIpwV0toGs+UaS3z0KMgHYaUhhayZOMzRuv8tfl8PdZEhDE+rJAE4zzdV8B0Y1SfGGDl+UlAi
/0OtD7RMqEKUKi+8F7FJis3r5XPYs1PIDokDlGV9Pux0+gciGdcJMNtusrWmcpBgY+BAhb1Hobzs
kU500wsTKBHybzOKjP9tsl5VwqLEWLeham+9oYQyzfyCC4KqC5KEcD13dhN7tG0mtH5uOA2bCNlq
+5I9Lqm71qgCf3TaSyqUuNriF9Eg+dyGFHYTAGLGzTntvhUbRJpm1bXpInfiwJ9FtvZo2QY0OMHo
0nDRzlgkAUWD4TcVcrIcSNJguTUsjl/Mhf0Ancp+q2i9zA+EFp2cwjrGFbdfQyzxrXMA9Zur9nBi
ABYJSR3cLXDh9dDrnIfXuvyqvNwxAeHqEEFWxUiehz918xwN7cPLB2FnATiW+oPLwFCPddonXqRv
POPAbHD1p5GRjPjgxSzCvb7UNkeLMZpWY6EDAXXMI+SG3qdRm5bR7Km/qt7g9hqn8TMNXXkhOvIi
BvSt6U/eD8N9hFWHXgkSoozlOL4cC/eimiDpoqBx8I4UoO6ye/wl4PYQl/SZSQd7gZWJmDmyXMjV
nVlJRnk6IEIpjEGuR0bXG0+ADq2JafBxcORBGCF3S7kvLD1XMNFSu8eK+P8SPmqkdBIkfeV5IiLY
NpCpi6wYMlpZC2CHSzFTh1f8YSinuvsHLpWJcRGhkMDLzWC9tpe8lNXs3zLFQ9T1PKbwPNe/jAQT
WN9wy75oX50PBWOc3KYja7b7PrG6GHYS1UNUFuNQf/JReudcfHhPvspkFqgBZtTW9LeyeBVjdZOa
xg8gUoQc903MVpRumTi99mtfcIZvCyItIJ5eVOT0FdjBhGT36Gr7Cd0VRXVVmgqrVeGOj19N9+0H
F5C3BdFRT902nTaqw2Eg0c3PRruKjiYNccK699U77iycTCqQFbcmTqVaKkZjip6P/3iBB+iYH81c
Kq9EuuAT2O8zjz0xZ4hcyfVfkTg34JSEDgBSb9X8nZM/nWAaDcofzcbTw1pB/IfkXAHAs0D5OKzf
oy8oI/DeRsojCf3tfBnbqivVzwxReoGgHL+KsoCME8ECKXu5EMPJIBoOn64YLGIKvsUuvvHZOS74
9pyC5fBEgt/ItWDVbb9yrFBP6ukS7Yem5Cm6fXsQrE7JEEQPXwPSXQDLDh9tnjgmbjcqEcfFh8Yu
0t2Hn4XGAtg/gI4csyn9nJgqVgpzdC2gBXSho86loIjzFRbcR1KIUqKftLxJoE7OpVggG5J3Dasb
DzAWItJpjf2kYLYqiMtq+mvfl93yfzJWtc1YOUcan7lQaJLdN1DOkmInjT0P/GkS47jqFjY10wSn
saApuW9hMJTBbGdAOvycidH9rL7SlbDqJTkD16Wx7zCfBmgPIYESfTNtufTR8+YZGhfZANZtZL7U
Wv5eH98Q/C1BuqqNT+cPtZ05YSp9ts9e8MOmfuK2v8nUTUqqHHqCZT0+pw0GKLwg5CjPbAO3cMjo
r+QcNyWNqDZ1/9XRb5gF4K2PCcjDSrGdTvTLs0K9Eccj+7dRsS8hNJLunoV1iwngCX5X+rWyBMun
zeXrocVk5d4ZBoSSZokEDrS8ngYmb62aL9qAasJZSl42zGWpH420fAkHCntTa0qZH7TBGO5dO3Py
YnBBlfxYyFM8q7D1XpsRN73ekJja/iaLU2hYds6LzT6OpNABdXbkcWenUM8uqFk+kULb+TrroDmx
jurT5IL0UzlgV9smmnUsq+ZLYFVGXgDft6cbCpkOU1Gx2cvgd43NEWNry8HDA8hT1zpRjl/VU2dk
b0EPNxMWiNJLLJC3Wlu/BeTiKUDJfgTjFyiN6TGlD31ZJueHqynGMaEsi7moOG+xYXUY4/hTX+NL
pyYFBDNstc5We0IivWBcdYFfK9RUXjllNFHcroocAlhSh+FR25YsfdM9L9hMh+sJgkhJBUGXlUg3
z7pKVm3YokydxjBzTuq0TbfMfbBn84nNeSGFB3HochpdawC0+chNFt9lUt9Tc54eazOH0+JF8EIX
13WtafDaWbwj2DbwwLXTezlWxQOU4yAgGOiWYStWlQ2engrrpn6OP4vnnf12RetykCnwB5wmokJM
NdMvxq3wqX4tWJyTO9C5nMq9b5XAD9wYvidHYgUMBnUX4pnPoPZJMsQMMTdckSSjmkOLMTmTwRGt
hhctXgf+eF2PGAU6zykeyLDAXo9TroLanhDikYIoC09lqDSZSUROyvRY2GyCaZZkfQyWNgRLshi7
dC3hRCAwJD091FozH9UsaS05h+I4kbzWUB7p6Yc/e45VqorGcSr27nfaBBEkTzDMBSs0ErOM1B6B
zTyfYe661kupeMlYO0GHoKq+TCMUoFqDDKHm2Moocw045D6aVqr0T6z+igk9Ex4WcJwy1mrVgrtw
tLWdcSXllYS9u3ylfTB7r0jaX5obCc0uCPEyYZJakWOHo7+a0HEvoiLE1p1VehxwfsqLeXpTyNX7
5wLPL2yT3Ab5gcMZU5OY9fK6vdEOAg2726aZkuno7WkSK9ObVsv9RfUA3uNhNCJs5YBDGFe2I1Oj
w8h5iHmgMaTufXPAjr/cpD1EJR9pW4SaBDyHs2GSQ8rrMur56oninCqnq03bLg4A4tPUjr5ova1f
a6oqbcvQd6jvOJDkxgg5e9fP1jLl2licGqWoVn8vfFJM9dYSRlEQym4Hhp0YyAoT+hVRIVNNuaHd
cgh2JQtmjJzfKDjlf9lxJYxlf/cG9HqPpXRb6hRZIjL0/EUwSA/nOgLxxGgnKuvJwr0Pg6sgWAjd
6HfrZLev6241UF5pfDPQYK/URxoc0yTTFI6skWbRW0R8uJyOGVozWSzc5AA9BAgRi9ycIvgVaOB9
Uy9OILHkD+lXAV69i2vBZpwVMR5L/157NwuEJB3ZGHC/nqhikzCgnqaDBOMedZUtZ2+3z4TINJJy
fbKnchmrcAsiBV0VVWp6fC01tGKRtAeumBA4ReeDQ9LpvYyi23F+ishsdfXq71oY9ZD8PwkNwifQ
VB1abuUhtVnn/P6U8d3X+fJqgCqvJtdSWKxfKxL5LjKu/e3DA0P7cBVDagEPo++pflvXqopgiZXB
K3EMZ9+U7ec0EVVPqjyf3W3M3Lul0GBv9jLRZAjSmv38c6QRUZj0Mm3VzIBqLpASrc0dShWHjyYx
xyZlzzfF+sRpQxSuxc2l/UcNuB08eskopQSZ0dgrR1LKm8v0mObexu0iEX+8we2RT87HpXDXFDf3
WjvqUbDKSWe0rAdsId4iK9S+wnAWRfI27gpGSZZ1qRGGJNBs/ty0F8knxM8oe6mEDDPLTUFhPS1R
4hp4mfkWAMAJK/woWwPm/iaRgareXy5uE0uE0z9Issm5F3W4WIBbStRKvX8OfNbyxk3VjZ3lSxxE
GkWZpFRd2F35YTk4X1fzMglw2wHcoSUCSdVjOk1xIIwgG78WYhTWczwqF3EV5mu8a//IJYD6wHBJ
/z4hUCbBpsVkKBkKPfq+PyC3ocyovYY2p2QH/NX/9RTGyyAiBngw560kcgEx04eZWfR4w+ZYgh0Z
sQOTPFBesvkkPuAYnldsoYIsWlIDru1uCMyY8Gt472U8X1h0OCVBE3K1wTczuYxflAGoPCv+mQCn
5SzjNn+d4O7Kg4QO7qGVn7RuxLmkHxPR6AtXaCP5QvY+gsL4dqqbLUY2pj7Hk73WLFl+dBfjoS99
FeNgMbd78MDCVXi9AxkPgM4eKI9MkekG2YGaQHg+tmsVJ9G/2cfbF1oDPhgsoLHV1amYBZjhUTXj
Kp5QyghheaEb+GRr5hbTQQOccaaFLo+u+tQeTH7Az5eeDZ1JSlqQ8h+LMU7MuzSGKwpxf2TjssCj
57nilPHZCDtgAp0KJHB0rJkUPiUilO5al0W8LpjBLVjfbJnguqPIzTeb4MQ/Eqofg8009jVScdyG
sH70vZjjJwT1j8ViCHU9F++6NoUFa81V5vApBm4YyJOvryhsLSFYOhKF/1Cn/mlcsNwQx3Psdxfd
10079IGACUGetApUITqEUWrFl4XumvlBagXdhlP20F2ewosZKPH0O6b0M/N07BHeLBeaNSRLmQwB
58bgNfLiDuOj39vYBfWgybZEb6MGtgmCv+x5VGteT4nk6sZYErLFLUs3ioUGuyvi5UFq41IFCm+v
Fod/mUenrNOjCVdvQFeSOngPf+Dcij5A0oqMPbgvh9nemgSw/+tW4YfyQ2aUuydc4xZsQetqfZeu
yY2spKS7fxdtqWjuFqWw2XKBqLte6dgo3Nt0UEYj80LT2Oojx6zqzy24UGyDBcSasv0knisKrLmA
c9QI+RZmniHni+cgrkD7kJ+okce/CsiAPrXAutWYqb+HCCgZu27wAYHsCuXowOExa6z+3/gs3Ydv
4mp0wnX5vipjbwi45FD6ZylTcUb7ZueN1LYe/CTJBh4q5ISTjSe5rew0Uq9cvh2useWgyA0Pvq4d
jS/s15nbLfNfsp7/UIFdVDxRt1onqh772AtHVkoDUJXlbPocYswpo8C1MG6qGPFT9ARReijIUyxU
jB/1mUCr4JMq40fL8JvBhkGad0PQU2P1MQIZEuRClsSpD2AYKsfPAlB9DF4EeaHtFGQWkgx8Lp1t
NjVX9/UMsO7pnNe/wV3LhqdaVj9gGFmv/Cg0SdvxMk0tcxhEk7IPxhuyKPIC5xeK5nqiRIP3ais1
sR41t8BjgmOn0AEe37zv6/1ZdWa3j9paesqpetDpNveLB5Z/LsbZp4pCTPKTr9Ldgfi26bfE2Sve
KRKxY5KlhY1nSBI1hRhPyOLSPi0TGUBVvPaxTH0vQdGOhRUQN44nZsqINLGTIF2SkPBYcPj7po5J
PpdKm463NAAXB1yuUDbZ81BuROsJG29y44O+r5jEdc5SBVGmGUxer1ECsdibmQy/W/J66mFhsmRc
Tjf4n3n/ERh0lhWFusw5t1DuNulfmVOhIjI5BgYx59oR3uOOHjONzLRccFNdJhVwvR//eRMUWf/Z
DIJDo39oV9htvklbqVS00lFWP65BNkTADbCjqDo0q433SkK9ewcpXFHzQlUb6P0SFZMHCEQF8oJB
fkdn17slnQPmy8B9EuaYnLXx3QVqqOeiZ6SJFhiLkUWvSBvPoFuGpaxEboSVp2KMHs4s1GbhNW9F
KGYXFUkY/uJH6sUjFYeoZzT4BGWEmA/jcA0QW5t+i9Ud3pp4jGfUHN4azUfSQ6RtfG2zT6fCiTGL
j73bdgsQ6S3X2p1xK3WwzCoGtJetF3pQErt+7Go66dgiCMfSXqSa01fm0vkxKy6jrKcL79W5vwOv
pxBV90pbqKnFhOrkNsDwdJYabi71e8ivx4XX6sSQ8X6stbrV074OyNUsuaF9Db6D/lxa8KqY8n8m
lXZzhOBCA7qixxrDYoCasypR3ehxuQhyBCtaoG/LVgARai4+JaQi+GuocV9aEKYkNSF3UdhONj0k
FzpQ8s4dhl4da1OEkPybwM3xlaDtmfMpyqsbTC5u9XECpDx+YmCbwvhnajekarMGZh6SLWnW5R+H
0+m+raM3Y2WOAbLyXMXaZW1CzABNGuT8zeYAxYFkUXS2fMsNugoTAk77z/HHXgKYABXsYbauBKfp
uekpyRKgSb0svsu5ARhICE2Xe8R1go2LrWezLB9gUx8L+Atrq6u32vkn2wpD1gRNkf8wuspG9dau
msfylWYV8jeR3UZjaMj226l/653ydyUF2gM+ldNrLV0iQAYdOuN6wWwB31xE7vgBm4AWfYaAZVvP
yqECDXxE3NR8ZNOaeuUGfqGpmPaoXdCoGk4VK41yAQ8UksGan4JEi5+vMjN9kR7OUId8OPOcIVCG
2xrYCCMav22cltiDyDbhB11jVAvZbiJUi1+Z/C3CkgGmhOtnT87i6TreP6cHPr7bxdTEaOIrqhvC
CxC42r9c2a8lMdRbj3veDW+UuWKiZqDTGg28NUfA2hMkZAFG3HAlb2yGNyJ3zw65Q6X2Hm7LeYw6
7WCsm6XejUby0HlTWV8HhsgrqvqFyK3C+GNaUuJ6fKuo0zUDk4iGOjMi+i9d89tVpAJuZbpbapH7
lIZO2ncnGP7HgXSFNHqbiJx3Pciq6ZllR2JmUPe3NxFAQI9HT2yXyMz0yUC1eHRXtLTlCmvG8qNh
1lXbiTPUFRDhE8/PP/2eccg8FvTerVIWTY+vGr6DtougXu/eU4oQwqyaNOzbcdch7FXiWi7ALGrz
SPFOwqkViw46C78+Ig4OJXXqEAqli8hoz5tQp1i/zOv0h6KS/U6PAkmspchvTQFqFqXEza89QEYs
6S7BSfn4tNZHMUzciLjhSFR8womfde34i1RVkCxmdwhPOjEUSUP8S3oG0VGNmIZMlRNHMr9jzyU8
k8cdaurFHqAYSESwYw2sNqoLwqb+tBQBeBXCd7mZK4SCkPOAAGTzZKl9F0cWQbhnem0nkw9PwsvF
2JtC6yHRK5FwpMTGfTuSio06LEYqnVBmlt8wSJtdtWybg2buf0p/2tef6E2A89TD/YZoovD5jUIm
jViHOriYfFEF6dbP/sFalL89rXI3rx0uPf6id7BZ6yIFV88XmfzED0mdnn1ZzwYFP9XLBRr2/PZy
C9V5zwDStx1wy94+TCBpPqev7LnRwL2FR2XHuuqTd1TOQtNJqHNVyrJWW479MH5wLzh+8gqzIBCd
nobKQBygrbRUsWRSq2jlzB5roWrujIBe/2nNtZ72QMcW3yHo29q7I8T/E0603duLtvsdxFVq2LaK
WOxyQeafAAPrAaA8YkTunQS7hFHVwJc9J/ip08d/zNJFqJ31gQpWF98blKk4VRu0egjlaqVgzX+M
Pn6O4/4uwAv+qhacgkIfEeBFfBB2T1Y7muB2GlmjFfGZzxVcSC6no0vljIajcqAdWTOk5BYalc2k
zQ77r5CYqvt5dLE2xoyOLv5r3iFfWyXlgLN4OIwcH8gYI7qFQsbZTQuV6RNfOtqFThTpTkyoq7fC
Uyl4RDsubuzaVa+9Ek8qbSjA/+1IywRURK8sPr9HYPf0fCNd2Rv5aOrNBXcuz0UY7Q73Uh0yxU+C
UwZ0Yo6RcWuT7oXd512SK86u6IHb8fle/qFSDkR06pWhLtPxFkJTMmLG16fJUHSI1N8GvdJZiI7n
NwrxjAfkb+H57e0fysZMh3a9Q49dyiG7CNtbAsjbj2WcoEXoBucmSH2vTxOak39K6bur3ViYmuIH
rDhIAjf0mz5dj40+Ut1WWaQ89LAb03IaOY/K+kf9IUk1PzkaItFrXrRKhgyckXjDFPAkyyakEFXU
gx4dmzxJWR3m8hOUpw7MbtXSRZbfCHwINUmSM3zw+Ws2SWHtzXd0Rbrid9nNILGCXCAk/GCHLFPt
30NroGjXLiYp4swElhktNIJqFnKRudVXlMjDopWSSax12oBxGWlNZXuBcGYy9Uiew5G9YtCihkU4
eCGfZcFqIb8nV/suEm7dLf+06kLoG44Rr99ZOXUu4C4E905MivBz6CSpVs/wCL43seH1yVyRrmC7
VOOT3jamWWVV/8IjOY5Ib3R7zJf7TgXSqmPrLXAryd3vD4L+W5WRSf9JCpPArZDpu6jTTlOT2oFP
GicVV4IiB7OS0oV/X/YyuWH6/8cdMKknN+i/maefpAm7bgPHJ2Y34KgKd6hcDmkDzgEsqkjNSuzC
LgriI6blOBq9TijtEdA4VBDUaITVRVvYhoIorRH45mBT+xDeddQqxd+HCh9RbGjNP4iZZyd4QTFr
U/T9+xEd/wT+R8kJH+G+ZvwIXnGDPuswrZDe77apCMCtF/t8xcN3bb9Wv7NTrULoTIOBO6XlIKhC
YhQ1ba7kpGlal7KiSKJDAcaanWJgmuz2P64k7STvhnwmntkpxMsonWHSPgOiFS4xv9n2UII51AKX
Lh4iPInFuM9E8JfEyM1YZ20coJqP0pw44/zguL1EL9qaDOD5BWKSNxuhdsvLcBaD7v6pwkAemGLd
fJ4eLjWduDqChCKbvRj81qXRSDS4+GwjvHzYf1zF5T2/lULOkIQqe0Fj6lfC3GIEVAmvT2JKGxow
vxG/YoFCy3U/K2gXAdZ7zOZQR8t8ENOYYAj0Nj8oMn5mONYq99pFsOwHNejJaPwLXkYN3S4Flocj
XSi3BdPNChgGJ7vjFd1ZW6bn1UxuDeatRFhQ1Vm6kA99IwmL+MVlu9PDIp0basXu5tbeZEBSuLoA
mVr4qu/C2zihAetEb8PztQP2iwP7Fe2ZuTMHTv4vRmaFk3vXvjuuvhj9oKFKHqBBbM7E0t+pNij4
/NX9OaxXNSLtcH29CyCQfVZfm5fMNI05rv69MvwH3fNYyKuzsV3gs6j5olDOQtAkLbg2FESG1n0i
PzYU0G4Chc7JbnxUS9yzcNDhXjVuquVg8m4nqJuG7rJyMDLQO12PpkFjoAwurmzDmXLVllvybXlt
PfZMTA5CEaRGSKwCSnyPQurVhbOppmSe0nJOUO/mYZ86LiPisDMLZC7+gEFXpgXItIqLOnc+NBu1
pQf29xKjsof6xyxjjXlOZCc2JnJupf1n/c4i/snCLhmad1NF0N083ppdQCofIrTRMVWuxDsnlD2L
oXcH/n+VLqeeNqXOj9T1XQmMcPAhz+qEMYb2pD3OAmjfgUpN4IfzkCcFPHcaLyH4/kPiewoiN4bt
WCEKvXGftz5lQJiQshNVJ+y37L7/BqdktUXxAyIfYVyfl/Fl1zRPnOgDNMcj+Y5AxHjQj1/aXLgm
BGxBRSY9/u1LoIKmouXuJDkBvkT0ntDwDogAroj2Zbvj2HpNfvwbtoQTXYKIB3N9JDpFBSYqiZ+r
X2HS1HINii2UZYhR7PuMX4bhvRIG5dCL/tjr1qgAnor6w5U6Pb93zAqdWABtk20AW8jrJwkJ91cH
qBj53XBhAAsGaCZ4z2XY87cc4fV621nnDRzg/5TskB0DHQx97voERiZhxqbqQo/0Qu3BQRta/EAF
yPhE1PIN1vZkOOmY7QPu8uMFkXVAtfwpVbv+sznGuRhTUPPWBKbgDCXNbGS+Noi0YMUoa54Tblvi
o3Cnl7QAfAwwJzdo+mneso3L56QBthu1FhhAvFicDYhy8ZOIcvdLGAsv8xNG0AmpIAQbnZbdyBft
yOPebXN7YlNe/Y9AS0LQRn05ZOaUhCt8x09kOrBC2CV/0kLXQiwUsXSzoLulz+Tq9Z/bp2QRxll0
Hn652fS15+FCcuip9ZR+Om8z8m/n7zb2VD/YDZfhhOb4XsXW7LbsDw78SnsNp7QDlDea2lc27BmO
BoTSh2BOcSdXqTgzOUBGkzvp1rf7ZBEZjE0QBWywpRGA44azt+9LlpojgDhgT0ETJ5R/sOevYkEX
9ZeTW/Jn+9nLaQdULb/NoensNwGWkJj7ozQf5TVCFiI8Cpm++m2GEeisTG57qrLAYYc1eldzgWI3
sw4gYpLFoGz2P0ACftRVDPArZfGdNHL2holOCnOutO6rpB96DGGmogFlAugrpUQu8gEQuanhRx7G
bcKHQ7QLNtUiOlSsArwsS3q6Kd18sMx9eMrRUI4qeBwBGzTWjtB5FpqQY/VxcyA+MQtL+lx9TXK/
8zARYYKaqVPpbuApSe8VA+Bj2KukUNjHNWBUP/rVc5c8NR29c+aPxlBj2Vd0pY1gAwRG8yuN7HP/
VrR55rz1eZsYQ6mztNANApOioZgoa6pPwDahaxNiho7Y/y6VurmCkTpiVOeBofDTNThwSdUC2CdA
eK/AmsLg+GRkhULc5c8P1SoqcjhdQY3g9qiQMhm+m4biAwVqfuwuKcR+p1YfLrlT82nadNWQ17mx
hRXAH6xZgJKWiGiLVaY7ZF8t0kVy4Dru/+KyBmRaFiwUtJEoOSxbcsCFt/R7K8MrXhfJAcQB5lxo
KVZ4bRQPhC4NCSPlCduWCooY2HUQacbMloT1MIrZXBUpLnUBr/LcHZ4jf36h/p8u1xyRB9w/XEEF
APuxr6Hjk6qI3xo39DOi8D1okdMF8uIbmpY/wc+GVKXWCIKBeJaAkbc77gTbOJJmDHmXuWZfHzGM
Eix008+FfFzp6t+TA7nR3Gh6R5m6lgy0fiWjzSIl3jHNZe+dAeXFtVheAJHqsxq914fk9I+a9oCm
oqjE76kix2bWW+9Yfb4lOIkU26sQ4vYzXK2C8WHhx64zAawwqmGrRExfEgj6ygQUrw2i9H8VFQIp
1maDxfiq5JysZezBkmWAn7tcaqKAcc3qxsEI0rvTEsdT0nUFurO1MFs1ibBlnEJprLmEShvCr/gR
cFqDJdwlKPy9ZEp5oqa2wdY9jtt7JUYKCQpEk6LRLTf/aBAkqeWETg13trq6ZpgNdWmnF0Daj0cu
HhCGri/UdPkdQ+m3TmQ9OuurcOdKJ/9+MTbeKiDsCs+cUXykshmGTV5QcOB2yZtNNL8B0h4xgmgt
81jq5aA7WtvrlncF87PAe3pXsTvjsbRIJXWjGI6rdtTY5EiRaH5++CfGMM+jpUfq0/qsaFf2lAq2
ZcagiAvhABkRph9w8PBiEifi1AWccBFNimoQBcmB3mm4Gs4t4giAEmw8sMQP2fbOEKnp3FUlnOz9
whPKZ5LrpB+S9JxZ8j5DS34Fw1TTlT9bMaY70i2QbC3ggHDr6jUtG5AjJGU6Omipa2SGVsjqXPF5
tVH21e+WX5CTxoyjTLR4Q6PdBNNGw7LxQLTDccuGfQ6o+lz1jV/mOuKb7BB1qyz4OHDeeUHi6np0
T49JDedM6Dil5rmAKQkP5H7ZDDVBFtE6Kz8ih9p7TeSTmWqXFzf8CwgFr5I6naQgqn+J9hU9gPrD
7tFIWTF68zkkpUkyjvZv4TFiNSZIkkqtJvlbJoLFaRn/nnL0wyVJC5HfseEBu28PuiP+5f8MaEwI
bB8EJaMOMQT+hGAN7wlG5gxjdSk9DdpJmCY2jr9iChbhOW6rzHR0q0P+8z9QGtHig+i3Izhvz8VK
ZmLcABlIN0NhqZ0IZC654fIz+65SLLu+z6O0o+MP1HweuLClIxEar8al409GLDlO141aAWfVY3Kk
76ENdoPmzGqRNJU7fm3Iz1lsgZSJm7uBEif/EcEYWcHH28zvdih+eaLmbquLdCm+QsJanfo5qEHd
o/LGHWaoqVIOWRV3sO110ABFph6jdLRzXAU3Lzrng+N/j+V6kQc6FUx0EjLQeOhqVwsyd7jhBytp
0PaMz/Zw0HxR/E8ds+Lbxw+Y4uX+VTmydSJ6240cM+lbtYOrCR/ThHK+u1bpdwFX+CdGwIL3k57N
QOmX4bZhtTS8oPNJBd855xPydzujsTZFj+/0S1DjmT6syQ4IlkA5mViJPHopfZJ4jXdXGDen0CX3
1cs4+P+ODlReo4I0iys8ipToxFnSZXHeNYfXZfMi9BWjotVMl5bW2VY8FPZCkjODevWsZzKYSA2n
kaGk306H1LXYlKYa064jPZeYKZcdtRHvK6Uo1ikUFtThlCoV5krkoVssp5qxyj843+3ANGQmNxH4
4PE3Emp+1zgNAwIkeRojwa8psxPdjPvS14WRIxvtBaN+PXuYFoUWgMH+2JMmdlrlNE+E5c1xQP30
sruIiZFwZ0hacxhQXSnfjRoncYItdOcFhO2DXvi4NNcem8YHgwHAV6GPnNdQiTbymhUR4MXTTjyY
2FKRhwNz/S/gAPsAu24hX8Jh67IXeA4jzG5CmJ31EpK5vrLMPV+tSVjRzEhcCiJWxuRvkzxJm69O
iumZplfMPNJIjdHEmodkppphGbJEpUYwwdms1hxnnGI4dghfPBeuRz+FHDzy6/MJ9WFsLAcA09K5
N/Wn1EllkJjj3Im32uTl1HXQYSskPqWOfHwaPf8EzXkZ++VvSXAFS2yWX2aaNMjcWiq8jIWcbrtI
vvdJtIOdkgqvOLH6uku/iIW37PufZlepVwQ/QtnK2IRHWZoDgpddsA+AcO1pesx0CUpLgmArHmNQ
QoU2idP4qAdEClDo921yBGpIdRnqPRYPAVA3IisSoF+HXjAZ7oIHX0zFbuaMqO8EXxh1Q510jUDx
ufqhk5EHiboSlEI+ggo9OJB6p7E2qbuRNJXeghC8fasTfXR0hAJL+To9IeDkvSEGrFLcxYDutd0U
Ww/hN59EWAkIQZSGZ3m16mxmYfrr2sgkzvIRUl5E6ysIVUN3fNnvI5gSIvxOjAnd8XLqVfk+rytG
AmkBfWEEv/4N6vcMsN4oJqAaqFvZbewLc1BTM6w2hqjk2gWArMU/YHBshVRhfCC/1knvvm++79Pf
BzhiJKwpwbfoTTwRKjjbTql5uDtjP2lOXF4j8He0c910zg3tiUfPKspwRTw4np2pJpkgoQPECeNs
wEPbeq2syLXOLuWc/7SzwC1F7k/FKQ7Yb34ZM3Z9/QEH2sMT5+2HjfI/eaSPmVKCbfkRjfsJItrv
x6dkWFZ2icnz26f/dllt8T2YHgFdS2rRiizSaXSr4NiONtsKQekSpj+q25TeH8LQAUyQv7gS6Aps
8xcitMl85a8yg2z/ewkU2V9bJBL08RbPQyronVlsdeaY4jLR/0omQTtilMsRMHuESkiZWP8r7tcp
DEQIvpbptFgpzW/F+A6Kxu2Vr8y5VsMRhG92V6hzVlJlI1uBCgGT+Roi+qPJ4bYqk4uYkH8ZCAim
UTI5JShVq45Z9vJKHkWJGsrkP08Lt3LtcakAupq0805FS8k9Cvj47PYVxHTyA58ux6zpurzhoEUm
84r1add3U4qDGRjyk4Mpc6Bl9dBdmMnz0DL6/bZl4dnA+c+x2P5sPsWNcQAVrofL/hrbRW40nsgS
Ejj+uUHSb9aNr0rcSuaJz4cTP2E9nVVPa3wrJLbJ9Vwz8+ige0l+2D+Lkw+xc5zJhRUtKTkxeMB/
HsYy9/XumR9rbQVhIFHgbKT1hPbqpoEquhUoqtohEb4Y7OyklisV0vwnLcNSwdMSTnYg4gfrlRwX
bw5OcQZTv+i7IUXziFZlFAQw+O8YtYW7AQzHBYHcTacPfm+pblOn1Raeg++GiUDIhDt+TtLULh//
RDHyC6T6quFZIdz9fMbZ8Ejvg78hq0QhUXVoNku6Db2HbsQAOds0eDqQKJXBfOEH6caf5ePkSNam
XGISVs7YmoPpIbo/3vcHUdwHV2LzTp6Btbl02TCCBug3+zBwjPpT1d0nO0dGMhb5/i2+yKK9v4QH
IU/azNO7paYi57kfNkhOJmhKQ9hoKcbQdGBTzvXuyU1hK472GDvfbwnwIh/p+EB7vXf0oUkx9o3w
COrhN2lX/tUPa/AF49Y3OwjmO8uA5LTsigHY9ycMr37oyGG00VwqHEOpJP3K0yV49UNGhpf7XpGd
hhkqhzx+NkRu8TFGaz7/reThNiCMI2+f6xby5gw/6KH2NANv+/RpXG2zBvDG1z0JzUGqLRY86H9k
bYGcxJ2Twce/xVltNrsAbYBW5z+d99h04KZtpw9PQN/lIOlnUvtBOBrjY1DSYwKxlw90Tborufjr
FhrN0CWhQx0Ee4eqITPdKngSaXxhUFrDIbluMybPA5CbFC5RbmkA+n+ORRGdGtFt0S7kmBfcT+2x
zvocc77jiKcgCPyv9GQh64StKYWACFeHP1zHL2S6y0fQ0LLdP8UqUeHHEUmr9b4nbUn/Hskjt85l
KS+xomZlEsxDqVT4lJ27ByseVE7XHdNAU1QXB24wCiq6f4nFLkGpZ04Y1XCPNQEJHDSzjgCq795A
7HMNSEbU/n/JUmD1dgPP2a+0FgZm46VTIis0MlOFQ8WK1/6Q4rf1D1vuZHdpU6VstvGC8iiMlJfH
K84ttZkEFppnP+Kf3UrZPyVqZ6NFE9qEQcaYYOqUUBqZYrQRgobU2ZJq+eE/xpfzAuG+6M+ykM7Z
qM3G95/1mgeNCTXXKRlcYNkS/mYycayj3ANJyAEd98JzJKesVOCG6h9KOl2VPs/r3PjHmv4Pbm0I
WjkXDFeJCKJFlXGx69knVDJxmmGbYwr795IisaAHmkxfSdSthBVrv8W+Rvy3dv6quQRoqBCGGxWj
ZH8iNxd9fSwTuAK3s1hPYSvtFwPxe5gv+d9fBkI6122zH2UVrSeEl6zNOTc3i0x7bKY2cFtwp7Ly
1vJ3Zw4v/I3CzgQPMFv5TMheKYqN39Xt8RtpU6hLXI/YIW3AonCkS0QJURhVND7tLGEH/maPby3S
m8cOFg8ol9d0jwy4DqONOQDgtfVR+n0TN4Oha2UN+aRl1ZlT/wnwR8ISjKp/zs+XtUj43VQPyCx+
aDYtval+P2bdV+e7UH3sYSU5qY0hWNXmRghtk5GGXFFJ6QChJNXYwwEbY5ll/mS6Qg208N0Bfo7f
jcU8L1GAvl4GpWPMag4jqcaxSVyjQtZioxrwaTGndHWY5n7Tp0Cp8cprOfXuxX0XEmbL4xpXbAxV
k33Spm1nqO3HqtvW4+RcIByuxZ2f/D/Hm3jXQgTRGIjD8Parseqz5UpekSIkAaWb1Ntv5qASn+pD
gYhYObdk7RHwoD34Gn2WRsoPtXYYDPb9Nhder6qTEzuXev2OGGgx3sKgIxw7F2HV1JwRjadFM/E4
xWpP4jbeZy+WoCUHYpqQrJZofyLeiflhYqdR7c/MqhVQNYr+L6CXMqKMI08Mj0qLzLlrh02lHk7r
cV3YaNuytdXNSozDX4J5dRfbyFZEZc91WYXhIumAQg+2SwzJgeFDK31/8M4ty4OeHyDd1I1JlNIa
LYE/4kEnZYx30T9Cy8s3gHbFopU8msZmYBOy7tyRYWmRDyS8zvQoDcIuHpxqArTaNy538DNGQTjV
98o0qG+MFeQpK8zdHyHJ58mpPGVusLna52adi64tIgHfMZ9bOkIuCTlVeYWPfazrWAO59XSDlW5N
H5A3Q3bj6Og5ApY2HHStXk9f+Xe0UPtXxeRhCtkl6LIbDe7alb4HIDy8YCPvysdg1ke41TogHDAV
cQRbZoopYXaybzhoMX+Bw4lIqY6g5BM+64YrVw4huUgvj2KZZrphIsemAFdbcc2GY+7nJ+9R0KI3
xkkqSe7bcZfrT7KcATvrnmrHInLHbNJIkss05InqymX6sOAOy0lw127NjU7dKY43XjyIlgZaAxab
xuLSXxcsJJeLyK2Ef4f1Nl80x8DedN4aGE6rggXvG6k3LAWPUjiVVEfNlaLDV1XpaFNiqLuoJj3E
tOae3LHPSXJRfrPqq0mP4gf7iRJw5fwQ5OWBSGc/SvOSqhYzMNzN1s2/rk2D3/LTiyREqDZyyGqA
ol9WEtGd3VNWcLHNjrnvydcpuVnEjZGkPp0TKLq5mijZzxTPqNSVNgGgWwvzFtRJ9bxXmZetP09V
19mpDiH6bNY5aRx8h5L7yoWp9PridMPKgRT57suYUI4s590MjCWVRe15G8VqBtQufAWXOg6Pv2/X
U6aFY5Vm0eg9ldfNQsHUyuCFGb5qq7I1yxKPLcylzwK1JdBVT8CIt/1mXNHHYF7BZMSiRQSWBtBq
IyFoUpx81KNxkqXE+XmVyKyjnXI3iSnqOZOna4rGXa4RGHd8f/6GtcNdecF9OyaFG/wFL/sUVPYg
BSWpH/w5MhUoD92dUAPHPG/dnB0VoZFNAJzlkorEx2BA1dtZM1Dzi+BlXO5K22hF98Krdl01FGjM
v0GDRFwH5uQA7wAgOl9XzJY+oIaH9h1uD9D1QdaI/cFvtxN2I7wbQYd1mk79tVt87AvzGNCjwoEK
a00FrBanhtnuL0wS+fe3C8u0yDu/frBtz6yqzElNgeqrZ1404YGjKGpV6wKaVnnCuyhPc2pKB/ll
l9skVJqLhWelNvmwBbrGvZlYQCyghulz7I6NxZLxoyDLnW7xlec5uGUSF+P9sz/OiWn5UgzxOEDO
r7fParlTCmgfDz13F8wtD+CYIaBlaKDxzVkUj+z7AKhVXqZXDSeDru78+tPc33htid9qcBb+okBO
n1zT3OFXnp2+JiROB3T7rGuQV8lWwXvx8uqHPZ5Teb+s3KAnAaZcGFTaj9L5WH16EWZ0Zng3Wt2R
nT+HdaZGc8YHnour4KfYQP658lZ1VynIeDgmEVE5YmeGwoS9BoUCL7awv4E0pkqqx0aQfhv9fDnu
oLj0amwoCpi/+Ky0nEYyOpWY+TBUHlFflKbfZY0DmNrExGanafQuWIV5QtvF/Wr3QFGR7l5NE132
0mJqw3y45jSeF5bFhrH1TvewWGVInF/RjtC0fZw9h3Gapdvxwa3zpAt/pdExYTvBteOkKCnPP2F4
JhCDPPjqT6IyDYjF/l2eA6Q9boAQmHPLIKkxxNN6i7d2VGcO+rUWEtKCzNpR3WiItZCZhZb2pzTB
vJGJe0hKfqce314aNY46aFvtlyDipOQ7fDpAaDIqHsR8yptzQId2SMwkV0dHCcUyvoRJNzKuhGcM
Fw7HPNewyQanIIGOSHktmQjHOzUPuAgLSOXlI1k5hlOaTChftT+vDoRyWKj8BKJmRgPTFjfguUOg
Q/mQJt58sdX0tHc4Fg1Y0KwW5+9GLiLJQVwuLxRVSqP9Qxl9tmJ8Rr3NphwGxOsL8YqiZ/Yg/njH
nuB2VGVKLgUKrPvBXjWioSug9Ztxmz/IyCKrqhCqsb5u/gckHDu6Cl5J71vRjTRDzI2knctOqesY
NmtRRk94BQBH4uRbNJsqFqhz0P5AhppoOdkAO1pcUQ4pQEDNi36wM5LFrqoWV3yZXO7w3Qhmx0O6
BnxB9PLEG7fn5FwOkuaVil47aErlHPkZTQy2p7DaJ4AvKgOTfBBvEKLueKkbksiSJkDOrMfD1wmE
t8d6kIuJ4mFaWDy4HNZH5ISoAHDm5BQ5d6Xzba7nUojXh//jbNP0Qh9zGYH56Ix5L7EA/c+ukWW/
yJYeII/hB1dajiahKfWm9L/AXcvReLAoBF/ugXD5PVmDog4gjG0vzcQDjWSqMq4loW1iilUC4iwf
kZVAvf8YQ0UO1a6/UtcDfaYDB7sPl633aqpnsvJb292rFbhLosNj1hCF8Ck38TMWDgjD4/Rm5gdd
iWoaDLD3YDGM6rZRdEaQJy4LtPvxOtnjtWaWglC7SNPQJrJvuO9dsZf6pTSpUQEpzw+WWYmbOy/7
THJHhSidSYGKiVTC2J7gfaZZi/+XDuJsAr3CgMOI4XATBaJt0M45tqDZ+uHWmIgY5dDtnH1X47u3
DSpptKutxisgEQCSRo469ILsh/eg9/sx/WPIwyOOH/xYqv0seRrYmOzheik3R3+vNQ+XT+/cYon6
3HCyZlQBIS3RB2Tss6KyJzXqdisvBJa0l2nqIR7hXlctktAnPWQcfzxG/yb/k1HrWYNAdjPB2hzR
r56BPPlInR01rKZFyyhHDAPzlctWSMr84YbvKnqYlx+Ny+0CjOPcGaxAuKTLL2XaqkU33F6OrzVj
knTSC0ckAc0PO9lN4B0WGG2KPArODlRUavne/ZRZ7j3whPeHZgxuEVLE6P6nGGJphWLBhG3ZCqhp
GJxc7p97X5mYS3nX0y9YbWSX6lG0IUIg33U6kIcuT9muOe9sXbW76j+Ii6toQ/KlV4anPmmHGqcQ
YkpExDUjPC4bM+rjKF6ULGZcqHKAl1IScEahoC+O5cQrPutJrndt/KswLMOq009OE9+qbD9vcZA0
9LUPCNpsb9QoOv6cr4uyXE59aPS60RycL+Kn/YLCcjuTyRUTUwB2+r6h19CL2HfY1wMLDk3xWyeA
zYanOPFwfrYJLG8JeqdFEmOH8YC7lhtawLO5eihehNw+oOBBvpsQTXtn2jEWGvSwDPDZc64pnQdV
lFvhqmk4qWDQASPSkJbqC6L/HMgYavhKu1I2Rgg//RWYatQ8tkHFgAYIzRWzJftjTai/EI5bVJe5
AAHijQxHBMMRK0fupdo+165K+ZKVbJDxlqKuXKC2AbPACTKmvEPFDTHjFL1SejdN6gRWTXCZiQ0b
MYqHZ+h3zGrH2sHjUGv8sKV/kSjSy+0QAarkHWONF9NTV4YAhPPPg3wQpoSU0lGfpLLwpjXe/+nd
5575nDKr+Y0k566bUOJ9VOOr5/Du4PBmsoo2U34bUGvBJDLPUDzz7bJ4KXRDY+EUO/gZl5VSlZTW
XbtmGdd+mZ82m4QbkFBW0JzABUFzYLIyJcYJJ/qfzkFc4L1FUThyZbutzYxB7NgqF6pbVSfl9UvB
pEF0CcCWYfq2xAf2+bWUQc2BjckAdgu2OT6FpCCkSEyIGbNtrUStw45ku5Md6PIV1CaN5w2fX4Be
DnPnPns/mioVBkarJUdbtF5cXTsnJ1evyoKj3SKJ1dwVQY6vSgjP2QvkAMHDVJ+/VtSrZIUW+gQf
lfwdAfWMk+xrC+fUfyK/EWIXx3MvjDF5zwMqrSUXEjPNlk7+cxDNWpSM+3UaTtLlUeh5JeDiFXcD
W3oUzoQnHJS1LaX0/gPsvPWkCXRG4AOHwB3rWYilXt/RdcofARTOtNQfnvfUB+6GAlfXejdG4lVH
QBcDvvupwiZIj8KJZ3L1nhQ0/Pbe16//j6cpRSxMqcnK+yOVsAd9VT/hjoclLY/yy8TzURorRLj+
8t0/KVKFDV1nM97PYwi9ijJVDAvScJpGFTJOaLoFFc5envDB2raG8vNZUNAmV3Lhm9oo9VFQmFL8
DxXwGGezOn/LQ38q2gQbQtWdjFZ9AMEWZqZ77wc4Us93AT89RGXfUg1nRGlVJpk6RCFb1gR2oIIA
aZBcJPFe1adDN/egQ4CUfHGSmto9OdjN5KYmfkSigkPqKsByb7l1Qj/PejD7I3RYL6TkEST3jfCH
FhbY1HpfoDE+CvQvzdjEwRLNmj8HQrEQlzmuRHK+n+7yVv24mboi7IDd4RavJjphnNc34SQuUXmp
JB9TPdF51Qt1rcZC4Bm0cITzGXfRK1UXkGdWYMoEo76wpP492a1d0mHwpzj+Sy+YLZu5exKvoO7m
rsqyVNbv2jwO97gwPUvuu/pzrwYpTVzZbzH3E7KbUxPG3W2DoUDPDxCsLTAg4GxrA0thzPm9CCZc
FjPkTl53/36N26AEcNGm3PQuvOJA0228L+96JceWaH0jqzVIuUTuzDvHzbi8Fb0AQ/hJyTdavKBc
kJ3NCp8W8WDEOaYSxHpvCjHpOm7njjhGsqJt9UxgpyXU3XCkiI4jacpsnMWeJX8FzvWfWrvOt8JM
8QIOXrGqSRCsXb+OULIm0zTyrdG8pmRVFF9p4j/Exlj8AHWwZfZez6vHR3gnRZA5rPz8nHHA7OvF
TGw7NUhoWL4QYvaA4yghurAVJM1w3Uvtha2ePtG9TP9RQcbGBro3YLPmpseO/ydWspcva/2F2Gpw
k7FM+wP5EZvGae9KGhwZ0j0nypI9PdzeujVuTwNLZVFGlxZf01iC/gx+nM1B90drVM4AFlluMV9w
JUE+cRIVtHJuWqIVo57oNbhaMRzjsGBzdi6DnE7yTHTWxUDIIKzX3MbRPpUld2495Jfe04i+QQ3K
4fDUyjkTjk9IH5QEoOJC0gaNCHvnfKvIbCGR70WO9VFksKkhXU+1hwyfXr5muMVeff0nu/VHaAwJ
OEavo656vLW9M+QoK38FAr9RYzZEOWYvm+5Bbjkt8l5+Ja7h7RyBFQG4/URY0l0ObSVRKI4+wDsp
MbCC8CwqJtgiISeKcpYr9X1Qdyh5m0xmSiKT0b7v92Fh5ORJIis6XMGsb7ZVF8TEhFYikXPkmoLl
0E4Vy2UkQ2yAoLZlZq8jdgZpkyhalVu0+6RuZspWh9wIjyey8FYrHWbNangJqYAITAD1ijCKJa7Y
QKTi+lDVVx2vASnSTi8a5g9M2G0Vjm/mlFPCRhLkFiI1x8Up8nln3iybN20xEjKmgRA77xTWEGVQ
3c5U4NuliUQMeq4Y7yM2LUx1cnty4YDkyTRrlpVpWdz6dLvUOaAecNarxqpEsY4hcoGwR88Dr+lt
zTLzba6O3eyTYem73h2rd0vBcpTDUufQJKNjZusQd7N+zUNTHULp/AFfKlq6m+avlYhHzwIyIgcp
1GdcAn2Rmx4f9ljD3D6wkLnT7YubrAveyilsGY9G/e+3kk63OFa4bcDkuES8DDz3kXB9zpPGyjC2
U0V8cVa0Oy00aMRTM0+tZC8aTPoxbq193oPSIctmc40I7lNVMZYRDQKKYJ8fN0agJnoHanuszmPL
RH47z4w0qyJ88z9zobuMz5T76Xq70oaUWpuMpq6SaAJZ3g+RW7N/lGogVTT49Z3PoW89A+FjUdZa
Ihj2TsfYyWdQ6rNLfx0wgLv2RWB+QZpS5aSuMg32uFr8ut3rGwiXxI5VrIMKTK7iK3j30jKXyq8l
oEFyNw9AbI16UiB4gyUbp/uill0p6cjpC2q7fRrTEbY7t/jGzL3wg+0oKTAlIqnJvZfIzjq6d0Fk
hxpXrmOoletF3mShjsBFkQri2SoZtwdXzOzVx5h2KcOvPtxfEqgYu+bePE+rph/rMSdx3heEKHY0
SvOkKRk5UxomsldjLip3pFLpFINEEVteS9r17oc/+mZRF2M7vokLEGV+SdFwRFYB6b6BFFsKYwy6
2J/V0j1i3T0tOcsL5O51xAtf42gKSev9Q5/EZP0Bp+JcxmISuuUmuCRvM/MGC+wserXiMKXHfqyk
zRegCZOMDAizISwPdYn30eeNZIR+jzE9Iz0lBFlvgoNZyudThnrGiaMInboy9zH8ERXLQErGZl/2
SxEAgEzu4YtzNtcmAY7XD+4mB/DwhnHeVPi6zgHnNfTVvGr5v516r/djes42E2oNC+RqsUuNJRJZ
x3rWjXR4FKvPXrjP9Ezy98AL1mgHNoiiqvkV/uwWk+VjJaCIVujWoBWCtaAguYmepUpnZwthUSIm
NQly8hxE5o6fzi9eYw4VRPhIgEWcl7G/9I3u/1/UmMg1eT0aUwJOJsceEx/4489xw/1azTUBtOzF
w93r93+S1xDv4rdCFNaBU0Ya9ZeYZfxyJaIpG/dOyjLNY9O++38F9Ig94q3dGItO2rlPuQwg4DAK
pDWszwfEs2widl4kek8I6WeyRQ6+cS6JK+YcBM39G3943r+3ahfST0B02iovRr0xNZNOU552JXwx
BDHJrtd2rWWDEAVz+omYyJSnKFMNLYeGQCfJV9+NYZ6gHzcuCuPsrqV+sjzz5OSUmiLVh3Wh8Sv9
zCu9XyYN84C6856S0sceTGaGsuS8i8kIwywqmzYBprDZyB0JMfG44ZWBTR1T5lA+SxB9Fj3+sqyH
XxBpvKm4nINggkuvLnWKnjnn/ujM0sWTgeHDgJ8Jn/EnQaB0pHitq0FYcH0fPt+sypdE1G5YCO8d
dqhfoAKN141Ljsr+8Vwv/M8uJJYUUp9Em61WlZ62mJTnv4K0f8LXy+nM8QqDvAujawp3U0fVIkMl
PaUTez95iUFoDdppWykbyeKNsmcRn3ZctWT3PaUQM6p2SroXiUk7TdtKUoT9KfS3VfUGST1am2j3
Foqjn+5rjFWTXKNd5bs69LnCVdNe4SqAsDR73aeo66p6PzbPgOMZzf+fwWAiyddcM7tV2BjzNB24
JhI4DAm9w+pWJJ4ywtFA0BrlK6hdGBHCnvuDDKrq75F02XvbTwTajZUX7UbdDg2SI9/Q3YWFZG2c
c71/gDGihMLNfg4I7+Fc3XknDL+YfZjZJG+JrC5NGkTkOZL4rEMYGnWnFWgUhcVtwZ/P0YA1cSc2
79ek5rbdB/Bi7b+YMcb/kGwtom1VEV5ZVsxoigLT0a74NxY5qoO2F0xURNqbQJVVoOmjy5CgVvwW
ltnYIL0VbK/ha9qCJO690IbcDjqzSxpSiTusZT+GCuu85m6XiR3jNKKIud24f3ajO5w532zgGega
TwWE1949XXjEQ2ahTaR7tbOmaXolRlmMHmoLz0LjqhBX7xaUfQ6m9TFp6o7/neX5FIi7hEua6Qdw
4mvYhQ3YVtRfGnCixhftL8q4+3a1lCbEJPn4zmnDrfRH6pkROZw2dU6toHU/TGhTdXs8PEu+5BJR
bxRiQRoNDi/voYx6i8SZUzwmjjwfHFNuvxsoNRIXW2eNtV+eYs3NZgACDoNEJ0Lnech7VcnpStcK
/kyv6XhThSED1af06klRQROlCEZImXrYG3kj/zz/hzHOYYK66zd3E5OXnzCqzsSX2Kh3mZ0PrFql
xiLUkGxom+y6By87gAP4BA1u6G+c3OqV1xZnWCLmeRAZCnywRlOy5hQ0+G+DOsdsHTdcHryrkMNy
ArAXcH+/ToePWDcLQjW6lS7afLjWilJQKydujwf+MOqrwhXMmXsA0aOCLw9OSAoqxup/b1/BfaDZ
UamDp3VLNLjm40C9oDb2vh93jr52Z+Xb70b1eNrwrZKHkEvQ0PFazn3vqOgd1bT6GH8LkkAx2cYn
lSvY4bQcqK081htEzwU0+Gk0lYetZJ/n/ys1N/I24gEPE+emt6MZTHzOTbiilAdsUfxT0+81ALzs
kpbxIF+MVp02mc5BhQNpZs01zqaukaJliZrLXZB7hB44Q5oZFoO5Ksg1uaOFItxo0d5e4fUHYDyv
qI0SynGZTwaipf3y9aSzVOYMUVmziEy6C5+2CkvGutu7N1CcmVtbw53p+R7gYsrz0m4kbuBSui3h
9Sm/8xlT4fZo2TElPXhzGczbbNuRNZZR1G3m5jLiWsKiwMn2FsqSuH8LBHxq4Q9OvPeXaZtHt8wi
6OG9lZwqnksduKHNMqlk5PthKfvHrJe3jcL5uwK87teVGuv4iyNT+CpZ4eX6bkZQ9ARvNtR86U6H
8a2+bdg4fFUMt13zexBHP2R7TDXKZrmizRxSVo8VV7JyFcMg6fVZVbcXEW0Iq54B4XuQ2SQcbvPR
68xBgfYrv5+cU658/ygG9k3/b13TZyjHXcrdTEMTC59DzsAyWCtHqcrGtIlRAyt0mT3pE8H3c1Oh
sk0KiiHVSIpkhGgf4IAW1yMu4ZwuQxQf9lkweRwdCvQOQHJVtTYvp6fQJBcbqIN1gajv2m31GKQR
m0YPTRn654quLtrWGVu6BPQ8m23ffpY03DyG4JKew7GrL83KmBais3TkmINgn6LroRxXMwe5MJFa
i9tpE5bMjg5jWwkDzniPcXjm+thcFtcOe2k+yYGQRACDKsoIn/b2bfwAs2iWrEywefgFpJ/gwfZF
sQzPVlLUS/Ctymyf2K3pIqqR80ka+p5MD+RHZaWM8nPn4172SDe2jeI6mH/MjXeyvikVPBrAgD9e
wRzsYobK39nBTze70NrMnMybyQy9OGfzHWpO7TeR1M4G7gp8yA+Buy7co9YjK6sn+TPm+nljTJww
IItlu+TJn10i0/ZJsgCQVCu7FLu+i4t2+JrRwA0D6HosO9wtjGOe+TkUOqK2HRKWa751dqMUeW8J
nYU964Tyu4Y0E6AePAWszKH5ftaT7A/U8f7USresK1Yw0pNEiaYgdwD1s3FWnEJ6iZUVsfK0n1OC
PtZdnOr0usXCGtZwmTncgDcKfUfhrBgqHN3hR7CasLaJXjMQjkFOS+OTTh6ZJUtn5v7RVYKmSkSX
oH+2qUfihG5NYcUr02bKSOTmfVbqM5fOrF/DwFwyQwR4/PGciQY0kiNG11eogLMYDEPXSwHZQXJ0
OumaZ0Dxt94cBqfWNt7EoKdqIZ5yDZd5efODf09n/yx7zzA6fWrWtJ5qe1bodyg1MlQqGMiScyvB
vMzd4+0ufOxEIS1JPnwaMzAg2s6xWSGHBf/t78fcyuzc7zeh06ioFJt2y+h2eL0VtFx0jBcGz/kv
clhUnI9WgCW5sj3R7AKm9VHndsGxK0oEOJK6/ocfXA5o1OQuriaZTe9mEVtp/E+Qm7w3GF5agAVa
iXri8p8eDvWp6264RhvQqdJxpLap7nHrfJ5EneIlUgV1nkC+6UZutilXDgbGdf9o04n92rK+qEdY
tXfeAL8h8beDRnA+GQkctNPoJnp/iVgVOFad1qxj4eCRrC6wVOBK/rB11jerPZhUgNJyCXQDB3Mk
LQRDGh2t6Ck30DPxHDFNCIQSsEQQDUNAzcPYaQWLgd3zZlQs19cBOmcks7y1oH4sXMVWVnt5pQsy
Hbf5OknS0UJ1QzGcDv4KcSz+Y0SWZhSZU24cydTSd8DxuQcpHDG0S9tRDo/nJwJzu0hZMh+9giaL
RzZDRiLP6GvETMkLwk+SD+ukyiXLdgG9eylCZ5VRSsaJOOrEkiXMDYtHpF9LPS02VrLjbFt7dSKK
vgAjCVe7agrY3RI438/lJm//hI5qdxk63G2UXSm+E5LebsL9vdQgaknGDBC7CKbWP/altkNGp1hN
nHwE0Shlrc5/LmdMXxd1GNsXibuJ7PKELrsvnQP9bMb8mDxad+Ju+wCdz60GmkpkU2VAvlrW2S8u
AMotGYgMKhYFms1RFE0Li5eeX6qFXbP30ErTwO6n34wmxngLfg2ZGfXiLlFzE2HhxvSjQrsgywDn
EkjIXaFfv9lE3pY+f09C8CZ9+zn6Azniq23G8g+vQGeSVSJQ2V6uFtsAdSBtCmgUsc8DS2F9XjjO
V6dIT+v9Bn7cgHrIP9Q6oJyDEzYRM4YR60MbhWM3iIE7+sl0DIHr183vT1fycf4V8b0FXvORlTPx
LzL8eKMxmletvdczqTGcoRjvA4y8+ngUkwigsnPN2rap2KdniYPsiOVkS28gfGA0KAPNFkN9ESKd
hAFLQPmxERlo7vyZzofEKCW+Xd74vX+qfsHdwBeirI6rLvlMLYPrgUdixPggTNgW8SlzbYaJEJyh
L48MUUUVnMlkKvrwIZKz63A0kVSp80jx/XYOK4V+oBfYiQXDztZ07LOxW0REY8DgeTn/MfT/sFhC
kWY6AHUEVMfPESvds/dfpwOmv5b5uRrZvWwOo4veMJlR3ZvuOb+XIERLRqQjjIPMLDAIPYlsjKQV
AIYf+NXnNxw664KgpmbLIMDmuw9AKI9b5QlaRpvY7oqI8d7xlWlFGJPLCScPpGDJjSRRtX4R69DI
eR5SZWrKVvKnl6rCkFYT2mCWmddFXH565McwElIqPj0+GiWcn+zsQ+F8U1bcIfNr/34sbD3/Y4+m
9yDzf3Bg9hHuQRRI7K+ztK02ipnAbLvWXYexvVWJ3f/40DiCJnnw1WYtayBQdBx93ANPEP/ua1Sw
MwFBRvUQbHmrOmkgH8Qcwy2dsng9d86rVaRcI6y5L5KyX0MPs35Xe/keWz4wwz4zard6soe59etG
7SRsXkppvlMftJq396KfwnU4aunxLkY2ohSfyBmoZJ3zJpFBDFalWhkih8vTm7WFW9muwzUd1hL/
/cekRzlVxdHQUvG/0Myr25pDDF7CCo/C3pDiwt3w3ETF7D9hQ6w6eaw+f7Eqk8oR0L9e8QSOT0kV
sJi81AHvEKS3dt5/ZJ1gqFapMLGMeUUhAnphE/5jhahLhYD3F+y3g0fqG2El8uOmXCZOQmSFLuQ+
hcBNFlg0yeKjeISOUG6R7XAWR8Cp96p6jEBXQkgltUWQ0wupU3Isgl+et8CIARLuxy025ZfHkQT4
dHpy/vxnLssSv7XfDn6HAOCxo4VhVhJb7fxKRcBmPami9E6jewIdo0U97ieqcwqPUlfz9Mq6xppb
5qwZdmnuQRASFIVRv1k2VxmjbBRvl5PfvA02EPx5r6M6FAGnocFtN++LSmKy9FSs1DsqKC0AUfYm
YISWCDoDMxOzbXbsigG9i2x3s1DDsDIZfVPYPrlSBhTBx0244cwoyYjRRo1jPhDXf736xHtMTJWt
7EGXh67j6AWZamNzD9qNTem+qI0rZH5UEEOMG0Q1fw/ccHRmMDUmSsRk1THPpcajL2elOlBUydY4
HkCn0uBHYaWlm0duuaJTSzpIFgoAcIWvQd8bNCfYoqxm+oj0+n+ulSSuPVpQty9bJda/nCn/G46W
ycEFHpJ8vOcIg+wkVPsKPiXCqlRgahD20m+D6/c/Kr0ED8qpwwpeBijRhAfJKY2W9lyS/YtHp40w
8xaD71m265dSiXEae1+ungiIJHL8hXuT+U/S306QMHXGGTfM3aGBHnpah14mcT7hnSfGUUhwRDRW
P9WCUB0L33Oemln47E2BknmlkTuCBC6rZLd5qt1J5gLULljhcOWFAP8iBxgWTOG2/VlKgnvbG6/q
8RlE6zLpIRiFD5ZRAb7pEzdfIzd8E1+GTnsjyli5BuuECYCWk+GrCB3c1GVK0AwrTo9P+P6ZSah+
xm4kVOe/bI1xLWGJVHZFeLF/b0V3u8hNrqHr6wUyYDVdeF0bHkCgsQ5vXzkS9ikiddrNQ4TRr3PM
Esqn2Ui1P7O3wZsHxSgYiuENU37o2cJLeyQfTrIdPt/Y8boWU2TGWWkC4CLPgduPtqmyLPbwrSip
6WDrzsPjJZTHY/3Rec8h6iDTewDTKhdDvg6d4Jv/yPoxGU68rGBpz+WBp+VnxoyZ0XTbW7AstXjf
Ltye/1hV+eG6/Ib/WeNNIjqMTab4Nf9m/8EIbNc+Ylmjy3Asan3ujP3xmlWIFwiOlfOphCBtIpFb
z5kv1AmwIr3lX4VU29l+XkdGSMV4HbuMwmdl/NBU/sR30vgDn7PcD4GhP3A6+d04SC6bA453bIuz
S85Sai1p4SDn1cBDNI4vf5QVgVVNjKGirYFjnBSeEAPm+VffzToBt9wdhXiaET/XMZCZ2eGXJpS1
daztctOKndNG7SRChX3c8kTCFD9wwSYI7MS8cyPxf4T2XqFH+XuI8jg4hBCEeZU+H50fLY7sfMUr
FE5TsMWM4/7H+gEtSyl1Ke8k7fpzO0+jXGMGDaFOHi64RLKF3SBTiEVgSnPWV59neRrUNjEGF4T6
GKk7SX+4LMoUKgUb8ql+ZxoxKCoNueaneFv/F8sOTVTZI/wz9pPFfblzvmThkB/r5MC8KUjRWAXH
QXxUAlseACoMk9OdTk48rZDQh4WCoSf/nhR2JUJf/e1S/sHwFZxus7KVQ+lwoaa4G8BIZBd0/b4/
8tmCjwYsEKjjfVNrkDW2xW0HrVC6yXwhjMQWmWBQyE7BAD7rruwaM6KDFFKQxnNgZyMGRbjFABRI
qHXzZYNXzCoh0vBfjF1XLY4FqyaWa5V+DtyhGcocTub8onDX+JLU548qqNWc3+9C4PCv4yJg0CME
1izHAfI/3gs5UwZ/xZqvnewsAua6DeNavku35N84bVNRBByKDYR1uApS4sVGn1TmVmJcbR71bk+p
WXyFCbwL+GeqI/LFMmqZIUswsgwt2JTEUzg9xwHFAsaskwvqCNaL3YvdkVsc3jlzBpg9cXm514Mz
jAecvmByNXw5C5+PvI+3Xbvlql3rIWkOsdRfe9vDMHCijUFkQUX6CayLHlGaaKUMYydcUOQG48jd
7V2DFm3JGbnRuXef5D4HZdUsIcVAbwSVLfq2FFLtdzpNiAasdfGT/DT8qCh+XnzEE38/jaB/+5m8
mp0Ax5Y+MD/t9UQHw+fvIId7DLrkiOk06qqtdceKLTzTj7m1HQQEBFE2UdtrszxmELKt/9454Ve5
v6njBR1ROSX+OlENb1czqo5db2algBeh44AWNjjhg4zLjVOJqkMJi1aG7PGWM5pPWxsvvxhJz1wV
vNo1eExaDYdxI6QANjkLXDd9rmptgexekxJYcOsvpvOhI/hFE1YXCQv/45d782mT6tWLjOIUdFND
fGscWH2xkGgJXtr2Wg85fmb1uQhwIIuO47yLzegwU5/UQ//EjF+OfI+iCKiq3++eu/T1+65Og+/0
ucsj3S4mD6oXLbW0DBDcUIW1IiWWrzbeEd2JZCnEtr7T+yjHUpT5cabaIE1p8jjPwDORThmr8Btk
v9LtXur40Ec3mvFUt+EhvVjTKw71mk6BmEKBi5eWi3HzV4JAnyO9difV8SVrA2tA2rWYe1Gwh+Ua
uHoh6F1z1Uq+jRgzVM2sfRlymdkUgxt89NOgggl/WWezT5/g2Z2n3ttInV0QUsxjD1z8Xmw4NIGw
dw5XRimqN0CWlfA/hpq2Ish6KDdbShJYw0LWxtLr59304l6P7T4z1P5Hz3EsgffK4ZwJOdoVRU6a
AJWoKaaptxaE0SIFJriXvvVNpmF0BkBQ3Xp6kXJ3gUsKM1nNpo/kPy9rlTgvNCiibfRg5v81ftHB
49B8nhUtgJHcF678RBmx+b728/Nl2t19z9P/M1eAd7hv6H/9EeGewd9JoWCgdFMAGn/ekX9YlxW2
2iU3JV8dQQkADl49Cmv0lq1XUc6nr9vnBbphUZpu6L/ZfF4d6W00OW77FQgvqYw13ij7EGA8IS2L
LnsI1aYD0e8KTZdP+fRuLD/qn+dmxjRP/kAISLkigDQ9LRl55nvDXNIPaLlzJ+/MslVVfTTkJs0D
0Fp7z972bsyZr3zGfcGQLLAiO64dO4PtlQwDR4N96xTKrzgk4ZeRBReqA/9xvTCOspTItxC+LiaV
mdj7dqokoPrUCUNZq+lVHkYBTSYmCbyO1u763a5kBHNVCVe3vnrk4fs9tagcafQFCUj8ESVJ2ov2
1Ff7mHAKcsvqpIPATnEohR9Me4hMkFbJQ94uOR5JTzzXYyGmtRUuiv9yUHUC10MkmO1blicXrLNo
mPmXyBo9DrGUif02IfpkTJ24RGi6WakMOf2zQCvf3oIXTalw0czZS0OgrBDVCKB/lgsNHfHrj+Ne
pOpwB9BQJx5XZ7EEQGL8Nmsq7z7z8Nbsvb8QYnOysNdkb5wQFNSMmp3LAAy+ecIEqKBE9wYRFMye
/G5aTBTQLwAkeou1s17p5J50/XNxnrJdYUzUzCSMwrynnYtaNpupTZPJ+Rye8NsUFowIW7mASm1A
F2lL3nXdtZsntmfNM1RiauFoX/fkrG8m0u7CN1jqnK2CjDVYpMXHufs0VzKUpf9jptg2AmAXnLs1
NHyEjWdrIIAemQHg1emCgSMfd07kAX35/HdM3qnSwD0RDrgw6ELrYdBHomnhO4iXlSdEucIP27am
zRdD9EyhVOxIW9VNh2VWNzbNUQVOSCJh/0ek2jcukqpWxO+D4gvTyun6x36W6qg89NUKOz1K6Fjd
KgcxpmB/0qVVZYqP4ZVGTRyvr8y42rXK/YRX1K0JfnFZC0JR1HuE3mhkw7aee0df2b2WbKkvbOHG
ApMfyimnNuhxbG8rB3NeIBWkk2ku0gSCkUyXGFM/nUt1iRUt8KTbEp+n9S6Sx2NPWhVcSCKa/nsX
VWmouXXOzYtnoPHSFPRVEF63xKoq2aS16EcXvMObcPWP3YRmW3Ms04hyhZMb1Jjfkx9lx8d53B2f
Qb27OgU24Ieetr6J8wAoI6n9kZYxgRb+QiN1qOuEgM0jkmBky6E70X6eDeXOhyZjeSoaRJHIkN5R
sS6nd/uo3piH8zy9NKWi5xmKObw/JjB400OwfpFFUIfyggv4pKXWUn/1QNBSwdIvgAiZFoXH1b/M
e5vMO//LBiKL3Y6+inx+FJtMVM/c8dosp+mzSRIJefCAooX7RNbnTNn660NoDHjckpeX8+Z+YHm7
QFKzhkny4ZNz10nEV8sMIt4cKGsUnnU+nJvvISTC7LTmbJGCbaorVo2PuGJUWP8G+5rCQQllI3p8
cSI9HRryIVcwjt+JBEWKmaGQK/KhsAJfv4wND/PWgTRi8dSgiawsbgeAf2SVcRfbwhYSRAqT7Svh
FvGpyIyC+m70VB5HT4Uuv0RuhbvrscLIeluzdaz9Qnb8MaBkshdmZlM7LcFyzrZemEFD63C0URQf
IK36AcwmMJe2CMUA8sVIzX3X+DzTBLMTEoIQm3xgsAmP4VD5sJpVA9hAeSAAvPcX7O9WVBX+s0Jo
T7gJd/ZimJhgmTk7rxT+YfV4FEkcT3BHNpEgN/co1kTOeu5CXWl1vGs3BmtUvnKDzxRALcNl7ban
XFzJmXcRx9RKv9R0eZY2susf4hYGZDHU6KccSysTebZrQZD7udfXdCyN8bGQpc9bwiJy8RV82zWQ
1b3ywGrWqTvriboSVvs0BFvaq+E1pwnBl0mgP+CYommJ6roH+7+8uBl333K8N0gFHjOVCfscGNEf
Yobe+Ud3Ybfwb3YNbbmx9b+aQJUxi4A0muxbCd3n4Z9dhzg/NBKsKWiaKzUCJhyz1XoGSWHdjqED
/YlSdN2NnT0BybfzG8gXKNnN8E3jZcjYniG9znL3qZc44c6iPLq1iNaXG0p1Mhfl0ucRXCuWkziD
hg1sLDisqgSeJsrDmofu55fynjl1VHvc9vhfYC8GkhZnUK/WXRkDCDSKaDN3YvjPm5muY+/8PetB
OHmNgrTY0n1c3ItGj95xTz+agK2yA71ZNyzVE7qf+lnBwmuopdro2FLrs1Ze+j7FfyMUeAp12Iwb
tdBbasbmISMjrMS5C8TpnF1r6KxWsrmrnRh66jZ0+SFGGZLsa1AV81UZdhNowGWviZr0QFzCEXn5
Ca4DbOK4LGBWJB9Zarx3aYradwkiPvJtG64QnsybFtTlnGv1Pkk2rwM2R3VJZpnq7CBzu/nupCQn
RuaKZuVRRYoPXrfJruEwHftbxIy6ev1V38HhKWAguQEI7Kry5Hk3jgMed06DyFp6k71Ro+dGz3bD
ghsLhgJieeyN+4gBKCbgvSoqu7Iq0VyiETfCAAsMb5dHWHKxrSme/D4hwgpEFQqqSA+E6Z8VMCJm
gK5P9evpymvPsytdBDILseUAnhb9txtqEUWOFrUDX0QbYxcQJWNo9f3qoWPCH7RGKXxsdLYE0L6T
Exj23molNKWacYUahGlKQLOAFEfQ9Aj62OWJCBXj0layBfsEE1IQ3aeuxB0VimIzXL9+iap9OcIT
uVrAjmYTTTAmrgyCfp+OQ9hGXSN9p6WQiKIlRlIgSwan4yIdIyyJw/xif0vqMDyrUsnSsO1IIZKS
RyJ4Z2pOzyNe21KZq4oNCIHdd/wpSlhJbjcxORJo9MBhZSXbhu5D6U3T3Yj2QgxPYBrwqIURYLnw
lFdqiVIZnpcl0fWQSecpxbfn2pHnXVDOnM6kWycu+vlrrHCZrK/fOToqnOEskPUmLENWK/lPIzTc
Hhxp2x09VJhY9U5uog15/JnkTvk6go5Cl+LlFYLAU/zCoNnNeGU/pVibxU1TuswSAB+SAwkPZCd2
wPGqw/EkHo6Fl3kHVASv1PnUKBDA/E5jukfOgkGU4jI3iQLHiWt55Eyp5oM05+oKFk0FtfRCkA2c
l6PQK8fSJCPcn47JvdkYjonxBD23kt0TX9zPVVKVvg1AJky/8mff02L/sHQigNFsmVqw8AP5BhEJ
IQx8gUDJlDMJH1dkTgxn/mC5gXLIu3UlWrA7bJtYbhixEP0c+0PRdiBEOEksNn8HZtmenaud1CV2
rw4lUz1faTT5u9ZzTbSPSpFnr/R+IdfBXKUQgwtY8VTuP34llIuAdpASIsXJMtSy3UL0cGbmE4Z9
4yFTV5+HZayA24JkgbZDlByvyjKAmuoOHTK7iQburYwHKg0IjZ7S7e314400k8KfRiEurtNs9+qd
Y3kuaT0W3Z7X5z8C48yE2H58zWuQN1emC5pwkiF1VuUChba1I8MWFPe+RZBMjwIF+dvttEYpUQhi
027UYyKTsLGngEPOwqq8Ld3U9HYGvtG+Jo/5z7VF5pq5aWZpVTnIoeRxB8QBDiHoqd23X/f4VqQe
649yOCSW333gKpF92zDNEiaXMRVfIIDaMuOSpk3FSsM7wAYFwVrgNCugIYFKad1RnLac9nk3VOPq
IpMqF0afXJsM91Ir/sSwRkGfGpi82qsFHEEAJRvu7TOlWKc+8lQhEz35wS0/wHvgTBLs/Jo/v+ZD
/YLj+3wSrzNSy8tvgHQU5Nd419NQQyK/ofHqnFMrS/cVActrsXC3/HNVC14ltZdoRifobpvU4MvK
k3Kx/vOK8aKpzNCxBqw1/8xRgswnzqRoZSAenLWFzD7uyiI0RpXv9lCFZ1xdoCHNv4Vls0fjsZSs
J6igNB2XLnaTuyAYg+y2ecPLjbDXgIxBqgL2EsFelzM+NYeACEjuhYiEq7ETljGI7TobinSw4slf
/XO5l9vxEOOQadBhlIGjVkG5RxE9LMxQouWdtE5+q/p6L0RzuP7vwBcgXICWzRUYUswKiHN9W/y9
8IHiyiFDSOVCOoCeR33IPuX72AjI/RM8qL7QEwoOTNdjcMxapx5AIVlvpcp/fBPRP6GQOkzFBqxN
+1UDxaSFqhVjCSEveVohzA4vt5wDYmKcHllH/MvWckKEKIaZNaWzM7YFEl+YjNatKXoJV84GXPYs
MXw4ts8YTtM15EwlCb/a8iTfQUpKlbpsQ5WEmpR9X0qeGPZnmF58FN/5E2tFPp7a5iunAXBzfFtx
HxCEUbwBL6zHnzwri4kuvIUctZyZ7dWnQ47OSDfVgLRJCXqRESSUnYLDilkMUjlT2w6dWpzrIgR1
PKHddos/Y3Uoul8YoVnNmkNwdYTOkUYkZbmnJTJH6mmmf/r3fIXgHX9Bw+KiaDMkUU2RAhyRhrl9
MujoQqfTdx5PT96qlj+pcbuYtYKFEnP5Ie10YC0g2/aDkSI0R99aXMZdQoPcC9xfpfzxU8CWmYsd
2sc+qCD40ln3sry+3/WfK7I8uTCyxxUOBl++tgoHOZtAyfNFvfNI/CV7wOVmVLt1z6aodjIcbbtu
rBTbm3rMu3zMTa3XyxAIEMKqVTqjRcZKBFc0i/3w52iLjV3S3ZpKxQ+/wwo3yby+z8PFA+WKrYCm
LEN38H+7QOwR+ed1EgvxpaGVNGQrLb5wWo56IN92WgIQiXhdMm6MyluKwBT/rSk/O1vI9B966U0n
oocW4OFg6CdpYAlWhAHoNA1U8XvSsyjm/vYzNqKNtD95fHH2/LkhEfp/IQAIUHImpn35OjeYaAaH
4RxWue+Zlj/f6l/QZwu7D7s61GcFWW3tgPxpvZybybS8JTfdJyMnKd2x3GvdAclt6auJKzr2ogNF
ubHoUijAGnxfDwH/5DwE24tyyWfTk86CqnA7SdfGXHCNhbopuRCJw3wHORKioAdnMfSBTe+ril0B
676N8bHHErSq0d7g7xIDOiw1L2m0DeG9aQ4DX4xM0qtVvjkpcEeSBaI0q2tNP8IL0VoTby8r4T9t
vsFl5qPeS88hnKB7Dpx9NxIFawquX8sLg5NqrOfsHfwD8UI+8oOGP3aA7+L8O7pvlmin9LWflh3/
G7IjWh5uUcWDDhvrZUIXjQqXH5JewZW3nDajttMWR3ztYY7+io+B3VvcYf/TKnVJ+tUY9v3Nz1Vg
j/wBrLIWJ+ii7rqwlNiG7jypPqTFgA5dOJlgspaafmluEnOqBWRup44gxI9NBHsd64QSPpPmkRdX
rEU4lazQGbtTFOQSZhgTeiELzqRqbQgHe4xYl8tqLHpzRV+nT29GBJmjtTRwhw7VJLrpVWkPdYjQ
qGdxGuiv+6A2pPktak10sb1FZgbWRYvPjuOHa/3oV06bcvWm+Yy2xprGuu6RvKF/3PCZGyxsSZUS
W5JiuOhcJJHn0hz4gHilqmaLX3b2hq0XQk5eNDUo242D4jEXW1Etf51y0XwftJTqLaIDZJhhDH+N
lus/W8+++vmEzFYCMOVrzKrb9r+O0zBHLIRLprTMQOjvGZ5I7mwjr4sdY2X8jCgy8A1NAFnXjSNf
h4+2QovLsBDmyFX4J8b2/DS+BYHg/d4sq7FVgP02Xyx6TTp81tvvw5cZg4qg70BVL18gDbySIKyT
DgqpRzKjdCGXxwSSj+mUTXwZ97vJyMEvtMHJbR6JACbFxba6mscVhM6B5oHIfzz6tXpNMqZoPXs2
7dI88/8XPJH2NvJg6q5mSb9o6FD8qf4JPSPZbqY72njMdO85yk6wFzDiOFpirD1cxi/5a8Nhvo7X
YZatbEF+qi3jRNMu+VZ0sGwvGk+JRONS4ul/BfVbgt+8nf/qoqVQhCyoWOnipCueJGBgWkOr5tbE
A7TXWpWz7Epze7k6sM+abk7q7oOtFb5PiTBKchxC/aI0ywVFiaMM+f1ADLVitKpE9fDcbKDZk7eb
rm+8mMRMnRDJBaxC2B2wvEYQnk8HEAokMtvhNXWE9T/Wy3wH2epZVPw9UY2e6rTsbYXbpyNI6rYf
r3xGNKaB8AkSLGrUN2jF8hey6XVDsaegDpuz5ci8nFoS9GNt/ylv4urDIYETaVNqD9esyMRWGTJ8
9gBsFAlYEYV+vLWiqDhwVNkZFBMWL4F//YsoTp7R/JFpnU5EBqPCxPxoJIK19QhYlDFvVZtbB2sx
fUNHVWhj440nQobhTCwLwnHS2LjixGcYIlEaFmGjN3dhh55Z74X/Y2yiD/XzgR3QwZFDNfsy3jPu
zwCyAT5Dp0P+6FKueilyhI36/ZRflyBJrif9ZY3fAPPe3F0IxSWFnourBNCyfLh6WDFYCdTcOmVQ
0S9CtVz9ZapaRi8KpS/11GCk/8yQl3v7UptiFzf/fijqJy8PCbdn26sWtShD+GHmujyANiC7DHmX
yRE9iFe8xq3cJTQyPDZPLd2Vq7bKdfxCHZTn0xHnd1xyWOvvH/bg8oQ6TfgNi8Vad/dpoDfAnhEy
jR1YFk8r302eImnQpcDjontbawwZa41eZsRyoT6Sxmwm6LIkjgf/LkEEck/FL57pWbBWM7k1q53L
9RQV/sn83yZ5QpUjDUXOvJ02Ob7OpBQzvmReaKblDSg/QOFgg5oOtlFihO0/C4BPNTKWD/lJx6Rj
RZ/yTAdqt+39V93wMyWJhg+plxio1T10RHgINUirdxqRbBnYstbFYGlX0VcEwCJgVj+nrNDXnhW7
kk1ur3OxYbHfAmDQ+Fm+LJkcWZZEdVmdXpd55ZoryK4tfs0jw0UZcfuSEhnOMgiXTNbHqhu+lnJ6
74zpteaggiLHb0LwNZf91U+r+Cz8nxBMtCeHdXX8za3nKLvuE3Cz+ba2Rxl4mSXcg5w7SxCkmgRg
sQ0PT6Wf6FlvycXQ1U3GT8YEGRlEL/adwE/gj+CYXLdewmeLxr50ick2FPexrzELgzsfh4AszasC
rS1hH0WAhFj24QUrWJ7wICl6FvVOJwTKCLuILLRyd0V7AUqvXdwF5OUnC1VIlFD6ZsejcalJvaMS
Qvu0wJqpoDpukfCJ1r/cSXfs2UgfRA8EGTJ3LCHDdYKzzUYvxqUDMghreQzzYbjhHF6/Rb82THkA
U7LDo/YL/7AW0zJw5RX1BHaGMFevT8ut9xZyB1hIEjIvbrmVifg98Rp1ZIy5YlVCXdKZUrYPb6u/
3QyxZrIBRTulPwEs701cj/TBXk4siAr7UpDUA5XenOK/GEMSfqu7s3wmOkn7BTWsAL8SbXxkc2RL
pY3iwJ3+PxRYpBCPdzWqppH9c9WwRZo9NoMkTgZYQ2YdGUKRm7RZFELHIgCHwv00YvWeHI17K638
wO24lPNgzjM6jrv7oUrbMzABLjG/cLqcxsxrmYUR8Gs/uLkm+sgJjF+Wk2bAxOFjvfRrAJPSra3g
GN72vdLHafQPQh8uNLKtFvYjbG7XwMUYQT2yNgdA2OINy13idAaLYz4DU1JhTq2ZzcrBkMlF3B+t
DwbkEAFBhbyh4qu+p+1z3gRXqtKaSWxploRQPuceD56GTZgBm9G+EL50SRYzKcx0nnTMGJEW3o2n
+/1x4NNpgSOse6Xvk5MeXZX8UcUvgP2Xn+MYWL6r1Ejigf9C7JqK9KqRd2dEb0FChTbTuuTVTdu8
IX6Gdit/DfkByM3QyBpi4lxKd1VUoYd0jviUEhFaeJSgIsPXjBUAHNOycHnRsxnTXXMj3Hw8kwkQ
Z80gYx0X8CszWzHqjhp1oNl/IZIqrzMwYuHDvbBftJ/h25pfq2RfczzmKZug4DZEA8iYTMII+hSV
nFzZabXwMkhzq/WeL3utQVVy+ZHeJYvj19dzU/MmQ2pS18I82eRytsl6zCQzyrkM0CkjAcmkrgWP
jPgNyz7adX0sVWylBMIvF7xJ95EaWJxRl1eIOvL9oL4QCIozCm2wpJPNkeO3j0/m4pOdKs4ibTQy
LwCSAdXCUujEJNGNW3mTcsTpNiZwqwB5WF4JG15izX8tlN5Zm5fTyoVC5eUUE1drcTeQ8O0lcS09
xCcQjaEk3Qf032ShV+FZ2HAAQX2xUMrWbDZYjLp6KMODQkBGCq8KmATIkIfxovWNF8WmLDneSojy
OHeUKhxrSsNLkR/yhRM1qOW6tuBE9GvJHno8qrYN9BlHZJXd+A8Z08Xde0oT5okNDKLLiIyt612g
lTCqoHogzuNZLehkyODwZU1SEHK4X/gmSnZgqsy/pa/Z1JzATFzI/Pi3EODgl6/vqXyubHSkX1lv
xtWOh0A2QQvdqFTPR18s0ui2ctiJ69S9xIfFWW/ttLOfMOuevVAy1CSTxp2hkRFrQEJe5oq7Gq7v
gFqgRVL64U8uE/W15Tt1vBU4sl/RKwFzqnasUlEBJndpx0ndAnCTnvafi/8TwOyIhNzvSRyrMb6T
dk5lP/tNjGxbcszuzUcKwDxHFNqgZkEZ/JqOt6FAdTq1Tt+0Hxl0TosCK5kMOJs9KVCqG4jW7kri
a7i22Aoi8vx4aaoa/Z3Gb8YVaxRDlikpGpZbXYqoTmJIGrfeJtV4mYdeZG2bgAQhcdkyuIthac3U
di4b+teGyFPp5x1DJaQj7noghtaMmjFThFFqbfMKjYSnWrG5PJ1J6SQSyOft6vZpZelnSpz+666f
SJWDTQY/CSSw90mtw78+cJ6vFwuawMgKlPbW7p2SRm3SzEOTQPihMGS3xMSmMqZfucCg2uQ7blBh
tWf1oirQjfTYuFgSRQkea2pAIo+YRa2ZAviMUlCYlV9XNmcarpp8mabXeIbJzaySB2IltsfJZEYi
QaRmPhd2U9YjX7EI/JLxGfi/2DTiXKm72nvVZACGCfMvULvCfOh0k4SzHJswICaGmzMF4YCNr/2I
TaD6AG9mKR5WZBV19irBjwgzbs3GPP3EwIycsj2/LpMgZ5X7BHxZoPgD4RE44sxqgGig0HgOJrWN
z8CwrmWieJ2oWuSVvwRsolCgh0D/H01HFuccbggpBHV4qOyAImoMvICa6MEHqh1ip4+OnLP3qdn8
4POwnMAPhbhHq/1zNiqayWSomGGna7T1eWY29XRK9QDvfZbDk7EL5m5c0cjJpGHGUISc3o+9rLiD
ExmudltOYbDblJYE8g+Cu+X9yTQiPcHA+AyS195eehGJyJlZQUJ537VqeaMHQP9OgenFT0+/AJzC
nhNwAbRa9J3kqU8Iq60yszTkEuyfM1+EM/Q7s0axlt0CgTmSTr+DdQQdwsCN48egWk6rV3xkC87F
tArvhL7fyb7pRGvsHgWz0MQh924Re0hu5rrXRKXv1P+GkNW1qXVntNTKFatYj/SQ99WhgoozJWIW
Z/WrcaXwnXEgIA/t7pzgBq3JNyRNMgMkS0yJlc/Xu9fhwOSGL/RE43tw6DhnmYNQHJF1ujyrfSUv
j5+y7XxnmYV/0cCZReHLs5oO7Oym2fT2JFKW5gOe9BFBojUDAKFP+b90+cxgxbVsX0Fjkqw4y43F
vO+xqEf5OvRWa5whJkSw3cVndEVH7jgnDA+JHdwPe3g4MBTvFzVbjdRodT7pLY4BHRNkZftiu8fm
4CA75BI8V0L9LyRTYr5GLnGuQNLH91cklvK/mz4EbtBe9FKfmxHUHWV0qh3o+h4N2GUFaYrQoTW9
kiwuQ9B7Wboc4sgB4UA1M7bsuwcRgNO3Udyk/tJ1XtAv5PNgjDVBiNCxpY9cS/XY6tC2cmin0UJj
kVY+e/h5pOhrHUh6bYr+naKG8NW1cUyQEGPRe1XEF09WNE2mpsPZaw/x0lXFkZEVsAwO52hKgOqI
8eq06YSiEN+B1gRAVTGKr/dh03af3d4Epx1oU5SoxDyvSu5IU6TGaEbxnbFtiSoqK9svOVl+oIdx
h33p3jFnk9VeI2ZN7zlt8oc+aSJgO7Kf+AZazdH2cICLOcvv5vm/QEPTtoprM2dL2BueZJ0XOqNP
rHdjYDiMjYhQc+agFTU2gb0lV6B4exeyHXpzj2tHoHA3mKYAGlPHSE58bTQuLYzwabeE7cQfk8sX
xQbiixGMzX7ru5RyKXW+xMnHsDk+ZI0MUhfTLu78PRK4T2WN8MkU3XhkWYHyw2Y6IbFnGa8VwCWq
F0UakFqOlZqQmhFZnvr+gKVn7z94MhaB3qW2rSiwsrdDgS5aGmuoAvtE2gd4O4n4AHnW0oEmLhy0
H4q5fCw0alb7OdC7/2KPkSC2b6IBLN7i2LqpeWiRk47h9fV4m7/iQvWZCn5kcV6ZGkuE6aFPOcXm
Ny/ULEG87Rla6KKEbLu6QVW9Op9QlaYqbx63FGdLBFIdeZ7IOfIRW42fA81EG4IVC96Y8iyVE6J6
gfCuHHjOpb3427w7vLZvfve3fWIHQB97d6dvDJYZ9TYFrbJe2BBMwLPRW6UZP1ZdYjjkBdQReVI9
SpKjYm6yQr9xf8EMCLbqW8YiHjZvoBACXY1QweRhwMIBH5/QnPbaKJNIUz4o2DqCaU+DL34H23dw
Q8mbacI3v8AW9gZBxo6f74Hns6wgXwXXHyU/D6AfkY8gbps4+P1qn3a8c/oiDDVEWwn4YIzBxtHv
cnCh+QqgO4bUsoJ99QKy4dElcDTdhM1ITaXkcvnUGvmOoZNVU8yXy6z2YNcha65TkLJnDmE34mMq
6VZ55GHum55tz9Vc1zbjdPronZnT/CvSPjN5pcEaQgQhe48DtzX6LY21cmk24hh+xKeP33kbaKbf
up/d6dIjPeDm+jORmWdMRwpEpwE7SdzE099lSQhVeyhQzbicHIt+Ya/KIynD1m9FM5lvkZvoelx0
J3wJxVAFHjzsiOvMKPVaia6atKEvFFZ9BfxEH69JwBQhP1zIc8TWm2PHduk/CrvIA5nlSXdT4tml
0FE+7ews+MFGwoedpIjSHwND5zRQnhtnc1c0We3rR2B/FXLdRSgldAW6FafkEsVWl1r36GO89UjI
p0g8faKxcPILtZfsJsFvepOUy2qsm157IgkvZkvZU0XmlSUgDbNGPKgBHQzkE+P4hkV8O7eOWTOb
XBamNUg5u4U/0RTKtwXhePnpC6KNsH3bTiJ7igiBLhGKf/X3rhBIlAuwnpoldWCqGe15fUhtNoWk
FKGL20H4u2BGBd+XTjp4z/8sxXd4s/SwGmTuFTcUoQopODhp4a+5XuBR5LBv7A4zhEW+ARjeYzqt
2vg48B+LZ6vKlNkoc2re1yNoGYg26FIc+/EbSYbTUTAC9+kkKa7RzkJnmtcUHPYdkY9CKMLiKv5X
6dby4NGY9riGqCoiC2NM4yuqlWrHtt7Bi7V3juB9wu/9f/pv/380/53+s5UZwZShBys6wrA8MDhi
DtgKuzRcT9Y7JI6zPEBjdJX+HLIR12nZHqgy+oqu+IX0k3O1WPDX7cs2s/i2Ft3wnzkwZdGmBNLF
bNXlPmV6Ru9fdK3h0/n/8jv9w9ZJauVC6Tm1py2HjXgXc8BcvWHows32//M5aBCZ8lnyGrvM0PU0
vl1h9B+lehMdVt5a7lniNFkdOPDTGwOGb3fusQBND3zpMRQ4vTxeBeDGunBBCG6G9yeHDaf8Ios8
l31wPpCY5q3AUeOS2Tz10Yv9w2zIhnqhkyPSisW6ucorIffpHhU0JJZEKg/HiEmd642wFVCygn0w
iuM9hSPwyDEVJSJ5mna0Ehmt4Da0lh8Xq8j+WWGJieFahLZ8ARVXUgKI3oHkmWTA+PDt3u4yTgDS
T4TX1S2Nzjtk9wVsyN/1sNmiGIitCvye1QPzN4dPr2pf5o5v41CNa2OYqpxXRAOAQ1533FcKEGLG
YP2O18IBcaYn0eeWN+keij1mSvHI+OPgP52R/NVAErc5t1Mxjj4s+ny9wIyWAM2kC6u+B7S2nwJx
5i/0itpYuKBQK/AGXzcPQEGRnyeNBRHIU5jjI2aU1ItPUadu4EMaXvgitWKl2eBcE6d78Tt3JyTs
S5BxNryE5DKB3fT+eB4y+ou2C09Ig6e4/DDHKn/T40+HtZvVdnz9E4Nf/QiyOvRpWQKkw16oduDm
Xrbq0AP9z0wYgOZLsPzA9V1fxm87vw+mzKBmSmJ4oLvNID+KbSE8M6L7jzaoS31K5QX3mEzQt+i8
gl5qRls8umPQbXc1N9lHGMH+X227khpUH7VSTBYx/CxHyxf5pw+Cdi11pHQuOv3NGx6upvunGPhD
ajPLv+GFlE4ZTn7r8FxM5ljS/D1VueMsMY5+0xDQW4qiw8m/jSgWY806bNDnqn3wqR168M1ukOf0
fIVuNf3uAwNHk65iCGq0WOupvwsy9HgMjFtSqK0GbTohSd+mxnE2rEOaDSNVHBTXGABj6V/OU3aW
HxFSOB3YrMuzQ2R4uTXJOfeHQuP5Bv2K3QGE7IXNOdelndh92P04F+TufB+BS/+EEHlnmsjdKdfB
oRobIIKAJaFJiq2r4yGDvCHixIaNMBh7G+AxXdxBWlKkH9a9iJin1eVWG/RmlxY01krLTEc7juWw
oi+Ba+RXuCwnMz0b1FoLjcfZtMDNpPt0lzxWIls6aOlTlTc0nUzdMqZJKnq4P06MpevD1rH9lgSY
X+y+DwBJg9krJJtfZYXtnfEvK0TB/Rmw/dXZhG3ZduXQeGapkHaWR5wn+ibGSUY6nbjBs0Y0/5s5
RWQzbuGBjbA57tjz7deN8RlrA4xcm629DpFsBpnDRas4eUsaXGBLggsDdTJ1Pc+p9hoWm70QGCl8
N7AyeWHVhhUUc9vXe7T3v23wvQfRITHFGrPLKLxIJBdmp4Ay731YLRkqSTbxKs0M+uNBUmL65qke
CMItv96lzXqe8Eyn2Vj7Y0XFpooQklaTnDaUYlcoqz3IIHlp/1u8rCS72X1d011z9b2BsO9yZvma
NwP4L844hCKUE7v2aES4FpI8uP1kwPdbqiyN3yo+XYleK8ZaYMNqjSycTP2FHdm8YFVzUHuIfNX8
C52Ch39Dpce2GHp1qoref6ljiRybcZSVoQA6/s1Hg9qzWvyfHnrFZsaQNie0qmGby5A1xUWS9oB/
GP+7fwFf565hiiL0FSogdLCfKPI6T1Zl/AMzYnGRFXVa0YLvp5aBq16LEcZTaLFdu4Gyp7747fCQ
dviaJZhNqjz6jcLaIk+1H9d307GTiy5gjaR0bfdlOsp/6875fQBOgBzoC+LcWWa1ZY1hiED/+D1i
FF+JkbnU7R6LnUFTSCput3a32RveMLM8GX2kbwZU2quohmgX85tPh2r4LTZYLYwcCXtQ+pL9AjAG
Su2TGaoKPRRU+GX6z/jIVXpzinQnQZgMbtdMuWDNxySVPedSN4vHYiln8NFBjnn9tkGbE1T0hoJR
OYJulFPqj1ge23KpzX9I2bTyk+QppWA+l72Gft+G8n5v3zCOYi9AeBWgUbT+7n8AEMDqaDUW0M2L
nDPWrFK9iOunCxrbVFqKmrXd0eE2kjP2k13PHaC7EarrAZlUqpuxikvsskdfsJmAc9ubhADNDuDz
bxfabo8YsMrraiJM5rKv6DZ6LWt7CWIpruBrev8YPLS+9Uw+/rjd9f+icomSH94+5bc+GjMrpyEe
R4Kc40fnSFQqHpUnit9I+5c7dFTv5BN7KMAF8JUyryQWNWs18GfAoJQ1zwYZcp4D31v8N6Bm1lsR
Z78XHqReFi6KNrwZo6JkzSuw+70xEk3TcKDlKQbUHog4+loFCcDvH2FCCW7dY5bMbNwCd/l3t1jo
CGk+9SUlUj8a4blCKwHVP6xaKNth+fAie7VXdTkd7ronAQKQtZJOW5r04hHnT9KVhf06Melmo9I5
1/9Id/gegS6zKWnRojSdz4BDXmLN4oXQ5U/tasNvitCjtr0pvxwMMoKqGQywBYCb1K23OGd/J6Z/
TMXD2y72nXQ2F8twWo9Zm+UV0urhZts/BB0VqQUc9dtKwJsf7/2mjLHBq7vvpHH9Yrt00JyeGrGQ
9JOMEb0pzcwYSsPYgfdZBE3odkMX+6LVF0GLrWxk1aBt74soU4dUUjzEmG9ctMQQ8WzUy/azmxC4
PcL7tZ/V3YsXCpcjFDHLD5v9Do1TvBh+U0gqkzzy7kgiP7NR2Qs0l6ejBmpv+DkVjx1TFz71E5xt
/Gy0pGrqfMM40nbjwmvr8mfRoTdkAJzc4LZ8ZrtQ5gRz8yzctiNIQIyxQsHGWWLd6C5XzkDZTwaZ
Dn7xLRsc/n5mLbp/jzuB+1Z1McTH+OjJNsZC0Sk5QWisuBuAsLGN+LZi9KlMRkBE74b/cyTaRpTU
89mswyZ9pVca5JB0LTsT195EexhyCOGoqrkDstyn5TbwTIMRrm4UqqDb4KnySgcpYOU3ZWsxLyFX
40dpVnMyfJqlJCEnNCMCtGbovvXwo5SAlPs89/pMKpZ0cthVcFYdcvLokf1VssZbLzyZszYXpAdu
jVr1iCO47OTZC/acTXYISqzzIUFBe4WrpkCSGZ02kNzibH0BEuAh9UxNrLlblax5Vh6kQgBUe8cM
s+wB1/KsC0mBUAszMtBLKBmJ13pNftSaBffmHtQ+EAoqztzBePV3uu0AyhFvMdu0bD1PgSw1enIy
jHbuCIkGmnbIh9DozlsrgmR+0JuvdgfwoDf1+m6YfuBFxRmyWt/me8O9vsxB3Ex3CfA/ZlvEjEMC
26xizYm+kpAvEQvlM6kkSJrzN7h2rFQKWmsog6kkkFz5QMkWNCPg19h86LPnFRt8qi0ORF9MG+oM
xGo7k9L/QIARlbMjXecELw0ePOAhFwb4XVgh+C3vRERFXRfgJmPddSLWlRLaSNEPSZ/v8bUkbuBD
JneOBKE1G/83sAcKOIAExOg3isu5bRqi8Nx17FsEP+DdkoyPRa2N9atQ3omVsF4JyrmUxFpI3bxN
3u7cJYwiSWqRJhSaVkVQjREcHDJ53ZisXgWVCf5XSxbNv23SZvEJ8IOZei3N0PSbpwzgITdavOMD
Y+Qq6m7vc+U26GlqffFcmqOisUxKsHEieZzfXF4WCzmUZBwgGDETzydXwNBBL9qSFyYMor2+H+hu
fOQle6azO9JrgKjq0HDl8k3bdGKvt0+XbWEvfD3007ZXEI7+HJ1+bE8MTUVkYhtwLXvWub0ITfX3
xclsFMcoQOPCI6vvhrguwMBH/iHUGKoKOrmQS++iPbuZ0/yBim7ey2R7cwXbEd8pkoyN+ZP85Vxm
pkF/RcYocAZMICNibs9RsffSinYXiyRYugJ+bDhqS0hGhfVB0orMtNwpfUumHmvy55eaoWTTzcH8
zC+2Ysf9tRIWVmcyGSO7u4EEjDD3rgNdv/0S9Q6wiO+RWnyi1SC3Gfq8sUj7G8tKRdFixL3MADMh
E8JZGNZ3l0XKfbF6H0XV5CsnQthTQBpMJdwcDCUCtIW58as0KeKY6vEOj3T9Wse4Ir7EsnSPHsI4
D+pzscls5EHAUepgEH8QSQshlubobxnAAzPvZ2uMLol5qYN1Yaz+S/hM2mOfCQikrBmoUlNBkxJE
eK65qeyo2cS6fwHL3Yzxpv0GmttoeQP9gJa7OjY2w80Eeb+SGWnSdvgninTtVzzaAMQxYnl4J5Xd
GELGzXofJBUNt3wRSqFJeWXwBEefs5QCsI7nb3c4WFWJ59Pk9tdDCsTwOcQDE5NNUIWyzy7EnBHi
I/K2evfzbkkI0bLebWvaOYly+RVQaxi5I8BGeDSW59s9zklN4fYI740PHado+YwzcGBj5TY9cozY
sIZkJ0q6sM3KtsxqEr8nxlFT0xdZ7BCZcqV3dgSbq31D0QZbnSyQOOTvjTaXxmuaJpNUBCCxOg95
Z2Y6wj5c90IxROk/BTki14gQcqtciTqORdkJBdiRmAY5xwmxX3NA4gNpcBrlDRTbhAjmX789TbOQ
g6yUvLfqv/6Fu8e0t4GrYyPoFrtatXJWGJSfBkX84UJA0LxhVdbaq5YzmEvpFgLI1BADZF1+I98S
C8V5MwtZH/MYLsvA57d8Wvwn1S/HHSor2r2YlqJHZFkxN8W9dV9QiELVyOaZGleT9AAa7fFcZyQ8
K0ZtDUytn1AxBD745WGmh+FO7Et3/7RRMrFRmErViliAhdOwogyh/RiIn2BuS6D+eBnY96rgFQLL
RPNensSWnLWDPLYrQnOrcYKBIIDK7wHZwX3yl91W9J6uy40vWA3veqc+qH9S9tyxUnS/hU9Jcj6J
JGDZXMMwm8N/qpVWZO+Z23FI9DlaBIq8njdMntKQAq0aWyANjbM6GWxUc3bzeF2U8qjih9L269qB
4fsYHueAgJkMFhZEryJp4JTQDGczqA/M/gInkRGF4jESCkusauCXBsO1jx0uoTlaHs5epihzisBf
0yGonDWEQQq41+VR4rBw/EPI4xu3cI4fmPKUnEG1opaUzTrynLcBJrPQbeS4xh2Y8UTiMa4AdzbB
y0EuQy9CqXUlC3Lb8jEBDcToOaBQsSxd0H83REsJIOL5a552R4/fLNB29VY+YG0aRdxUr8uWbkZ4
+LeLhpLpcv54pU/3tXwO604PiFCZShpW3V8Izd9eIuE9LigZlFKA+yboFykQGEEkF/hDvtRtZWgD
J/Q0bJNSdJGCEntNqFIScHxyQ99Ao29TdheRJwC00BRMiPYIp6l/XgmsPJEapEpUTMzGLzLc50A5
2J4+6i8E50z1DUtlswVABUOJ54xJIhlq70eYp7w8ezfDxs6f9hTs9P1jt3kdF22mtQCp44OYbyE+
Y5C5RAkeNfRb4EGxvedkg6X3XEUQOjlBsLXGY8e8a/ywIIhXJRxYJh8YjW+fnQeuwcIrMapDp5Qz
LXn0eCt39gFmbhli/arAXrxsfSgO9CKXSRLQ2Pa/5E00fLFBtMm9w0NtkkJ1lvwWaWgOo+AIzkPB
akBWsWR2vDrUwzjGkSWnf01lNTPfqRnCJGKAbFV1SL3Q2XEtM5ihAv/4Hbso3CwV3tMeERI1R6cu
FVSVExDB0S81Y+qV+wCxHFshoW6WXx7dG7g8D4aoAs1+RBD3GHwRElLKC6GW4Y5IezO5/0d5ajNv
gS628wJJ0QDedpHGTsIrt5W7GZHJcBS7aQVrtslyLsRL3MudcH4eegSJXcGmfJ8zW8zeg8u38qUF
YFrIchHqbYfQw+wXIZZ6XO9MtW0S3NRZxwjaZg85hdTLGrMLmYJXJFEGK/6I1MAEukdm7r2/cCp+
OXWZ0FR6SmG9gyGVEwrp8809Ec2GlHENRpjXAK9ZNKWj5bgZE3s04t6JAI7xE7TsAkBWCUiskWHq
Q6CDzJAV7gzSOEOSc5gmECgG/rkfvhNHvwkU+gi5Z9Ffni8tt09SdusdNac1O6qxAh5xaj0L+5QS
WXilNkAgFDjOJfF3crpQnqMS5f8B4A34CRC5Ih/iXyCo94NLyOPm6bPS0LWQXM3NSY74xz5GE+WU
FRdR7kepuy7LafuAEbrw8lgm/O7Sn6iUY24q33Q1Z9Rk+RoIMUAOieBWkNVzJsvubn9bye766FLV
qloW7fyNkuA5CGaG3IU3up0hqd4aCPMlkzV/Y2V3Wsr1+575/6Ad/f1pcKooqV1mN3go9WV3KcJK
wXW4Ei5a+BEG3CUR99LDbyPnT/eW5lZviXwRJV81ww8ucN6dCwluqBk7G6Cmvk2EH3BmUX8gVlOI
bPS2Y53SXnwp6uUVk+safk55TLWLLOPCr6eyjWGWcL6i5TEcBh/VeAHgAUii6s9c/hV0WSiy07o/
HkfvtwDYTGHlP3CYqKRKWEZgDggqyewRoGS3TZwIxgllIeatYq4BI9JxBS2los9bvoIlIp2VHDQP
uWyWOjZRAomx/+tcN6zyxPfp7SrOBjFfD9xXXzs7gRMo0stIjE+N5mLzmiQjVAWstGz9gXNfzqHo
8kQb9M/ivLcaxKvsDAvO6KOcZJoQHvmfEtvQsACN+Tiz1h+8fkn32fsV15VUbFClo+79pLYWwFvH
fFZ3aB5WFOlT3AOg+4IOjZBttQL2FE1JA+ynchudGDticcDD/u9JBbGYcsz8/m27MtIDzXMj08N4
ySfgIoNyO2NLJbolLVG77v1Ely+0P9rSr/lGPiuBGXhLZUKr2RAMToGB44BVLwZO/MnWd9ya1+Pm
bYv6c7QBvx8u7QikKtwdCobqSfHWaOmwMU7FF22QFSZogLOMTJTDmTJVMTLEFRbupG12c/qKognl
xsNE+d3W+v990NZM24tb8FXajU9aBqjouAF3UJ87BcA0yRNYq5NqjfncFxEQVyqDYRi37tsggSko
uQSWLQkNE/g7oiku3KAL8A3DkZfD5Xn6MqR7nWXeIiFh/TZZ77RZuWrn2ixAUgF0izFE80u3MHuG
da2ViEcboCmDLax7iFyb+BUIjaGYFAbqO7Z8ITSyIIMxO8lvpiXAXy2qJxKBDb6VsGzEqGwLiKoW
bp0LrwvV5xI71IKkLUpAYYGOwppLjl5YejGQS8XCRXiPN5rf09A1IRcZAlJsdEW3j/yxsbybij16
mf0Ws1KPv4ZBpgP7A1gu8307XeVCTo+HfdJdXzQPx61EQwIOyjkpXgEU9CHmXEg0b4Lo41Wf3zEK
altxXE13oly6ltR65SRQv5UN/jMwlumjP+vK20DiG0uty4QQBhWQkTS272s/mJZ0mbItbnD+dXFN
mLNcK+Ls1g4H3pkh2si5lfEoH90i1hKaTANEHEEput5Dz78xBt3KZcBKEhTopM3O8MLIjxzQj7+y
kV3XCOjaWvqVHQP6JVLyALuhvTLvVXfmR40SqMX6WERdCZgqr6QpoBLOtUiyaoOPblt12MCXsNGT
k4oK4sAE+wyGwLLkiix0HCmbPGebFl2DKGlMv/Bh0rL3HRCTTrGQ9Ib4o62imZ6tj3heQ7qxIt9j
GddCmVF5ITC6KVsOEvg4p7gJEv4I2ZVODwW0Gd/r3EfORp9eLgc43Vb0OyFg3PskbB/YegQk1YPg
fR0gBF/1rlTCX9EMTFOvWAilkqYUXtTx3VWzD90p3HFTKlkLrfOnAfkIy+rEDn6QojKc3cu/oK5C
wLn0dQaW/TaaBuLX4wskFTPgnRHala+44j89Vj3SmjB23r4B18yLKyXibDUsYWD6GTR2pcun81H2
tWqZ0Sehtk7orAmBP2Tn5EtJfY/YtmTEYALwh4c2+0fkGYPv+uilVXuKZPQNZRXcbni2efmwzo2t
u4NtyVWL7NiDN53KswVSutNkBw47v+bW6vHiS1DyuE+x06f+8BiQv1SrjPEf+9/mQNtpPlT+LR/d
7fv4NqQLHOsI67FgvRqSrhxflVxzGy9yGKHJbdWFud7QDP/Nvh3rjwtQeNOLX+HLG6IWKW6BbuWK
/7mSEGVUwycHofL8H8OphH/7iIURPeJF0kgM10XkofnBXndZu/pkyNXMQEwv8xD4/W7NyTG2ePwq
6kI1SuuJ1sIj4Y5HqMvsik8xRGFB30L8MPhHkuBiCzLzWcG8UO7RL2uWDBPz7MzRmhDfTHM7S9hd
L+wJGfGjz0bUgehHSX0uJUkVxlPEtNh+UV2cqG4+nOJHZ3Q7aNJsQ+fafCsrqDY/1Mc5vKNV9tAN
Ptg6kgPQTZCzKEjy2mLptRsfPs7gPCtEPjUnEHA/vPIX8O5Y4y/nCfYpyUeiju6W9Vbm0IlrrAJ3
gyh7m3ibBxqr9NRQzzj6x5eSs0VDOCkkqaJYWmJGqNg7UAahZGon/2xOqXgscG0mM2w4npVoVCW1
t/ig8mtzTZGnt7TjmAj5g4ri6ciOhZrobtbmkoxgtfe95X9ffhXzevvhAlSnwbUMDazWfPpCjIAn
6aqjgWb5yDQfsB5sTwOBKJ3KIF4PT0xa8ljHgTSQ0sW2b9IEWKYqY9I6i4bwYtdrZgQz30hcyG9b
uYCriumqA8cuwfxTZP3BH5xIzdB+njK1maP8FSvT86pSFhxHppVzGfL+6TQRHs7NlIGW4PYR+uOt
MrvzkGwlRvRw6jUhdOcKDnsbZa8eejJEoPKLLV6jPQHKjrFkcOBVgOs5NCCZ8YxtHiGACAfXt8n0
nrqPlOLFOo9iumoi7DQTS1gkTYdfYhf8DZutnWTUIhhwoxbxmpUG8nRxtaEHAP0nCXA1dIaLEPOC
+6pTuvarXWq650Bp+tyyng05R6WGKPdMxmmIh/gsKRnH/CV6ADTs4lujb9E0ooNiZNTtm+HURtKp
2uhTIPLabzT7u0DDd8baR+tUa6D0yytO24K9aF2y/DK7nTC08aA1yYpPyNo46yOs3ek6kni6rzEd
V3hdn6abAlqbUngqPQLjuxUe+tHlHT54Y2Z83x3kWFnotGZku5Uoe1KFbKEilG7NSUNP5AODZbJK
ir6/VZtBgnB7GMBW3700FzhBRNKY6s1ucuwCDTHfU3VOUoL6/kRccQJ2bLaxoIIIQbeCeahoYuAE
B5Lb7uvSDgARS24r4UMlfWlUL9mm3/R9J/HCzR/3d20ZByWZ8pnKcWD2PP/VKuIAu0RlihiEhTRI
zrV1EqEw6RsO4Ik+3s043k5DM28InEyYkZ3TSiz535s3T9E4Vp91Y5s5F7JNjnwJMXmH0fOF3P0I
arn90+1nLacdnO2yQ4dx5JsNuS5wdk0SenhRASznXO7XhDCUUG6H5tHTm5d0E6Q665rrRZeiic5m
d3lOx8fkoZ2zQkI/qdHb0HfQt0Ofme+pIjsUsb30oZrLcAjbBVV7zdSTNI/5vuDDba2PioKkkPMK
X1QmizEJHEP8w2pipc/TgHBYbGFghjwYRrFnEzbfHVU1bFBFFSz5N8Ex+1edzqfFc/E6p10iMEeE
a8oCBd2pyj+5UB64/gjj/ZG1mxPXpzDsVwSV5FR1xzrgjSrArJWySoUlGo9263Oq4wURKglwvrMU
oXH6GS0y3jvbd/B7VHlXeE9jI81TYUGAKYHyNhBkwurc3YhTJ4+tzac9fBBSjWRVRhC51IqQXWav
hOlzpj0KeuVf1K3ZJJVe2wB0SUjCJ64gYCDNxqgwPf48GiQQIedCi502z25lAhQkV0dj8DrorWFm
k50C7pM6SnbUOligLEXl9wp3L4o+9uCcgnSymbl6r53AMh2ezn4/k9BxdiB2ZJ4fBtsChIzLuH/n
rsow7T1IHTMumahuxgoWr4ROO9+V4zOUO1lkuyGMbSWBD/W5JtPFpfK+wrVQObBMeU1tiA6EecBV
lk3xYfNnYLSIJtmaCcJxg8X2h6Tpl/5lcaxLJIoKrFF9VOjWcCpHNXPxJFObhYi61AeDWwUh28LW
JcsXhiaSiui/dNL1+kxKKujzalPNPsvIPpneH2lA0YG+3wyIkYIqiglpKQW69fKT3G7VsyCIdxXz
U6ftxSiMdiXiUSS+GbeuUOIYPd05ac3XZhZgYizY80q/SghGjueMUm4gvlNBKPZ4y12vAfcntYdM
dT+kckV1q5K1ArOVylmYZ2cvuYPGZpXFyjuRf9hs/cu4asE2aQyQExKz65NxcAdHGdnV3Zwi7e+1
UKCZDqBo+GvjTQ7hclepBRB0fJmc0D8aOejHcAGZhe2XtG2cJKPTKOUIefUFfstzEyq70Yh9XpxZ
MFohdA/oC1gL4gdGCnVsCfvp22gZ3yjUA4S8Yxld9G04gZAwig0aWUzSStiSfeMtsYYnq/vysgQA
nkigo5UFLR1U1lwtFA+Ab21QlA7QULtCl1kkSVPw2jONb0xknm3u4DVinNyLYCCvLH0vkngvHjw8
WDMSbSsGgeNu7RCsnHYlKRJXb7/ybfJc2pR0MEWPwQmgyKgZGZJuZIglJl+3sxKAeNpRx0puae4g
fjpE3nDnaou240AFey/GckFgRTpzhtrabrkjUIa/d+K+eXO6EFfGPTyATmx8pnGaII9b7hSt72Gv
ua+RQuZ02UbZlgHLGKaNNOnm661XgFMm6h32FShzfHiPBNP3TDjGTu9xiyI7w+/7wqBccTHX1H31
q4HRM2nq+rYDGsLGvbmHlkJxMj13AkKSis8t7hOvBTySlEuGViIx7Qu3oiiyjsLfHRGJiKCvNNNa
H/BaxON9gFQjNYXa72Dkvyne2FWZx9QzQX4V3vKEatZMmMgatHgvZDknEQByqWYxEjS1ZSpr6fDE
P9qJF1+j79THorMZCbLfdbe/l1JYGOza51X06gphNSuuxyt0bWTAQQGNt75FT034o0cmzJdThruO
S/eXb7y9DKZUFMIKUw8clQ6mLFoEeKXsfaXfLOHEzmEJFpdV4X8Kq4TTcoRLMa0Quw+IM5vAOcRh
03/cENijTVm3TFAzcsDONxOWoB+yp/W1sXq4JXWh+5o415Im/0mHxAqqGjRqN7otF+SfQbdYHlBw
pQgmZxR2I2fB8Do8NZsQdHxDgsxq1O3hdf6+2zk2yhtHXvQk37to0ViwUzJkUUgCkUayqgg9qOYd
dliWWwCMPYwCbLn72+FT25CoXM/wDrd8+aYlgW9rsU+3HEnv2E1nPtvk+EpYgAQOHVdJBR3E5KPe
hCch+TffO47JvbhPnPc/Ie/TbvcDZhu2narBcdbfS8vfKdtxqmA+s0QxJevrC1bDfFXgNwPE/KzZ
sXqzMjna9vfT16yOC2ZfgMKmwP8UW9TncCtj3VJdASFyZCyFEkmmZwxZwCUqOrvxuyqxslAjspqN
bk4Ld9arX/ncmo3QMppYLccM43PYf6cWOgVpwN6zmeHYpgGyHsBSypL4UJjEZnX18rsDl9yzVhQ6
O6Fvyu0pUTCeN2tiE1Ze72lLpqwEJEHCiG0S+vuTfHbq+g5cGie930UlQ0h/ejtARh0jEN1qTf5x
yT0Beb3xvp5qTbh6hNPhZHeOiW9EUe4ggdK4NptjlnECgr5sf5twdmuO5nECjsT5wO0wcTUAAqiU
gVzZ14mSGF8jxdOHGM3nOVhXRTJFwSooXq4LG2Q+baWIJxDkY6HPm1fGwPziXMhKmJKXXX0Ml4Yq
0Lpqt1MQZZbSA3+AWXhZeBEOVc99WVrEAARv1K2mYTvKuKflPRxKp+FPApZeOGJWsuUaaabdxl/y
jJ8Mr39OU3bgfCS15miiEM23wlvO5iZMaKBPYo6Qd0E8y2U/Q3fuYFYivw4gA513Fremrji5rPOH
Ae48U0+gQfIt+g1NtAQdCeqZVMzCY0+ZhC4+gi0W6eqlV3nP7rTFEYSSX+nw24nakFD6ggIzjsGo
F05zYPGjvlPg1lBmIrFuMwKFnVFrtkI/iTJDMzMFFr50b3cJzIVS1F0fHNnpmIlx+M8l53xTJJNK
NbFAknRjQVHwUZlfxy39Eajw1yhhLYW4AzYrcmCSFtQtey6W4MbkWVQt5xD/VgKK+CXGCgTexPUp
T4O/pxMLbZXFPmfECJG4+vBX61bYs19e1diXgqpNsV8CISJQIICvrJ69ok1oMCu3sAyToLT9oAUu
GlL5u18afg0mzZ588kAJuMucOq/3ipm8eqUqK8381WmpqXnRfzDidzSGuVIph6aKXcoyBdV1Uz9i
i225TC05lrm5+GN7tw6Rlo0gJgRrDs+ysDRQLq4rNTL3wm4dDfXUjLpM2eqAPqE4cAwLXqqxrCyN
uEFNEYg91kJabLyyp2ZJoODyTNfvgXxPpbZhHgnwnYxSP8ZKpVzMtwhDucFBOycZ48SIxxcNK4hd
bzEJiP6+WYvqAw4TsstvMTKxDgbUPH55lRcmFGE5PysBPEbURl95oEe6871gHii45oVA87/u7gzp
qPgdhM6MtCp1D+hkjWuvbjmhtogXQYihWOgKhcTSeGWmJo572alljJ4FMRvgfI4ykQaev9OQ1BlC
tkIbbRSWmiAdOAVLJwn42jDbLwfFxKZw17C6aoc2MaKjyB+v9XogcX8NfycWKAepS2d4Cqv+Ahfj
W953GSLYMaHbududZoWZwWQBFYjSCR4Lt+/nbgKM3r6PaW+vGYguNvO+nJSgSkZxLwOvX31Zy1pJ
+UsJqREOPuGcHCO06I5DXRMu2BkE/XAIE1Lo0fLpTBGGPU9Vpx+DTjU88hGmbJ1sSvgIPFx1b9qQ
mjVDnd8+Y1MPhlDXraAFTglg2H1goineYmu4Vn4GWm4rKSgnl9zaOMEkOfP5KD62mofwN010/SAX
RBdi2HQoDUePN0tjEKfEmVb7ipGnmWk7jXc2Pu630KcwvbXkOwDe01XpFKD+bjC91gqBndObUIO9
YcsiCvQMpW49PgMx77+QH4EmDjn/EqSJnW9gKXn+6YG0jKQUak0VRNSOaqS3n1UhoSNsacfPA1+/
Dm5luufYT8cVQIvTqkjD+j/vKSyZJgj9/RIl9NcxPxO/kE7W7ymeJOPPYycLGHes9ddjEKml9m2v
fYFumZtiGDyc9P0aDXc+DmkGmJwyIzEcAiPElziSB8aB38ArqO42q+jjoKT4BxiREhQrj5Wz4nma
PJptfWALHEX5TAr9mW1SprViCelptBQu8xSNE6J6ZG0so2i94SjB6+PGRV8BgqZbP1E3VxClhFL0
Zvky/eX+1W29ALKigCUSSqY1h3IdxaU6JjuHvT1UMtHCWEmexed6xbT5piAMQ9Ib3kzs7y0A5Q2Z
HZbfNttgIL5hSmA434q55/LpJmW15JJIEEvfe9Ju8jHyG4Cc6RdvhOpDiQWVKrYeK/uPWDQbMw+M
u73XJqyKLVdES6A0rjWg1UrZz4xGZJfKNIP1RHr9EPZYNvGJrp6R3Z+woymofOUuST/ruWlEYlGD
ZsVGAIbDGF/cE733SOug1cO7bPM0i5+ghK7hIoSzONLJ/Z5FdoFkvdVo2ICfm+jT03O8DsAsVDuw
lwMXh2MM6bKUJE1Fe7FWRl06mRwwTE1KLV7TB9fuI2HyY22McDy6/vEzNBUq98eMZLwq9hBLUe1s
LQyjDcknzFHEhZ9dUV8VqHmjO02P0FksFt6kuE8n6IGnTmh+p+2okDwtvEHYBWBW6+jinDw/tIgM
5tR46SG9GZJ6kXw5auIjxdqAmy3iKPi5J16e3FB6du6iq8GI8l+BUOlm+v0RzRmQsrBI8CZgg/Fn
QpJjPl79aT4JXDrpZCKDUfgX6KV4upb8hENJFTMh+hAwiw/UR/XmhsE2BUBQQPE8Ux+xk0g+aHhM
jzDxXuRSFdftpTUtIqyuRTwMsZacBJ9MrETfl4SkwU0eDQ+ALju2gep7Eo5EfymHMupez4OJMcrj
U5XzO+C1gcNErhWkrXvSrpINBujx542ajliXANk2XZ9CVxwKMyj3M3kcEofbNWuqvULoIgvkwNsM
qfp3jiPhPNpX1i33JTHlJrvG9KODjiTFFX49677qjljVPqqsYIVIZR6a3/f6xB9CXqilIJiHfdyH
qRtwktEBzL+vb3GqkbsISbOIK9LDiTO2TeEJ33jgrN9UJZrtSQxrOY3ERdNM5eYaI3zbG1N4UrZy
5chTOR2OD4rV5ENT8NlOCJx9292paNIdZBEJvcPYp5wHscp2YCvnP97g7M46/3xtAJbJMrFz3j4V
9n+20r+fWSOGl/L8Qk3Qc2MZrAGBGeyLfEzwl/BffE+9O6D6KfxJ4sFFL00IuVaURbL2UfZa2jWB
yD73H1j8XwJOlMyYDgWWlXgKw5VPq+KEyS0h5MRaoFCv/g1oH8mELuDcfRnpOx0PrX/jKKi7mE4i
9QYj/7s8I/GRQ5/L4T9TAGTGtuduaucWX+Dp/WSAjuYuKf1FMt+8ztLJKk6CzfUH2yFdaG8eK3d1
VSw12gkoL5weZ05AuwD/wl//Bag4rcM0ozmTGsY/LOgglMBRT7yLzj6/+o048BL1j+5KDt9TIZEF
iSlRRnftsFn+YeCl+g9o/jcxY+kt9GLiW2QiaRi5X4o8cb31A99EW3vRk5m09WFFfzf5Y1p+8zXR
3Bfggexy+t+iaGau5OysqxbpDN4Mvv7vKkldaUd/yw2HztaW1mHVAdqGs3pgzgs8TGhMDQqRw9Mw
YhgA8XZJzgraR49mpXR9ZGODDI4nXwz7EJ3g6oW516Vs710MBz3/lReqJt6lOpY6VXLmyYnlbBc7
iaSOsd09w6IPX1jxb54fuSzvPnFEyoWHsMVLXWdQBaowjtQ62PnhppFgjnLKFAX/i8awyfFbtLK0
JkIxp+TSkAQRaLCVnU/7c6UGAikCyDwm42M2d/APlcCm9YQMp7Yrp+dsgUYzBeX+OcAzMzkTyXVt
vk3XDk7KbptffHnx7zPXZt3oOUeebavbkAuOAoCNuye3HaMaq85vzcCnmWKU1Ks3xZHMEgj4Hl8z
hQuRFNpgGE9x2OybxerYVTTE2hT6tkVp/ZU6o5NAzhr7llWoqHS1U6FxRF6yfvgwvTBLNZYpymyF
mDR1zm3TZj2nJtNp8WEYK3b36+5YYCfxhWmf5p/2s/yznC26QcTMnKEuNj3JLOKKBdJvtRtnU5aX
d4/gEYc72v4TOLsayfSii3zCsvyJcw+3E7+0UWGISwVZztoQJG+jg0zIm2a33pgCM/NGFrYypNAK
FdDTV3JNC0IKWbWSEUYK8Rg/ILaKvz/U5l0OMnSrNHW4Bf6pJZ1x28cp0iHbbkv40eF7YsbDGpEC
RTlFQd2hLqdm6eEn/YvyLJicMda++dQ2GCpM93KgxX08rUfs+BmfoOppMOGs0Wc788kH9Hy/79Mg
tz9NCnu6qu9cjfD5ToiV/QmvFhnPk65VOgmC4vtRWYRw5wnaoc/F3YsnvUfSamQk38oim0BDDipO
oKcZi3aVONWoW73q0I+whcIeu5V1BICX3omgSY0rYowLMjUpp7qwWTzJBQT7whPEUDMnfZz95H+L
WYUc1K+2Rg0A3J2Z0xL4AgHiE4nl3MFu+cKce003sGTnaipfumKM06G5ecY2JUU9lGdaaucP5DK4
TnXOVqzT15plilOnBoi5CU/CIESmF3eoY0ZoKI5ojSWl2USFY8tOgqYcaevn5R+rzOvO0JEX5xZP
XRKsxc9Sh2GooOQ7DmU8rVek9CFMH2WDAerG3qSvFmrau+nIdF4d6nFmIh1S2difUKVOsTB3UgCB
7o2nRwEc/9wlTsbJnCmKrsf+8KBc/uamFD5EPgjupaZhhgB+aADpVmLZtAdYLQTZu/iEHDqvPLkX
LcwPQIbiU14Ufdc9zNTvRslqYJWQfxYp9soPeVkagLIgdOsqp4OrgTnj+Rw+RwbtVW9mLajZuiAX
HtSNgzZsXZdwiPYxq/DgDDsNifzENf2MJSkfDG6UMn+O3MEXpamdpLVrsX5Z9N3wSvHvniUnv1Np
HmMcycnvsswVG2YRs4kz2mIIBEk3twIbiBPxncRqjwGBpvFKUYqgEnoQgpnSooQd4Blv6rvM+78E
hR3bIrfVnwGw1Th7xzs+FHfQWGqk6XSmYXur3GAAzp9T9Nfcnn5HcKVl1RAUHCXUmjKSabEGC9Zx
V1Qhz+arW2c16/jOUzc+nLCzF0rw/5CFbWgmd/2I+JlLzkJU1V7BgXAr44H/ugcJG3MIXlaC9pgs
bZBK26B6xEtL+ZOx+NwPUdpQ9ahbhh8z/EdRW1LNHlCYUP4J3lXBFxcalSJMa6Y4qUtLBaqu+Hst
dxjoMqOHvuSh0UPFw3eC8ZuAXy4H7srEisJit96LPoarwZR+tJofNYWaFoYdMP9nSPCm/I9fhhYx
E8pSKO55rHixL39Z7esFJ+geRIQ+ztcWxxLJ9MGwLQ8YAmhWM3ZaLTFkfJT7Y+n5H1JIfOlCoJR+
VO/1/1krSMZdj/Lt+NPq7GX98Mv8g/4OrUbFIzK7Ax3cgOiNOcj0Ts2YjPlOcruEzj9Xp2lfHapp
7FdYbFBxTEL9gjAPmwwxml+My0H9J2qyiFtwHJTt7fthLdWP3ScDJQeT8lIVjEzXToL2DY8cLGws
lxLAeGrWStKyx+NKjRHgKU0CQBOSlRO8ly1+lGySwLsCHB9oF5Eobkc69HC5fNNmR0RIK/eHqtwu
LkT6hgD+IQWRlYao1yzoM50hTV0yPkdcy1ClHkK1qCdZSAowYMCEbjdPZ8brFfIDYONyLh7faauC
wVHEYB7fqGMZ03Hbb2tRDjFxBRB9FYYRe0/nPOi4bYDTy/orBb9FtQsPgSJSZiduwoN2Pvse06x9
nlj60YMagNVeqLf1gjgofXVSTnHuX0oP9Q61hSa33ohAYDO6fJO+LqthL1egyegNkmoWMfbi8lTz
iGnKQjJxRoOzqMdrPvyMMd87JeLUtAB8wd8VfQl+J+AyJ+PLRVbgq8WslxF5wtZogQX0JoecC7un
LrBNkAN9egKL3LATZkXrXGf7DZOf2vorAD4aw9M7op61Wsh3uq7AaDlv7hsL7x6BmGKTJaal9Knk
mwR9UvtDkewTYT4hlQ+P8WOfRH1/E8SuiD9id14GDcew4qb3eTpqDsYEPdyq58pDM52qNQk7HMM5
pXSWETF5FXlDH3tSEMBnflyTZ91X8/OU8Fsv9ycGqImLwzctXatlRuoAC9CtXHvUsxEW4tfo22E6
mkt83ER9BwOq4BEdBW9w+nA6ZWPmGkjppkfBcmfbARO54T3B1tBTHnME/X24V0hNhOsGgFsqVhoe
J4psiUlS1pnraO/5mgRFUlkDYVLCtpgL+5fpQOI3mGRu1ZftVUNGU5fQ6nABcxUpJCbTHl32Zn4m
GnPij5s64YksYhsEXBQDUszqQhJle0hL0aMqKoTgtAR3jRd02YiyTqmFjWCdTNiDV5NMMwa74LqF
t0niEdMGqCpULESQuWSMP7SPma8zVq3ckE9k07pyE8ivO4FpoeBTLI/inJemkUZ9I3ZDt1NZnK01
CmONl98OITQoyF/GcLy0RNuZPk7n4fgcag4adoM7VnX2PsQ9rKJHuirYPXmdeIgO3EEgFflqUBj9
+IDfwnZVS/dv13cxSGbHA9sn9B39WNGV7UQD6yCPQx2M5JoY5XWQGD9Y//zHRWvQo4Gb+NtxoqKT
s8vnuLqKtMw8gx06tQ0+cHCSscm8Fh1gf2eFVfbf4Yg1Iu8v1YRzKyhgKKIZaiyFuNbJI1wsxAcw
t+iq6ybh7t1uUzU0cDh/F2nsF1Oh2VdJ/ZX6kOofVTqahSav/sRLmocshaOKDjex4BWc5Bh+FlEh
XeoN0GAFaJ0eqHANBnzXfQE5A3Y+dDH4Aw++dZIBbX4drSYm3InX9KZ123TChp/04N8jR1q2i48k
PwM4erOXjwJfurq9DihJzAN/SB/hWIO2kIVB5DFm60SO9pLNMt0i/kYYo7+o9bFCK/3EZvhsJmGS
+XOidGlN9C7zmGClE03H8mL4IFKGIA8kMI23FR+YE5WD2jXAlaBOuduG/kI67Dz6899iPP/Scva4
rWKC1DaQgQxI0lpC6/FHtHPAisxcCFB+PCpQr92G+M9R2PQRGbGTcOLNdG1fAunH6TB5MNFv6c8K
XMgzFpajNUPxxgVtpKAAh6Z37akJS2k6nTt5qGOBID9dCjyuDtZ0ziKvNaVV0ohhEwmR5bhw+MmX
7nnuYN6IeCnsQVb5zUBRF8liv6QpL00ptNlcxwd+ccxCKATV+7scNlhrPce6lkCLrg0OdcKXc6Av
e6Hv2uQ9lLW/m1se41Vf5DW/Bkzqnz6bHIVDw1JBw9FOl4+dyR70egK0BV2Tv4G3vEVPrsRp0RP3
0EyMeg1eawGZ+IxqLVyTGZKM2Ilsx5AUkS4Pq6npGLp9XCgUBolWuzKdUH2rWT2NLQXtRXNBdVw8
lLe+lnDvIhFnnZklZWBZecm6WLryJYneeLyFM2yvXa+1E5M1mrqUd4vORDeY1XTKRVi34PhWFqxc
CA76yL1UOcxYxcQ8NkkL70tgTn1wUK0dAKLZzqvjiMut8vpG6WTxr/hS3k0wNvtljCEj1SpDVgeo
tEgn0InOqM+E2Q0aEnqu4cxh1ARa5ik1ksmL1rHZ03h0AmixvueQOjmoKzTfE2SNLc97cpFswmSs
sANPCeE84+bFpv0egSPIL4FBz2K/ab9qWyb4cg8IRCk28sHUaj7ABlF8odGRHecAI7G3P7fSkkAK
32G6GO/mmZa02vnSGyrSbh0SpRwk2XH6F/3NPz/dfG3R+byHjkPQCtVnJBIfhHPP3mz4q+J9J9My
R6yRWJqM2yRkEjl+lO0mh2Kp0KhoEWquKEwzCLGJHqPrymwXqWQkPjwt0mhraySTzIBOERVmXin+
5P59eeblAD3Xn0qq2cQwTiNQSkch/fn93BFkxWjT6S1hx5FRyx8R28302+RrHfYPx+RkP9ulnP7n
63+0SzyrEC7Bmf+FL5s1iun7+R5v2nflXvxeGgg1c/ldS/V8j8PEv9SPXoUWH9KL8thm16zCi5dx
zBYDBI2EPwowNX3jTxn9dlHF/BaWcs1k7iCUMxg2N07BQafdg5yjx7B3EQh5cjVyQj7NJGZljGmg
GKozKZacVXJmMEvlfpvWQ+KZ5q7RCnuUTdCpTF5mm/4k9KhubNs1bU/w34JO2WKgSHxws+mVfbpS
EUM6Q3kpxMcrCdSjVjFF7L5tOyDy5r57Vax6qPF6LWhYuPCDo9V5+j2kg2Mn2Zqs8AsjhHXnngZE
02E6dE7ui/7NHxb8+w8cmIaC18WAGqpNlozpJ03lrxIE2wdj/MH+Tdek/VTX9TCTfF3Og+Imz4jR
L03D74luKIoj1BZtzBhFfkh5GFwVV3agipVW6iaEW5S/SCRhy42gb2T75xGiRgoTQPGHG3F5CGcx
EllFl9Pu6Zq2xfnXawoUssG3wqddO5QCGuHYV/206fndq6rzWlkw5Ps27sLza2MFJlfkZCdb9ZoO
FO75vEQcuiBXG6ltoDNfzW3NOaH9VnhUFCS0iL30FrZMfYGzXJpo98pyXU/Uu3Gy8Efv9qLZbrC0
oZGURNI+TbfmiXK4zHFhbNGNt5cfKv31y+U622H+L+FvZq2ovkamYD8VOpv+1VXgow9CqOQc8C+J
pR3C2XYvkytF1/F4cQ2EbxHSzvI7xl3OQcxCQjCVXIbtXjih35eOVwsDz4ctMLB+W1TcQt/FkqkP
2dbbe9H4Ghj5gEh4vewvLsCBXqjv78riejCl5ruqQZP7wHDFDxmA6fGKbkBi/YvTVepwNty0Xt8G
ocGWN1Le+blfotwGqnWp6mv42Mgo7uf/hlAjXYkXQlIipL99F6yfjg7eSRNg2SCPGKk5RQ++hrFe
xxY0GnhpVllqyKtB3VugMMke6YgVYcWgDgA70TVvExUaOYUXCWSNNoRSuecFGGl1TZyhoRaeH3zn
UBYjBJqzXCfckvVkoXjKzBGnHSeRy5DTcRVI+OIptSdlVlclXvQ9l6JaooeD14SovIFIIR43RKQf
F0mnuLXkvH/0UNbD9BYEXUYTB1eSbYjySsjV9sDirBGJAA+BY+5FxG9vKmeRDsdHzRZKKBCKYjxO
LoDXW80YHVt2FPq/859q1RDO+opnK9HXNvqaarTdeEiPYY5qgBc1Es5pqI+2KjfyLkB9NPQVrZAV
ZX1FlJhczlIT7FkKTdkNJcwGVMtUK3I9CCtpGsCyd7vMJcShZhGrH5dXoAniwNk+7kPWOtl12or3
V/0aTLx1F5Zvxd31r0llEI7FUBNZ2KUJ7Jwj/8FPCNfzSe1J8kh+FWOeqnJtiTnVfjrFV9etoM2n
YXXyU7F9cojDdfWzkGeVuiYveJhVmlieiGPPFF/fCWSloEagsl4S7uOrLSL7uawedsmjKv0mRHhY
igTwtnn0YSp5fTuRhMwoF/LSFi8sw7YG6KddxoaPR7HiG+WWBMMtbkL4JBqYLqbC54f/cYcu5T6t
xp72Nu18qbudnDPX4uVzQhdcukRF0AVKdjqo867C2REbMmOLTXtm23MgAHiusxRPn7KtD53pFrgl
Auo2EeCbiRQqib5/V/7iygMQRec7gBWib59PGRTUgBWExNKzqXPKFLjUYYZQfpoVveGcIy7qo7vB
9QgNFn/FhxLRls5dgkQfXcBmnqHYU6rwllogQUXLM4Nr7HOomszopt81sQNLMOa+Jm32bD5pjiHP
dml4nMDbiWK8vsBdB+UKAeqZ4TE7EAbdhPLaXiBRtDmaudit6XHWIT0ZBRxPj1QWmX6aIZ6cKhZN
WCYWSpcJa+QuBrCQ1LGDWZq8dr/0jNcOgSiHVvKmkyR6EZBXUBsJHlbXZFZWadwldX97vZ5c/Dxb
D3mhJPk0NWBDsqbSGazAoYKegAv0h9Vlg0YTdyF1CLfx3Iu70qJw867ArlCYqU/D1uQzzGrKyEpy
JwYWFA0vtVQbNOHSEyKV6yTvQzWb5tuLX8JVu1ALjXHnDspZUI0qO+tH/6chlkffcRj+uPDqj80r
CTmJFFu/YDjaQIJcWQU6jWK/2v9GvcmT7i6A9OUCAnZgsfm6ySK3DLL0bq/0ADawontUcIElUUoq
978mXCxce8vQGXpmnOzVaWLrFbeTtJ3+w6p57pToTXYbJ7J7noJ9vkwAv+/VQ+vJ8r0AvJVy0pAh
jZC6JiUT+HSucSHlXJkjxYfLBd4oCHqBZSQ67bmy53Yl/TsfVciUhQyz0k8DIuybuN0y7/gv9NfF
k/FVTSOIf4eQQ2ZQFvWA70cUDwnJGLUwLmcOvqhCgzBJjZR6WE2Zh0mpqJeE3M2Iz4Fk3/UdoWgq
1gJfHzwtuwdibGq/JJr3vk/5rXgtQPEybj/+Ws68/y8jcuj7A3FWKdHhRXujB0m/ePw/y/SgT96x
Q+bhwPAfNnMdFGrfMFHjhc3+rgHhhezc1qj0GIiOYGMf3k1DyxkpeaRenRqIFy9ICO3DTeOKaNlb
IUihp3cqsVT2YtR8Y8eMRbUhXeOOJ5Lf/f45ky2m7jxIcsH6d4l9LS5+Qixy+CaJFKC4IKiobdxT
ery1Zu9bBj7Rqu1li2tTHvljxhsEiVu3uwumu38uxlEUIrsDQp3S6o4vCPcR9Yx25TQmpw3rIIXD
cNZvWxLvxYvgvEklyTC8J/Fp/v/TLreBUP6eaJX6YIz31+TcCA7pOkP1RYNkdwK66IV7Cv4vltsO
vMWjzWGdvGUULMOV9AZ+1db6bW5NUQhbM40QMkQJGSN2Y2L89sSUbICABmvTYHoCFqV6WgzPkRzU
TCrJxIuTQNCkef/n7Pm/MKM5as1W50z2P0yILf9xEH/A+X5zfOWUqGhaGm3Twh+itUbtDpBYTIDX
hjjnVllRPWgXyr/Lf0vrylA2oBK/R0k0MogIzeYeHEqfWaavB4C1sJ0gnDUjmsh7GzFZL3ElLr+l
dDHjz5I2suEEMVYlNcTpd6UCIyAYwZ90pq65Iv0kzL6EFDUnOBItHeULPsUSwwd6J+WV7ZjGnOib
Ow5HL/533futnT02gSwowuHVG45b3R8pbpjeuWWOhvOnBuzHX2X1gc6K4w7V1yQ9i6fON7WcKUEx
S0YwqznKAQeUg+Jj99hxET0dfCILbR/9FxIWmq6+fCu+14PyA7WFHVCSNyIUTfoGlToBr3oihPXf
3bJZZJRFhFWpP0VMEegFy+dy5mw2MO6TjthiitNfjo1991gIfVR1dJXM2p6S+03Jw7rWkuTov13z
7Qf97fzcsafMNnkH48Ni8rglBWCXy5tIsgk3AAqu9ibJ7DmvK0R7nnzL9ymZR5ckOecWPfXUapnP
JvXS8isCQJc9B4CX+IG0219+DK5Q2WGawgN1X9+0BWcbQrIef49daH0gc4Skh7sGidX04ftjXJMz
4Y6rAzeyCjZCUfIcUCdSAfVZecreWO/29VUJ3BeTA9v3kV5KyK6Np8xFKGmz1zTZpHOywYUbVMz1
gY5NPYE4PY8Usymhw4grCE4p/osBvzgteLQHUAphMaD7gLqUH81ULjIZ/vxnr8/oTLgfWllNvmw1
m1S7Oi3EUGp/JV26hXCC5pG0sP2XnSd8gLuyCpMkVKLy7QID3UhPIAKBvGc7yBL10JUQgFB5y+Gp
NzqENfrk7grreBYbey5+WzXuTkgHAQjZw6cVsgxD/zDUGyLLJGvaSke9xLSv86xCrnC1hDWBPL3X
it/OQeCw2XYKRda2cTL2PxDx+gjG6nlw+mDhNakhG+PtoIsreVLfHGPD7v0WX/7Bb3AyxVrGEkof
Rgzkb4V+PiiNekT48b95XzarGGL9vlSJX7/GIPbdmzRPeRht6Ha0EX7m/yWjfCJSOnlKeGocLumF
q0GH0+0AUxHz5GaBlKG8a90z9vsoiZFyTxnY/UtfPP/5CoMcSN8/UDAISeEIi9R/R2ndFZvFoujq
q7ocesilI7KAy/WEZlRznwkiBvYJweMxatPygf8sRdzWQMCNXYE/i0y2vAK6XUaHo4we27q39GOP
R7UTpO0OiQK+oRarM3Bkxb3lhQ6J97K/jgJhJ6GcK4LJJjTMZ8OV11T77ak2Fa8SOaWAWjUJ/3dw
ZfEegSgExcWYYh5xjaqsqLY8Irx8Idfcdw+iPDQkw74zmfa5e1tx/vjvxbN4QBocyHjet1n99qYS
EQqO0PvkMqmQehZ1HmqeorLxjnk5B7BpVH+gwxXgsnqWPXXOvca7xAKPly59u6Rqx/kgUdFpctko
FuRnxQpjQKT1SDsXIOlPMahFryAL5N+xoxPOx2LTduabEd2bTp0Vde7Pz9pr3IZ1PuX383aQEPKR
RsXCeWrqUEor1aWU5dy98/MUmGkOLtZXbHHWPSDnSF3Riy5yUBIeGNcpYuNd+gNfBvfS/cm7ClSX
eCWrTwQs76i7a4lHSVwBWJGSaMhlMVl2RbaaBR94dVOY3/NWSS+GXEOTnM+VwwIP0gq2BkAIpBdu
MWRkzHipI/uYtsVGvP5Lvohx+vxdDaWbf+EtcBjQLiisvYgwU4b2YyVfI6uuB7rN0ckNcUYPCE/j
Mhq7DPEji0ipqnVvJh7WB8bhXDjY6rHPEwNOd8SDOfykcuG/WWke/8m8FA8P9hKbElN8akEutmN3
QXLdZ12BIKV15YFLhhfKgcyGXd26R9+f0RNjvtkL/mqjFz57UmEoR7EBTzD0mqZoz5XXIfg9nNU6
Qtga02Xpskdjus9Q/27V0oEYgHj+Qc5pzDWHhLy+nKB6kX4HQtM2Y9V5KZKZJUtT11HV4jhGngsq
Z1Bpu2P6KBae0cmEsxJfe3r8ZkOqK5RM5j2LBFEt46BxEeFyrhh1386pYtB69TTP4SiR2NqK1Y0m
clq4RuStiXbuI7eQrtFRV8ix/mmoNw3HCaVD4gzkqIwsrS70fgTPv0FglaLTbSy/RZRhY9TRYJdY
icfPRlKGmnZHhnqtr+vHzWRo5Pxq6mjxCpcc9eFOqpzbQhjiYwwdzJLc7lQhDzoHv2nt+Rsqpqq8
VE1DPnquxSWirEdCkg5DEyhlrf7Fswu7ihhKGe9JroVoxZJe5ZGzbSaVZtruAbLYEavePTznznuB
EK/i4CORpbxTAriQkWFCwNcdY94HaKWPRIx2QMIih0ocEtIOZ6sdicwYo9BZaIaUrvyYPfAJS/fs
gLAwYGF2DG+p5LfTO3Mi5qcZpEAQAFIUHlUNtf5OZyJHZyAWNSM/CL0+/cwAkPijqsKEYRByNszZ
Z4OLtXe3/u1ZKfa7DcR8xr4mXu+gF3f+++DFR/82MmAar+7xlWGeprzXBA1/4vjJDkAOHVsYqzqS
8IRhayXODnofM1Q2Av+73JtlDUQRNrZ2ArKhMb/wAY1ecz16n18aXnyyKtbOqEleswM4tfGgfeDm
FDjbCBmEh/5oR8TCASbQrcvypzw3DjhK5k4NiboWe6zbAjLKkORElpQoWogW2e8zu/89mPSlCgk5
heZxRNXQXfTOnkGe1yUIwthcerj+3ilQVf+FNAcVX7inXr0Y5xEZ1rB7p+osk46KWa5lhrxGAbMa
5rqd4/HEt5E7uI3RKCvW9RvWB3j/dIn/ulkR6ezSE4yqoh3lZtHfDtwMcNHjgXBlI9A6EQX9HNoy
ErRtxVrpwvwIGKKp+N2ZBFC/lAM5nYHpXGhYULZ52m+tULdSkT1CEPFpJejq2dgIp8dMoTY04eq0
IKliPZVM9TxE5+t4zUdsW7LxHht08O1eWkgz9z6v8qYobPLSUNqzOM0iO10jGY6LuMh4pOwgzMxC
W8WOquKvMhPahaOS3mhbS4lHQ01LWE96ybQo1JxuVD2w0m9hSyjpBKVnDLZl9e2zWBVtSTGr571E
zOW4VKKwG2AmH/8l9eYX76AEOk+mr9rxbTomCbGujxhfmCjKz9J4fV16EJ5SRFF+xCZtTva5X4pn
SRalMpNHpRCNx4BGeTUHdNpOouMKpIkamgVXGPJQA9QY4WbwoxGIHv3E1FDq3WTYaLtrZFbrAzkb
NQvul2ocnGYBKD+A7Rth8RaFfbVrGvtohJhV+UGHGgX1ZykL7Vqya0A78uMHD0qPajH6+//NyZzM
/pxJuxqnkl5okOAsNljiJKfxUEXfAM7WMsUPQ9B4ZqPc5MkJ3VF4SrQlLEmkEdm7GaAdFGSMKgHR
/YA08Mv03p7PfqNbQHc8Jw+ILDImpFWUmPdOXKaL+DDIk53SJ21ap1FRsGqSx99o1wWvoNZVRvQh
V8Tf5+3vSTI8v5lXCEuP2H/pL4hIrXaKmY3FEgZ8Qk8n1bX0PmJvxL1MxL36xLZI5EcIdT4PHw6x
VW/MCeVmsWZ4xsPTl0SZUiSCa65HsbzbgFRKAmos9+6+cB2MtknCOVNUWenthp1UU4vMsQAP706K
nIOXdts1cYrphV99SI+LJklhErQu93eYfJdEI7IL5Jd9bABbQXdLzxZX8LYO8egVYwStTl9Fpdhm
K25mTLwDGmoIuaHK2tF1xX9QhN9Ber4rxXBOtxjVGUHJvHN6edRApALhxSIMEaZY5esyQsNO3rQl
ROrvjRtJ8RJ1HpokwvgyyP7g/oz/wAOIulE8eaTbDKUwpBXWZqEcPscsMrDDrHT08WDfX6qgz0Uy
9vpdLgFjfw8iBLL5Fkyw8KGR9XGOFHX+F0aTDt12AujnioUT8L38hA7hXCtRAGU6kYpoGOQdc/p0
VuUK4aSxNagsKeM80oLHQfi1TIxBfPAtP4Ud3S15pOfh5Ikhl/KQ0om9f6GrsljFFPKk5Fmq40WZ
GjrhfgztFfDa1FyhYIoPwz3qsKKVsbDH0Q7ES/OzJw0hSCv4faiVdU3FqYtYztPDiuozgS9+HnEt
M3wH/ykn0HQel9nm8HP3wGjfcO4qejIkPxu55vgGLx7+z6olgUV5X+TUo5WsLxRHp/pPfB96wdTl
v3HYymBIg/ujYQS2LXk6/vXFuN5X8fXmlGqOC8HYWR2Cilb+VNGCZ/30nby2X2gwQBKw/0f5ox0s
LZ+sB4TYsmAIGPI0ASv5Zwpmd4hxJurh5u92Q98bUXn82HoE9WW0jgzasWCs0zz4oYA2D7BKvD+u
ap199OGee4k5q6gmDuNtmCNnn7qZcL0XLSYel+e2hnNhPGks3FmDiXwvFMNzH9sHX9Mpp8Act53a
y2HMvURdKdEHTYaMyR3gG1BHDmO/Vvoe+CxFGl2/+cLS3OyhFLpmbXQzEA5EINGSFoWiKivpA0cc
d7EOXcoOK/HVKncW4QkYbf8edT3V/Dlg3zUs/zpMDnflDW+DYqZGsIWCdb/LJZjLCK8ec6haFDLv
ggL9/u7/QtgvsHOGuVHu9NjJehtzw+opu4f37FyureIUOvDuxxv6iBZ6zzXjM75Hdce2SAEqT+Q/
BPum49fMsro/usTXSiobPs+eW728rgRwUlMKzGKlYkaa+3lhm16uMmlxiNs9hdTrqoifLg5rVtWb
+H6q+FOJS8RwO1z/IWnThUgP9jUJOoLg3M9FnzFK3rhOTKpBSHoF1bwVi25nXD4TPa/10wKMAVMZ
py7TAbAD67Uwjh9NWFbWV4xzFnbOGthtGT3F6qkB54wqMP69QbOGGIwYYbupC+F5lS38WOsLJ0NW
ZzuuSHTwLgbRFTrGMEzEJ3/lGvyND3kvLvxL7Dx9iMdhBfnw01MZxQC4ItKdBK31FH8JJcJF7Ok5
HcqNOrLl7XmfvFHR8iZmwS9DfzcrzV/beezZqrj9NE77E8a/WmIzUiEmU6j05R3V6yxH9ffM+ImN
gGPq0KAO+VPgfTWa3oGDXHw1uNpg3ZAjOnyHyPKg/IbiFSYRICv1T9QNGEX8wN/vE+okPztQqV5P
QqlYRxu1mSF0R1WhZtOmQ6eWtxwVs0pj9AmxqzH5FhXp39TZdFw8hCJx3GYYcGgykDmL7cmJWaEj
jZ0fDyHBd8MA4+rASJyjlrgfrTI4zTDlklwJk5qiH3fdqoxW4WEijDno6O4Tr8Os2U+spXEQvcnF
cohVqRmh0yO76lyJF5hSKZ+MsWeDNeVK4b64SJ1G7///3HPmuCO3BmhfT6Pcha0WZMWYyHq8tR1S
A5Orh81x5OzIlspZqCei0KxEdekVBtlKB8hOu6ZdHKZuzHWuEG6+rNI0QB8tSIJ/hnlLOn2JUUT5
9FIHbLksv60/3bOUQNIMOiOYUak9/TSA8R28YzNQ62CybgDTZX7MhOeVqD06vlR0o3WrFLfawYr/
pHup/yE48C14zGdHkLJH2s4lbUXOGTl0ta4MhBRe7rY58uHN0djp20aIBYzBxaU+FZvSujQBHG7E
9U2wqm6cHMeGnEyVTnnL1h1t6WGl/Gu8CQrviQDIPqYWMeBYMbkyMR7H61lQ6qCKA7iOxnX/DOXT
lAXr9DOgJWngatiWo1gQwcilqAMpy0F+JVDpFYMHusNlZV0sLsiqOkfhckPRA52zZlIg07X3f3vQ
MIRCeOcAYzvlnlxtKCX63HLelT1SB+1W/hyL/eRMzQKhV4xjYERy0pY39lts5pwo68NLvJiqqOG8
iiu6MOrSj8c52qDTMBbaW+dfp2zXYxU1a2zhnFFwAkKGf7XU05dbIXgfcFTUev/BJf0SjMhtbOe4
QhChgLUDEc68WFruo4ahVGbVlgrwxRaKonVHY71694po3Bmg8eB5beGEveHXRNuqzpdkVtkintbZ
81Z0GfDE7IXTxZPsDKE84WOU4A8WxacEn6dHbZvw5QyJRWwUoQYOV9RKhxhEjhXGbz+xa+MAo/yT
XunRYeiHwuTPTxda2FgRBHspWD6ndxZM6JgtTB804H/b3nS95hcFWqnqdMAwUasv+yZSQPuuPmd0
AuWG01CqWpp1tagcb/yqvX5WebF1ECy9/1cTnfMtCUKDzMrqQLLQthrRiQW/6Vn7n3CDUI9b2+/T
NYranhEecUc1RWXqVoOs+0c26AGEIVk1DbCeYfJIVENIqXWkatxgmSC3nBYIZIROikX2fVQJJix5
qbPqDxds6d/CpOqJvf4NTeHpfF8mQrDmkRhLpNSvzBWi/VIl/OPVv9YN7AQfzKrhPWpRA+yutk0M
xZ1zW8o/D2LfJjIk/b7BI2sj/ADIJk+QgHmU038wdRcbE1xEBqvpOd1i3QXBwIAdZZfFMB8arlaB
lzaR3L1sWEUeUOLUdkY0MLIH4MJeGpBfH6TKechduDLa3v15gzXzd9Kk1hvvlMt/eAWyB+6Rp11Z
PxFFbN4ZsELFzV043/b4+jmRxUEwNCrBPx+QxCybEH1fAH9HF/NRsqL6eA4fMP/b33PnpfAuoLYn
4oVAF2KUKULsb3Ee52bkvN9i91Hw4cS544OBXgCzmupTZMwdpwxvifmXb87yqH4dEjY9e52qIP1x
rxp6ueG2M5X6tcF/QRd0Nvws0dQJyNhbnotC55sB5qe0zDHP4qHnUzcAnzj2HNQuVqAVZFfKLjSf
jyVj1IDCyxrkb6RC7XBt98hj1vnctYeNb31DcHl+f00ggOIvWTN5e70q8RbJBxsiAgwEppLmDH4t
LYw+vZjJc2lgbVn+YXm5ay9iZ7m2z9eCpW40e4814Npi7nwnAyYYibbQjvgvx1lRbPwlFL/xziQj
Py3aIMeRNAGhUV50IibLyuwjamodaYX41x7CyQRDuXBpel4OFQj5AHZIrAGoSQy69/vbbizL8ulF
sxEV7s7q0HiErCCG8U5GBS8tOu8jPUtjUxsNOWFK6YYFC7vcjCzJrIpL4gK0omD+4qhDeEhjtD5Z
KaP/mp+ljctSF2FcSCfTx4U6rl7WGHINRQqBbezFFbY3vwxbS4t0exB5fdqgmFWCtszaHqYx2+vl
YjnDf0woPJpIC2ww3gzj+mRGlqZ/AOWoE/eLcry5y7urEqNTnUNQAW1vbb8w8kiZxFKNCcQIfpPj
Gqbwlt5sO+k5lzHEBp2eFHn4jJDi4+smjU2PLRMX2byDwe+nF7l070uVkBwS46YJQGcOzQvsIoIB
L2Sd7hs3SwEIN6O1+rmL3SDVB0J+UvNwAySHh2YCAlCuvA/z5ttWI0ZNmpawSFUfQDJDYI/4QVUf
GTmbwe/jVt4UlYsxnxZ6KnICDNIZLWCa5hgFevmKLIL3hCNuwju2hGOoK+t0Mffi3J6GMoDUDMx7
a6IVpE6WEU269wx5wIQrQBYxF1CnHLXK1msIzseyYGK4F7i5woz9ACNe8EJ1vXUlvHuWTskKJ0sT
OVMw5FWpu9EXcIjVAPmNiaU9GSXczwN5uqmLCwIBU8yLrEr6YsOabbAb3hdRbdGNdDcE5UXXL+E2
QpXVR1ywElcm6DQiiygFk6VDuYrpC8e2rCE1+W1J157UPDFEJpT7+2m2jCMOThx7n8Oin6meFHww
To3ojEjgQOQsiJvWSRd9pQtntpeimmPn2H6PDwlFKh7N37mTpLarpdep5Q/I2dmn2vP1AvBWma1q
Xounl3Kubtji4QCSZuX7F0MgQT7V3dqBwjuykyoUZsMxChsOJHut/Priroh0AHA5J9v/yLpoFhbr
+vZDmVn6CMyrRQjK+jMqOJvUWBe3gf3ZG+gs3z/oP/g4L+aylARzUYoYDDeHvsNwv6GohQoVPjJz
35vCcq00JCNYYXe5aidb3xQXZJzTbmZ0zG5VOc8fxdtV14yJp6gtbdgijc3EN0e38WzTkf12+TTX
DtyEfP/kuMJWfegEWWYT7mEziJsUd+7K+2rUczpIfKuQsGcu8il9etqu71/a9rqko5/s3SpqKXfL
M2r1880h36sPGfAKubQAs/Os4MM7PQN1+sEXCf4Gs6FQytl2mcGw+WHJvNFgBIfkmCvGc6dE1H5a
O9gdFqHEoOBYCKgzYlCRQYZUkKXbg+BKd9sOPAVsEix5ZxJgzJHSDKdAtlFeXQcGBy3U6MGVKlHl
Pz0JYVXD+ASunkv144LVBDB5sfwHxiA7jxXQwm0LoTi/jZ1skB1l/rSuWiGK8L6UqiQ9DRqCIgBC
IWvdz1hqv82XQo35tr4DaorGd6nrkEEZU2lmoIUthfDSaNTHcoYmQVgTINHbdkiK5OKeLd7GWIA8
+g4vlA+RatwcAitlemzoRXOlJ5sDFSBIOqBHM8Shg/g8tlUJ8H0UMkGV8Pm1M4NaI5R62fd9d/9+
KQeKvfcEFYSau26KkYjESxxjg7lFk880PdWLJgTc81jIiuKNqSeuctyhdwaz3JY15FuZW5AZaa68
KTgMeLsef4ir00svab/KCvrk2Lsk5XOrV94xfLTDuGugVQZM3sHPmL+EccJwiuULrbBsmbtS1KGQ
Q7/J39GKRf2Jbd9Sl7XEIcwE4iTbvVjqzCdu8B1BHpX9N4iVBts3bDWmap5VWUafJYTzD9PJvPI+
0j9Ft6ZQnDcpUJ10o70U6PpwBNvet+FDZSfl0zU06lC9nSuHAPlg1yGswA75F2oDza8S1eBImOm8
hTw1QmTwqLkjwWyf804hk8t0270Fxkf5MFQh2QCcOYMGDpbqLLRwOm+f1crknrJq1CPZeX9b7CM0
pU8g0wu9Ml3fSHWT8Uauxg4XtUOLCiG5Y2O4dptuA7z2Ij7I1bTyrVtfbJ4PZ/anfghhyXXx+rpv
05KsgI68b+o6O0QmtoCjieSNdLrotNHWc0Q9y+Bb+/xlBuNdGIK2Dm6VyhGWimGyESu/4Z6iPl41
NmetDBgwjmZbRBwmhHJlrvbRyx6VT4pS3tACyeMkUibUN5gTYohYIv1DqUnE9b0OjxBa9SFi/HwD
t3JH7UKD1VgoFDdsccs/AApZyydIyuZeXq5Pw9uVqPOkG5LpBjVRZS0kOlTmwO/tBbMwetH37ZXU
U24wWmd3yb5bLp53AyrvUk5DfuMHTJNBc1WdGPWmRNuvJ45eR7sH1hLijyNxnc1H5Ecx/M59MWHy
hjeRaaR+nbV4MNmiWgZsMfqIR8bJ1d+J0NkqQcwq3qoslLCAbInEigT1NMlRpuEYEGrMDr6zdRRI
dasPbJolXH/blo5QneMyRXdvwyRlDmmetDQVqRltYPWgC4Hvr1V3jn0iFZSyc8Ax96RWJgREvAuw
WNHgsDgvp7zpzcvd86gyonO6XH5B2mKIHIkjv9w4oF3b2cMcid2p0bJKC/+HgQxhFxD6FR5csv2S
+8e78hRoerZS6v7tpt4hAK/I7REjeU6dwD38bu5rrI89kJeaxPkHpnS5wBRDqN0BCswtfj37lsCs
oG2eEVc0I8eFf3Vx76Qbdwpo6nHm1jVuEcRJZi9soKzT5qpStFijj9VvqfDAznq/CQi9OY4NlFS5
XgEnROQ1Y0VJzIQ4Myqg27lN0f+nF3AKqujPPRB4z9EsE533Z8htAYNHGtWPMQ02gXkWGqbpyumF
5wj3wC3C46E+WF3De8Tiq27yCD7kW64AcI0ocr6Ok7cUL9bkOdhzqkCNZg/YBxmPk+0nnstxGnkO
Q+zEBHSewtQDhbfPgEGGx6dBMg1C3xHqcJNeqnNt+vF8i2dJwIsov7um2KXJ4AGCJucAaIcJ3YZD
q6cUqALJQwaBpeYy3kClHd/rJxipV6cu77ws7Q91AOJ+OjJZOfbipAht6gqdR1wCveAU4v4b9eAv
2yaYcLUrbqjHJ6zKL3+iG9wiO5eKyxAp55KXHVcOROiXhQhdUaMwFFtSXazXyBQEDFn6K/0sa//M
YPKzG2dpuV6QcAigmjb4oNykhVF/uDGBx/0tXzemTQvMjCZJHKm5T+UVkU12SKoKxCfoLipD75gN
DrQdEb9xbhqNJbMEWEV2XUcLCZNlValeNZkh18f62+WOKS1fVqebRIUq2uGJ9HC9FLLr91vJn7j6
WyShpVXnFUy9IHch4Vn3JtKGOYezbDKOLYU6W0MxfcNDsCKn4WhJA2j35SQPNnX50VvCCats/2Hu
OBY0hMtb3o+2gHrThGDSUD7kFIp6a2lnoNuxJsb4HKNARev04j/BqBKgHmQ2wJi53EyeVzri3nSZ
15BNAoOgn1SLA1X7v8N2sJFIuSJZDxGDotC/WnbW2yvnntzka8Hxi3JMBuWBwmo6O0bgD05ox05z
FnkSSwm2i/VvZoqtNk5ZOOylwfotDRyTTaV9ZH0aAjHn2pwHXD+7YsY7aKel8c5/xPHcWhK3RVVk
tknZOi67v8ynuqmxc1312uIkww0WowBxAWonDrPjiZbu+QKCrEdVkWcrJX7Mipr2Kc6nvnGkGMXS
3uDquIq1TISPGzDAaU55vKLZjKUAXODkcgm+dBg/xvId+ojROr4Oquvq0WDatRMDs5alPkg41kF6
M2M1M+2dH+pNrRpR09em2tiLNFXxCu2NG3g2LIOVSZxFgrVuAXtovbXR74RrqCAW2UeW7o84HEO5
cT2g9ZsgG5GYcrB0WBWtOSb642OWcKHct6CrUAOiD6FHUIoM4xkGkfzZDcimiRVTw4janiEQGgTS
5WXW/d4/EJx3Zx1F2sRmtHi1pxzIs2WLYzhyq6WBgFrFQjITkRHimyfQuQuDX5Nkiuz6GkDxjzCm
kAoiQVwFUs1ZlrkOc4EirtDE16OTTro3VB+DmkyREypyWF9LNKwGXR794E+AhndUjtIShJkxvaz3
XqS+qGWHnpyPIq9nQz9gCf8p3uohoMp+KNdS9xrwS4rZ8ClPGzXJQUislEVe4Q2AgJKEqRy+bfIn
N2xthwU5Zjrhiwa/HploXywUPMwFSQlhsCa+mMP+lAZP+qAHrNb3vOa/g+EtJipr0a0BzCRA7cr5
VjFipKlRhDaQjoAqLmRMt9PyVBV7dPTo7Yt1SKYgZPDqc8UOh1XwJDDp3uET+Fxqx+FJgNWNyDqK
PrD8nIpgVO0JPvTrpe873VLK0nfb2gSiUMDI1w4fmJ2pEyqkPJA06JXF+9Mzbv99aTZC44BKA79K
TByxIjrVVQY0rDgVk42mdKcPzCqi6zB5Ye8L+14Guf3Zb2InQ4JCRerKOHdyP37ZH6a/AOkTfAAC
pDFFIHui0U5JVvPNYdErOXOSSL8J4P3M0YGa1DAqR3xdUXiUrVpvKdVllDh5mVAds5NsOcdAiaKq
auxWN+9ZUe26M8ioDrdhIXxI6lnkXhKardSfounskqOwPcrhqwD+ev0gSY6QFGOIA/DfEM6bXLLU
hl1zxDX5TgxATsv7vM4+RfhwCbu1UQ782Yp+z7uvKlf9jewKUDWaLSkv6eG1gvvkLoH9tuOkjUhY
VxqA1mxZHSEdxITZpMsSSXGMQ6uOjXpOGkZxihm32u3zWHbnV0zbuiw1PFAPNjjI1EtTUA/p0GmF
d7VnzTICwpoxs+Db86smxOCoqBXedQTQvohjusw+nA27AdPuCGQbZuGmtw5wx/if6NS3vXKoPCdh
vxBpYGh6LYLwcXumQN4b7FfmUUCcrXq8aCxzj00AqlGIqgcqOtoLmuX/bv91zC5gwZ7D2hvPMavJ
cwFCFHGmbK2GIG6pNagoFd+inSh2MZmcjbmDSjDu7x06yGEGa73vc+Nby36c7xu1RiZtkqNyHqGs
FooVM6g5hXc/oYfAJKVeKRWWqJVrYpXAw1WvM06q+Jpjafxj6J1waSkae9/VBZ4qrO/hhdbP8npY
aNqquQnlq3mUHozHfgViuv7DFW/tpVivnhZmuPTs0DOpuT2Wi8B+ZzQjxecrKDWTtpHzRIOKoeb+
4MjkJQqn165z1+GXyHXnNYLI7NYd+knW6sG/zOM5jPhqC/WhYqxx8S0LSqeHxQEBSmah3lGxc2OF
2XNbqdV3XoPvX3HUglEgJdc4NzKPqoK9Yw9ifyNPd4je51nLoqqy884risNctwdJ29IA6/XmGLjS
xioZcBW85KvNQfWNYgKey183umsXrEX6N+F0ICqnzmplqTXLQf3oGAO9AG+ttNGzjvPHMc/4zigu
hHn/0gqxn7GGSITfAS91rs0xX713kppPU5xHnX00X5wbeNM8CYHC2w/v/Wl40x9uQFTQqGszrgnc
j1oYlWWOqs/h3bix9iKCdY3PtsBdbCIwgevOxsX2ji3W8Gyg93CEunMQomTSFoniwrSP6oPWms3x
+s1CmfasqBr3w3pnjMYik0UCHU3ZNT+Sl9BIdI0NsacYxmpwcQajNrHx8KU/39qqN5smOZj8Hv0q
XuV/V241Tn3C9hiJ7p37ewvT9LkMHh00eF6Dg7QCRy5rj4BXjp5VilQtD0TEr57iSKVS8O+4UNQL
5pzB4HEcOUA9dJUg8sRRGMm9ffPPq7LfhW3MsL/AxlGqLdMIEbpfKnL+VrHNrxxA1sGQWb5WtYH2
ZER3Udl1qVuwhjEO8713N5T74dzbKDEyWdTGg8nqcjv+rIUN/diUIoyJrWynEwhzNO3JlKnQAF8N
84eL1kMeY4ovM3ud59hhVAp8hou36JHxOUTrlb+xlgtYYSl+eoA/fCTpYFZ5DUjLFfULNNtl8Z6z
+CSI88X/eIZ1j5VL0vHVz/P7Q/9fcjVioqh57+jSGf9/Cho7J3ikiTGRxQZAzH0ADKkeGzO+X2qj
7Y1uyEwGsQykUpxft9evVHVB35sT/TpBKFKxHykhGBWF3IAKjQKR82LlOwzkuHog9/5Rn2daAClp
BWZ7EgJm3Yw9sd/J2k4l8WyxNcjkWOUVu7zPrGXhLu/izMiAIVoCF3sqM0eHF8mDwnwgoYBCQUVp
Gcc2eiw9E230pDMLyYf9BIbmss8CmFDkVPorun5jq1Iy/wRs4uBGmeBBx7rAohUgGnoh0h029EHN
KBCcNCo/FAowN9ZltNdfq1YCA1+oALYyi+jE1ycqIpgEOYgKkt8U53/GO6BmqERk5w1bKNRCgOe7
ug+S4u9zVYznpuKcQUzMfBDbKKEmJStCkv/h6tK8oyKKX4UWWTHMvbM3q08MZTg/O560rAARZnMW
wZglb5FPixhgokdW9tTPFQO2wkStuHJ+Sr+lzc7D1BYaEugyyBtXl4vqydGYFxbmcXbR2+uVkgES
q8UJaMSLzTCNOHaYGAZjwWSCHXL7Uyyq2zlrW7AUHj+q1ebqpIZE+7NTWBm+aTXvFgNF7IMqjSoY
DArmZwCMZ9TrjOnrZw8DhLnjxUxXwAWpo3BIuLFJnV8/C9s44OCEMdoxmEj+qjApeiq61/PxljYm
r0yu7JLkARyT43YNMPLmwhAgUIMSqE52lOGcDJw5CBael2oFBI3cRjGrsOo67VybgOKjMXNiLl0M
EAS0m706LgJH/Oj76e31ZK3k0V+QIXtftlyZzNPDUkk+13F2KTHrFVgPQQqCbOC7Rno71UPrC5kP
v2ESEI/PszpyFDFzWluTgnxkUT363z2j/UFGGA6aYLX9pzqBztAk3nJljsbqX40Vtp+k1vY48x45
XJRZyJeH9S2GwDOoZ9PVPm09HcKsGS+UR0ZdZce3y5eXugJadkjTEyF/Zqj5rC9fWpmjVFey5lMT
PaC9Wx4MFMIe93QaqEj5+7gDC2ntcM12peBlRHIj9l7jbnZJ3zsmaR5pBJ38iy71o3fa1wsQEzZl
TIbmZwshdtMAYzyCd0Gu39WfPdbKcF6Zi/eceWHlTJVnaHuasc6knfV37R0PD+ywPsmclJyQ5Mga
nWUL9Osr4My4wOcIsA+cP+mhD8c0GqtsiMs1rJ/eHSA3T//Dwix/0p1+bJS/iAtLFFXx6E3F/ysh
OSTcmmfuWle4s9Ye+nYL0WqL7YSjyh97yphX6N4aEJtNuoFI9yF+iDeW4C1PaLji7W42WW5Z1QZj
1xFdBvxaZacutv8Qse8FECLbDWZJr5yEfevldx4D1aTLa9BthEj/shzhlfC+PVh/dXMyS43PEl/l
oIN+Hg/+9qdEwIyPNdV8rYrcFM1QkMnZBLGpLYvp3dhhHbwS/PyLT36yWei6YPNxhr644fqvrBSn
Gmapu9rPH5vn9N8WFIv3pjBv3tdSQnYd9tDZFdE5hDEVTzoAZWxl+deX8keC+R24blXNU7BIisB1
wPh+zkbeL0rra1aYI0Tq8NONGwTd0R9NyAaCPVYq0NRxhMvxi7NOpyS+jpudGOj0FmBb+ZbnFXWm
gHntoqzG/n+QwM7JPSlFWMkNOxuDSHJjNPED37OcfDXN9ulfOjj7OXCMqj9ubBH9SP/SkMA9pciy
JJHS7iWq66TaxYH3W/eFXMAKPShLFOX9fP4jz9BRgdLhHJIyLdaa1E/WrerHgWBNHI4SEvpc7S9y
6s5+sXKirWyKtRpl0UljNV+GmxTM0lfuktlbqQOmHOYx+jvUyCqlCmMwTF+i4hiOAPvWohYTLrlX
JdA3dujAxMi5KqekT6qX6L46lmEncEfA5VudMtdqad5pvajfG3YyMB3bV5Y3e2AUqSH4UxA5wxhw
tZwkTFbJeN+x/Rx9v8hfKNnnV/sHN68Yadtpkcb3+w9lhGf0Jh9SCVP2KQyBtGnf1xsUixUT7M6q
8S+tz0UwM2MvBgCh0VU2WE6YRJqpm2uLraiuz2SWxISaO1AlgAc/hhzxApjYgUx9Sn0SMmVxUTXY
synADgoueMjEyZFMcOh7HX7vrvRtuT21ey0TZ/vAV+w3RHl3/6dEFamcCIfHRPyrlCf0yPpvHGp3
eestbQGa4ZoX3pPsB5HaGtUaIHpWDhFWb7lVwXXK97cb8MYa8JoOzqE4GQIkCWHb9PDEvP6ozWqs
WgAN5l8uswG/8yd3V2QZLqzYJKP4lKrollnFRaWQx2nkqzoMsfcO1Pljzk9wWdSikqKfaS86q/Tu
VHWa2Es/eLtE8/331PGdBxhiX74FIB57AkVWug3BZFl5oOHgFh64HYPP/wF/Yp9m9WDI3z8FkzpG
1Kta9TIZb0ipulVc5bM0lcy75fhuSgLtATNaxQ0jfTGwnEGiZ1xxfK8m/f8nAk+MCLkfxWyB/qmU
HiizrEMYQDgmd4fIIE9HUyKpQ5dV5pj7DUbRd/zAlfhwTYMfT5F+ioh2wgkJEoYeJojpE3SBWEKs
RQ3Wv/R0HYoY70YT9Aqowb6jqha+6kuQTKGzrIS+oMZG/XMYdjfPX9W12SuZLHrENWwFhtxuhaOR
AErbfeL4HOq67KIZ12CCO+8iz/KOmimRX1Vc0n8c15mN7QLZObEFo1jkXNDnkF8+/puVfKOmQNQr
2EveTnvH6y+BrJCFpaQadWqYM/e6tI9kQkjzuoqyAPyon0BtVfX9KslFH97gusLAD1ZoTSx6Uog4
mLNbxEmf87PRHkHnu9s2IDEV0vrREWJr+K1iZqRji1UTsU5E0uVMYt4PMBBE9bwJONvIbB1WJrQZ
7Ta16pR5W9tfbInO8Zn0ZLkBODOOvvJvDuanAWhBggweWly/WI29whHvEI625WPOr84qusfjOxwF
IWfrbJkXMp931+DWcJGQTE8PLCSGT+rfKYEe6gY7E6y3KCgScP2vvdzaFd3bnrmivGLsgcOe3mSc
WtTYe4Wdy0uGOGwagQx79SHBK/dswc3TuG9EPEzkek1swyLdbMvMx+JgeqiVRrS1GngxNSeQFlYi
tT8CqsVJA6xc2k6hwNCzfQz0Ptka6sBwpKlC1vSukGRpZ4MAAHjhu5cBhfnkaUXjPnU/ihuyuR+2
yog1up7vEdOGCNNMrYx4/RqtPtGN5pBznfPj0AaMa0A8rxXot5/prLqoRtdeeAJzN1DT6aIkEB8U
jvdoEaHnenI/EadYHorXtahVqyc4/7uxOecB2mKfM2z9+AZqscGQL5KRoVVET60oMfnanx/YqBzs
yZNM69u1m+KsDBbHW0T0EQmrNNdzMjyHPnn/t2rONoVz78gWPZPCxLusLOVms6BPHYhAkK2dJhNe
1J23EWFbUTqpHTi8fIC6HMBhq3+hp3Di2eJoI43YkyWOZdnvccZ2Hc/8qkZ0ue4iqxvsWQ3/BpN4
7zZTA4r208tLmo+zAQL4RNKfGkYEOSBlB3RVEMpH6stf9jlKIhfkOL7bjdE6YKvRbEKO9LE7Bgrn
0/C2hrH91WSsytSYyXD2sj5hMij8811LVMV5TjPd0ZzUAW+c7Oz1ENdIjgxXfxv4qHOnAkUHG5fL
au61JnRsP73Js5GTXwG49iUB4d1K6nZmqhAQ5bw/7wdtUdgnM1kQARAxX688EyhKZ34R1IGN8L8M
Jmh9jJOA8pue4DeyA08kLBGOtJ43dvDUgJXl8fYUq+eK/le+8ogdmWlpKM/zdjPseEk0n7kkq4qz
UxtPPXXPJuuQMJNBfMVPEp8yuXXluHVxifXB5BvKA1D0/a2hy1jFL1gRjbbW9ZEt71zDfYWvO1Nq
GetHs5I7AsJ+bXKCG5iRFDYsjsXNda0K7twnKwVDDMjcHoWAIy3S7F+lNKG9Y6iFFGrlSRgjHIJ8
RkhTq6Q43ZllBco0p6A4J7WIw40xbiYbJ/3/1emCjAE/1btNr4ayEGb7sknmx3IjyxAXHUq8FDkP
IrzQSytHhEowsOmJTdEQ/DUMJj1pTgDkvc345MM5HCUg5fnWhqIA1O4i6VOSKxO1B16EzHztDd/R
IGI8fsacambuKUGTC5syMHg2w2RMgqwyh1cU5pAbPGwz0jGEnlJ8ZIVKYhLNEU31gmt3Ic/utzLf
FAGeF+n+p+81A9urbcNK/TRXchPTB32cXrX09r1nCliY2bIGdB0wmYwTaPjHU9Obop8oP1NrfCaZ
qTncerEHI5aw9h5Vbeal9uZo7DfcpXiANBL8UCuvsisQ+PURfcSslswmplz332KKFKfqulUomFIM
OjcDYHvwF61C28f9SlIZOs3ixWVfp6HJ7/Bm9Nt7IY3tvKfN/TzyR+fYu3NhQPcpnCeqwgT0eFmJ
YotiKWoQ2DY4kiwA6jaOfCgR2JJdAUZ0+f64DNNQW8wb+/Gc3iLv7FstAI+T77VHLA9EbDx8jcdt
x4+hZ5oxFnI+ULdKCeTGRFXQvC7KPuvq9cpMuYkjW1CDRxiFtv3vpdJOJ8N57EebtCUyAPMrlAHK
EASkWF7y8gl80Xv7jmQpRFUh3IUUr6wGvBx5cuiQ8cIvfkp+3Xr4FfxaxMccqMHLcPuhhb0eKVSQ
qCWOnrIB27SaG38EfSr+Jhpqh79PYWOQcj9QXdrXO9chHmbdK8gYCatbuTjXd8P68AucNz1VF3PF
T0n4ml5Knb8kcrk5RWaBsHDM+w7LwHAiWy1D3MgsgTPWal8h6fTJiOFUoMRXk7f1/CY9bHwX2ieb
yE7yFYaowfj87xu37GylPhAlE/fKegr0r7/aSkoOrKaH/5MXKtUlDgJOl0pUnN1wS59v28d750h6
czIZmHTBk6BeQbcG8Qq61EJpyLx/A2fRlrNJXpDjuQ32lHIFsv8/OdRrqmpkZp9/sezDpHTEBp6H
uq82y/e1tPjAqZuLnFIuEJIJbUC1e8h3gt/9tE6kV7uUhCBEJNM5RNUHVtSfkTVG+Sr2jbEpfWpf
e5n0ACHhPejQ/8KNZyN9loos+YMC8aLAgKsyZ7B49Fw827a4leDoJoUAV7vJ2bNHOH/jT/nT73Ba
kyOlhgKgSRxRd4JDIq/a+rLsVtf148dlGeZvdHFeWFTz1I9n+DEQNCos+dW7X4vGgcw+n4isyYQ8
/+Pb46QNuhOHsJxyO7jLzuJr37AfXagQXrmKrJA9MJcpOYm5UjyI6pObRk98M1ODSwLFHUyVjhyY
+my2ANKhRlzT1/iP1oRyNLrSWF+zxp0s6/Hp000nGiJIKfbf8fIF/tUn4cmTfVgDujXQyPLF7UFF
wkJht+m6XC8Bqal7y6CBd17E9WJUpleHxAJhgGTCTYzICYrgkFMX3Ln2Skwc0/hdbBYbbmmdqNnb
sqOEzHoy2on/zIjN65/YUukVLn4YJSONUTIzToJmuT+2pQ25Av9uAOG9UXYN9U1H/1Wctq4a6RIW
UFgGTxl6A9ddtQCE1lJV2Zst9P5w5vXQm8K3WqRG9owog4bvNITdO9UNQjmo7MgniLlqReMSEHFP
31gl/Mun9wimVCumGj6S1mGDFWsJ4wTzFya84SfKboHH+WdsxdkIMY46cbEsfgjZoHIbCYaujPt3
5D2pnoM28XolmTCFOeqyhEm7DhjUhnvsoTOMw1dQ1vcPhrEam+6oamSIJpk267R77J/CMoqhkOix
kY5lBOms0m+/TG9rexQIMm4vTGDx1Trvaq+R7EFgxwQSZ533DekVwA8Us7ueT2QZyw+mwOLMTAof
wjGi9VsVba5sr9SzjwgTCnpZyrM0x0gvHdizM31LAav6wFDtGqew0bIu2gUq2GinIhKbTbUtnF2z
Pwb8uj6U/leuVnQ0z4sEyiI+LziAayRbZ28iajoPP4F2IKTfcHOvlAVRQiZR44NkXQCUI5l74TCQ
KddY5WuxTl0MYUKRZMOMN8ACpDhAcrrhsaTiS+DSQp/K+CL4bU4+HiGPP1CMonWG3UZDPz54fQpm
18h4QD7Yay94PUJXUdNiwuxdg2sCVhP3nmnp54dD/IhIdoCRK8hbz/xJzr15GIMsVShKjhDll4oO
4dznNAaih86COrxtTBTBSmAmnCgeWp27Dq0zFkPBJ0rOIm+ZCCb0zSH1FK/RsjPm2lsLfCUA5yiE
xR7gnIENgjRPmAhppt0c+Cnha89VikCHZWjPmbE/Ch67zM8HvIrmW9QPBGOY3QFKRnYAYLRzRORs
nGIq88O5SY0couXmaWLtY4XyC5CHn0kxSpcWueCOI9HKeU7oHctX5fIK6U/iyGET81DAtsfXw0DB
OLoKm6bbcv40nkep6f8R9uMj2eQ76EvU33LRJThgp1mKqxEzjd8oxxxxeAb/JxcAYBn21nRj8wGe
3lJXQ5zvMbkZZ5umXog3VLvJoNSp80qDN3dZfiZ/7OBAnpePEav1H1yEQM6q5GKEabv1kRd6MrqN
lR/aSeVqBSmlAo4Th/diGl45m7vdE4QSgzc4uaEDiJJvugBBp9lB1HJriPJnGttSdc6EtGeQdT3M
79ce8kewXyGFwPNlDS/90wolLoxv/2na5UrgE5ZIIraWpcFHDt75yasy6mHgq6Dx5zMKZ21f0oCF
Zugz5FrSZjRMrrTkqEzDzMgHlhWG3mjUHZGa4LPNj5Lh7AY+44NwugY8N/7tyyYF/71UZbtCEgq+
VXQW7t1nWxT06Yn25EZM9fjEuqEUcV5SHq4S8EsUv3WOBM3nMG7ecNafRzIR7KI0Y0gIKbGo+egl
0k4D7W5cyhCsiwpxQjPRFkrUoJH8Lc2imofolKSjQnR1p/NwbAsAifoWriSQl7JTkoVqBJ8a9Lqw
cYK7gocjrjQuVK6HbUr9RZFwKXQSA1iRHPGBM1l5pyd0TrX50LPrx//qIx8wb3N3nyR0WE73uKMl
aiSUeyqrVL3EeeYf7Qh1zwPaAR/RCO7PNKNORyOK6dzcKYkHZ4DkdlgQpAopNmofLA+4qiUVaGxn
POHvcbA0GLIAGsokQNKTj5Ip4LAkQS3WH8Lv3ESaZm0wYO11pKw8oWQ3YoFGkvijs0Ch58Yij7OA
drmuQCW+UD/n362DgXU4oQgcAQkoqvwiMU/z9I2BWQ0FNr3q3tGK+h88mYs3hvcBIsKXyUTpL8Dx
Sem87xRdl6mgJkR6Suc9blX92R+GHcwBrR3645j452j4NxIBdYnkGVrUpROT9klhqlgNh0iJB9ei
ejxusQ9gNYcIoQcWN+kHriQx9Y1UFgVwnLSUhQdyCV70wNGfGq9Fogslk460b2davIIGUPYGlAzF
trjqkyRwJEsCvQ0zRJMe9nMn+tAK87XmKQJfyNagb+CKfWlUuxUtvTWmHEA55MvXVASEPOUULBJW
tebiye3bbCyBESQlwNDJO8ZSLsJ3VzMs7BxSIE1RSh4O6JkOnpnAKOEln320QVrS5YdsWB7vHcB1
E593BIit2C1cMW7aHpdul/lRtk0AkKBUepwNLhpR8D8HmKbPY0pN1GwE7qCgF8gUd9O35+dUCNWv
Z6XTL/vsuHBojr7WWIVpgnNjyI9MyOvepqYR4VjN15yZjS84asGP9koPUs3HPvpEcgEQKlkEewEd
pls7MvWtdfneubEK+/B5QBXGBkYpCUmbQPRAQhrRLwFpEm8bMxuteCAhAcxNIkCyCa+tb//ji7QP
z7uEJ9Wja5uBvK4SrpHVyVgKXgMYx2z92vvhNMQg0NpA3AbonY0qkdTagEVU8iMMDxVlSAaCIr2W
G8SkQ7n5rC6OEzNe6d3eRPtOEQcGAspikrTZMGAHv8gI07CKwbhBjfCOAct8LGHUvxBsbx0SYI5B
swlrf7xd8Xn4Vh9j8USvBCGk+JL48sAZgvC5cMpogr6UHqFTV/Dj+xBiWCpdY2rjhVTeBPbc3XeU
p+sD0sWBgwFfhm9FXpjqc6tIrtQX1ts/BD/1EhVRLrxvg1sL0Mjo2QtOmueQgZgpJ3hi6sV0RPD7
U3y7TaPCxp5u3AQBtmAz0nHJZAOBi64fkkH5gsxIaIcSe2wZOVX6XCeHnzDHuQ9OZxVAI5BchJDI
1NqldZm2aT3P3ePyLUM7i10A4ew1B7NxTwDYhAeW2bE7jcioKel7odvdAvLiMPFIF9fUR+LPZPtl
ukTQN+zG/O+BNr9HVc2tJt9CTN7T5xCQ2PFOVW3Bj4srYAJwrFUSoDE8P3UB9kJjcohZWKWO1nxw
HnkFmFOzrDCZqCl05AkcG6WblvjbOJoxtRYs4l3nw5fJaRp/x/FGoxeo9phIJNXOoldvsapsMXH6
DdRg9/BmhS6BqHxGFV/RmrB4LUUM0I3jaV4wCEtIwapfVUQVSn/Q4wreM3OryVS9yz9WWPm9Ocu6
h8ZChxERnlHffNpGhSHKpxtimWLYWXiJrqK60/dD8HJvzhdJQfurYvujlOkSSov0RCBcg2CWPjxk
PW+KCeP+m6lB3bFyTvBsolwRDrcWep2wJnuD/uzmnjZmTUWNj/Zg+n3jierdJ68xWbA3PjAJ9ufd
DnzhCnS5hMzmzHbIDvba57WTS2RsWwCKfvBX+HcsiGjA07kOpt9c+Ma3zj/G3PdEdl1mdZIpC+K/
1b8b3AJHkRpZS2jnTdrURKqr9G7PcDxZuXusVUqDwi86CPCt7l0YLCaoMhM1DMsI/Mpug8gYkYG3
ObDxDQZaW2EyOgHN18kbaBv+/PesXyQ/avjxDElmtuMOnP2RQaLbRxgHNvHgcP+CjIAB/YOvxFJX
9dvXRenhISpUPT+6YYLkszLfM8oApnlFgmSjfM6OMWJjo8mByJeCuUl22X8aNM8tQMuFTS1PFWbX
rUzR0mK4SuR6nRVOuqCpi88bGHgQAFU6xNjJLIIHlOF1ZX2oF4foCHdU96qt1rs3YJS6Sr0vXAVw
7IrBMVknGycZAfqhapzIBU1YDCqktuB+t7goaFS1dMccVZzV0c2MJm/wzWYbMTmznWqUUyxJNwNX
tvPc2EjfJq6kJ1n32HLc1vk7AmvAk/+Su1WU5liQyYdrDg0ZBJ2uHVetGC7BXSefPnAFblDeOhZJ
8MmqrdI+xSEuUoQO/cf0RNSMwNSO7pWbvmQqt2eycIO9znh2Lf/ujOwDQZOVBaI/V9vOaWsJIO6d
NVpNBDtY30V+AjAPZvAMsG+UVVqDcE/lMgXWfpx/iqCdd+1611dWYd+YF/eheCzDfChM6i0FlUy2
BpbUGrhXo0YGNipKiE9PP0NiAG/16gbcdtqczpTzyb3v9Gao5g8Snvp/2ERdBRHYrD2216J4uNlS
XIF23Owi20Qx3dB1yqPuQMo+xzKDMTsIGQpIOLKN5Erknggq7/IZQzJVydLTH+UkE2T4IIvAyH6Y
D7tbRizRuWKCAeI5OGx+0RjLNMgK3SaBZFfIAuaBIs246fZNssOyEbERzWnE5u0q0fTeF6U+WyAx
PCC12kDXIFzoFCbaWhoZAhRMVGc/6PX/eGzRPY/M84NvyQhBkL7h2wZsCdCqrFDeSiJW7LhULQ0I
LUkLXpFH+q5zteXDbYJi2uXH+CzeMt1J1X0JYC2jYyf0W5A+ETqNKrCkziwSqrTVKiuQW+Q54gFc
Tb5l78pPXEeHSehPsCpn34eQyq+QMRWrP5DUKPj7qsjebr4MAgORQvfqmUOXxvFqKvdWIHZOhhS9
TA8LxJmkyz4Bi7XHD1+rI75Dwkvb+zb1+Kj2BKyay30OT8IdQEb6qIVn9T0As01lhs94gmfCH8nl
B2775IygaV7TB0aKY8adPNSV4OmCOenLI5LvHofC2eXQey9DqU5dfNcXqjU74RbLO7A2XQYOM3Zl
Zgm2X4GvEu7oriNppidynuWyTMcRNL2Du38rmu/mEien4W+MHy3G+bcjPt1dZE31mlI6j/uT1Ny0
3+xfJ9547Nf81xOgnYUwda6WkOqBhK64ezYAuXpb/tEZgekv35CNIkNZsD8BPvliKI+gD6S4Yt9P
h3UvVVycNBOJNDdsrACtq4WntVygYTB6I24I8jLeAJr4MEq8an1GkFDYkPn1yQ4+jFdd3PTB2qEE
UNZW/fuvuliLhrwC2uHWmlJT2mo+jQaAt9Q2fvAkPZujbVz39UL+04HJz055CZz98twAMVJRs7ps
rHZ5dL09+AAkRtsGgBSPvgdKk94+qIfzu54o+WflE3OQktVm/i6peH9rSm5WveQ7C5ePKl/QZznY
SQzldSOAkf/Finfjd3sLkdjq3KZnzLd4Po6WP0a3lqu+6sSq+WDcvq1WS+3xvmnd6ryVnEm0OdxI
0DS5teCqx4CtJ/fen0NUchb/eGf16cOzB2rqRu0SjkR6NQMRNJfbD6FxXEKAn8fUIb9qnyjJ5VIM
DzSkTj5UakteybFPqoVx8IonKwNkM+fhjCO/kQoVMVbtaOG4apip9q4g6U6dEVp2gUgKCRSwEDNl
W80/ksilSKh+MCHgw+VmiVd2sj1sYXQL+Lv8iMT7UWbMNGY78qKOJf+F/QuiXyuaIPPbLwtqvI8q
4bEe7HQOW/DAtjIAkA5qn0yR/qQn7AuykCPsp2tyTFFyj+cMSU9fhMwU6i9n6Y+7u4rn1u99B9p+
RLuyWLR+LxK3uOgaOYC1W2vEHlZfwwrPHz9skRmBWposH4YWbrajorQub++EIcVh3SydRMxODCW2
p7wLMAbGWrNTHiOfcDWwcimsB+oj66v0HvK0Il0ch+W0dTJ4yVRz+lRQs0dWyGurdw1dX+TgCYqi
6zSIuy58y9XwcGNGTNdjIlOtCoLWETM3wi5vpYXtQ7k8T1mbLuXVJ351KyQJnKkUq+poZr5rNM6R
sJqUHGaThNWX0ZqjiM6nRXDNZjgHoEofCA7Qp7pwgRdTdmppZ31GOmXDH43r8kPrCTCBT4qjDtPc
7tdPoBaAt/rDjBmWLH3iP8OlyaF9q8F5a7X6lBDlFWMyG5NfEx7P3LPj4ggr8NyfWw8H6cyyDf8G
YqjfqbOtcNkLXtjsxeO1pOQBbka5nl0IJaRZBDmK1KDQVpB9fRBrmxTbtGTT9fmmSMcutae3Rl39
4WpokKmO+LrT7J823P9X5kMXHQy+k8pEejk5izH6Q62U9JWUuosj5484ikpjCUU6r/R89B0zr6QP
cImGxY8qWWAcAY67RXOHP0a1zQDUVidueBll56g0cGrBjMX2fu/wFOyqLUKDZWgA0LbQ1P8BYxAl
yRKoAmsUEoDnAr2L8pb9kQqB89VIsoTJDwuMKJQ0rPnNgkZmlKyDf66qoUjUkRwiCOEF8y+LjNC8
NX/iCpbR5gVdt/h5u27xD6CgsnlrZTfvSrBI2IlgLc7oRA+0ofBjjojYHJLi3RvX/8gAhMvAP4g1
pdVy/Xi1FZJnQjc9cB48gphnXBAkGyDWg3JAMpHzYzz5Q3BHm715cdmluoxZWKkhnYl7at+7yGco
ShLosCGDRp53bm2+ucBGAmPTytix52O8bSeXsKHfis6UgtSxU9BLk8DDNzQBBhC3sH3gBX/zB5O7
SHRnqPgna7KsEr37fs+CCcSAXUutTWWHWXXHrkS0r9UwCBjOFB5t51XhRdMLYcW3i2m5z4vXDL2M
Vi+daQqxKqAhNgQPWacfqUsAT2SXuyjG5imaQZQQKmOnZmLGBjKz6CKMFBrV+Y7O1Ri2CFB4zV4r
XUg9r87ltUM/oxf2pgKtnw34fMBNVjNsR7W7PZtPvKkDrZ9cqc42auej38hgi1tPVfDwo5aEhmdw
F47JHgN3yznj5vwomMUa5VdigZ3acxVyfyTi3HwmsfnQYEjwZlyyvLRLE27GTIFX0erkxyUXK/xN
JEjBJS0k5mxCG8oVVr0jkPjNqKS0CjAbs/vHG66nGg0U8owBhk018znJhrW+sSrffDSUeOeBlKGw
1qnnyRxOW1eVHm14IG25Fj7Adbi+d/46oHPyLkxHCMfFo/KWStaBVIHOYD86g8nU7g+z/mpu537D
vHKoZ3VBpiiWVRrTeeedWaaDTcL0Gwkj2/QQDCGExy8GvH9xZc0ZWm84bfi8CUCECb8hqPrlLELD
9fV7wmm2L7thE4+lCaQ7eqdwQYbIEJKuVsDy6KcU8O0sqQDYNg2bvbPj7NUJGGjYTrNGPl6G+q+g
tlh6KF9wBI/wTkDLV/uht1hU2PYsa2+ygAuSaXmFeqrATCSW0ZcMDt4y7+ztopDPrwmvZbfObW8r
jvyiqedxBGXwUrlNTXG8xr1M3G2HjtMx4XWhVc+o9NIWn7DrCBwlR6lzb1MqZiv/Moz7v2537HY2
AgEglbAMisy4a6e/QzD4I14sAeOiEwilsTun2Akf7hTzAsP8HaMKKRsIUGzHOGIlVN8svKzP7A4s
BdZiAHKDQVg4GpmH4xWMk8NlEdr9rC+R5c3buG4JFsVXuSB0GHSpL2wrpoR2jQOqTWQlpRLMj2Kg
YkGrp4Mo/HG530k9luyQI6QGIyP3F9TykFooUuvSMrUF2iyl5+rYZqiXSiwKFDhY2x0hIWOVB+OX
l516/Ucg2O6DScPx0wngaUAgCpK6Hu3M11hpgkHyk41+1IdojUtDW3+KN9KU3nnN+ahmIcWwlBiN
Ge5CHNyrx+Phv9odOfZzQJiVuXoPhHxz/9lAamUCxPjDqZ91VgpocPi5kauhd/NgkhOmdqqqs/3j
tau0MxE7zsb2g4G7LQxSHNV+106NLUMogopWjYn5+riI09YfWCxTVrnTl6PK6mUp4zcy5z1oL6pS
jq6MkjjCOgLM3+wulLzwNLcuknsDcAGTCSglN16UN211tlWjzVqP2LoCvTZkDGFZXrgFk2xFXJlK
1OWEhhcSXb9vXCadU+wXS+cIR/0IOZ9yHhHoK5ROATF7dL0x4F4ScWLFJogu42/lyn2vHKCEZphv
o1i+Qekj8LBsrz74eks7oqEdGHzdm8XeSpm3CI8BJGNjaTdYLgSEAGLwYfNmkI42IxCBHYGFDxUF
BFVsgN5HUgLFT55iBT7u8+De/kzN0TXX65wdeW2wPh++/sIAl7e7WEa5AkivOTrgV0zCgB6LauNR
TWLpabj63xaupMB15ka9Lnzv9iqd6uwaCyzOP9p0+2DwjshedKyt7yuHcEyQOCmfD31jJVdK067P
Rv6GATrPOaynRpe6OMc08oQfHvVArWdi09n/DnFaI9z6gMYIEzNp+bBxw4PPQAJtzhLrPBhRk4MI
0Xi51kB0mDy/nP6+idyVgBsLhk7+2mlF2LZ+MC/AVi8C2BBz2qqi49IqWJOt4AUG9ei6fLVlovdT
h1/kzZtQzXHeU5t3qd3Pc2b+p3JWxxn+CQHTAcI95RX4YiQ98XgUwnU9zSTSvyBTXf2L+nkejOQt
+VriTO74+eJT3RxSn8NDgc5equDuHd0dPBwV1eirIKEztVtyFZxxxz8bwf98DHj89FMAsC5ASHTU
Y3D00pJ04WQ/1F1n3L6MoIPkZcHwNK1CfZiMX5i6FhyYI9vzrUcZjce7yg2njpkYuySJshD12406
t7WFLWr2fG5UQgwUemlVQoCqgLbRs3LlrNs2s44KFk7g/sib1WWyI8FnrUXpehWcUctSsO5Xn2pl
znzEZZ0Fh3ob7c/MABG6MHPFsWl2kDwE8PY1VaGcCePTB1c/ttWGRWWHmVEJJHI9m7v6BmrrPFr/
jN81ctmA8MIdcHnCHWNv59IETZnqnDLClhrXFuGFZnW0SyuEENtI00XBaaMSMSGFX8tjKYBxYAUB
3tScbZUQ4Xt+AzSnB1RkWTZd4ETK5knD4Xsz78z5cwmA+1oi7u4jp4JMX9tQ+nV1v0TI7943+h60
jSDxKQEhf2640cwEYP1CbG9x52GEFyNoXGqjqzmm88fOLMGaaHGNmHMs+sjx4Ovjv8MOxycodUwN
dY8QBmIkDttsjOThmqsaMd7a/0zesqx8W4YsGHT/L4TTBdR3vweXq8Q0WCd1xMBQ646Q/+RmlBwH
bH8Kut1h5k9NXXXYU1XtjA0crp1hBy9yS+j4MA8KQIsRYMb+gfg98XQW/PMkm+n2KegxKm8VU7XH
01njuaXsA84AvJCQX7M5ZTQ+uYhjm37z6f4hjTLT/3BimHc8ddSdXtd68CWD3OgoctnmSSATJ310
Gblu+nRFHgLEqhHGskjhuaBU1wXM9/rDxThJ0le/8jUW8YU0lvRmHDGf3utED2T+iOJ8/CE5F/nD
W5oPkta7a+r078ESgO6ha8faNnc5FiuO77yHDBhNeHWQCEwlSr3IlAQpY+fTSFw176aFtatkiGwA
oXTvUNI69qtYlfchQLQfEqMdud7eCDqIrfB4b9NiSsIifzxld/SymxZzzEREmBRtIUNPy0mVFTZ4
+Dmq4Luc5WIHaWCPfUBJnklk8vq6zpEDDbta+cYYZowEWJtQJirMpHozJgqxUoDym68f6RTjAyyq
DTMc3nwnlJZauqxdcBJpICEpctaZ+Pac4MySWzfaM+/MFQznjZDVOYqavrzQQGZL4Ggt7/nR8TpR
hYRtEiw8+686DLnKkbTiodMnrVIQSsIqFVK3RrQ4fhIVGjxTL8FrQkHaC+Tr/q1mOpIAk6D8+xDo
tyImvQ4X2S4cc3bn9x3Uy/Qq6RU/sBqjcMYdFEIY7CeytQuma3iKV8cwR3jsWyCKuQGSI6AtRG0w
kR5RUOjcH7haMTIouk/ABOnWgN14og2GQdLAttrEdTWRpxJbdlSXisDjmhZawY8HqkgeLy9kbD+f
nHsQ+xuPfRR8GAA0Jkg8dmZ12T6X6DMpjJC5fN4oZ6d7YNmkWdDjYFFP1oiN3yTGj+y7paYlvucy
UMI0q0E8Fo9tKGo6+tvXFk5SMiOgIDGSyc3ho+zpgi7gmmIfH7J5Ph2Erlsma859DFz0NjNU3Q0V
EIfco0u8h8MeLkkYbmrFzsFo149AvPBkVoGX15Lxt+De2DAPdDz0TN4nIRNoOtT8pdW7NnHjsEWV
BpFxgAhUcUgGKSLudPZ8zEzdBRDAd3uYifC2Wn/YRSGMK/xjE1zgFY9zd43BuYEhYA8ohC85/0qe
OXx3TnTzI2v0OqgFajxAdcD7JliVdDNn5QpDfQoNVMh8TVg5lh2cafqbpATshJ9pOWtIUO6TAnKE
Em3RV6ggOlUx/+Wsr/12kovaqS7A0MrmJ0eOeiPifj248qyWdjmDrvVRvDcKVA66EWbIV5RawOeY
h7FMPxyJ2TbzE2ItnDvBPpISXWpFcxtjYw8WSU0zeeLQtNyrCDAGvdJizes6mnO688TYYjjcnBhV
x9iz/m6/EJRtMw2ANE53ZII/686oEPursqTHImOBpAP/uiJg7+UM1ZwCJFhllg/MMBGIQ3DaJoin
hQcyGC692pF70IjUFu6NjIoxGfIsgx/LeN6noB9PuahkTzxUmQmffCdB+L2YlwfXL1FYJTX4NxU4
VP5kHPwdwXtQmZPLp+20Ze8IGu9Fo358v74HNf+X+Lmxdivz/SxCNNduEUPfy5TWXjxe6RmDakir
HO9fxEuz462S9acRP+wXlDf1PZlZ5/DEpwREd41+7QoYwjwq+EbqqHQn7Mu3zI/rtJ9ICphXLMBD
g39GBTm/miU6RS9/ZEj9RqKX2Q4NZV4Prr57LasX2yvbV+1KRWQOvruMYxJOWffYxmpGGLZOBYaW
8reUf+eEcdcimW8Q7/1ApcezoC4hDj7UPf32UqaL/u91F+niXPRf5hZ6LJVC4QLcD4szj8yCz9zq
05yRo13olfvzigBuMsbNyfhrNxVElwUYp50WBtDyBO9O5YvTYoFQUVyxBzJee3s629SC0EqrHDgM
q1qLRZx7o0x5FE+fG+gJuSMeQSRBGJwV4GYRcOSWQOjJOmHKaaILkUZZB3nib8h8CjFOSa/bd4hI
xe277V+ygcb89pIHZqkf5cShxlgOld9eA69jD76u7AH6+NhYXhBPWvoBXmW6UxPleWxPct/kfe9u
rIb8nFJAHhghc/hkvhKzYTEklhejTfHWedWY0ZWnrwZahFqQB98vQkstpXBDjfeA9ta2s+Yxvrvp
+4n3DVxY5jpWt1DOVlTXJVMkmN5hu333HIN8itn+rEqwW2bF6BEA6Cx9fCZNTC+e1r9y91do/fKI
73SeAtyl/uGDthRM3sAfzmEXFQCYUb+0cBedYUrWTQWKX91+Wwzg9H2rOT16VYeyvWcwPwwYVVG6
4iiSPxio9Mix/eXI0hjxiMfjwWVK1AbvvUDk7/RxrpxSkkKSECAI2b34N2fxtR11xUhtKiUw9bMd
GYRYR6FZGqNOe37C5R2k6L1/XGOVCPX+29jO8QAxLpFFYpp5h1DbVNNWCQbnR5CGejmrtc/xNTqx
aP2lT2Dm9JY+L0hRA+sYkGDCmyrDrPfz9YiJC0d7Gl2YwrRVhG6V3FvOe1eK48DBTknyulSljiAj
CSq1SeMB/4Ri6N9sZ+Iyku5toSmIKkbaLSJBmCT3WiJul4mkTMuc8QZTc/tMa+Jldm2X/lhofAwt
qEQ3jrGSqmbwWUhFEiQ08GBOI9bAY/oqI19RmWxBTI7qeyjAarOUhnKT/HTdxBfphEAsFrLGHAhs
D7808OuW9lqQGXmgnjCdVpL8YuarXl9cgoNIjddzlOM8IuzjHP42+bCk5nyohE0hWHiVWgj2+zOS
43QvQbbY3bbEWk97viau6jRo7fQoAQrQL9/TeBpTPHeLOSCAtZmFuZecD+35yv5lxjU9kEDvOnoN
+d5R9Z1AFWM732rH7fkcUwoRodTFe0XjLIIlMX1Hd/aE+gOnYZoA+q6CQ3+t+MOeoBvOEO5PZkg6
OHM00FhKm63+BQNsJFz/Y/4kIbZACh1QItmhQB4r+aIwWY6Gi5ZdpIrq98p/zrcc3ALGdFGqPsTW
w9qck3mDk/DRWyMXVbh19pwlFYjllqHR1COQ91VrlfixH+s6Op65QAE7GxAlj5J9O2t4nUmBSZ9H
Q9/DwEox2pd5LeZ8HxYQrRrSGqZvlAELvXG6AupfE+bwLbi27sbLDFRtEQyiVsR4o3nHmceSFPYn
Z1D/DtPNsvBE+1DWmW/5riKmoTflVjVc7IrXVa/Vy6KR0Uisx8oCBOpiiaUiodNWpyLXHcTgI5nZ
a6Z4Kmvshshry+Xt1Azjd9vR2w2JGfY678ipeeJsJefKg2a5bRivyR94QPuvZhEIrVUJ+T+L8Row
gSAZzjHcNurGxOZGGKqkkPvomNkHmsrEw5aETQ5BR33yLfXTwxZOMLGoqakzlw6FYdAMMTxbj8hR
HxHutVIIOuEcfCHvBuyU7nkDW75Gn4lveQkNd/3Febk8sfKTtXYCayKFjuFcLDFL20uC+9Eubywe
rCwRGdPiV8DeV7/zJhENgzwc6N7lkd4BoXXEg8mMZ9lY17xDrRKpSx5GiYfpRLteAFg2taTJ+V7l
Yra6BFVdQvvtUF8G/vUISlUFr0a9IYD09Gq3q8yPC+phpytJKY4ihpOVITg68xvXkREvwxIZXgZk
THYN7VbtuyANNIecG8ez+EVTWjqlVhQolDJsWQqS5mG5SkUaptRujmEksHQru5cfuy6qR3mUmnVx
4++ODTBcDJ9OLPtJ5FGB9tCVauKSwEqJKjTW43yiO/JDeQ9q9JgeR0qr9ufXkTxOKZY6dqc+mV0j
bWQgYau62QjiAulfOh45WgyPhihpMe6FKlQigA/iPw7xVB8cO17yDzalcai4HpwUsJXfzXiFiYSf
dlc967hQqBexuvVF9qyM6J4C0OJ+u8JYwRPZOR5sjgvGmfzuu1pV+z1voZyXjN4NrWigmr6uaRoM
cpicpTqMHn5ypBh79U1cXxU1zLxQy+SFxAl98btqZv5bD6sRHMG+mZPYx3/XLaBBRzNQvbbhzkrk
+N3rOE/tkyH3t6e444qDl8O/wMXHzyo44yrWUe254TkHchkrwNXJol8blghWmVZMS/lxLD30zU6X
d+sPZkwpU6FUg1+T2XRzbDON7jhrMDvvF8J5ySVb+gDWtw0bOEIeLu7nJHqAhEQVW6MFZZuBnBWe
3FzpQ+Y2Ala8o+KhMY0yif2gJAd2ZsjQBVH06ym5ibtl4jeV11Zs47I2QIPQcJzsYxruDQpmoYHW
78z7UXYOweehdhBZbDB7xVS7EVvnMeeWLGr92Ia2bPmxnD2ld3SZvgsQFMHjAg/QFJesIobmP3K4
UkTRR5PM2dIhZAMAds3vZEzN91mM7X/ytbUmhISDJN7YVawvBIgU27vjONolzoUuL6+aQz3qdzld
q7XIvsFZkFfY/q8cw3nS/Pks6Hk3LmvhB7oRjWs3oIpQtwI0htBFB1nOjm0YxKU84x5fJ+QxD/YX
ZR7AeW9aHnqqhcwcClwcAHnPqDWjPC7DcqYMmfjjjgbSVrat7dqybhsGUDLysb4fw/XITU2ceeMA
8Pw8J/FmvqPOtLVjwLLvCNxz9TywuUvQZZOmZ6yFrbUxOotGv6nqeVS4pi0WRVb1+Os2bI4REBBK
PRWjB8rmC/sifHVDR6eJm+abuQj5/qnEn5fCZCn4D3Gcwu1U30mnv62+pf7yZgwwS7oYX6FgkmgJ
cvis3Hsec4tGpZo3TL+SNV+T/1avQXsypsz1+rwYEWi5KdJLdmBd608/cAkbOhGA70kCXmqYF/qp
aBhSdfQgTkmRym0Yodh2fcodObziLiayq0Sq4UmQAU1pAmuMwX+h7G6F/YXST13K1IR+5DKxaHsd
Os4XrI5STVWWOOsDte/nnDzUuIWzcLIwHWfxp0gXINXlhLOwLZnHEvanuFGz+da0BItyS2yoOS/p
Cw/Ydpz1c3aWyg7JV95VB+fmgtNiHW+WkWx4e04a4jbLAvO4nnDITho4TXSeQmNxY86GWqM26eg3
3PEePwBV0SltdLFUDUjA7WqXWBCiv++2k2g3F8W+EXTEL/+RU/F/sK97IvL3keVM08mJN9GigiDW
DeOSJ+qxswuT8GWT58Va26g6dL+Fo2ETU/QMZjswc5spzSb24kU5DFhchStAIJ1i1FihHWRprnQp
jEwvrbPy4nEfV8Bs4Pu0rhkmWKhXgg+DRF68CMB37+dna58sa3WTyhXmZqn8acjuqHPX2jk9mMvk
H6npy4KKnO8xCJ7jvWRv+whfcj5MrAH4HOhNXhkRKO/UPd/l77THLU3uVa4pq2zJVbyCkxJThiJe
7iYDOWFYwcgEk5xQwz2MNvwGC/0BuA9jO8NXHLK0La9UqSJf//MVECt7WtPsNetTvZVs9xMtkI+x
ThsvhMZa13meMr+FVAmyHJRJMrMZAx69Vg0Z5zPggHIcKeDc4AcSlWXGWnwpR604FSYy7Mm5s6RV
5Bq7U7sbPw28No9YUZ2yopw8eXS1ivBr+AsNhUcYzV2488DhSD/r4Cvyji+xTuTMK2Q5z31AwY77
gnfDmuR7N+qGXYmCIf0bvh3JB7uZXlQ+bGj6RhTFh7/a3xSBxqMBwu7Vvk4E9MRjJ8l1bm/cH/hc
W0lDrGXwYzGNczuEMnOQp1kS6iQfcae7OWbtmi7A7ouIde4aFgVMEcl3S5U3IrQKRSyFuyr4yti0
USzjMvZCIzpV/dIp1GxmryGxgvU0TrndagynXlR5Fuzpmv5rIzvQXUJMn+3odEajhK8tq/iwq6ND
hRAoPgXg75leeSSQ+OaQ8N4JJHfGr/hr1T9DGQYArPmcS8IiUDYXCO7TPC3yU2dtyA4Km1qtshW1
vJeGr1VaFTkmUddyiHfcKzs1dIbfAxNrdOESjPS/luCJjZ7PKZ34L43J9jwMjEczOlwZBU9+465g
QAcS+Ckwyhy1Tm4wkxNX/KyPVUQGC3fkT2aqWe72iTi5X7y9bSL9G9RUWO14BeVu0OsjOen0EcMa
sjnSSqjfi8f3IVI5Gf8urWBxzQBTP3vkM9Naoe+i/AlXHLZpapyojU3nHl7yMb0X96XGc9Ifct1n
SzPdfYRGqhu6dePJ/nn4VIYFeSrghR/4jXSgHjwY0L6A/v24yfRE6m+taETbtmeQm7pzowgE3b+y
Cz+xBHqxGKE/0qWcy2SpiKM3iCfHQjwzKEzka9RyJOeqOjv6T28v26zYslRjOEYZD/09gsDRqbTl
3mWg6W5NVMd/WquG/xRd8ch1hpaFggTzamBA1wfv39ceaW4Fh0RhLcGAfsorLPe+0bY4c3r5sN25
wrruUEdLOzxAItRbpzbM54doFvRnAnSjng7iBa8QYq16yYu1P4eOuIXobluindVLPTQI9nLeGIcm
Nl1Xq3o4OL5TLzwI8WrHcKM4Meuvo9T8OfG77ky8QOwwUITbBknO/xrYT6fJkovdx6JuCJ/5zl5/
ER4xaNAyGzMYuUnqeWB3YAIH9UpZzS7Lo02FsSOOhsjNWJKsyj6WVCDQDV3yQanMo4y5GZ6/2q90
SOFjy3yFZoPVGupvIvbf0dnvungo7U+2d0c0LQble3vQECeOo83lCFpo0RUf4wbyp/pCF2Mk6xt9
r5oOcCmZpkLzGvW92uU2w/3l6HsHfOPv857wY9ZJ0jCHNmEQQTlU1QoLsea0UywKXT/kRY+rYuly
1BDF0AF3xMKXVdy5j0c6CH1XF5DO8IV07afbR/pzmBcWk9Vw7IB1v8MTkpleuQM+isQXhSfWTPxM
vpuJ3ypTjtBsIWpDEC3HXqMLS+Ye2PCE2nIA6kwKQN+yzsOZYHxeQ6x8n2gb7oKE8+M8AuSerjTG
egj+tnzW+IhaYY3DWUeoie7zrb1nOsgjYizTf9f77TUozuMvZES/cM3krkqsrPkHenutgT80oA6J
zdMmMiAU/1PCSJk91Y0M5XwqnoQ6b5Tnmsqp7kJsZ/14kHPeSfT5jiB3c7Gr8WXUdr8Dluqt0jpK
NAjxz6Rlsf5lRTq9yE7P/gjR7h+n8E9o8AkiY7aFr5/w+1Ysu0jVkUhoobJyVIMImn7NMQNRVS+y
7pKNKzwCdt60Fb9CvYJKdb/Z5NreA9nOLJ2r9htdymRiJ754sBK14OTFoy0EOLBQW4Vj3vZD+uMt
8H2ND4e+qIgrlUIvLnqvUVaKGMj9yJDINmKWJKkGwTkHlL2xz6ub5K1UqGFm90kKinbWsIlQo/Fc
aiYnExTB9woUGs7jeGIYX5cGqDh7mPYmK1+FoOSwHPb2JrOU0aWZJ24pBe/j1zpC2WfyTnt+22ot
FUsr3WduFBbfVAXBE/Yb125LNs7HTK0obqg86AQSllICb6hZKa5KAhjrmYKydiUTLp7qPUkml/A8
vSWPBh+J4odIkczXZ1rZPwSA2T2SZPj2+NnmHH4WUC0L/kt29waFt1NRpipq7bKADLgKxjLbcguT
18w0t4P5Ry4xQOUjk7E1326OwHgqi1dirc9LjtdP9zJtK3lYWrqPmlB6uGEJHFynWATzzLcXg7PS
1r8orahNQWI6r4QxbweWiCRDmQ/QkX1sbgSc5Izu3COeab4uryMmWcXYV32u+1ss6MmsMNQ/LXyv
Vi9Wa19uhyFSjGuc9gj9hC2BNecxmIdZflhmBILkS7TdCJs8si4bKXQhw6B3Hb615KUPGlQXw4b6
nf8TVens0nnB2GLEeBOL5+VF1rJaN8GMl+nOYxJH/SDdU+1hm5acJylbBx3LHFD68y8z0pOzArrW
Bmb+AgTfdfVwJqfBUMVaXLV2CAAuQkOVWjeYUiQGgUEMpAEjikOIGNIErtzCtupqrQt1j8fO9aoi
qP4plxEbo1jD6JDKUvWvfLGPnK74d0OoDy3TCYu9sICdxXe1gAdbqttPM1SkhLR1YZN8ORsv40PT
rgOSPObuJBKmgc/B1zG848WBglRQhNxYATgcrITF4h47lve60mZoNvyn1BXUH2SM+EEA91bkq4Dj
lQG1jNthV/ghki9wk5Dpk5dLmgs/Kxma2NpUgBUiRTo9R5djD8SeeO5P65WQwSkptyRImBkGAa+k
b3q8/yk0K4snMFNGUG+ERKRGJf8DH3lGpiZcvJD7f4B1FW/wEdOwXNLNLvMI94wiSHqsjkBNaYeL
EdymLG44rbMYNG4MJbaOCpc3U+OdIuWvEZzuYJZ3C1oI6ya7KwR/CtYqdvlNtNsUrxYD1sHHfZ6q
PeKREf18ewNsRxS7LymsGdBx1ofeM7rWkwrZL1roZa3R3opmCJl337/EITl2NTqsYVw2nF5qVYVY
OB4VVUcs7NONr3nYMqg6k+CDBEfCgMNQFnPjxEKFtcDBBynvx8yD/8QT4eJDJjwocu6r4qWQRO1p
thT0lCV79ozZlRb9RlGRCdN3HeSr3HJ5ax9dTaWf7aQay4H3r0GkkJUL1RANbLy2wY6nkWy3rf4W
jOWV4IYGGJhwKOE6EZuV+sO8JgxxaxmjI2YcsusPKjQN12t90RK/6Zxq8srbBiKr3gzGRQSsiJ6n
K0kmVqalMrbC5Hs55bbdCV3dxmlA89mQqU9oZk98xAuk4JqnzH4OQtwUlZVUEjkxkig/eo0BTXII
fxzFje1VAU2zLwPI2/LaGtBtx75tpxC7O9MPai+5Hm3ZRPBfVv2+GUs/V4sRByoZF8r2kq+wErNz
frPqE9sokRq81iqYVRCpQQ/N8L/6PC02aF6D8JRyep5ypskG4DdhfiGjCynvkpTUqOjzkfX0OZ5M
PMZO+RFDfKZ8xaoY45xiRkVwho3m/BYFM0G9zaDTdUaUwyUXRV/VRwcGvVrMyR/RiZB2cqq3PTm2
ZshyMlZFHKIrRFe43DkFebRr8Hsp6uvYE82KUNotbuDrZm7WggwCfyV5taVUgtBL0tU3S4+o6gJY
CSY74owxagkrQhpzdhCSXg4AzJlpygsVI6U8lHBVjNLAllRQv+nmDA98dSpd5/zhPtgxXlStE7i7
Iqu/uuqvfykt2/gqE1byLC84HihOqvH91eDucfLeAmQtUpIW1M6sc2UVaF6biojfcxlk5mSaup1c
bZaYfOi1lMc9UsZO4XhDyZelS1uA8Rzmq2z713b/I/JQcuGCImhkSwPGVD4jhjemVe7eoaDbYR+b
mE7WHb0brHkdwuLxBFIMW9hweSPl6p+K6hITIj7Q6/p/J6qqgPe8pNONEx6iYZqFzxLZ5MptL4Ww
+8KS5h43JUYJQmStTxbNpU9mnRR9AF3NJqg210KBe0WK5Ki4vL9e0ip18hEV5L7H+7f6vNud/Nwg
7y9w7gzfRfLQNLUvtoeYrsMbHYJQso8vbSkaDeaAMA4zq/ipQz8SX5qaC4T3H3cYIusO1SRdjlFz
ccM0Ym4TOs4kmeo3VFGB1NS+XHFBBtHF+qB8F7ZlI/mV04BZpXef2+11V8yKMt8e7oqYtVQExxo6
MgMhgdhGR/yHa44ZYj748zBvUlHMgYuDyNMDlyig8FGsVIvqLKWQxtH++QiBTDOtLdL/0eOYKG+O
WoIPgeeHJj8sk6bE/jvbsQG+HecNT3HB1Z5hPP93lF7sj1ZfWa13KByDDD6D03ppkxrjXWIr92Jd
CmzvlPx3ByUpcMvamem7VFAgz0lB6lS3C9U1r3rHRuLEM8pFt9QQeqXqzO3bGyroAGKnG1qh0n77
SvA+9soRFsSFh0ZnQaB2RH08C8V1SAANaJJo5aT+itc7Xh20kcEinq/lh6lV4MxhpixCo9ItJ1jK
1feY+JD4CgB4HXjqyjouU+fqxxQ0kb+jJajnZ9wbH9dAwdzEBU35GSXcP0Dj4JwSqk9joh8YTGC7
p9Wotr6cEX5+mCNEDPs8x/c/UHq5CQVzpWuf6nUj7Ax1DMzRHiufaiCf0LmRCaQe/HaI+4FD2Ail
cbmghW2ttzN93Cz9w0RomQbdIgpDMSWHKir2GBdF/om5VtTU4Uaj+X/3u1w3t6baKRn9eXSypnSz
U8FiFiWa6Tu+Iiu7k7ZjZratRPwGkRv+mP4t4NrLzfijdXWBt5JC9+KfOAqrt6lX74Moml3efHnK
J9n1t9HOr4HVV8rlK+oQe6Pc8Rgw/CWpuzxWzwknovvoVdD6DxMwW1BlvCZIfbpW7lPy79kC4kTD
ZhKwcqZ93HLT+7eHX/msWK9LdVoy1c1aCKP+mARuu2D0XReipWaFbZVSRFeH8O0DQCGxyR0ujPOw
Z+xk0Cysj0VKWxITF0ck8Hs52oifriqEzm/8E1EO8eaxH4//BkssvE0ox5adaFKngiF0A2X9lNZp
N4suaLEQMTGsrajRcwCoQYz/IbBkUku5pi1FFJ7AeQKNZQlGUU1HgpjC/nMadoeLt8nhE65EXtfs
WFZHUiQ2hqcVsYTTiZp00t8DDbidHaMSC5MOjqmHi+ppt/Qy/Om2yGl6oiGUxOlag7IFdjWfdzcL
GHi3aDkV1u0mdL1AN8CY5/e/s0OrYz7GnCpugzKvarFrXxcKxwC7OI/dyQ46Fx7ORL3PH4wORYJl
w2Zzv2XBGno64gQGEvNE68iQCWKAvRYP6/4rCIDByJx4yHj4hhLVZbt7KzVGoYyV4B+ETVJJ+Teb
sOiIRxDm4iKRGmnxQWg9pnBsKaC2Zq+QheL+guIsoEZzpCYDu4U9AvTYchUdCnxl9jdp8k62+e04
g0TCw4mM3+V2eGjjwVSyVgnErCl0nxFO7dmfbZSf5EYeez5nrXCmBPspK/o0ZUDGlxHCTcN5dN79
/lyxNfML5mPJixDqYfOP17F9pzxZbr/amAl2SGFSy1iYYdktjXPjDlTrINrzx+EjqhWAi4dZ9K5o
Rbn+huFURLiyEb0sZF6gf8rkK5l4hgHZkgjbD+s6oqibAh+oknA5gYBiuI4C//PlUb5xqDH6rxT7
RV9o1fIKjJ0uDYPHNBXttEHOqpRbs9KfJJSciwOvRvupJUmiwORg5xanK6OgTxm5eOHcZ7SM5JrH
6IClHwnec/gWKK2UGypux/W4W7jn/88eE6h544jyvQXUjaAYx3Gwdlt5imgoEfrHdHVAkW/0AMV3
qV3hyu/JuVbV9JLQH8z9hUmY46bvvOpPMBDGOW1Q50l1Kw3cMabpO350sc6Ysk1XYiXpLA9dbXRJ
6/T2fXeM9CAAeVsWy16odz5Xcgp8berHrAtAxr+VxMhqe4HXYHrPwbebHBAwlAQakiq/OJtTnm/r
S6RgQTOE5kp2R69ohu3oylKywv/ZLOb1Iq+B2qFMBZ/fnjM/DJBzw21yRqxvi3VRY4etQDlom7fa
cXyCpiT7WZiHKxZhmqNNBs7dFsuGoiHuy8BXo5flY1tPGYCVA/pRmZ41i9u1zanTUtRIHHrYu0RF
4kIGHdaUaxvPMCIHYQ50rty9mQMR84Gxx6YIQuZV76H8Cfx0Egzbi6xG1PQnr4iM9dHPjobJh9Yp
Ml8rwKFeilKHhyg85dBWoRYHY/+c7XaG3o7kHGmlecWe8UdwrARO4CeJcafKu2uta4raKhz8wd8M
sLvM17e9iVMHjfNKX6iu2Qq6bVbEWn/IwGvW0SVNmXU2ONfZlxUKr3pRbGS6i4c8hIsAsttyLO2e
EOVhXD3nMheX7A3bbA7w9aoVNdCS/tAJvvqZimuACSZIYHihRxmH38w30hr7w3umGwa704/65rk5
BfZbv1HxQtGgbYWybZnqzcJ5V4+rgzQct2F1bqBGGmAOcIfTLbLemk+u7jkcsOQkJ9NK96pstB+x
jjBSPU0sWq9h7tbrQscrJGHcZkfDy8UqTBCcKu4XHDEd7sk80dD41oBq7amASzTvDcKLS8CKxMaX
4YhdoraKSO+VqTHuQt/wC77aePSvODaRdwMJFcymqqYw4nXXOhmRM54d6WiNyftmOMcyeot6TpWF
NX3wcV1lmGurPEw5dfS6H7owdUeTwsUya3ha2L1+6sJhGdd+ujKzcXx72voo28v8KLcaX0cBhmUW
RnFwQ17cEvYOtTS0HHJcM1W0VLz5BJEvOT1rX2j7+cqSl+uOmZ4JZTXuch8laTGb5sYhKj9xJFQU
wZNZ+XvkeHKXtvCC0ZpIUfPXoGNYPxKCQr9cT44M8EI41IkwLALZ6OkT1jTYrfKFdAHdxC2AfrPH
FbXQ4qMSncvnKdun0peEq4MxmFR5MubRsu+kpUX+Gub3xh/sMi0CU0YeqOt1Zyl3jcVm7jfg3Db9
+Pl3RAy0bdtDzeryPP6yszIoJ3AVPKC181XX5k5wEtovqchzP8BbPYD0E6YMbIc8RXDbPtcylK9y
vm9G3H0Sc9v33EKCD8tidc17l6FfOsbVsttx+aUiIVjDPWgrKVvCW0jmLSmUNF5CHlHvgM4L7iWk
dgZdTG8rKadG1Vp7+E/58FH8Tv7etqmywkLw7A1Ry10yTgPr+wtmk49PWGHLSLRdZq7GUimagnTt
H17cMdOricGKJmHRpcZxbvsz1yVC2RyrDh/2k0wm+cd1eSc/20+bkkkNgFc/J5lzIbF+1blNNHBr
rfzTX8pHJDrPqzAEUePLtpMgNIhGv4qIJIJNEOmilKkZK3EZTDlPSfk6B7hRsb4wGiCcNm8uEUQT
n6i9rmcKSDBJwYf/k/l3yE7WO05UAoresYMKiCzXkrZnGhUsq1LMavHK7+dWlMyqQ3PEmAPf9Yfb
dUDpk1zhiPIdbYpYQtW3upww6l2QLfOp1/aU3onnrQbA0wUt5I+l7YWto9HYyA8wL87EZb+g+wAa
gjBul7psGI9viiGH7DvZZSKd34ZkMfmtEf8a9TfbLWocF1thDEIT8jX2kP6HAD9glgboBY9RYFYH
uoaVgCRjIJdp08B4VK2kOi6NZGSOY8MyTQwLjPp8/cvkO5+lAzHoAJ4qd9npAXEmXZtuzUPynbUS
nkffksmCDtl/5yTJxGhNG7OQn487v7++8deudPJxETQHOoxf96rMRZv/alo5bqfge8dHeGsMSBtq
84LDUdIJw0D0hp23zpsM8Su3ZOdrpR1uvfKzdS8cJNmJaSWVWqa8lcCZu+K8h9K0TW+3o7arTvUa
r/5r/tnXyyqDeJkbOr5+vauUc6+wgR5R/6HcK78nmdjRzjrTGKIPxi3MHX7fKowm4OXgsuUTM+Nd
TC7kUed+aybaKC+DM0EZl4mk1+LPQxUEGxHLfoBCjbd5jkT74UT67WLD/AD/ij8MAVgO++GR9fFt
lcatKo4VoDhX0jr6bXCzVR5Y6SN1AP/X0WJGR5DC41dgo2QYxGGsXA4K3MPNsE/FOnzgzcJGovg0
S5UjViVOhlA3mX5JjMW9Q+aGsGJuYsCM9jl5J9vETow3Kv1v26suZFuVn+2bbKX21qTlPucqGupU
4jW4qTd6LSY7Br3ULQNuQrZ+v0LckeJSYIgm7S+9eAGBYc1k0B5LISAq2kpy+cFy2n3JYO23z0eh
r9oCFv+NStawy+q29b9VKkV4BYQNys8hFqjH+trc15ti+fjGFjJhCQjJXzNJ5IlGbmqZ1RZ+QWVA
efIW8l/FCsOJISakmD2sP9jSKq+SxGZ+3sSEODcyP2Gr2uxNF5jblGC76w3B2e++8z++mh68nkTa
XnPKZezYyyYQDcAYB6zzy/Sl9vIaFc8KWa8iWj3lcoy55/I9cjlnpvKr+vCuAnGBw8xp98/Jvg08
LMzhwCy6OG6J5irmU15qB2G2Dsst3f3mpPyiaotaP4Rd+x7DUIM+z/FAWBJ4AA45GwRp5YpjI4bi
rBBdVVLzYGnRLrckiw3tbu4pzdSbeow05iLDifb0PIlG5yMSPypZBV1qS7h/BeZqXTSGs3ETU6m/
4MZCwtlsAjhlQhs3wM66epOyopmEdQ/0Pqj2uEZEt8wGgpRU8DnwUjcQSWNMsyZPyyexs9YN+gLL
PUb1die0WpVi9yW6yaaRYpeP/Q6WE8kQEyunjUb9YAfvAlJuhubKVGh3Q9UjQq1XULntNJvw9a35
PYOUMt8ad6xTH+x0XLXlydzXy8KWLZsgg2C+rS6XUECGYrUUWsF0p4UaHoJMYloO1o4uYGq3ftAY
KSJeH72BePYzKWLBYqMwL3tCXP7GqywkbJ1kU/I0biNFkhEf77M51CRZr/U+hPDoZOX9xAXpfyre
4/Uf6DqBhMFcFFZRqQIxZc9uWJse+nfdpQLVTnPcFrNtgE1kqC4KG/Ceyjdqokv7SUlyn+pest+A
qmX961hBcytTrrSqM/qFzuMKhJg1Avb2UChG8JEOCEZLFiQt8VH9gprZeyKCQ99H1QCLBgaa3t7O
KVjqufkAlWeeUDANuWLnXN2oYTIeWXtRgenmZW0rKENAkD+pnnitvinEteXoF2rapcK20MzB4Iqw
F1RQs4/5tLJglLjim7CTLUmRVJtAwMDFITvgsKcIQAgBYTxouWGvdFXajCyYPEzs7i6rDbiy0Qdg
5km7AUVSw9vlugPxN1db0QMSI0S65DBQU1pwDB4M1PC1J/SioU1Cxtm6JtTbcGSFdTWcosbH0yLL
610FpDEXX7gt/0IcRa0NZDp2giPpPSplgy4NNMZe8r6K59xYHJ5+yVWtKxzmVW0lGI96AogLpxHX
x4XuozM2vYIfp33uLyl2HFpmIbQuI6RDjJxwNm0GwZuZNr2znDORVnCtR8UeHhM3u9T9YHyt3amB
jrzM3gkD99S5MgOfndbVyfmmzhNsTzb+8NNWJLbxVKZ1vUtBa/G+0bWibRVMtx6uQxEkcvNQWm6F
2+Be/b0LxOGbAiw/Xmzd/2xu4Kq/Qow8ilXaV6kKIbi7z+xanmbhCrizkMK5n6MwT21JDzq9GYco
xW/Lf1BJpsQQQZlNFkwNBcCXHB/JpEiWuCJMEOU+jDDw2y8Q4yjeDRZPAooegWmxEimh5ndsxVZo
mw7cHdh1Tt8otiJ6YxlmG4kCKa3EsqSUUzxqVGRF+SRzTuC4nbKt9KZvFNAkgNCv/bMxcGzq+5pj
gkdFE4sbyY1xKx77s/BIYw6VNoFreJ/SmjCUKBsVLUy/Kk3QH8bIOSSP8RgLESG9ITofeXlU8RNg
YL8D0sAEOirABBtwtvAyQLtgwTFGREVA4Ve/ysv1ktonmHdlPoRI0oNqddjz9INpCw0NO1XaYTvY
5wAL7TBNSCNvIUIhielNoL3Oy+Gqyz6OuyKLo0KvcLAZxC1rGiXFwGwyEJgBFBnQ2OFFhDgdRSOs
s+ltkYOXqXey555WDa9euh2FpESOk3t1mDZagRi1xa+SVqnaCSTWT5ohpIYA5caH8eIpdGUvht62
ctRSlBUvHpKvjeY9l6WvvWE0Ij3B6V+J+Z6Li3MsTTulSD4jwGCBvcJmxTxRomGMYulm3mF6vQzU
VHh9POp7133T7DF+WHmCYemke9AiW4GvtjNGvzBjp/D4NaylvVGO0Dtu/KleU9RsdCKiZRuT6ytE
DaQnJu56yHEVvfAkk4xoaWmIzea426FzQUxH4pA0MXyoYTUuGQ9p83EN7MIVLKIP8fIJL24Y+5lE
NOrDBJTPxYJV3BwK5SHa23nbIjzHmUiQ9yp4lvX2C0ewVY/Ny178dQqZ1xASQUb1wW6BrW7jVTnf
TE7DcTlvubI57JsLzKM5oWvFXl0IYp4cHYBWxRAnStGfXQKqyjyN4H/npJUubbWMfUpEY2s4uXfC
Q0OAoYQwnKmLQQyijvV3EQow3oGJobggFmBxcY/bhXuR6ZBsmIGduww4Bac1Zmuwy4e3x8oyoE8K
5jmy9MJt/0j7Tj2YqDLsma5/KZATo7H/gQXRCUJz4xnhHfSIlf7bPcH3BDGNzEZqN+9bx6HL0Pch
bEvwAMRVDGVfnjQd7LHpYgT5Cw8QK4PV2YwACT69Zh8rJ0+WMUJoqKjnSGgkXG+z/dJSmK89ZZi/
7buA5S8lRcvPhYB+uaIuLBTHxuT1QEYzZKinmu4toIUYFx6KIH82MBzbiFxhw4C1rOSWohTunVfr
qEEtWxG8wv3fDwCTZm4BAraPDfpCrNX8zOhf2mt7NSQnKKZw7n/ozHHcqGJSOYQ9SarDNEmfZR8p
LV2r8oUjvvXJF2M7gqql/Fjf7j83J9mx3gLKwDVRek2AdHw5J4VAVW/Jfci/wBiwHDGFrxSkTK71
PT8D0GADpqklg1RPz8vN1H8hXt3D+mkPGWmIHZiqFzOZBM8fqdCO+kbO0ar7RTe4C+i7ESxhhj+P
4ibUceqRRvE1mt3t+TVwH2+2ATxQw04PxfC2epBbFmX1tuQN0dp2z+pcaHvaC36zJGrrawUCq1MZ
SW0hRGLX7Sw/PNwkzDSqD9/Cj/5ORotILlQC8xabg6MPB/SmFrbu6/D4lCWZm9MVxi45uqvD0ySV
OkmpIV/c8jKEn73RfTMXYxxTT3wkVxq28+tGVidtyIPS2OefP5WKQ7UngXGWik4JcvIyGAaVg19z
yC6fz1S7E5n4r/aQ8fbtMHaeTk6e3nbIV6cMuFi9XGT7sMLo89iWrrfgfEUnC9xrY1NhbvyFvTa1
KWJ7whNCE6+Ero67aBQ7In6wTks8mJ+cymSpFR/4Xqj2DWihqBoqmAFp02Ki6S+F2gGfT6xkPSQw
Cg7skYsd85hf1fP/ti1RbHVooL4cWSKme2Puvyt6KFK3lBcoQaqNGz3H6SXDg5aaOPj8N+4SEvDn
5TyyEb0rhW5Admzg7+fhPnVIB8x7Q+rCyRjG1Z7/PCRbOrzh3QIGD3oBAHy1+UtTybAKnSIBX0rN
y4AaQW/L5ho35OhIq8WBInWfPX+NdyCABmDIzVr9/WwXFgbJbz0th2pP6+ADeARk6JFq9BSpvwJd
sk1ziVnyRxr8Txq4hJmXnFMGIJDNQxHAjG0c2TYBkFg5MVBKwd3zcxtOXObSQZYyMPhl322U3Y85
vVA8HoIWC+z9A5K1bFqhZetZP3YSdIaIeZtGLvW3u2u9IzIHS05LjbdiSmslFjtvCVLlGjz+QI5B
EO47pdKx56d7gVJWKVRkKjHLYFTcgrhWHnwkYzvKG6eV97yADT4UAlZGUgwnftyUD1YLEwrtj4sM
GwoQKXTCJ2137GeMdfEhL8lsLFBWJAhy8Uod8+8BC3msFERlLk+4Ptc0b13IY5rs62GxnP+/rZLc
vw2zTNK3MQXNwN0GuckwbuJllQ9JDMzpQd5LrH82M1AuiaaXXjwiyVkGavnRw8TQ8hnFspcGevTq
Uj4mUVcyyu2y0fqoWbZKrmGBrvANAWLXVstNGFConjtoVOnL37K1LAf+pB6TmnPVkEPv/1PXTxYq
3jx5xWC+5jPi2KCUkZ+f67qblHGgIsslBYBqLartSXcVe12WccF+AnDJubDh6PslLCuEjwc3YQ36
xVisNRbExM+j+XbSLFH1+LcL5aBRudMshj4AvY9un2oEINDy3NQb3upsUv6RTMCDVlBAKToND0UL
xrC2dWpOjgfZijlzabQt83NYagmIX6k1OUi7t7jEMnE5XosmNLqVZMuGOSZ4XUHPQmpWso0H0Dqp
uu379PWVs10XcsLZoaaO0vaWtTANXrD9hqOg4s2axyBbMMI7pbwaXax8k577tZFZ6J8WVx1J/fjP
6ahRFZwXfPmm94PHnTD6879CBXdfG9vvMRY0eNYX48NOLdMcmNsh54MLCVjTXCjFBiaEmTTSyjdk
iJxq40OnXOXSsUjiEga13Ptx0LiUmwH/tstg8vfo8K7dcIJ/sgnqDMOXSgMHXLn1o5aI/Q+FDf0J
7zo623WqH4aZg5RtujqYecbyekFoRysJq1fz9FGvSJaZjAUMKJvgm5tClX3IE3SkTCbrbdo7DMjP
ukGyI6euMZD3bWDhPkrqgW36eeIKTXqigth+hyywDF8R5S8lSLVTwiz7mGtbqdDcbZxEQ6QrnTpH
O9ah2NhyE1Ps9+XitmdyDVwKVAh6NeybX1yHlEk0zR77GZdQPNruE+m4DAmc8WSTTreFGhUkQi6F
JP/XhiKDv7yJEcVYZriWUChifuccN2NGZUmRccrdlnNun+VTapfllw5VVr85Xfhdcu2L+d38bwgP
qryNUUIt+EPGS5HLXZGUjCkQaY2mntwTUqd6e2dH6gfl47So1OxL56L4kzqgy9HUwXnfzNO4U3E7
WmCY2Fgki8qAdBRCOB1/XJ+jUflvdnYpQEHdUx68IbeJPmI6S2JszzUMtXbMk6xcG/O/M+fEQKbo
TUGs5NJc2iBpFhS25+LU5yVaSiubPP6TWkqUSvW5gIH7TP/pzGp8JTodERWM4dUhNt+ri1Sy7C0L
cqQbYqQWSwfCGf1JTsgTD65BstYnutE/HkFLcZtwtAfhkNXpkv6dSnULgNRvQkicRmi/GAK79SRB
s/gF8OPyAFdoCA/47kb2s+QV84C7vYHegFH1XndQqFUsZ2RS4p7H4nJpwC+RJevDssn3DOsVOO8/
Dl7ci8gyljrqKjMDSK8XfDXfyl52+dcdn65LBgoaodcMvgodL6SFwpMH6VzuoCBVo9ybxMXDipF0
cpwCNfaV9/9dN2n1UHnHjv16XmlDOV/11/lI2Df2nCRCNHLRmxqKJwOUJQXhROkeLsGVkP73AXKv
dpMFwVuqf1f48TZAx2qyfLEyqt1wl/JpBasAr0op3wBDrZN8rMFpfQ+OeF7F9X4J6UgXznHTs4mg
CzZkYGjeaVG6gHqV5hK9jk0H5Svl8JqEXPmzFk1GBUOO6GUT6JYv/vFg+++WoK/5B57Ma4CrvNe9
PfdsYIMe5Qh2/DLz9RgSdv+E5Qq84Yzn3rZHz/Bmqo7oytRvn0fWltTzDFoecDH7W1/VYOgYygL1
vOknyb5viatwdTJhzYFMEPCmXNjxazFnkuDsGOUbYWXzHrL8QbVdyx3eJwVyYRAW+yVcxvB89FYi
VdW3sAoJJL4glReriXD7lDDt6XxsF2lPLm04+ZEQs+E4Qd1fQoHHhIQ1JI6Ojnetz6z5rjSCJ5ax
gd1CopcwpOlT8nd5m2Ye4O2ShREhvpnpoydHxfjcv7QpH4WYFUbzBnzUAPxHS6S1/EZ/7jb8J7jw
rN/5NPmt3Ll7ae8RIfQZX1o8W7iJkn4sP8go4/LtsKXa0knmLytx4EQiyEryzWiIHYAYfRLQoDIl
MUEdOBhdcWhujlurzNGU3BOrDsomo2yljySR6ZRT4jF6OEd5OtBv1Ov3nj3GPByKZr2S/5i3uixT
ZVa/mhi59vviqYGnqUXG00qvtfmIhpaFdoyb+5FcBhDg9q1Cp00BcGUzOonJ26yktgw7vJqXI+Az
gZuLBnFOIM4yXjJ/sKxFlpoSUBoOKA4w+hK0GEFFWAOIChcETKI8P0fCVivrkPmhGr7RcyGF35gh
CtoZB3FdAQfB947PSiQKz/OhcynmaJOtye8sGwSZvPJZ5Ihe8JJO65A4UNnVIUbZbaUXrQQozmZq
9rLqXaUMZPmgDKLBcNWDoym61tXRx9UrnInAmMFSMToodvxcUDSe9BTlIEDpo/bBJSmDBiHVt3Ic
GdxdnPS+jZIo6xJfSz3+3Jf2OoZlBMGfVFUw+y3AN7yrcECSHxz1Y8KsuRiGg951uGAH7x2F0vAu
fpdHvYK/2gXYHDL7TtJXkEuqROPo9DWKXqzD5yT9x60eMYESkwgkATzSOuvVP/BOVjXCgnX52HEy
q+46E1L9fe+dY4FYer93k+s4rJfFlnvdBN5/ThNMsTolUn/p380Itch3bz7SJUwP8Ddc5HA0PHQ4
Oij0iLiK6ifOzCcydL20Hv+W0TpURSjKa7TdajYZdOb4wC25Nt398flXORtpxpLEcC7qCMF62xuE
XZtaThULhVvj1KYItQqg7EGIo7VuHxB5BRWtXz/niArXQbSh1v1tALXqrevrtqiC+wa3vsp7GMvq
Z7xFWii/GZqaNvsi73BIa3uvsL4r3SXWanNAMeSljfErGNMnYrqMVZi3zg5k3ZYmLezUFMwjLIci
oFDSJZ6phFrWGRRv7JJW/RRgJN2KwNZCmm7xdkIJRD1R6yww1csVZN3e2zr3tL+XQH1MjzT93K5p
Jr6cJ/zlbr+/010z4T+pJgi1pbND3NuQaIpAhhefvyTqalxUb8xhduy1wYWdRjKynSP1LxSsbBYL
apqZR4Enyo2iL8ohEfJyzQxcCaJF4IEnK/mGvtytxchG9V5z+rcNNna11cb6Hx3b74wSYjwi+mp7
CbS7sBkkpnk9OFZyzPCL/23fLFDMF9ivUc90sLu6p533LWolchv3JJdH7JmYEgRLS2b3xnAYhf6e
Uh8w9PfqOpPqx/4Lk39apDYiK9cdPCgkfi6IYgZS+rtXMaaF4CIGn5gPa1wkLzYLCLfuO8r4Xy8f
4d07I+8FPatJ3I9jDGjn5HFQD6WOvVJ5U2y+fN9b2yXwO/Yy3HnTarS/gM52TdZQPApaodGOIfc/
Jz56OlblCVCb3oq58NJVl17Ya9jINOCXpu3+TJawYyqg5yV3pV6hHZTLa5DGPuZN5dkjJwZxfdfL
DYFwZFtJQ8iRAxyXU4l2p+8jxItWX7WQHBCjglysdWBS5CKHwMLyZS9egAUdckcC+99GEnvz4OWQ
981YPZLFcD1MIxfJwvIStrqs+BMgAAybNJPJpHkWwdROCWxD+L3YCB+uI5NMRuJzgU2H989FYfLa
hkMXwwqqISkrszfQlLaXqyLhdI8XsiDzTFnvIrBFWvDsIcR5YQz9AsyflpdNJH3ggg+mRHoImfBv
OLZrgRVU6oJTXk9QTGvWVPDRI01rSw9vDIski/nYjdwfOgaTfBfE2gobVaNQd52i35FyaaTimzH3
vgC6KLw6xNgQI9B+i/ztF6CRJ+7Rq4NUVqlJCx/detTTRYkJ2yezqG+hgn+506pSIsrkwt8orQm1
Q4v+xcgL4hiuXRIrwnqxyw5YR+jH/K+8EvRed4PQ0dwBXwZPEhbDeM9nQ4R+Ezj3uzwOXXkOiRud
iJYxvtVt40p6WAPlsL7qfEYybdVPjCY9b+S8HoJ4V62V7CzpjIN41WK8vFNMqT9rGzgnMpQTRmCo
i0cWzUyBDu0j1zmwIHaVLkOTbu+6q37CZmnIWzbK1hSqarp4maOIe6723jXQoV7taNJ4qriWAQKK
zjEUdFid6RdtWHc1ZZ5f4BZLwi1UHsrULS2k5x7eWa/Mb63+Po6kex1BgrYIoAfIMvO1a1wIujh9
eFX/lvuPdIKa0pjXvNp86ql1BpKg2OQqLI9GZllwzKwgL9wqigYCKOS1kVjrJEus6SxCzzJiv0iu
zgiUbYLAscfaky9z1AFVJqs45OY/OybtLJSjHYfTkGdf+qngAYP5ey4LGCrZgWpXF/++Br5ufhoL
9nHVMZmI65vL2pUN8HuBq3mkmTBWRNK4RxZT0ktJKcUuIzJpoJtHw8f3GgyZXMUYGcIHXNWgxgvC
CNELFJh1Wx8oF0Bl9+xaeALQCu5ULSGacZckO1yLzl7O1yVvtbhBy3Y4JJGc0qmQspF0yB5FCr4q
O+YKwNIKGFysPwyr7B4BVAbWEGQaSoVejks39Hv0qYAntQln2UXiMzFhIKn5yA8kYKurzMrfbl0Q
Laia9m6WNoM1hhTUslsfcCNTv927vzUyJR1AaZWxKH4RjQF95B03+icnFSUAVnCh+kHRkxMFd48f
Q8Wpyoa7n5WYy43RGvUEDgPTWgno3RT5f329av07jIK4U4N1TSNowDqtskaT3YokraG6/7Dji88f
/WjaelARRUOiMB4IO+VJHJsmJrfd/O9ZYTtngiyT595zke1ErSuF45EcZV9OZE4BBjXStBd/zMO+
45EenzHvlDW7uYfvk8ko5a4TbwVD6Dcv5KAkF467UAF+winfJdKNnqUwYdNDSEVFhVMhxf+XHZWl
ZpF2Cp3YLzUmyKupKOZ2LEWlutYb2ZS0KKWN8hzMYsztGvBQ89rtEya2btt9Z6uKp/fbO983HErU
ui7RZuAUC52NYvjwhjSAK+rSzs/egx/vAfh7rvjQgh/z1c7Ui02PHsoz4ZHuAp0CNTCiETN7L/Rn
jsV20RxXvstJobl7zgXELDc+hss7PsfQXNKHwcETh7+mAAU9lgiyeJVOR/EMqv4RXop+SLz6kY0z
GUVuVFd2ts08RFlbYxuOaKR5+PUcZKA1o9UH4PHGB+S8SHgJV9gFNBn6hsphy+pWCURkBPTyIbDe
kJov2s8IZdW2Eh/n07NBdP7ZaTLzJVG7m3FuPdrOzQiBYbHV3b6nDAxD6+tjvQnKn1AsYIgUMduz
NIBxVuwWS2mF1v3g42BMa02a5Ryp/Um3IEVHxpBEOaSTCQ5ijE4ktjEr5RxZwTy05obF1eRycrTT
195t9ItUWghCPQVTVi1gkDijsOnZEW6EOvl11i3tdkS+SgwdqNI3z2cfhHxyNjzV2GM9nKDPoGqE
0WvBjBLsx8kIKrHm26B2p5Dbhn7JhOJdT454Uc91O7vY9PNvzkPUN6ozF3ZAZpQhVKNsD2VqLn51
m25rv78eeHIidF0TdqCYbDWL+vvrnHoiGLd3IW1RB1Gm+8PTXJ/XcpTp/ukVMPedmdtw2+Nh5Dzd
8HcqFtGlgNRbPIfkTgtRbCynMMXNpWun91i0kSeIEw/uxwGRiostPxZlgU8Gbc37xJidbvcqKpKs
C1HFkJRxqKrW1jhdOljrwJBvft/nQPSclryTmPMGNL46LLGsg1e/h56O3MbcXl8iWNbKQ3QIfcJK
CgxYxGyc126U95YaRSnoqiDXyKq9NxiZsItel5i1jNI+TPw4NEWF6UqO2EpURWwKlUxJ1Huim1It
mSLASL1zlmukcnkwK/MNdQEHnfnn83b8klItGv9Vjt2ezyenDjeQmbqNm/Jqw8O5kiLVHwX3zg0h
5Sv22PHnHkkgWRaXajzueb7EOu6bCAc3J8ZS6vP8zFG6HVEv8kMf1I4+6pcUnHMccSEmSUKxSirW
lgsa75pnbUc92kbbEa4D7GELwcW3b/lVzS8MX50V7iCiiQWI+ouCbrRaR5KBw5MWpSU6gQ1yei7M
EfLURQzvUTHLP7rti7a3btOisyiYAPJhaV27T5uG0rmSvdMdHwzXErE6adF6d66LyJhLAADnx0q7
wfWpyU5iDvw5bJiW9XCIQ+orWFcW07EPdYdrmLUrCA9CGYAMSdtlmzC48YYGoeB4Fb1UrRWkwGHQ
xTFk6VfswyxU4hOsO1D+/8dg9UcV3rDX+NRT1k6IqC+xxWxuGr6I3pGj+F83YcbzXywRiY40PhcZ
BmVvEWrB7nPUaFP/vP4DmDhOpPRnpHrK2nmfJwFhaB7y5XpUvUdNdoCttN1C4kKCcrC+88azexI9
tNMWU1dZwk4TmzEia0C8ZiIyUhrWh4saIYDfby5oVodHMYJFp2IA42xdPNy/GAwt3iOHMLyr7d72
/CF26TM9akjsjjFL49t0cl7GyYIH+6nKiTBFntfiNMxuaEMSVxQiYnGnbTELr//Bh0b5cpKdnWY3
PR11/dvGnFAjRQp5owCjhfpbZjHuGEY095TIY6i8ooph1UVzda9gwhxLO7pYl4bSdBWy5Dyu9lkX
PVF3DHYNBVKfuSoRvvEb+8rtS5psef5WfHquwT8ZNmp6MJQrd3E+QPfS9aq8JJFTxZNRtNdSkv0b
xnPh65aVkLyNWhOaa6F/rhaF0ziovEh6t0QF0/9dR33TYB6KMxpqCibj+rrQDinInsc64A7O5/sj
Br5u8+DmwdRXld/VPampUZrBwaZvkC/eOFOQi1MyU1TSSI73+OOFkRAssCkFCeJIoLWnkSjOMhsC
Wuf7DyNswUE5nSyKBOulDV7oJjiQ6y/FT9vYJvibBOKxhio860xgs/vrp1i0iRk3rek5H/93T3x4
X+DHAg4ILOklWSDZ6kB81a7+JVoV6qbNZ6vkPa5o614HtbUZYWN4x57VufQbBGlQrKrv7t0c80HI
5msq7HoMMJHvBYt5/yCiHxq7RPfz8e5iTBhHVMDdloMaNHguqbFGLtH3eQqOlt4MBCBBYwcyyILv
bbdq/e1nNDDfA/b3d7+M1RIH53GxMr8mABRIFvWGfcHbUHyBv+EEuP8lJTCvlCezgVzM04xaB7XP
eDss0YoZNFXmuHakboFIO7pdlZWWyhIKXVd2FIniDgnjKeWVrdm3b2GwCjwETEfn6XRxY6bDeC/f
u1fhY/hPqZM9drHATCs8VvQhRxA33wUTFsujKTbJdRl5a2U/HeSClq1z8CCG+/1bxZblO5JJvgyZ
zcdbeFARcJccoTcQgl93bgdIeUgIJm55VYESn+J4pwwP95rq+i9oNcxrjUrkDcKw6p+Aqu0dein4
WvhVoIDDKWU9iVbb9LQlbJDabnUq1EKOmEt5CnXtemWgAOEvmj4093jSXpt3Sh1zWlgEVYW8cYtu
yymv9wrwTivIGUPFMICB6VvA/b4Wvv55mwjJlzZd65mtDqnd099RxXJ4enFTYiJmRIWOSxnrLgEB
QSDvVzRBR2TFf8ulcMMYF2fOK6cCzDfPXxGhwltKqoPQiv9nVdfqMCZ/538Bf2aLBF1w8GLx8fDc
/R+aEo0ztirKpoboinTd5EomRdGLGq2Vt8tO66+hGsWJ/eHFbUyENEEUdoOrERAuhgJ6DVAhI8kQ
29A9PaLdldgUVqAXTPvzMKEKcK2x0Iyc9VPWPizbTobnvzeNPO92z0wLE0Q6uU6EWTleuJ7+eZXe
mQ8JKLu+7JcF4M59TzyuSsHnuuoNltPL2ddMl2SnJrm7SchjNpCpY4DA/EevzXle4iBcN7fQuSDR
+52FGCJwBEbNOd03W05rNtdn8rZMAWOPisbWGOGupgd2+talAORvwcT/Bepyf4tQF82p4nKh9sRq
ZsWgi9hJ+4vT6ReGCf3uqKw/44vFqAROXMrpxoRvUHcLty6YimhhfW1xWcYYlTapQW2db68f63QP
Nk0kKL476GyjQz2yFP64/sMbaTsIqB9E0/WuKDBSWsH54xyt8rhcOjez/We3wOskvoLoFlmQBGoB
9ClK0bFVs5Hz2KodPKDjY4XQ0cJBO+hFkqN7/nV1CdIjxGpG6HEFEV9FKsyeccv8T9M8KdHYWrY4
fIDhQPTKgR3aOZbu2wLMiXPGFe6Iz8v8SAKrqfQjhZ8SB7MGBjQtqJusXj76ijlONcgVS/foAEbh
oz1UkLVjgWIwY6kyo1IoFPoHkkoBlwmPh26KiQV4errXCThVopm1xKbPX5TGs4fwDQjr2Jc5BouY
bo82IwpH6hjm9czeq2FARQfvOO04YIJvdwUQeH6VvBfiwMyKQz8BBvyU6hzFSVscE5IHEMDF39Mk
wdF6Mqp3QOiiAX7STUocWRvnLfWrPpBIgCLjE5gpGckVW7I9/PR263AF77m3sFpPahMJgHrf//8R
SPBhDSPaTjtJioqMPqbCxHpEI+fJzlZjifb5lVihR+hSvNo2U4w9IgqZdZs869cvhA0bzyx0c0jy
f8YCRrC27ss0IgCSZRmWA2nOB1I5+ncfLoIIwwSjQXjuzu73i4jEF99nxK+FEdXHr89LjNKU5u+D
Vb47vOsjA47UqLrAkEJ8JGx5tEdqq1nPPNSWBIiaEBS5gqbS6RBXq5eigFmTvNZyBg+IRd+tZH5B
1hBOQl/idmCZ2t5d3eMjAh3f2I+DLqnW3P+ZUPm8TGhzmH0OigIWuLQ7Q1gwp0fk7NcO/3GZiGby
poEcVfUEAcVd3wOpdbckqndEnCa1bxnfjZMMtEv97agXEYXR7fH5xC0IAK1HcX9WIaWlAZZbl/83
DVhgCLpiHu0FGg1YWgMcPdiY8tSgylyguQayYJUrHd+/fL4IH92ZT8t7BTTRGj3FiTIj9kInZRez
/Y0g7IEWQxO11pDiTQ+OUYawXw0DFzNTG+OjLpGjvrv8LhzO+nSFlgmwFXd1PIQvXm3baNeJ7DA+
VIhzSReOap5yN+BqpFovZznaafJgoNVpheQzZimnnFBY7nF3mO9jv+ATiwSfLcsOZcUhH4V1dQCE
iYpFHfAdIuKt6KVvSaGujz77xau+52E8R5GucOcMUV3OESup2T0LdYASxA2BA20te89q/VHOLT0j
amnv6SXKGqgNErz9vmWIvP4QGs5PwoifVR7BTxS52KQi4Lhk87mG9E/cpu2x8WGszHS2SZDsqq4l
J4gn5LfHt89BYeNObtyqKYAtCxlc6UN/01hEnhAHlzTPVIDq4FQRG5gI2RD4/O+kufqYJeEA3ueq
eszdqkc21PK5RReCCm7JmJu/HNsnuAFKFcSXZO9MqtOed7GLf3fhExUEL3i+rSWMqa18H5ogvPTX
xnfOAuZP4sjjhyLDaJGHt2bfBQpzOX7ko8cypOz+SoZyJt+426ov/8zFl35MHSorp654pmnY95aP
08bXI+ffI0bwrVAcc+V5ZreQnexIwaSgq8+WJi992LfB5H4QZg4Pi6jnTXw+xOFfWmtnLfTbWAC+
Xzik0EvoQIM3D7ZvWQ1XSA7Af1TnlKuBC5kXDXWMliQ9j0iEmzGXY4PRyAnpkXMVL5mgOc4JppyF
V/C9olPlYI+Iz9VdvPgrraPz0U8Wv60vJTrsYH2HVSLEnfoIta+TH8vOLfNKgf6c6lnWXNCU0Zqa
1SX586HjplQQWDQ6QhXDTDirmD2nkvxJqpdOErgyAcdeErHZIurZooRZjTcvJpbMsyvpNHGZAyLq
cOoZlyFeHI6awByjHA4BqovGO0p8eST8IgnUBIXnw/cYu1+QSRlfhzvpkkXZouSTnO7+TovTme3/
GnxcoGJCrr0KUixU2w7yaCX442rZ7/pTvE2e/bZ15V6BBn5HWMBqrMeBbT8kFDwB6Of/Djr0pDVo
itZ5agRbwV/soesc2g7b7ev5oCYajNimLUUN7SIOuqs3Gh1y8DBdSOJPaWeXhwuSgQ+ug5cBLD1y
ca9kOPHmR77B3j1qB4DGPYnoqZVuCDxiIguETkzdVsOC5b9Vkk3/en5tlwGq3Z9z0RzpMpIH+9w8
UiykdV+jwbNy73MiEOS58z77bJ1P46+LFllnD2EP1+YtjEZQBfJSxJJmJGej4BhOxu8tzBEdQzCM
CcKQhgWOj3y3tjbrXrsZ+Bs4R9UACyDS3+OtwYhJ/8wGsKl15gVjCS2W3ZVlba4sls87PWLUpCE1
7M0P5736Mwwtly3FL8sccS+mZoHxkxKvEuTYH+Sx3WLBFvqsZfgjnwdCGNXkLCuBJadcmtNCnQC0
yxhVlpLgtdPwNWHVfXofsir8WvLwzleieOXpLxpVI0ACVu1U4BLS7SZDV5jWl1MLDikIOGgj9HCj
AdTdalGfWywjnLIBFOucoMKv8I1awNSNd/wLBnQNbTicksYRrkIFR5G6TckmmaHeUR7GxG9QsAf0
LJE61dW2X82Pf3mcz+7wyK50/vYd7ThoE2/kwsObsNDB9uFggBblUMvB3v40qxoN+F+IFx6DahBn
ZMQOhCEX/QGYGPdiSSyTIM2nfu4XRDdK1Sns5N0MVyVnzE4aHT1ZufuNffyK29OA+ZYL/Lt3UP8f
TP3+cODluXX5dVA7wiZodj7TQY4KhVL41VziFR8g9NX5NBBhidMlbtvZdpn/bQ8loUzTHM2PqKYF
VAmLv2A9a7af8QtFATzQgiRGfcRxNIVhTq5rbBIDET7QnZWZdAL6eaJF1WcvLyHOyOPq281Rgz5O
t0XqXC1ZVpkC2SfX/hcmx7UR/ycOuUjC85efxrGYaEtePlnR0O5JBVx2A+eSBt3rKP0/X3TRerdM
J0rYGFC6nbSZfYk7Wmil+zGZSXs7Ts6TD8a5ohdyoex2N4W4xyVTKrqXeRUwapVaMI3OrLx80G4i
kljY60nTBgU3JA54dRwR1J12MiICA+8F97ahAzA2ujRZs8oYA5p5nyu6A6Ez5DLg09UkLsYAprIZ
IvQ7IWi9I5tx3RXMaXg4jwb9QNn0z+OwlnNrfGTzKNCGs7E809YgnLReEH1j4mkRLRHdYrcRhtrW
JOrijFyB6GM6y6Un0F0D5yPWzq/0gC2uYTpU0skjZvviIaxkRF1HPnZEck8lKefTyn1Cs2sS1/2n
kb0MBTWmJVJNBnto38J+FYupDjUXtVVHQapeZb3jehTkN8BTXhI8sEC1K3L4mc2Wm1Z21nEVPCcd
FFqHpc2stgM638j+46rRvFmhG53+m3N/KqWjuyaO5qFnylGX3HIxgZ5A8ZNGSvUtnLHiXd1gZnKM
GX1ts/ynMAWS1kDs10WfFAauTL3JtIQ3+U26By7sHAJa7w5pNrHMpCkOaTORWUuCq2ozas7OEbKK
B8hZGFXXVbJ+ZkH8Xm2/Om8WaBBmEwahiYguQtCkN8C/zM6DfBSWZueaX42A+8T6UFVnhNsRzjY6
LE5j0CtAzgUy0+UHbYCZUvi+KdkzGyAhy6Sf8elqbLW3YJxQwwBkHBsdOvY+klpmCy8GnIghIX/r
C5IKSZZ/8qeqQlyU2m8l3xbvzevKr+xDkXxeATa52ICBLE/ryhz8VehytOXiQEreYRafjRDe2o34
RVl9CsVGMMIQGLGOA1fmJxOQlrm9LMFP8WluyCSYPAKeimahmelixiasmF+TV5jdo6KykPsv4hFc
ilyJGeyM62HjAQk4kVWLi0Y1IcOyNKO2/xmaP5anR8rkyghkkbPW2TbD7n7wVqiT2RMeeLjwg2XR
yx2fYXHK8FlnM74a9uhgk4ve/5JM3188Wm43lT/oi5VsDq1SjsT3J3Jz1nxRFU+ME4l/54NTC81Q
+M6B4p38A65JkIZjBamoczxVNG6DW8UpjsK/gd7psLiywaGaE6LW6ztpQ7aMXsociuyenkW/GdL6
F4Knqis+qAS3vSVxKnN+BVHITr0G/x1Yg/X8zViht9KZoVP3C9PfJs20hBLqMUXZT6cZEylY/yz6
mNpORfBFwqh93aTDA6LsafOLWZiGjSUrutvkcfnC/A+q42Xjmd1PcoQHVBS+NW/IJYgvS/NInn4i
YkvrOC0Mv+Cz9b6jLgrXBbmCHc5LqqtrrBX+0XysgqB2wuj46FT23aTUERaKjn0rmQpVpMFKLV8C
0FGyoQEr9OvGjBQiSwhmbGHqCzaiam2p+sAL4soBYPZ9GoLI44koWqufp6f56Thn36uPHFcjgs0x
ny5pq53A07uGIzNpz3AqZ33h9xwzDWm2+l6c0HAT5EYoAEUlgzs+6DZ8Okw9O4Y/eBGvPVOIh1uc
9UTp3qC4Enu6DleWrAQum/tyXa/6rpNFa28smnDqMvQnXzYTX0xYNebnKrs+BRauUxl1pqt6kpvv
vaXpHF7LP6iKLRaYpLCDW7dKnXNwynGSzoRkJl5MxKX37AdplW3Of0+cvOBLpgNS+biqJLdjsYfD
462p/a0qUO6JefF0TzFbgPCGsij4RHF7yU++Mpqok9NnXYGqnhOV4N9J0l34ZaqpVdbN8BbGnEnV
W/dWp6wO36GrZhsS9D2KonoflJ1IlLIwvuOJvBqLdpTFQnUP0ZdaY2p+sEr4W57n5CNC8HehEyS3
GxhFhl2kv7Hzw91k9sxtt/EpfYS4xkaipypC6bFk+p0GGMZBX9pCHF3qh/SdDcUWYHUhqRavCgtK
g9B7vLNDEMVf3ywbSHXEVAy1e4l6IecEQiOvfc2dUXyIH9WSVoqxgp9EsK1oauMG3IRjNXHXmrM0
BrHRG8/gd4RHtvrCTc353MiOppAG1b3VfI2BUqyYCqoDaCBKNn/BFMXtt9MuugODA7128xBb4lKW
9n50Jdh1AzLQuLDBjsjqhvp4YiQ6rs6E6dukEtXjCzhCZIuDW2lQG9K5dtyWstLmcBO6WJE3n6CI
jRh0XDGQ8uTriLX8qbdTx73rMGn79M+x2q+pzHsvXwqya3HHfkF0ScVfHuIY6mp53OiVnbdo9VX3
iLPuUjMe2mxn/1ljHaAg5EO8ntfDyraZ0n9wMwZYCEyHrhKFrkOBgsFN+t4CtHF8Y+0srH3twTnA
Giw13fr4WygSgMh+yJWxQ4oZXh8OjN1EFw7YAMED1Ob3PakDMH87O1/zlXBp2DStzXBCd6DWj8gs
TKSumOkxfrS3zANLRFb/v4OqklZyXs43GU+n9113+IljjRXJXYV3wGYln0kqG+dtlZWOvwFKaKDV
0MbqxQ378i4m+J59D1W+NbHUZu9gIJQxdUeDEukR2te7Qi1W93SLmnJltm0WI/rpYTfhmVi0QY6b
n0jxi1gUELNesxBWUXsN79RVOFsPJbDAZxMFQ7aiPdMjwil6yizRFqr3hcy5p0+PO5Nihox826Hn
WTlCHr1k+Em3GSRFXvEb1WPihHCaAiFGfZ2MkGH5aLgzYWxje33ZVOynW2y1YJKCYETRDeSWI/a2
PqAri6XSjIwiEQrbhZ8XbahJiRb+pdBx9giW4QM+rZvTyeLovbvUXsI1PCFDeOD1OHXrrQEmFP7o
t6iu7SEhBTe8jG6rDa3qXMwerJ8xmvagr8oX4NlnjYaupKa/eLklmzSkJWKXS+flgLrQIMuDm3+v
T43PE6CxBvUV+2BYx/UOF2JEBBnAN/uw9gw+SaPNecAaOiFBVy1reyJM8aCPY3/rop2qFhubO0Vo
camRPtyiJ2NW130UwFRjmqru/8eBo8dOXEIg987VntyboZEn7gsPU9o7vCH44quH9bxw4mM287pQ
x8sL+86mio86ZeBUA0DM6gaGhzUoNvfj7HTA7Y6mWU5cpaZnfQIXoJgFmbb76ug0A1rVc1Vr6OQ2
XI/V/8oCQmUD3MNToxFR4aMKUncfuMWD+Rxj30mFhnEMUwuemNE7kjawS11hP8m5oL0PLPGhE01S
nq+xMLBPzBLRmNqP8yjwyFowYcVHQSe2elU1iufUjJxLKZpJ1KKr4N177FT8zbN7R5CXwhbCWpSl
VClhsZOBBRutKu8ZqcMyowe9CLHEJR7cDAYdoSI3qDCtD/XsKZGWly++sDXUwBDM7+9zSpQyiovS
u9QC1hz6VYyss217uB79ZcYRzi2P70c/FmoNJEfUQvv5fwHRqVjmIGSXNF+NldYLQjvA2+cSbfmK
EnBJLNEbYwlhaGljwcCXjLKlddsgNDfx5Ri3h7bQy7vIuWGKPOXuK3aj1kPJFY1+RzNn/NnIj9A4
CuLEcsvJRQh8ACFKfTFEAMjQPLPwN2pIUwGuFm5Omod3jehHDbP13UZ31zApPjaeHMFBgUfe7SBS
KZ0aw3l6PASzJ385VjDDmNK0f9V9qUGxPlTqY/H7TvA+7tUHck2HjyIGn95JypgjfJ2qBjtSc9Be
zN1ihKLkuGk0rBNlv7VYWlDSEA/+eDpT2prEAW7ZkSD9DWH6BX81PuGMqXqQNJJtqKrSuxjr4RWi
AO2pkjnomVuT0jpInlZ8/hwRdylcYVGHeYuUACIsHNslthXZDEEI9PFnBY+5knUK+OukeXJPl5JQ
Bj1+6HPi7x4rf2eZ5r4hFIaLi9GjCbnTfzk6K8OL7NIk7xYOxq/ZoP1B9u5UsJn2c66r3tWXXnWK
vOnunUKqv4jjsEtrUw5MGy6vle/+pzQOEPD0eLMbKSQ2CdsgogX7xXZgLZFYpq1WAxGcr5AR9jLP
FgT5k8c9HxjkDnuX5UXsIyeGxBMunutf9ihk9hGwLAVb8h3p3ZpESiRrg/rarCblMr9l3u5ktIY8
l5fyp3U11I4zurICeyHroRVjrYuw6IK/dZezK5Yuq6PpqHGZRWluM6FeX/fQPDp8oTzxmGznuE3u
oVz8H8MofU2cYoFJyd93zh6HyT1sItHOXjFi/dKbkHpbuJjxjgxr5rExzNobPBA5lpGgS9ylIdPC
FUFvREgoCnk3dk8urg6BEIYO60OPHmsFjIM8qJv/389J9ixPTzIOF2f2knZ6sJjTfOWiI8oB79pg
p2cMmOWbNlzNFt3s+dSFTh6Z/uYRLoN6Iuynikfd8UqBEYAR2EEfrrlyY1P9mqeDhd58C214LjRh
A+FZBePuUbGt5lK+nkmZoM/Edi+lbmvhwTylH1dWqQ1BhxUFqPr42Lgz/KaQXZCsWz0jzLHzWILi
SRnJGQ0RVQ70RGNLsp2li690ein+XUS3jhYd43oduGoxlEn2BBCUtphC3/nEtQ1a+tvJ5Wq9uE15
49I9vQPij/qWtlpyCIIlEm+AYKbTPnrIqjEFtOUEObSMPbOiRthcbuQ9R62NTRx1OBBeg3wBV3dw
9DOs8IoWZ/5W7TWrXLW+g/UjbA4OtF5LnaAIsqPQacdjGZzM48LgBMdAsBijMM9YTDN26J+bf5rs
uEaIbeDuJ77nZD9oroU+iPvFdGoBRkETzE9gijSMGZ+mpncuQkHYM+xodJgSTg0EsRTeBbXurhL2
xBKnJUOr3xlj9wDCAVcTw7jDEcjPg3YzLek8xyLGruBAM4Qv9qnM3M79ctnasn5QDFgoFJhJM6ZH
DvSZ9ZzjgkPLjVPy9S5cNdhpID9ubHdo1xA6VU6P9oXt4QYltrOtOYHBpupOKfm9t5SZeuozhdhn
YsFftAcLSUNIG9Jfn9v1uT4fjewkd0fZaBzNgVyeSwaTHFNqMozGVAQtJkHrHS5veIxMQxXo9aAz
EPNb9EJyG3kO1Q3+hrqgc4JJF6Ryp2/FH+U1QtYzgqfAo6CP+L5EAX2A9DeVXrm35xaEjGVIZ5jw
uEqsor3ClfG2oe7UX9vDdYbAxvommoj5RXactl3vh0eQs4yIXe7cTO9oUzbLK9Wcaylto21ZloN+
s2IAheucaJZAD58yLznPa4+D6AXTirI71sXc+39HFfWP1T3AbuY6HGMTqSsVnIBmDvDltU3zScNL
BhjwOU/qE5c2f4GiZkt3dIZYndiCfSgXolUDh7Rgx9qzZZFLiWoAOcyodN37PEIPBmEblZf6syXS
6RNTR4DQgaGPUxapRI8kIZBB42HI/CvTESiriXYWsx76C94BMdrBMtpPanUKKu9KAakPl3dCxUei
oRfj4Gu/sHCJDACE19ixZNq6QfmsDkzGj1VB/t5mTf1dTCCnaZpv5YKTa91gUeBcwo83K7oEeQdl
fZNVFIdTF/MXehE89WnCWYoXgL1/lp2kdkU/lCUz/oaFJ/PPCCP8WokORkgeSQTGIrYe7Iea9OCI
O16CTOed5psAjyD6MMY/ZYNbyfAJ1vcC6rlpJmXZDlKNT++4g8HsP325NYXYbq7AatWuZBl/cP0B
rL3kZuF59wW8nGaNv6yggW4Pwq0q2K0ptsACUY6+JLUPi7gQ4OdFnBTusWSqmPBBakun9i0Q2sph
OZkhSwdcYJZUrH7IknU+k+C0IpsQEwhANh5Cv6oaqnShQ1zneLCVLBOU7m0uLEAcrr6BamuGchWn
UYo/kiTT+0qoTf7Y75TcpA6g4RXTmyIdPf62agw6O/xIkr/Hsm+ltjnsMJX7YlbpcAG0J9QpZ9k7
4S7wd1M5D54lhxM2I4CE580xhNr/rGc3+XHyPnmtLUwiY55T7TsAb4U4y83XCjI7ynxS0kkgL8pH
goIqlZUAJPm8gx1Ln2U3ST7SriuByf/YHhERDHrOdLyY7T5YV85Hx97oMFmE3tiXr5iXDm8ordWj
HL/LkCmXCBfC0OzpDfe8bwGww0G9Q/OXRXhCv+g41FVaGcQeWvch9fx8bn0on6ASVT5hsYR6qlBO
o4IS6O2FO4W4CJnZw+tQECpzlt5msVYpxQnJiKMU/Kqiyu47hxriyRtKBkXeOgPcDQ3SDojL02LT
cuuGpHxWwld9JwUUhkWcdLff7h7nV7z+UPW0+mR0VcjQtzdTHxS48U5QLRP6GXHYlwyVNcC0rXIl
wVZTzlCUR5YtkMpFoAxhXwtSmRq8TtZyrhR11U5yMuapLvAi2+4zMxnZLwS752NFFzcpYe49eVLp
1D7rqQQGAU+2tgWDn5PAIx6SE0dl7PfT3St92J3PVm6r+WOYcmIAjP8pPiESmZrW8KdcCRXqiiJH
O6LtvQZqY2Jyusi2bpHxRYShGhkgAFd6SeA0KfVjDWsCkEKXpQ0ciSq1+72eYnRxpnsXRLczMcFQ
7qORs6PVgTbU4y4S7mwXg4mELibWxtNid9dSSimEDDgCA8nS2lAQ/reDSAxYkDWgDKZH4TTZ9/8h
oaWt6ZNXDYkN4sUS46Ksmq96OKNBejQ4Mx4H5Sab/5LBb4bdlf4bXUtJaeW01wNF4pmsenhHRyM9
RRwH1kf4UTuSgIT+Twt/dhW6Nr1hAA61zZI52Jq2ITX0c/DnXQcbFj8vt9HAFAzmaEBqCNzKlMJa
62IKUwjl+1K+Nr2+gaTbwd+KRrRlP3UIdOO8S0NaqNHM93v/3WL7Eyi/8m/ZmcYV72Bv3lINZ/3F
Kh4i9elkl9hvoD/xqTOoZkodn1fo/Inb/x1noa/Gi3JiyyaDd1b9ntwDeCao42mn3o3k1A7dC4lU
2s4cGmZgeJ4DdVlmnoGQt35mGJNEMftrbDsKRZ00Gp9GDj2JkSwlA7pCniCqfplp11W3DBpNLrwo
UQHH8fsoff/TYXHjTr0zUzU8tWh1vYfGDiji3EruIyMCM2nzwm6zVxnc867S5Uan1SSwTOJiEd+J
cABX5OHWkaiAA3dxWJ4XeX3KwUpz9nqMXyhBC15MlOSiRgODNFoLik02PsWCcOuZu1blEPHAnrhA
e2TvCleFcntwV4diLiE7QpQus8ySw7+EkU0wLgsc+hZiSVtpD6hQ3ZEeG88383dUEPDT/DS2dLfC
t+/sd6a7EhdlhpLh54EWPt1aE9Ho50X1EuuCv1osXemD5r7dpDinUL/PY4tS7hIYmchfEAI6/L+E
oPZ4eVzCGOyBsNcUFxq7Itd1s53hWmV+LvGnZa/yRSk7nVfyAYJbVDsy+IPyHREz6BARL74DVHGz
8i5sy1bsdWFHJNjCaoWzc4sZGexA4F7pEgU0+YIP2NLutK2MfeaOYTqiEtYgA2XMvSK3r6vOGbaj
d0iV+wXH2TbJ79/V0dJQWDgLoQkoUUSCCJvHodIcoVzYor9THohz/AdWOqgqq7cCmrB688MUZC+3
z9MhRHxubfOT/0t45qQK+dKhFF8hagmoDBAv60RZkcY/1SfPO/fC8jgAqGGtvthXOf4SJHpmmIDc
oWWyN6crdAQPW2pLLvNLMwhU7wQBD6YCBd04CyrqwUA2KyTHOeaSOgoooVeCQuKhqWBY4kYC1OIY
BftBJkTgAHt3g1ikzPyCXFht3NUcaJIjHdxhsFfe2cNnq3rp04aczH0zF58HdZzsku0/y4/Uqzsu
wFIwFqgiVaJyQz3fbWJ6Z7lmmxWbUoanhn/dZJ80AP91z+acvPgvWeXaqVxuaRCKz2lAQzxvHaGQ
0XaC2HED83SvhaXN0NZHyuZ+r+3c7dkxjSiRY83srWnKY6/8J1bm2DROf5b2i9eWxOE+n2kC4QVi
0zbJFwEMPmd3A/PWlpNhCy8OES+HYNof35pMJ/6oJbYJpJpBUXm9/g2Umk9jxooFK3qZmkj+wmYH
EmWt6dOSyODPTtGJ1v44WabAARbJDje6kQJoy8TQ3NXn1xACBJX8mL9SyNYzIR7/lI7Cu0GLifdO
6mU3FxZCEKLjn/QUXO44z/OY6qo9g+GEWpPsdFq7eiB7a4AZS7mzScUl4p60cm9Cow4Rf2rHAs0p
ZI982+1TlyoR0/3KxfnlS6DnNOjbld+vNmi0EdSmYbzb29YymioZ2GnjWq8tDcTRPAVggLFnIJMD
+9cr4lFkg15Z8KcyjdZEOhWJcj+hU2JwBJnVNtlLhSx4cFNICLSouYa7wPT5u5DphT/XMcuFxxl5
5z9ch1N3xFwpH2yJmRuqKzEPs+9idPPQw8i8fBEG9kHWamHl8QX6zuQBP+XYzfNLbiTtHPaRMcD2
epB+32JJrQPigutP2Ffbxnc4AicCM4X+qgGa4D7xYH7bI8hqA5vWbEjO7IUgnDPiWKxskvc5iTpq
RWzpIQ7mzjaU+UGLgA+Y0wAaRxTrbJRNXFp47oCOkMmjFRqSWtrTfmHuM6efxmfnOK2d5HT5RipB
gIfMD6x0uvo3cbsVVmbVtE+MtcJ5XpGd7aBxZ0b4/b1s3h7CI/AF7iE5g5XdVM0hLHJI6UpWDov1
2cP52rxY8/TThpl5NyCQS+drBVer7vWSUPC3So7Lag3EESqJbPeoN7Ma/vUqUwaF29mUAB52Whi7
KIGorzTxftbRvxo3JRuChHBU5P4O3CPhmhbqcYx1oxHQERGZ1qzP651rwdZNZC95UQJMpTBgce/a
98ashgMnimNk/ITdPUzWdJVznGY8WxX2fJHagXZMJ9F7q/lO+/+PmG1tDhZ8GQi31LQf0voDD54v
ercs5l7vqYG2NWzw0dhdlf5P4BV4IuZRqPStrMXQhHCkP3VaFxmTwxBHcgtugoQZazuM30GJPggg
AZ22rcylsyYyNHnEW4V9+Od4RXe9MRq5ESsHGSqkM2WVe1yxHUyF3D6/4NPZ2QpZNX4EdusRDWOl
VoXuNtG74a5wZ7Ezkjafz5bqkPr1geOXFS0O/TmQVjYOM5IaXfoeARU0H0ofSFsSzRLfh/s7NOW0
G1Xv748M5l6Vf8IEgkrzjCx0QgNGB16WKe6WT6li2AXxku6GZVNnNVRBntkWg1v61wTjTSicCDbL
eVsgKo1uQrK84lvUPFY8RTZ9XcTvcvAgwtXQxeRQOTIVyINx7gpBtVKiiT6wq20iEgiGKN4K42q+
v7odlUjrCdCSRDgmr+1F09QZ21DS1exFWSCYgn/Bc23Pt7FrpgGdYHr1BFRVX0yHpk5hrIhUNJxM
73WWjaF98My8DjTvhW6j7zKpbDG07X07Wg+SzuTjAB0QfuuLsosbRmTq66uEOQzlEu5+LWEFdlRE
eA6Hltc04gFLSU23j1Ibz8K5lsH3EKeUliAyTHzjx3A1I9D9clpf8D8nOw3wIzi5LOVF6xNHPcwZ
AZ/rcVOeZwD4SK2XafhAzKvoqxh1Z7b6bcDRJ204RrdO6X855fd06pTcWyeGq11R1d7qDGaaANgx
NSl6V4//RjmLhNGGn1vmpUwA2m8lD5RyjU8c09kKXZFKWaF/A4OYSDlnIKHCNrdy/KHaLSw96YtZ
0wuBWH1Vel4JwfM1/kw1gVDRDMA1orw5quIe4q0TeIrMLXucH2vt1XzZRb/OcQmfkW6X4hSraM+G
stjeXNUpLR2+FoPWHGN2FfONMSaE7qvBu2DqnkfMAT2WC2ZdpxH714w+HmAZ51WDPF4saN/wS3a9
sega5khfdi8+H8+rRbl307/YyitZrxX6skzHyQlPVDVE+wGx0beqU2EwhoAK19ckyeggzbib8C/5
z1s7fRQz0a5P3NY4RSkEAq/UoxfIC+TEDSVdMoFGPDZ6EIE9LZMIKJTbpwC7SgT+v4etnOxwpww+
WU0MpwXD5ZHt1fjCM01HBu28iurbwFV4XWAufGH7b51E4zkPjgLA82bbkQbUIjdcWZfb8/7h3uI2
dh46BCbkhMq7eKux5nuhBXQ+4CWEduIr2gMPsUc8dVysCmoX/ZIGPlduYX8/9wEBanskjrWZvTEx
zOe+npqRZ5lWhhCpV0rt2b4OVyn9tKec3PzDwo7a2pSRILBJ7SdBcOt4IK4yXu83AInMBAhq5Yq3
qM6x/TXVlIPJXGzhbvxfd1SxM84goF9S9ISUQNaZChdz0iHLZREWFcpYUwFmAl1mXGXI7lXXlnJq
TzKSqaKcJfixLh4W25h4V7yp57eIjghgr/Tlxooj0PZj5fD5MdPRfbb2CLEN9eR1/olUf1jVvkxE
001LTgG+XMyswBEaK9TmhMcTsKgzZRbZ/oRk9P5uP59M9zXqdcyv9mMc22ITbPESNtWI+QyYTY79
f7mvmtkBvRiF1KRZaaQJmQVHzc8PbDSNqU7jouGDCrWbxAqU1aoXIniEV2uOk4JXYey76AcjvbrI
1R2Svyd1p8qoxHG+/M2CVpTUvlEOjejVdhWhVeDiMQhRdcG+dLrHFOGW4naczoCv0UPoUnr6bt3M
nWbA6nf1Q32GLKUaSX4YxPfGrnuQlAY/l8E7lYaHZlgrQmSCQkWxuGcdQBozitCtYxP4oabEDLwi
NvJlkFUgHpXqfbSoWsTPnX8DvHABiR3r0HwYIDTHyA1+o6eQUpd8dlIuESzU6DX8BMPVHhD63Cmr
CB6i0KtTpo9Outve58iOvrGV+U1zYvf4cTgMNVL5GMG0UxsKIX3KJzR+11Y96xPhkLZIV7RtqNtQ
jMofFwjJS1ZH5dq+eUZ+lTi9yMZhSX/muACJThJ1DXNQXd151U5hGbg619jGnQDpGMAI69a/kOxw
uxPEALIarMEHRP3xldji9qGLYHH0BG5vhrbs6pM1Erkm62cg6soY0T6HadH0wS3PDmdmsLJjjfgX
J7cOT0maZgaO6rSicvqDbMbxk/lfN5rNAcMYwmISZm9DFL6BwObEeGFzUwae62HgVKk9H+RGJWO5
I9YwiwAyDFxXGqEDJPuF0834QLvq0bwZ+2vScBoYNk9/p6ueuWi5FUgud8OyhVFaoVJ8xs48EE+g
Xbiu8C6SJxYN461N7g1DXRMzrdycEUyw26iv5aGCKdcrDEV1qIx8v9CLGdwAq3Vcmj2oUOnOWbHx
pjN1kxWRojGtbHMZUyH2QuvIr5TUcaRrrZQ6EKl9O8gfsGX/+vQchcF6msSJ/jFpIo6dzeIPkxua
MouCkNptmirWji3dO9+iENZbiJ8fHbTDGpPt2LrzzHOpOGSmZ/0BRc81ggaTQqNs8FW9RyVDJ9hc
/z1jl9r25ckgNAOcspT/5pWWUfVma5t79eK3pGFE8XOPtQTJADXbheltIiDZAqjZu+78OOnUsQcV
dYV+wKMHA+7N0AfvpDwV3+1OKP2r+Eo8bzg/ogzS57ONAOA28IooIbSaonsWEnJRI7nAZSoboJdR
EwGx2wlM3GHwh3kSflLVNV6U6CdXyRC0HdIk8Nm8eHB6dXsq/lECL/ebQr6HWKQzvWIqZV4Xh2Qb
SXUHvdHlXh6ZKta5K2S4/Mm86ND7Se16cyEZVm6WMfOisxlUa0Hwlgn2XCswlczUmvQmRQjzBzYD
b9Kl0Gwk5vcv7vQFsa9hCCZ1SEuxYETpbz5ku3DI9TF5tKfShDCM3ohycIeuD/LttE0NPD/k4Jme
RYP3DxCvYJhUGrmocyK6vtVwCMDXFP+rrC0TWE8R0Tri26SQI/tVYTXRRiwbbeRGJH5LY/WtV1+G
AHm2tFKeTl1wSuX5F57OK+asPRFxed8krk3tk+EJt8+gQpmRa54tmXfwVVrzAHdJz0hpKSvss+WS
gC9tNeix3XKoHK4RbHPd966fDec1BI8kbAJPFEntOMS8NGDyjB588PV4eWJKetqvJU8rzgKvLujB
nGFOGVHg1T2TDOPDRjUnzVWF6zYqs3lXDuv+bOLiwyOUXhHpksl5SeJiO6m3PaopbKQ5aGW/31qO
wqFVEiu6f98eFP5tRv44M0XB2nhHvrCcnbVAFpKjXK50JHP5ueAM9hsB6Oyn0VCWhHYGGDn6ixQt
1bmLHn1C8offHHEpJOWyWw0QKO51Xszs6Zt4iXZWrptv8Q8cfP+ov5wdvf9uBGQ1kJS75SRv0geI
nNyrCzu5GiQ6+fNgtumZkYUbwEMBHMX6HrWcumKWAwU+MDkE3xImHYKEqbtpfuttEf9JdruN94uM
D+uSQykxO+DVf6iZ/Thkm4EEcllFrTm1Lb8ZcCf0dlIB5KACcR1RQGHKQsQPNZGMTsfsYk9JI2fa
C8tVN3pxMzmAuztlrDWGxXM718qtBw1IvYos9ulFevj0TUsvJFIfEiw8B3y4noiTF7zeKkfyhJia
A4srkRGeaVwVuMqT4ETeCfqp6aPhwKg5TsT8JbRAHKJy2kV3C6GahN2qW7i0dnJJ8C5Npoe0FE7n
hdgw/Mq2iS1HO/nHe1qVS8tyFd1qaWVPYhUot/5G1X3vjxn8zAOJsjKcjeyOyxMHRyZt2nknWVoz
83xLJaYOaewT0F3wa+3Bw3gc0X4IlhLVf8LKMnupPeKsyPdThbAQfnYv3B2bBTxA/DBAY//+mQT0
5g2oIKpPK0J8u0o4xWwzUQ1AldKtpRaSyxtKbD1AvZY0L8CTzeP1jytca2wuz1b43QG3tfYlj0//
ar7+o+t6/JRGJ4/8umDW53tY6CLiYNCgoE+kRKt8XQO/VUWleP+xBfk7GF79U49kzdY0talSoz4A
e/3SnqxtlVT9Lrm3H5U+t6SR2Ke4TbumTZ5NOU/fenRrKd3HUWaWnvGUYEuhF7ESxb3WgSE/5b9X
V7DZlYWgpqvSrmxo3PyOtdQR6nyRkZkixpwk46xVggTmq9wlnwq08OEh5FlAEoyoKgUvMeVyBkdk
ZLigsrS1ROrs++JTNGvzbCO0RlFXVSo0wSLFSOeXCkEFSmXxFizTr4+lA0rqORz0RI8/DxfEnlvW
8C3one+u08A/SZ/xk+bDD+U4xD/3RhhLrN6L2u34nb+U9Rx8z9w97bXyC/GqA2kvF2e1BE65uYVG
U4TKiy/dqwe2KG57oQRDDysZI1S7901CJGBPS+seDYCLarHF+GXZMHk2OuPPB5UPYlc9JdWEIyl8
OtrbjRWcYxHf3ajDIPEezdkfhrwzVWrWBiBaTYCe/vI08otbEG+hWK0B747cUDJpkbF3262TNmqS
RKN7PEgj0u7b4wy98Ia6ryfH5+fnrm0ukR/GNV49iIaDUHDsJgyZVmEXq14ZVUmSbeM5IBQhrvci
3Bs6Rc3MYytFmfkqPTlYxd8pzJ3d625qFRuudY0e3WXgqvPSPki8LjW1PLR0NmCg8wb0vAWrCVv9
6jvKCNYb1w553njI9YVLh5pOC4nJVJ7YpbJUTMh9wYIBSjyZ6YAHs/6Bu/QLc27IU/Ri101gHC3s
zUxkGhH7f4m9prcrE7Eljvona4hK5CvvlSDHdFzq8FU8uhY+D22oMBKvOe01+lODXNde9BLlSG74
QWu20ss3R7s/oRq/kai4rkfAxGhjyFD9jbQ6o2WH4N9I4IcuoykJi1qiIcu42ixPya3RDGBxdBiG
dJsiaMhrZZWcXVR+WnCQDBX5zNj8gZm5AvV7V55A6V5V+d7u6DYf4bnfrQC7JgSD42jWuXgSYYQj
xU3iorR1MNFUBC1It3mWcdTrol07NDEHDl/xZHxaBqKo6XXwzxkSHc8mqisXVoA5Y0o5PsCyrZbv
7X0rCR5BYN5RRa94besITen0zuckGRR31dPGbLu26JYCXvXlotfCjFcz845Em5xLuGZah5JRhZ+a
wtnS8XolKRcmogLwg/oyUL/1x8ICbV+eL/AcvHzOhkcFUISzqlQigY4QXtpl3GLHzR6NOG4a41yY
yMbVHBidmycAQe9OBlZA+2huRAMoZYoJg2lU1l1e080UY9LynJtEJMFMDiQs8wnPO7a9Il5JEiND
Qs+9NXDJdeRAQq+9vBdKyKG4K1hpHwTE98kFQZjgfW7RMVAP/1aR8e4saytpF3KYVIhA0gLfY9zh
RyZ5RIp70PYbaa0V7XmYqDrzKDKS6R6S8K/1fnGuoj2lcfmTWHcaSEa+raSjuxDm65iyc/ck3eWA
XrvA8XWUt4JeRLFMeOvKVi9S+bO1YsdAvgl0M8Hz07jW3d/7ffvJi0U2HW3E2RuM70Hb03HrSMmG
24fRxG6qWS43oA5EGaE5jCO5eBmIRu5ijLJSLcPCG/37KvrsjSwFq1pTpqlSNsVGpmV5EcRTRRpZ
L2W1Ugc6OhhuCN9Ak+xMn8VYl1Hbc3axyANS9c41afuu4/K1gJOil8B7fecFViZ5MiBlqPTIVgWF
o3IjPSWUrChpEH94DEXxao7Dla2DtbAlKluM5DKmENet2BNNGHX7K4tydgEdUKi8sNAaLEdw3Ujl
VSjUoVW4dKkmjbNsY+9G8VluTt+WRnm1pdsdiq2cNI+uM7Hg8zTumo/SH+Sb/qnS6eUE4d/0vP7F
WEtpmAK8k6ny6Oym+q1dtBjFxrUBd3W5qfvW6+F2LnAbIpJxLcAHqFE+Qi50XwfpR3z2qPPeC82M
eVDWuu3AisorI+CnBgrT9VzmgMdOrATVd18duTdqSN9yx5u/bRNRpWVrUsTSXfV5R4V4SmzKPo0j
qHIGfBUtQcRy3pHn/YnCW852lqi//Q55nXmzGgTzEoQmonFc1MD0RLFGrylLqvQlKw/zm9WKZPU4
UUk08cC0y2uasNApzuStZycJ+F8bQ288T//LJiCn/eBmmul3EZf/C7QtO3ZYCqle8ucwE2285hRs
gdk/OSHRyTIeZN8rk61AAYMKVtq5namp/3gJDBDNLOa+NGlY8sb9QXfUdJEccc3lluVkw4LpfeS6
nN/T1fxZ8Nu1OiCTr+X2rXjWBH8du/jPvx3RUa8KQzrXXwoTSGvSBBNTQkG7nQipCN5+uu2OQf+Y
SjmZ2Evr8m1FPIvK3a+PieHNi+9Qay719bplLMVsKCD5KpiiRAXGUGfil1dk8iWO0OWUZIUD95g1
v2kBC9ONEpJ9dETrUNvbwyphxYVgufnhKMjD+hC6MDjtM2eGSwYm5zhdmN58RsKJApO+GS1NsSKp
H3DaqG+6NgimwBK/BTUIUJbydaNOjG97wDmJKV8xTXNDrZIOs+r2GbEsEzRolw5WXBf0OKc4v4K4
zFd/Lw3kOaCejt5H2kCvRCpFFe1Kcz99hpK20sIQnlFcYZApx5rPSllvlSd+eomAeLf81XmriVG5
lEy06jeqp/P+TT+JDrs0dUGSKEj+pIty1cIeFyOQHUFmS83YekzfoTfz6QoQ8dTjAIYgj+RXXPLp
39Ud8ev1nsmg2ytSBepGqSjjbbHJbzkkaaz443YO6s9wZhgO0YxW1ExHweq35uLPU6My42T5A6ud
ewKIYoJj8XRMP5lOYfGW5nnnA5rkxfqD5fTyiKa3D0XMod5YFan2Hr021cQ+F/q5dg1IcHFrv5qo
R1otf39DFheKAfCaPdu+rHTfhNcRRdXnWugOUq/mO+R6FbwelrW2190Q3sEYpGIebEU0aKlV4N+I
KhEm5ciGEBmlU8Hahfz/5I2aV3QK5tuTKoXPnIVJidIkpB2iUzwOmr+IGEEYsEIYBQ0AT8TzfvDR
h8qhAY289OEV/jMEqeYqNW5WPdhl26jNv0LIl/Q0jgYVyC3P/KmHEzagIX01RpM5Ed+ynS2M3qlk
w48vrbmk0iktVtf+jcctSn3Ccv7t7tG5IFds1mXJ+uUPXyvlghsoAY2rDA7blhxSrRlAHlpZB20q
XICl5leOamhXP3mw+YdO99n6lWwG95I9tWgSZfh1f3OguJtkAW5iHYIDE43mzY/aK39GFl23s5KZ
iq2FHXPhcIHUJfaC/8ZKI19M9h8Nr1+Rfw3l3NrlRJVq75KjsNH2wyS0DvxCr4qy++GWLVbs0QJX
mdFtNWiBqspZ8UdUpUdXqpddvL8ZVIb6nXJM2UFRSfVQ9vIPZv1Vq/HFuAu4iem7nXkbilGQkBgj
CvJR4NrMWUgp+s782IrOfSpThUowc0T2uDd9f8VdEnEqf4lvAFNmGA+/EaIGEgLdY1d541M+aaBI
ze/cFM7kdiy4lcJfEk5aAGuTSBwGQRO3YxzY1Vz2g4TxaR3YXjQ/vH27vvsTJGvz6CIlfkQ7cy0m
z1+z4minlfluL8KCy6jBbLizn6EeOw/OYI8LT+LJETCjtbqj58JXep6sY6nQi7hje/dygBjniRGM
WFzE7Wt/gff04P+JK2fvbZhCTOVDRIM2iNooLrq/xtcNXCkAQwPVq/43KZBnhyzc6lXIDeURTDBf
50prXhRGh8c9bQgQnxMv3Gg8w+bpRjIlnZIjWNAM/7kDiQCfxccrF7Y2778mZ5gWcm6LJTZX9JbQ
qsGRLuh6ALhjXSYoaROvoDR94Wv0vKGwvJgy/GT0Aeoca0RM1PEZOCgVK317FJLMkqvyRbu2twKa
Lbr5/qjqns/KemAjJqVQgX78H4Vsi4ct0SOZfFBD01nw06TRkPjFcz/DMbaM5MRCm11Om302I4y7
cztXhAoP4PdR8Sp3K2G+8smEYqJgB4EWgnfDjnEXCyN2MjHeGSCT7AbQYotMkJi4aT7blIRARd8Y
Io7p0vjs+0uJdlai11npw3ATFjSqGLg1u18HYPKwB/n4Jb7fsvc3dj0vCeQhFLeKlyglZAvwY11r
VdfP/EQQUJsUFQMfIwNT9xK2Or6q2ZVS/a352p5vCtFKjc7g5tTauLk436rUnoIFAFcKTbjdKU+5
oqqnUplBja5Tk0T5sivdFDafbTjachr5eD6pSgXD/7p/ypK8L01yZZOatNCr8eN0IEaXLLu1nWd+
O1+z5A6qC0zNMxNmAYK97x9wjWsY97xWgXaIRC8vGuYhKtf3SA/eVZSCWihCrXyMW0ftv1udRU7A
oaePUWS+3GKYadwxX6TMxW+i+eo/HlPhCOHseGTHV38QYCg/3amaOy8y6ttb7GvPp3qcn4RnOB7j
J0pjSoMBy0nr4mhbzuktY1k0iCW5ms/4nvbA1c3h/sewt5NosljTK532JqHauwBumk2ldP1mH5cN
YdeDdXSxGyNBRW2X4jChtc5zUaxyD6kbw9Jy6/KoGOTMv7JEEpNOxLOZaXhMAdH8Lnxw1/wPFWcl
p5SxTjCeCiwPYXsXPQzTUhOH/smMiE2pK6W2YB4672PJOzTmlIox1AtusoFc5ah4a/lY+FRmsiK5
B39sowdARAHIDYcAIp2cTsEP8SM7q5/Zx2VNpHBR5rF63t8mqx6sbQYu33qJasbLgPfx9K9lnrur
fmaV2GrAD04BsKjXbCfalV+3b9V2x5azKHGNEG/RBjccsBzoFdFhwVHe2/IDozybJbawIvsA7Ce0
+/9sL+CDZ1WulWu8URTFhgltDP/bzJEnLSC+hX4uURETdu5dMmaZgS4IOHtpJlqqhPnHn3gAyAt9
hd8V+1lbDLsrRA/pnkRU9rIqxUMyXle1YWx75FE/GgT0AiJGx7swZtucJaUzAxZup83JIOj6CFLX
6gqNVhyFCqfVRDTgb+VtJTwXlPgjLQdKS+vxexmC68lsiF+mZ8VKR5OYVW4XKhh4MESYe1uta0C+
O+BLgRoPNQLrE9hWSJHTYkY+xB9v+tyokCu1TLc/vHX85QI9HSr+CvmwwbeH7zkvQfxu+L/KdGwy
fPdEsdKPa2uhew/URSq6ggwnXr5Mvyd8J3QA6fdTj6tDv0Dl17zJe5TG/u7btd9JNqKNmln4dS/K
a3NWTgzxMUsWYxi4t9pM0gj92MIAs/D/wwyepI2CvUjTN9G2SbGk5or/F3ubUNlnLGdkJli61vja
YvC7p5s/1KCtr+irrhz8Kr4uDi2JlHwtpR+baHAfViT4wj2biM3QT8+vXfdNeWFoCkX5//g+YbaO
hEOTM+6phTZ0OXXb7IP6DSgWRmVHCnYlsmv3QfrPEsCU5E6f9S929HhgyxtY3p7D3GESj3H1PV3/
7czhUXe7PQhQDPlx20KrsN8hsRQVwqAsiWYKVXCx0C1CtnSyEDQBlKqjOPCccZPElKGmKg6vUYGe
lHPQt68cKYiGObePaF6d5ThCNR+j4XhwXmA8iCY65ca8CKVSE2K74kpdO0f4Z8/CLkAF73KdBz7S
jTgQpTtPqLeaaALrA2rIqA4HDqI0jg8Ru8/31HCsspIQOljV8E2PyZ/RcFlM6JgGEGmw1VQgoKPD
lbe4k/p7+E/RscJugtDMqX02TLSOlYRTZgp9UEeit5p81JYLZPcUE5lrv5y0szu9GSDNy/yG/6za
Qs2ElfZRS/HIoQwRyiLRaad+ZK1uneCXHG2dwP+mikfMagsluoIK0fqAcyWOkmcpz1QdRprb2jEB
oBvas3hZnSiO5B8vj7TRdEyu/BE1CJIxtqKIam1bku2a/Quu+oPYBXmq0CIzgzZz3SSs8xghsZzD
622DYOmtf6iYbb0+05wr9QTdwaXLVQ+mzML8Y/LkpsPBhIlGoBeTIL3bkOHsXI7HDVrJhptw0krA
/3SmG4tbGbLdpklpmt12al9Vumt6Pq2neirZzDfHr+nVUs1YswnvDxZ0Z7vIigq9VelhMYl6IkHJ
jJWUNR5t+xagPMCVwdw5cuwLuatGazNl0uiENPwGhYdIdnK+EsVY/MUNclDtBMQVhqo84E/vARql
v51DzENO1A20WSH39ivezBPYiFN5CoNZjjzFhkWfCV7KKtb4SC9KO0vrmWkTNdMyYzeytuE4PhXY
BR1MHEHXH6v7b2B6Kgon9TYbM/Nd1gznmiSImVVQ3n1AeHU/KMAMKDGI4ziaot7pRgKgM0nmO7MU
7vQtuDcRunQmV5fa/jnAYUnp0zCVocieeSQWZXIHOzHRbvDYaUuLKIIw5K9w+dCiAi9S3U8Wxzg6
sZmcdwFucz7xs+i8jgZGJdMU5JOeH+m5nLFjNCXq6lTP1XP+OzF1E7c4gJoHuPk2cweqDIf5SPRl
PoBC82MhEc9TBHRxR6qRfDRm+kNFTHCeDXRtKFwew/s9F98t0a7crxyC8NQcWlixYXafgzMteIuU
CeV8Vxz1IGz+pYGqirW2matjGBhpvSpvZEQUlAOo+nFi8tgLh8gMj73olEdXeNf5w8kaisYgqdiN
EEk4O0mSsvOOMt1zSx3D5HPq+jkbJF0SqtCv/MwQYwDYWl8hO/JEEFOjb1Kk11KUbfHhueRl7qN7
wLBdEgC1TWHzeKr7tnrIywaQBAknAxLWIt87ZYe/cfKyla2mOC0sUwdKA+83n4wQJscfRA292IQc
+kDRfM+SZZu14g2ZXCjIS8FwzKaKt2lEC/r8PYNZ6KekbueSEIGLk4o8dSN8eMEH/TJsa6FdXmqf
sO9olnFx7R5lf1BK90RLbch31/K/iFYl9JIjIK2QLgGXuwbDHmSDvHquXiLk70kcDLO1X2Xxs0vf
vuTmqsvr50HI5WvWkeP4SQE+MbyMfAmLEPu7FdcHcGZdWBOe6kljZWkG6wHRkjfMFNoFjy4uvx3G
7k3PyFWuyx5+q5cuQfAqbDDmT9MXLez/Ra2j7g37C5IvxiOvqXt1bH8vQTlR1tFMwj8O3CuO39ux
929+ryF3e2mjqgVcGXsecLton8XvWjBnXuWDWu3y1pu0aQntB2e9CtVuhp4KeF67CMoFOZSsbgFW
zg9CbFyM/qMuYZWTRKRUBLIHKsfHQQqNYipZOHBf5JqhtrnbnmMA3P8JWVgKWNgZQzn2FzBixnqT
KJLDXplQAe+RSS13VaKe4TpM5JS43bta/oflB4gKFIyKwUHeTIJ7mAOL9hFOqSoHmBe4uod25oC8
SUDmu95kOOP0/vzGP5LAa3pKt3guazhSj22sxnhoyhaUxJfV55LfSKGphdp7+ivRmVo3l+w4veZz
gepNp4VYEW+B/b6LhXVh5vD4sh48ijb3rWX5oLqSrU/IlHQPl9QxKUXMbpGAL/xA443BT6TE/cO/
yfZsub7sB314VNCnJxH56xfrh5iJg8ay335adZ5ncqeGmYJVpylFOaGHUG/WjWyZfgc+VVbuJys8
2aVCgmigpCWnpROi2OwKsyAMbYONTatnLWlEJKsX00CsrOuiDO/RlTYUYFv782XKp7NU3MplfdOq
EbEn7rrJ7VMZKyPB/OxeYpDKRqA9MxP0tw7kBeSv1eEXOPw5KbJgUzV3TyxjgyNP3A/y1VPHtiLP
BPUL5amGi/FHbF6Vk7aE8zZL7owxV14YM0D4C2od95XtTK6v7Gr5fdnv/0fJ2YULWD5mNQZFDRbL
W7mSrpXkE94JD1w9vviXb91xv8M5RRhcuvesK08VaQLNNesewLxQtRGzMDLjdF8pOHvPbFKNBUVB
144pfGu1nfzMKBL///K3Y6fG2aKcmARc9UtL5Yu18jbgshfDO8jAEfks9ZGae4gynGgZQAi9aMLo
D0Rlid/2BpStlwfKaXKzHxTVWo1R8WhkKjodgPG48TjzrKI47E3t7DcUGqD5KWCEQr1MPnZJlfp2
G5mqHwKFO8ifov4pRS0Gs1cXTDbLe+UoI9SWwjpdbb87QZGXkH3OKzrkaZndACc8nuLl5/8fKTmc
+i+BHmN7TFEqCOf1FbB5S+6dbG2w/Vg666eeTHV5nBST6vXLAoGFjF9BuvC/akd5vPJvSovhhvo5
ACNMaCaFCAn2RxQ4k54n3a0pGvolKtNBwYh2TiWVmcs9T+iGm8JsLOWglGVygxd5tH2E194LhjVD
4Z+7UpHo0mlw7+B5V9cajHiy9WRX2dzCqPW2jC8f2AwgjMAqFan52EFZEzxcRfatDy7HkxVPHo+K
fYccMvTW4ZX2bV699GR4gxcPDySSvcfnFtHyEV271C5xhOu8v8TEFKwIiwDsD3HVTaATQUk//nYD
LK06jKnL1VJBZW+wo6BDgw5AsFJV6L4WeEoGTF/QvO45GA5KNYY/oaCCqbsvpGWHRbO1irf6U4fd
xUzvitJH2XtcXgrGbVqmQYcmPwvK5is82K77GXOxZ/Sb0aQbH6IWlmShss+VWQ4KKbo6WY4ZqfpP
7dwSwdwU4LovJkjguntg7V86S3ZgsfTFZCmdD2XM7It01MEdrFY8Fme0Qp/n7ETR2LUGIJHB1fKu
md7zS0LhUAFw48jo9O9tmFQHnH3h3zfx6RbjMIixs7XD2Ncq0Tqv23M1/ap5nK/moFCI4UAA+vcP
OSvD7dZYvlBcdDtckc05iFN9MnPlYYbRA+cc8uBFUh5j6oSwxP6Gf7X3tZlnP9rX5oIb04QlG3M1
MsPrdIokJa8palhMHw1q/fq9zd8LUpoj9V5jLpTid9uBf+rhEs/RAgd4/yuVmEBRyeGXhc2AkXK+
ZIwh8EDzhHvxj+Ebqt64+9EDMAfb1lzzrcGQ48km4No044HVO++G/dDuOufUDWDqBiBv1Gk+Rl4r
lFUQ89BC4b9YDZLptROUaOENQ4KqP9A12N5Ce4JClv62ZenYlPfRrGSuAkAMHe/yQq7DgvgfSHCm
oh2+AAJ/3oOYuyJaLqRtWUJnyJShMD2PcHEXdQw1RvW8WpEAoiVYmeDMbHXfXrSRvzYGRav0e8ux
QxBG7sYAKe2q9wG630LEhNaB5D0cVydQLhq/5MyqNjAbvk+uiB7XWJ1H9y0c/3ylyO27fChkJHVp
PSq1FVs29l4bR8lMWrYwrzFARf8QokvrhLOhxjPC/b0pHBQbRxsJgL7uAyy7O/4ObservpElKOhl
5yZEWyhTtESDKV15Y/knxNOPTLSv9TXQ89GkF8G/IoEbvTBbxCNKb2ofROUWvXLc532McFsenjFR
tixYttxq6L+hfnby2IIih2C/ScD/TLTxBkr3PU+qoL1NizX0sPy1gvnlDKyjYdnRTtjiIrR6jGQz
dhbEgK54ie9zqwr9JK0Ui2VUmXiLlZ6ZNORTXduOwCx8sSiV9RaBoUo3vV3aHDwHKjaQ9BjF2g+O
Lt8AB3l2D/xh809TasW8PImzg1pQp9urhlGYzFCyvLp79gRlOMA+f9InmR9MrgGnNgwa67sBvAAS
mj/rOmdoMeZiZI4NcTInxBU9MKtGWfVVDST0E8zT1lfwXY4XLhkJNDo2DcqKDiOglitWIdoGOrVl
0I+c5cTb13ay6Zuekb7kit6ib4qsW5Tazen+HDgLKBcGVVOyQqLpTTke31VREjirVnD4tbzZYjJQ
tjVw0CinqGBQl+nx+vjRAyL8CAoQHIrkdfPmVkg3zLd98J3xw6RsMt/F6pIvjuFzqH1zpEEoGJ0N
L47E5wGnD9IZY2Y1vWYg1HwoW2mwha0wmQmN4JMglI8wGg3TDd64yZzFV61kVeqm7IWXglpCIgv0
++zEFNrpN77qdjOwzYQblx6TviabkGn7Zbon1WHR3Vuit1DkLLCRcEM5JciqMbQq+Kb59YHrPI48
7VB+t49Tllfxs+wU1GP++yANhmVNFoBPBR+7koToDMPA4/p3vaYsIFUUW3TRjvLdzDdMqG/+8Vio
6SqjlkxsWXdWn2RVAAPc9iSmAHLONsmJriiKYD28/f5F3BlQJHpkseBKP0JJ09IBbUZ8LLCUdD2k
ANGIfUoq34SsQ8ILVUC1ikxsKc3sMKilyxUpLFYZ39f56cHJqJi6CzjRvCl5Mm61D4nXqatA6WZ3
uzjxrOzyJrbkKW4cBb3t5ySjBpbgt+jLSAbvcunO4nkVgkmtZvxUoBfqL1Rh1TiIVX6OUdRulm7k
kx/PVpaQkecVN9IZTu22du/ck8e2QO2qNgWPBz9TK2u3Rl1/laMbchFbH8hWMAFZ3qxsXFTIerOQ
MMrTeWIzHda//NMAXeONdzmBxcSRAjKJX10t9tH/+wm+wEB7hzv6CYV3FUbZ8DDdVxTS0dB7ZcGJ
7NQMmDp7Bohd+lyhXrSwuN45Wqln/WiriCOApuMPWqsoDmKdRkCOwHOSDKSn8eZjGZqTnA36jhVl
vHNffkppHEPH6FU69e7glELrhYY+qlKEljCC0OhqikiPP29pQSlUPPB1zbtnx6qE8cpR8UeM2azL
AgIXx8Q9BXEDOEf1f9bUAPPoa6nf4ewvFaJ/A/gdGuxvkbvi0vPqMGCWSo5SmN/GnLSWXOdi7S/w
4bkGXKn2PrIgTzeMfNbtEAD6dygncTljoY9dFds5mEOgXjFzqOBGJUYmvx3M3j4DPD+iq0Tdk1RA
aPVJmAuWjljMaH0+oj5VBDP6xbKOcimwHOuZ+Qsl1J1ksX82uxPrgFyG45SVgCQOwFGVH4m/1FoX
6w6WqcX/zl1p/jtD6frbQsOSg7C3dFOeRoR6+m2RPzhPt8s2fh3QrgssOWq+kM8V8zo1E3ZJrO4D
gkRh4PYgl2HJA/si0me+PUBr0oH+T9Ga3NVtb6WfQ9N/qUXbInM2cNfVBf/cysMdHBGoDb7q+rb1
16f317Tbh9Rq6r4FGef6iXzeq+kft+PcBcS0HZ8PMcQhyHmCizSJm0JGqAbGUl+TO4mWuARs09c5
62hKcVZkVLsYji51HX8RG24M/TzkjwinxCVJ+pYznuiRsGnpAuZG9DEJIWDMAgHOZedGhTHco8Bs
QAJEmJ3kbme+Ydf+k2LiX51DF9N7OnUez67ccjQ5AdbWv6iJ7xPK1tQHDS6zucE5CLDiH4D36np3
mVNxc0ICeCi+XciBasrhf6sKp8SQooRWfNKB9UxB7RXIzwxVTnTGp/cBZOo+Cizy3cJ4m1zLxvfr
abcoSfbXO/wns7XQeeoLmTdAuPLZcGTUAL4ObXKHLRw/CvAwIr8rrav5BcVKvObDvuRhknHbcN+N
n/KGY8MAQTD5TiCKE6+OZjUQC/G19fua2AK1WdEhZ2x7uhFvAz6PyCOC9BSFUwliAGvbsKTwoSvx
PsZzSWSvL4hiX6Kw7XiFXYDc7XF5tH7kXnZgOHXgLl1qaVPpn8+KemnKk7248JqwJwQSU+snLSCm
X8HYxeaR/EOevZbkk0Nl1GIzGZJl0e1hUua8jJ6UJiz12TEX3Vxm0G3++rOTI6s6Iepk3XULYGAU
09Hhk9LLmvTjDz6Dv2hrYsihnDc4Cd56YmWMN3Jx72E+P12GG6a4Ei1nzHirdeOhQwcwcfryxvra
oJDiXULhfwncbNdFk2nyG9JSvqYZWoFFLhcMtScWgtR2wyg2Z9t0K8aixKqEG60GjrFUDkzTDW/5
ZzDCZIOjWTQo9uJvCnOatonyOa77gQxEBjRPHvyUoFl8Pg4H7+x3XhsQO/A7G4l2X5oao3U++vdZ
BIUqn9jgkjeWATXE+xV0HL9B/pI9G6HcZdYi6NjZeKQvr4LSgrrTnvIcbI6Tb0u6nvScTb2VkWLJ
Ond5TH6X1gqyRpynWaW83IUNlUfnWxhIgLVUTQZgMReiu1S4qqfUXaT4bszXhXYcnblI8PyYHKQZ
KPJ8tRCEwkUqUkOezkf9MWIFHoUjlpabVVAQByAe6JX6qnMlTLusyJ4NfPCSA9Poh7AyNzCLSMWW
it2sYVwsMSaBp07g7XCxC5I7NCmPHDeuvrI8CPHPYHEYDL4wUxfpvwCHeQGTPoQDVBgB6QxD50Zk
fZGIhMGnQxbTyNk3zGs7FLgYYurIvEyDFHgI1QEYsTuUkS/nIPsiOpE67UAEbP6g4z4Qd0kIwlOd
wpaPnsYyq4FxSeRQdBzwdWmj7i0TsnJPaIdIQ0L3BfWxCoet6Br/tuse/tH991TuemPFmMd8JSlI
KRhn0bIbJYF9vVK0Q1thNAHcjaoyZudsaAgQrjeKm1M2dTRkaUV+rp+0khRefLCeVwIJsn2eGiUi
8XXOl+3MSsgcY3seaAuvzlIwkbU0fyAKIHirIiZhzMehTfWsckTHnAUOgjlsU6toJ2hqXMvJByi/
77gq6idJaiZmnteB9bLHmqFXxJFzYnbgvosWTY8VFj/Vukb2lIdGygI8VHejzoPW7S/wr6qwDiYM
C4pO6T1cbQ9cK+Sm8JyNrylDc3D89fTzCSXGTQTQwjwrUu4qkJF9KEWGbE9f+H/nDxBFooTRDZnv
CCC9KXAHQEu/5s1ckNIXmI/DQUYle/HmcWMU2gbCSf2CZlvmKMfUVISWGurZPKcGUxo82I1BjLrF
iA0xkLPErvZ2z5+Ouwu3gxOsH0HVNzTk/ft1o+28sn71nLIX7RafJD7BaEPKwIpOxUE194oqzooH
oWjDNvlqvN83iKAYowWaWkYZYel5PhZwLT/3SqYjXHgOzDON6RM5ifUOahoZD7JqYyc0A4rTce6B
+9GhnxbmaKujGTaPC1HewWUXJOFUTwImSMzkN2g0bSIObCH914NfxYOvL6Le6NqxmUCN3ElrU1NN
8h+t52SnGmxZrBugp7PqFViLNjUyt4hvreGLV4KqLxBbaWx7SsJCcnPUhPs50eGHK4d6AcvAVUOF
bS+bD8blB3xyqMuO5Aw7sxDB4z0jffJPG+pWmWrTEuFJOhkfQuQ5l5AV/26tBvJpALhtA3QO0UNx
mgrMZgiU1gVnVEwMrPsJhZxUav9o6Tw4u92oloP9MRrHJJ6OdEl8G+YGU0VWujutqb7lyTXdzXa6
yXw5KzQgjNPBXYUgQiAek53PcMSk9ykqDEagEU59jDQpQjjwYbXqAbRoTfhN5h9yfcByqIFB4i5L
BUUfQ/3q8qoZPo0j7NbdBAqwItMC5hsFyUMiH8JZCGX9h89/5KxRA9Hq4ZCG8rAmOwjzHcvt4wqv
80oJbg6/CTnTwp6vS2hwgQTQSfEN0Zj8CRKbWuU9Vanr46izmuNZOELjfuxaKhc/y5mUT9WXXvRL
tiT+6tdsKByxKTUmhOlU5DvN7Ktfw7i3XxtS0H71kjT7j8ztYPIKps1MlqsDXJ05HsMtytFGD08u
+aiUCxmuxs/kZNfVrUD9RLpaEWMf7UWD0whe35fo6Z90G/mUPpzp4S0VEjv31MwG/TCpvUed9RCM
paLxaWIAqktxh45ckrRs9jgQEvwK5RY4x3KojE1VCp0qUGx0A1WLDTvkylMF1ZJS9lN+uVGh6ysz
Gny6kUXlJp/ChCnNVUfCfzgMF6QQS1oYw7rQ7LeIZYioOpchcABAxTD55rkFG26LGKRW97sJJqdg
zyq+4P1uINQ0ZJGkNdvAjcv05NVdK+raqj0qWYbTzRqdby9Tj5l3VMNdkndPpFa5763FW242cv7P
cMwX79cKULVnRPnSWT6RPtL1sZ6TEhpLPLRQ4yFtrx3u8e8LntNurz/V9Xp9ZicYVRsD5YIz7VC5
8U4b7RXSByDz5ge6x2PcooOYn+GQDUom1Gqimx2IBqyEObZJSJz9Zvo+fegEa9Atmu0XRvvlWJ1i
oxq6oNBDplAj946Ih1j23rK1Jo5eS74oWhscGseOv44rvGr6qxhrpbSx3KgGCS4M0aP7U5SuMeOU
dSsj12iT3zdUg4UlrPuaX1Anzc6HkrUcMzkafxmGWLQyin39GZQjFe9L7arA0SpNis/Xw873Jz8k
YHvPVaHV2QL7GmE1Uy1zHeLHEK5trYRzaZBIsfzXEHkxOOePajAjjZ23TODIgQxrhp1VIzkIeFG7
eReoeAKZ2nYfte9ZQxbP+Gr7hwN65MoA8IJu6RitYsYT/8vXRgPjxRVHzvUmeA93nfH4ffPKVzlD
LlsbSrCJE75CeP4MHxWUuG8lhokxTASqO8br9LJNvJcl/kNraWucMtHRzkZaPjfUyNp2c61lM4au
nUmHqWpP6kHC1VNDHxZG2heycn4CuEKhYKqN3Mo6pgp5zxm1brr5F4nj1xYf2T12V/MCZvjrrwVW
VIKMyTE5cbdYGFWuB9ocAhCKW5eygM47TwXaTDhM9MbLGdcVP+KrttRAhsxYLrbpFkKvpxlmFbmi
oUChN3kiJWFjSFZbc+8H1di/KNbfu1Mgo/Q3DtyCHpwxHEPhI1KJ/aI6En9/v0o56d21QAApZuE3
NlrVNf+yjvbssHxYFA4R0+93YMUK8vh7ZxtYx5Sq78gVHP5aL/xmcH8XuLBkMchasCo6SQOOEH57
nTFKYRJf4rzDyYrPs0swxCo9TsRw9ZHSHlhweontVtj9G7aFMn3v8QZIR3auURI41vSvuxRmolCM
65WBDT6u8E80k1RC2e671t1u+xPzmEmOUxVT/NvlGhOw7tBhE4Wan1tCRwhUyXZ2qOqy/GUs/c92
8iA2DkHF+4hh4rzJ2eDZ7RkiT/MWsUC/IdfSBZhMcJjPNuHdrtONGTPS4lZBcKQrA3KdihwKqnfm
dlbzMRorVZk11pnEV7ha94xYdJF24wP4574QJ7C2wo8ssKa/ue1FYas4l5NjFAHJ//2vOE9qFRlq
iwElCWjZtwlBfD0vnnf2ru+MagVpp5FqHj81iMaTST9CzQTB0hf2fkdH1twevx0UwQjY1QknNh2S
jIouV8Jb+N19johiHEV6vTkrWM+seWJDxXtDA/B/39dxkumAUNIz4wfgAifa3IJBQCLcABra8Epg
0K3B+HWBgsjjoojsMJVUDbVIOARt1iX9njpTEdljsYmx3JOApN8QdOnXzF6FWQwExpCHlGZDIJWf
PhzjXQUuU0mvOQD2Nfk+6q0zA4+twK2B9F+hWT+pgOy4cQUvxoV5deG0dNXmYVh6WaFlbwsaN56r
8v/xY1Nb1bi4eUrQQj7+DuOjq+bw7EnXYtyiSbUlCtvRji4IBFcMmK2k/r3OWNu5hgnEY2VILdzi
juxfO5cMD/YowfLkbgTJYDyhvDQ8BgYvAf4NFeHpt6Zbrjv5PskSzsYr3uoSgMm17clG/R25+898
JhKj6ZTQJOoG6uix53oiq9PZeCXKB6kahrQS9D0NgWRL8ArqbWT8cS3z/Be7lTGnixF3dxf5hORV
Sm7AyzwTjuMkwBULn49mz/yJzh2W1u9sq4Mz2IyIKA82iM4fky/nBfExm+pBYGApiTvNk3Q6GGvp
dFFrEJiRaPUe9EdQ6H5OIV1kN1XMXxtDTKdoSBS8bWEml31FZlKe1insGrbvXoBJr4zYs7yXbJ6V
gHZsvQ7MsGzEZi3D5J+Vr8VV8+noIT1RtylYMDnBi4VRWtXoEsUXkEBvOi8f21pGaYaHbO56oyUA
4CY6GTWf5kVK+ElGc0131oEzdLhnx75sHNaUkxevAb3aIR44unprp+EE3DD7kHKHsrpd4TwtoqKa
YiWR6FkIbzYCHjKv7sTPWA6eIGlSCUt0k11sNd+8G6lBMMbz5RtxTvxoPmLz6PwnuEWfRUrrCuHX
MyQabDB73MnSb8hkf8K9NnRx9BnthiKGb8W+5kIdiySWLJVgK2zC9HtQ0UghmBupRm8e+1u/yfQ1
K+QrkOT3lPHsVgGTtfAhvVzn1p3APAjNxi4bobN32KoM9BES0XEhd9X8hmwlH2GrRm4zFrzB+CHs
hjIopSHWhZdTa3gahqE94UIo7ZmA3RfCSK+9rWg89JdC7JLd+wgrV4DTK++t+JO07vIl8mXAuqt4
kRT4Ndvb7tMb2KKG/O/xsfqm3XDlJazLb9+5ZYyMywAmUWmSYF5LLecJT2EUttEP37esa4gosb6p
1SG7DzK0/oXseejuPMFsvTg1T18NOOrKiotA+Jf2aW/TENRMatKTmxkOOiPTby8SQzj5O9dk7SSM
NaEO9L+/kn13LkwvpRraDzcktMuON38dVcfEbqA3vPwe6YRmtD5OK3TyVQWxXI3GBDUg400mdYO+
L7YZhot44KbbU8ut5DCJ0iXeaJD8wYXTRdA6OyYbm2ZU3kRN4f6QtTdijITN6g89zbxNrEYAUZeK
eag5xFxrN/uTUgDd5LZ8+Yr3IR8wRfqr8oj0ukUQFpGaqTMcw63S63Jh1f4sAkaB3dyDvWZZsNCN
zdZVOIRfWmEDgs85rjF2jQkGh8INN9CBsbMlQVbWfOWX4/lKl7JPZF1O9gnldCm3CKTc+cU3MnxH
8Q8rB4aOsMCmFoVJbUIfbibzxtVPmHP68z6+krWwH2bTgm4hYObMWDiFfpNRQP37LQP5wWbc2cwf
e7irtPu4JtB1vOeUSDUNVKXIVjz9CddfumkE4tPuQX6XLiAZDY49W/VmC8r/saZs0p720Wxg2jNv
EZ2pPK5m1NaU4G88fnRl0JAgHwIQfipT3Q1P1CuR+OxOxyGOMrZxoWss4dEFc6ptX/EX3X6sQ0ew
pVh4no9WcvHeOVtt7tq3FUwF0zdRd9laSZ5OZRHPZkvGt3uOXuatEmb35igAAXj6kHGzlPKoeyKT
XvlhLVKgMIdBhnRHWV0wAh9odsRoWpN0TVlov38y5Q6RhP7btjmwxdjdQKdgxdgP4JYcSS8qtp3E
QT19d3A3fy1dX/wf7sBQYIFEV47YGkKHoMcoqYVNF5cbsJAG4KhmvFIHDIcQuq9WkMIZhDTQq/9T
/96K0JRlRe+WXHnWH6sRuzlPC1GyixmHLlm1cAX8h05sNIwOYWA6Rlhcy4YWANk3IpHc1UmOrWpn
KFqQZSNCFG6lVxYlgUUDwoBWXID5GVPlCnX58SSWteNq5E3uO+8XDVE5iDY9VK74pS1Qgm/OkYXp
Gce+j/5C39/QS9JI/y5BKAwRFHa2au9eUJxT9d+F86TKtVepx9FFFpu0QLFE659PdxRqQgOqIgmF
aZLMDF5fpJAo6HxvS+pR6dmqoJiOHYhudnQTYJ8ov8LXFYCovxYHPfGREtgHPo1iESHZZLChL9Y6
LdiAQERRASX67p2uSh9dX01RMlkqpU0kgbV8Oo1VLtNqSMT24v1fFOBP1mT1K0YDu76Pes6sxVDE
RkC6RzLtsiShtGsDIEuMO6rm/QtzOZsTzmanWKS8i/xn5rATAGdHI7fRu99v+Azn8hJpghuEl5IF
k6s0Der0bTGF/SZMhihvK8+XgPEYJIJF7h4Pa3g9/dng0ZDjoaMMMJxlE1TgetSOPw62RiRQW+5Z
MPIFP3tFDlAjAK7sc8OPyXkjfBzNY2QqlPwkPiIq0Q91QqgEv9O6WDIumhQLaiLUoTNrGjOz8iDc
Q/lYkyRnxcQL1+A9cQt9XGRRYBP4v1YlYVoC4WNZAg1HP8exq1TXIFw1TLBM7UI5+ipeJMqXCndu
8sG2qsU0pGH/OAKFE/8zJPXXvS+AkfzBvWeAYBD331ntpaFZGtmPfpL+IIuQYP+LhD5ycH98Pm4k
XZ9yz5XYsaPHY+A1LV8TcgGGMunf72DhmkFO1YO8IIQFpmemvm+osZoQGrhXN8avR+BJF13mxyZX
9Y1+RJraxwEpzLSVsXB2gskD13wIQV/kVkm539jiCITc6tekoIdb5LlLO3DldG+JG4KwuHExNxvI
VHce1fZ1k2f9mzEtTFS9CxWx/pwWQypBgfiKFVb2MmCSX0cEmLMJTfSQ2SYpmhtPoY1NFo2OiVt9
1QgnTYZG5ByayoDcWskQZZBRPGqSTn9taqb592lN4PeUM2E9Msndl/LRaBUkgB0a+RPBmNR51Fbp
i5vBq8i3ne2Xuf5ttQstQEsfwksDVstwO6VzslbOaUK6PZzK45f8aZ3otILV1mR8vMZ8Mn+oyVMJ
vWMFo9hIUyspQaQI50eR0DqytkpuoAoIrfVBkhgKBH/cEjl5odvc9hrDE0Zo/c2uSoUhBk7MWS1s
aAPMMZMpdWedvzK/q0TFjqv1Bi1YaSf2DsLFTuVNmeoEHio9iVapZn9mzL+bnZ422WpdWcQsqd3t
VMA9ensbux0I3atcTC1dVyfO1Bjqf7xZ+h+51d085OWoQBz5xujFMSDo/SSJbLZgDG8edNqLuK4w
5N3We+h3wh7va78NMXH1ESur/n3cc/2RYpDf8xow0hUo8tIWnkhX7mLGe9qD76HFfgyclzft0TCk
pnQeFbwwMfe+2yvZeaa5rpZM1qCV0OPSOencPSoAsV8QlctE0/ucWhrLRaMIfiHXrLGcZV0duwsM
zof3naWYgysyuMd1AqG1Bs1UkxqwhZwDYlrTd2teTXN600yxxdKjzxIZaKr5GUHdrSCERLg83fcW
S1vQJA0dC1ZggFK6SySusN9anZpGnPef3ic+keY8muGsVygrYUjIORrJbFvhzrKcZT/FRNkfbLpo
tPXn4BC5xnXLI2ePxc3Oeq7KC0jV8rOQE/jOnDGv8yw+BlUkOxW6pHklc/tJIx01QVRCK4hNDv5M
5Xo3Xn4eEj6B87TGVfxHMwHn2YGPWcx3TmLP2RiOIu2dFnuglwOVWzRlqJv6qW3rb3Ini0RNtcp9
rYNry4r4itKyykSyjYSEuuSjlv/DDaJpRodeuKmNhv8/rW9G3JsGJPZJrXuNKt0FhGlXggwVLJlP
qIHx8eWYCB3y3RdNUHLuAHnZOJTQIZX38d+SLYNnIr+pv0lyOoYILwHJ8qq8qeGd4JUQYJ/hUtih
87GoTiKdXp8qCJcP3VrZd5l7XfqPzgslb6DvX9EuAY2U3++Q/FKmCVvbiScEDyxAi1TRV2Y9wJwW
nRf6OldoNR3GTR8CE0V/Q7bPfJ8PAtr2Oka6cLvE8P3dlbwKsTiuw8nyFEPN0vENteti0A9p6jGJ
SoQA9yV8VSGICFKha7n9jlN+nkQ+vWzfEj/LgW/y23jY1IkXvjDX3G5FiCIRk8nJlr5K6fuIsVwl
wo1rzTWBXHxiMryQq76RIxAvCRzyxLaAvWIf95TwJObvHNL9OvIS5+TE3gOmZacXnobyuqZ8z5N7
bgboKrKIGI0CratqLrR86G6NF5qE4WMWcSK36TfeNG2/np38gidC5Tjk/mDnITQ79/ooXeNTKnOs
BEn/7mjXERirUN2rfS26OZ16im01PRtvjU8tLrTvot74ONgSkEA2j86iF3ZSnE8irRPdEnHLCcm2
1DKNEqoHzU81o9iE7njZx/BwxNWiw9vgczeJov8Z36T4Qwr5OPoH88GKKEaQglBYlKAtwYKTkPJP
IPKxwyMXrEPNxauJ2TMCZmh6mnAQpv4wdgHhsCNcsHbN4+4nIWDaP3J0vLrH3CeRw/xjRZEF6cSw
+sAklKvbam7QxekoBENJ9UwNSAVBNvJw75/Wvo4TUnLTolyvWqUiX3pBbno2nS5EuyjpzHCUWcv3
sT9qj0w0SBC87GSoJOdmJ025SUtOyHRYX6/Tm/41/qhALjqGAzThMi7xKyuyNTNlbYpdye10rKmY
HFvlCmdZS68+/yyVlHsmyJqv0QGgOtPicLbZR51iRoHljEEXTuA87Tq+1mKsdE6M4INpDh1Mg5xx
p0CoaPf9AERky5pziZWa76y7e+x9Vd9qlplDqrob2969TOVFtW2f7ANFU3lpIgChzuXABbmEX04H
cMYGs4EH/NJAjY+7ie1vPKb8omnwaTVYMGIrXptGdTt0u/IY4METPeI9wr4cm68H8Ih9+oroJY13
GSm9YXcwPBkPMyIzbRNWwnrk8JNHrGtbIKCeAexaiZjkjjYn8M+H4uITpX3mSUEjyzEVzMFoo4BY
DVLyvDA/DxhCicT3PRcc7oahKx6oSCNMdqRSdXdN1+j4O2hqPFLS+63wAzy69dABh+yQy5vdU553
CCIfc2eROLEaCY9ZUmyTSC2NTQWcm4ugUKxiiwp340gsxYGlW23sxxQdtDVgg/sV4f26ESX5p+d/
BgQCwKVAoO+dSbIa19G3VK39PBvMFJ1nUgkZaI59lL3PgzA6eJbZpYHrm3bhf+oHGI14k7B2O1Ao
N+da8Rm7V/p8S3qWBRYj/n1Vbgs4NZuq/77CuqZCIAXbzTPrZFjwMuAiQKbDr0Qe1GyhNnfVt0LO
A0p92b0GH0lO/XWstoxnwIQu5/lopWVYAxaKcw7N5Vl0/1WRpDOTyTyF2EDHgCkO96UBSyF5tnxh
3AHrH9bQztZ6vWE9xcEdG+EHSoAR4B6SnNnHnMP8fbW9p8a/0hxePh6Nor98+I4h5TRiJ5MnFgDo
oOEm6ipu8mzq3JW8nWeAlzEITH2QbmxuQb4x0jlrx03pg4nZ6KuhwUT2TckpUQF33zGF/euguh0q
q2h+JewdD33zamM8X2UqT/4sYwtY3U6dNZ0YYCaWARtYSDKqcfIE9BdrYEZq04bdD8eONdRtrnuM
nlcHH4nZnBbogkvEjde5O16CBsN7znrZBqv9Ben0sRx4oUo8SJ0M8sfvhcH05hfqG/q+5i6tGQAv
+tKOAJrqwSxBfZOTZhEr7/FP8HVKIC58USGCSbLMqDwIlZrjqNbwRthSc0DWZ/+BQOvtGzd77/Ee
Fa4tt/Vc6hdhgRIwDOkteyW/2ZGKSAi81oG4E4zsxaSYFl+i7kmgTyzOkwz5ji1xvlRz577SBKOl
2ci1uOILeg3j7teCMFlQ1QpI4j0X2x0np7QPM7jH89BhTCRgIIgHXxtlSbFJYH8hYg2qacExMUlo
FCcOOXf/O2tynmBJMf+PJihCC7tWWglOpXGJAirfZgHrMcAlytoG9B5idHLVtv0hTyrnOzGoELAK
B41wiF+uRvqomBD3mgFJz4r53mPsjBuoaw4f+C3GEtC8tfDyC7ZyCKy8yI9umhCpE9Va4HGKW7vN
C9AHI4VSIkJo8dihuApEYC74jPccOBjCjLn0U8TIYkC8ocM0kEfKP4cpxG999Ubpv026MhynptKU
9M1wo2h2Y2QNbuBP0U2rYIj+av0lVdsta/szkt6s9s7UM1lD4FCRbonIxepc6Jw1kqe8yt9wE9mb
qinYLuK7ylwAs6mGlkshucVD3mbolvAnaHV2ZfqE6IPp4v/L3vULNrHzIyz3gO1ST1lY7Y7fFJHu
Ql4a1i0L+ShtiywZFL1pu8Qk5QUyLW/q5FI3/3KnHJthJBMq4Sy/LuvIq69gnhhUKV4HZfvcVC85
cBKq1Bk150xhcs1oz9h2+aY/z4XQRJum2m23sCa0Kel8REaudByk+XRVzx2VxiVM2Bf9a+ItjTtZ
qWq+bYP/Mrv88VWpDimz52F0HM+2CdUT2ASNF/PvXaPJYiZx7TD2PSsu7XHnr1OT0Bhu5qVt475S
NV/Abm4jOZgZSyIUKCGOgPxDH2ACHRnt5kY9MUuRx82nigl+bJBI2s8+vGJbcO4gVYSzwU3dt6nC
L509rwMFXPP+LzFMDYpKuJMhnpghK7osZa3iEF5c3v8UDnLWbMtngPDHYguvtCJ0y73wPgNghYr2
gtoMvQCjf/a8RACdqnQrhqppuZfxRHT545BxhtpyL7Fo3FiD5s10MWNtxGIy956xL+uXUUj5aWB1
Dyfq8lCrnrKJufDaQw8+Izzi96wLoDxspM8n95Z9ibgPLtN3dYK9CMiH7ECyyvTxG/aVyvI67Uyj
RnJGWKbCKtzpakKVS/30Bg5lWGNwGulqF8Fy5Z/eiJJfwRavEpusXCpDc95YA8HahwtfeA43KQtj
mt6sX5pmRQZYNLkMkodMEr7dcgwnVNx5Ho7ynFFx+xpSUFS4J2kYxw9/gDOjnLiaEZQFcuyOsazH
UcQDzoyNfolAuhgrYJfYOX6Vm18WRB/SSGa2p+3DtCeuHh3rwXdfqHdiUpm41Xn0mzXxEoOoKC8L
5UykmVMzoTAahaIoYLsJfzyBsHWWMjVbdCUdfvpjdPnmD38waeEFnB8fb1EcVHYKbGYKB0Ag2gLR
xWFb5keGkwSa087v39jhSWQbgfLQXT/bcrBXRa+WIrFgGrzb1I+T050T0Lkae5Q7hhT1LJTftsYt
T/u2C1Rv8WlN35M1NDnRnlCG/bH0/DMx1dHTIcXCewKBQjFEnPOrEMAys4+5gKLluLo/225CcxzO
+U4mmqoy/QFYvEnHvWskAKXLdMskXVvildWRPBBbQNQIXRnLK1D94TK11gckb2mBwO8S8aYy7vjC
K9NtOCeUbnedxms/ji1wY7TDy9I7lhaRqgJqg9vchKNtPIPEclBIEJfykx0bnKaPqc3trR/6xfMi
5ADMpTa2sQkMJrj+SNMJSK90zcKSUyaU95fl5ecclm0Rbl/QAc2cS84lKPvRsJ1zK+KElXikZn4r
4ejCojsSHupuXjedIjqZZrTcpfsVPScPfKjy3Do/Y4bsW4b8LgosLssaRTh/jeSQLZCktyS2NyNd
0ccnalB/2Sx6NQeAG5V0IFvDfQ1nlGPRDZE4qbOFba22AIrD6pxR4tZt676X4qHm+vA/aXlf1Q6z
nui9KLQVLUp4qYr+7+n/JPNreBjBU/m8C3Q1H7dYwAUn/dPhMUx1SXE2hpm7Xg7m5UvLd4JmojGK
2lGpIiOrsQKXnCGoM7xjl233QHzL57b4NLJqWUjI682rP0GTtIE4NDLITM36jJK0KXCe005c3Bj/
xXZeC+yjF83dWlfskh8Su5anQfhpogLTo6pZjupjaTHjR0C3Ol0sWhftnCmO9sKkRdqBkCzAxxl/
EaO7EyXPdqFAkkH2Hw5RSXjHaOaMEkm6x+psqYfTrncK3ibVMBMCLMiq9I6Pqjan+mk5tPehZK4I
Wn828fKql7KtWypyDXrWCO/PretOdnvTF1197cNH5dYDoPj9UhPaOT+cpAzgRMcwVt8yWg9RbU8G
rws1toECbHrtHApdBiaNRJh7RSiGpZ9/MgAW7LaSc8qfgYGPE9zf9OqFj8TivuO8gvewTwOFQYRf
lTcazVABW05HZGckv4Zb/fLM4Td7LcSWxNVOVDpacyIg1oJ0Ova6pZqQTVZ0aLYPRBUKlbpxE8WL
CAI0kGAGWQpb41IXlMiiWw9XRNmUbbkTwg9t7mzTO3E2O1Qj6c5mjUgDlwvmwEOnIfzVFbyPQwws
9HumOzc6hnxPekgtMnJopYEJ9nNPDG3DR/PcJ4NHGYiPTjeC1kvBrDk2lcXOh7gO3M59Fkba7SKY
MHsHmqTurEEXCEWc6Hi96F0E53wWh+9ozMP1gegO9BVGiMGXMZ/QSmEuJujeTdoGyM6lr6N0j/lO
GJd1KwOfmQ9WzaovY8S3HsWzL0e/UpADagk8wtt5FgHVI4x0fhatoHboamr+sZLFkOF4hlhninJR
OpGvvXXAsp4wzCdELS/Z9N2zO4Hfb6HTXjLp5Qw3adVFM2fzX+EJ30PHKKCMGxMGhmlw4xvTXk7w
8xBDL2Dy8Z4k7g6rN/uYnfHL042Jzd5n9v7e9cP7OpRacrSk7VbaHi4dpLSedHOutiVNixAs2pxj
LhKYxxuGDZOcl83omX7uWc+vko2V4SjKRKOJXz+3Ql+BcYBtobeZJRuyIifSYHstht9qGA5HM6S6
kEYuwteBK/IFq+8Rf2ml07jdhpssM6PaMPy6lqH62iOh5OPmR7OVGKTQom345j/sVYRyGhazjvEf
VAmxPwuscFENoCU1BBj8N+1uIpKXqn/O2NRzb5o0SdrVE08SNuBo/QraiUQEXr4nY6SWzBK0wZwy
vVjKzUQSyNUO4tnRwdXB9duiLpliflIpeFgwQIFeqGT/Ll7wkkUW1Vt5mZ660cF06qKZcn2dMDlN
jr2j3Ut1IhqMXByBTBs8pLrTZTuXxO1rFNASRfj9uYNBAUoRG9ICA6kmxP2taEMXEAFUjK5IzGTT
hHWjp0Hs6yA1d/63jCjZYfJtmuEIYkxMFC9BFiw/tQWDzwK2rN2LSZ0Zilu/i0JKy7+EbtVtF1Rz
oXtkMppPxBcBYrOoTL2IGOfbz62IBq2o+59jxFq3Ci6N4AKmZ/jcUD7IEq8ujWBMTOa44/VV5+yu
GjaHPC2uhSHXHt6wF7yDGrlgHsTNulMl3xyozY+3huaNNB8KbKhUgb6KooO+PWt4eLr9OR1HRLEP
s/XHx2UryjQMa13e+0C4pEXoziaOiABWMPSuxdfeGejE6m7zrGPIsH8djawVH125LW9Zkd1IoUoO
hNMKszoLcfjsJXJvGOqySBlCI5w1ojJOixfpd4GnjUAzxbLgy0ZAAZJ32SdrK0ifJivMoElN/km2
Jj1IGAJP/K7YV7AJs/P9W3c6marENdqunAkrCH5OphrshasJ9OHDCCSDabyuxk1lMqu30qFrCPNZ
h/PB5RY42VVPAJx4H2fhlksAklQi51wpm0uEqY66QrxLyp4Hq9RGGeFmHTUPh9Qg0nxebQb9T4FE
W7M1U/axkN1AJ27ElCI2E6SIwpvMnOMM3PvTETNTbuzGm24y9QHo/AvxDUzB6hKU7zqtNQMU1MgB
yyRt89M5qUBy2717NjI+iNjSDecFgn/obwdg6RHJHGUXF0NOPgmz0EGqOOEOyPIvpMcK9A/3Ghuu
C6lZ5nVQy7yIJCdStw55T+4sk/YTmJTfVWrYrhx79EPvskNgDmxVyUr1iOEWJABNSXmnJvpbVVbt
6IrL/OZM6YIBPuVsjmg0G+YXdKmtQ6wgy1ezJ84i4k1kZPy0yclh7YYUIGRPvDOynJ1542J+6plG
XpnYqToR3a+w6Dqy9aVxqK/DfIy/j2gPRhKWNyVphY28aJmIBaClag6KGRbgalrV204lZqQJ0Phb
GpSBb7r4E+pexVjPnZD9qsE0f2SfZe4WdU3PGr6DkLlo8U+2I1S0gR55l1wjUtYgreDiraH9yDSo
wzJQLtVV0SsCJet36fnethBssZ9YE5OpypsV7WlLT2IgfYJyqr5+L0SASBGa/wUIc3dO1zCpu8gD
20e0rqbmwk+w3rEJjOWA6VnQNQiv9TnGwu5EEl3NaOgYq3C/hzJ18lVFSI9ZmLmcjZIJOyxnXIlm
2Jw4C6A+y1enxV/OPiGuQPamybJMQMfF+u8D33ZOc/ccPdaYwJa0jm3NM0whSnrKpxHH29ltumki
kLlxxlbhH41DoSqcykyNMgZaETTjLMeS+mootT2UBSyPJyGzFYQ/WCkDfi68Fmca6/UDWS/5RcBh
ARCLvSrKk5c2r3ZYL0+BaS3SS+Rpnwlc4Hs2cPWVh2yZDMAwZbWDcTXTH2ncuQLHZao3zDKj3upu
ZjX5Y+a3TrIByyBRPWBzHhoP4IZV8HzeJ5KN/jH7VkjiigTXYZ5McqM+Q/YI5LCx8/x6D3fe3wng
+GuQttqS8YBypoG9RFgThfxiyd9l12e3yRkCLkce7ZrhNNphNQlnNq/dJKf3iiJcfXsMO3r+HlCM
MBFpTgJyCRYMMO2IPy2KPkCT9cUiUflk5N7KS9XyKf1ggljiRdLT4xJPi2pcsu6hWpBRKayFDiy6
59S9N8jyWvRpl5B1MReMqIX77yAPZ0M/jPWD0faMK2pl7Pxzr+7ZbwUNsqUM4u4mBnhOam995UZT
5bqGT4f5WwhqawiR1b5qUvfhXokjwUDV2sHi4+ZABoKpDg1hsdaY0ciAppogXwW0UQWYD0q8cjtL
/zZHsPYOVMG+34VTnf0PjK5dm1EcSH0R9mfjPts5GendfGtwzr09TEXX8YkUzW5lyTdcgGOoVVjS
3hjaXSoXE8HROAKVOpM+wGwH62hACPZz7p3xI/FJc52uOKuXEtnVQ/UYghvCD8Bx0j9oAqZJzvtD
ba9lAAY/pmv7jP7JPkKLWwR9iYoOqfOmiqnZi0jG1NSnYJstfy7v6BOumh9qHrGHOxPYz6cxVuy4
FYvLvwA0hfBdqYomGchvWnBbswRWBBNjYI+kz/zCE30AQvwIFYc/wPIIiExvwpIEWWbR2fwlG+E4
qBu8wckyp0QfarPyVIMFlHU8tk/PFujXtsZMcjGAxNWICgO2HWvwr+ybiRXc7SwmsKJUhRWAZ5pF
MSBYQEt8afBuw5erjULMW+tpn0+bfau6hLO+82n/G/GDe22q+AuqFXz/xH8oUSHTdf50EbKhivqq
D8lh1TtMdUlY9lgMcKxU0XPG0A8oe6CrpcIFtzlFVK6Tz/g9zvXfQ4URoYhxI3R1yKRwEJJADeSG
rek0IwOeD52OdTFWIaBqqNLgYrZFSS8KiiHqmOMRdW/qQ8S7uXym68h2W1+SVT7Qod/fBcd+baCs
grjJcRFQHDe5qGt8qx/1IOlODScq0H1JC5B7GJmrERF4B9fVrENl59+ILNNjT0xFBmRuvu678lAB
5Mgo5+VkEOsQXHJjEjgA1SIDoNh8TcyfzaDhFen13oF36ig7OLL0cJp39NpjKG783JzxpQKNyVVc
8FHuSOHBxJpbh/RtPSnXVn0Zaro/ZlkBVTHFIu/X4MXI+1/JQnvSIiyz8aWaQp3LwIGwNMg4HwlD
6gg70/+LMm5LV5RLLPh6W19TYNw+HySIROn5XXbvmKyPqugqT/VR/f1lMQnR3iPRUa5Sb69jmbMq
rbnvDKblC9yeAl+dl4lGTIHz8V5dTnZPLwutSewEbel1c4XdAU2iyVOadzu3sWSKdbMiqxJP7HFK
3sFYw1s3dRM3pZQCHCTX1Ti29K8O0WZYwCKvrqEGCp9L2EDnLz2VoVu9sXuycJtmVKB4et/w/ZyB
z6i0g7FT2K94rAXxr8kD3s7Zr8VKrl+dJW5TK3X05qbVLLVlNfiLDdtJ9hELwsoEWxqsqj0KzWpE
/sw1usIN9bkY+/TzUT6G66OHgWfOkiLu1EaT5nhXpbpqv23WAdsCJXa9JtFu7usrtrvfVI4yeVL/
uIyvkSeuMp2nhfbCWN8b6jvYtgnVgXA2f+spQMnkixbbhULQgPXOvEaMf8j/ZyBsPb7xBtcbU0PG
KNIevtxD20k50FisKZ1lhVx0+jPl3PQqIgZgFgH6AgPZEFr5zKLDFPiStVP5qkcLqGU3b5aCWz/K
mjyOiO0y39uMYNONEWW24PDaOfCN21MOJQf3xs1BpuGlJ5z/ulFT0M22r3b6hHq0MmNrFiAk+V6W
ExSPRjb+tbpfXP+ullw43xa14DdLwTMN5wGVS1V9PmS6vISeAytGtWs6fvvPf1YyD/j9EpgenJJB
QG4kj0ltmg3VIYXpcjzOIhdXHZhqIx9XXsc6axc0gtzor20FQRpr8Zw60ac8y+VW1Zvm4d1RNA2w
ZWuNJVclGpmBow+qcQpRFeUosikFT05shPpYeR0aQjiyWHrcSptUKbPLZ0hrLQTY+Jeyv5ggjlH7
YGSyeaya+IZFBFEAy77PiOkWJw5Iqto4DpJBJtljMbVbPeYeqB9sI5LpXJKtFKtjjRmyBhUrLATl
X6KJ+tbq7AqNLryWFg9Yw8IaXyzi/XGVK2ah3pQWloUaa3GlpxaZH1gwXwZtJ7N1etG0YORPJkPJ
ajOcngDGN73SoypSEnLaggfYRnxLWkAqAbaZ6zhtk8dZ9ivkmLZJpZ3EnD8NqjFQHImEyYqT4oXs
pSTju3gZH2xnjEoKLy+MNT0nwOktq5j5Frnbqi6dfySozP8nhVoIlX8OgETdhSkw8sBlbHxHXq4K
MiadBp6GzXTUNndzIyqRaCLGmsNhKp2v9Z/XIKhb/U8+nX4Z4rOVAmstw1+PorOLxQSTvryVTcUu
/BcLzG4b+uhCFgzJYrXJ7PI5VT66i1ZBjO7Kp5nmjswiUN8GGbf+j2OF2PFbDcAZ8OTqPN4SXuAo
O4r+fg/H5+sd+kMbWPz4CvP0rAhIsfuoIne4xy0cH6Hat9nF96XwJ651mrl7oMHKI2d+bDaQVHQG
LIAhixu1rsNp0pcO4hVrBoe3+Oqwpgq8IgJ4ysXgmMkUR++AVPqXNa+RitikSMFqeSe/A4oSRJwY
AlnUDbI4USDqnryn8Q8xDsAGPmd6boJUekddlYP0zMhRjv58kasbSXTf3oLVZN03tmhdWPn7uPvt
bniupz/4Spu3mgOU8ahAR1+A5wzbTCqrgP8lzS/I3QHjgmqWCeIx3DP/VeGTf+f5OUe6rdewQCQl
7HwoftprOSANv5m3hZAOE5o3sFO7q/6LfpdURUh/tFgdGJbgdwMYsfjcCvPoTtjiXmhjzxt6htRu
gpmw42qE9eXfN6CX4qOyiCZ6y4ZUp3HfhY2diSjogLJfym2/bQgPrfKTAXJB3pnt3XNJd2aet7P8
XnBNvKNszAUhWQA+XxGtOF/OiRNB/KbFZiMzIXw2vKhfPqxE8UowxYRHwQpeIJDcnnzgwxElziC/
6ORMbTJpk2fifIduHO21020XatX1ZsFp4RCfxoDzWw0aJZLsU/ueqBNiAU/bAufMFyb6TIZOnkip
nCHBJY5/zx/7gxvgiBWRlWj1jn3Bg3tRcVMUFd3UgfeJm3F4Nt4ViS7E9zNga4HwZOlGW72+xM9r
Ewfq5qAsDI+97M6Vb6rPMBrjRLzu93NDxZU5Y7Uk3tNeoWWgd3pvpKw4rDEVqQZAy5H2fjalzbn4
Mx0U4/P3/rPgpTVlq68aPgg3og5yPZqRWRu6H5GRiP1OL16l4m/obAJnfwC8CCIvFQJVyUDC/8Dl
khRy6ZrabMRBMsLvcvT5mn3Pj6zokdUcpMfI5Lc8/6W6OI8Ar2xa2HzVCrSzYNXxKADsbumbkFyh
372XzSsiHbSGcUsatPoUp5uMIQIB34ULuqYjSn1tJqMFq26QCHq08WX5plRjeyLqBNxEw6hG8mwp
dvezBlf8SL8hTdnzRNcubLol0IPA1JWaSVriqChVlxLPr2JrLttI22cXrbt82wIhdLLqScce2R+/
msSH0SzAu0OX98AdAo8D/T4RG1cVUxtBKXwW557gTG/5yrKSNM/YigqEHBcuZhalL5rj4EUlB1ey
Q2qcZ0oPge+rsxZjtd0V77lEN5LPuJGtSSd3UvigwQmMH702RUjyTIt5jmGVU2mVFx7GJCQApXvL
XJxAI2PW5yNl2aPkTbFZjoRJl4HUiJ+uFAg8DMbrH61l2TPC2XW7FdH6u5k3Dh2XV+wpaQX1/qdh
VLWiHMvPJGErOzK0eBozUduY2c367UtnW1LsOvASKK3ifQGW/dyC56sU/5olCkMzjIZckWfQRW/A
SG/onOf24b7WmpTNP213bH6Vs0T9zSw5GfJzVQHTGq4X/ctYdW257nF+Db5NhbA6nM89F2yLn7iY
jTwJep5MCoH5d6qIMlUo/bU3qhyONB1r9BesRKolBjTLdqQ3vNnGPePd11mp9jsoaqVhrJYYrwJK
nGdgfh+4mwqMr4iXGr0A/F8puqbrpDBwNAyvh9yN3ZltuMFuVKdHvki7u9aOZYD6BVyR9iwSM6ev
1twaRKUnrrCdyks9n7foUuh9SS/RPWwInqQoqsrCjmXtn5CXEpiUP5vjzG5S9EaLergDo0JY5Hy+
NkYGFK3XuOOjjc5ID6H1dnKdyfO/THcdXMg4wjfgnKxwIFGj12gZ65IvtpgsGFLoyD5YTKpQUllU
JiFhILfvcNq4z5TzXyg+rC/z6YOck8lhsY4tIx8rZMJs9lbcXTn929eRMjJv+UhJ5e9WD45GBTzJ
kbKt5aHoAdEfsPunjfwYYb8246x6++JojkijugyfvI/Bdvd4g9eKr3mekQnXejzRAQ73bsweDQBP
qN1XunZdYF4gHTpMQ8ZhXSjdvLcp36bVUPIh2ml3eZBPWkDE7BbYn6+trApwaCUJi6g3e659mtCa
MQmR22OTLV2VotntYtFQS+M0HG0SnhocCVpd0aPwnLHjfWUsFCCCNy7dASewXPyZFEoKZ27OdBDB
0U4NPv+tyOUIV7pOZUz0BL+VbyVEnqHJ66V1Qu8nSTRmt9CuaCy286vvffwHPuJdovqOxTcfEv3P
NrYWOaWgSWBIyxrHBWEO77Yj9HKcjHTZ2SJoRLz1ZSs1RbwPLlaKONpxTFd3odei5tOo9/+bAZf9
VKSLJotX30uaZJDIpcXB2GfhhD3I8p3wUJAOvX2y+UEDc7aR2sUtZIIcZn/AN9k7wQmydWEHz2WJ
7tmaV1YMPmBrzcryabjBi+Roa/hwc/bkLR/tuE3AvSkk3KxQxTUc15o1fEvsykbivf+DjhY4bNtF
xWX6TwdKWKUPzfR1yn9iACEp889DlVQAKjvZlwimBTwitKzTUo4RBx4taIbP5LmyMgSuhtWHAFBq
bAsuyoSr/urK+VkaleZoO2LrWp7J4DohYOFKx7LcQfXquwvIAWeMhEh43eU8LriAaGj6Z2oIbgGc
D974iCZN9DG5Lmw+5l82rICCMPt4rhx5I+IYJWD+aHUIBvH8e9aiXsLgSp9adJWigwNDfSUPc949
HRdSuU0b/DFbF8hIqMMuvXTO+n+qhGZdNjDKNIj2ojVtKAKl25wziGwyyjSD3mE+KeW6MAW2Pgpg
pXMnLOt8IrOn7B57qQ84UoSi2VlkzvxwP2g4WjCayl5DALRdPBdh9ku/BHdDFj9E4CuKhWbdRa8i
93wfTyIWSZ2H37P5DTWHuYdLquURseV62SZg/lI7T6YXxHQ7Anv3OiPGQ2fBe7elUr93ZUpkZ7mz
DLURyFdYcV+q7loraJS5SAObweS1R+ALgJ6LRgsIFEEmSbYE2vJmoDhLT1ZJTxi221MsEXbA/llI
J3LJOIW+pQBN8/AnOI+EYeiC24jZfVb5vzdIOkaz7IZA9L4UlqIUy2TUYxE04bMlvlXU0+wfwWw+
NvGYZ37Rqj6l+HA+dFL0qmzYchlCICeP7NRmfB9iFgA0Kt4t+2IRUWPDBBgSN1d3VW98NhjjALhc
FhkBNQwJ73rDi4VBHTU0yROXCnjOB6e9obEvBSXR1yGB5stlG8Ln9wkI51AGiXIi5/wx00Y95HSi
ES4H1evnm6nHW80orr4FjAPFTBV8SbQrMucsSx0EfFkhcXBHKHS4f9q52vEIT9sF1pUAJ9sxj1h8
+bHkagl5iaed6776D+u8qn15w9EmK5fIERpxZnxR8dZ4mCQxfW2fLNuvgFkJDJdhaRCeWjEkNPZR
avfXDwvMCkSgC9JfqtzkPtuKRCAyDWTxnQ1ag5mR+VKyCiT8b7ghE209U+OTRINvYiFlKfKpGVg2
URfBbZgXNNFYiJr2rIhUmC34emT8RaLRDOFyd90y3vf7hzlJ/Ll/XznGHMoBvrQF6eceYz99F2Oy
hi0nrxuXXONZT05lAkhvFul4Un+PA+i6AGsSaNjcPpbQuFeGoEmo12FLEiISFZMc5eNzuGPDqLik
bv1AzgPckTweoJ0skGJ8wG7J0kWKzoPc4Ak461xXssWYEr+Tcm4CB3Sp0hD/WWcW2mF6gkvbXy1J
RBzoEmOUPl3tBd16WuXMNLA4zhqmh5GLpOovmJ1ZT8OQcBjKRDD6QiAPrqiPhbEpcDTcoCdGMlWN
Qrdp65t2oQrIm/nZwjnVnqV05+DnE62QS7uBDFizMC09teGPaG02Bt8F6zVNAn3908UC+3reOiRV
yVePCQNbLJI7GbHNs4iIExXyq4qlVWd5hrIVTLOdOPsWKb5xr8BwJeNvUns2qQy0+JtujwPqkYOi
4rzs0eGWFvk9KWnTk6AKhfu6OEPdOcdhhffi6eOfiK4/eLfj73t089rtjgT2XpKg/rtAKLyCX4V8
oxM/RG9lMH5fUCn8ah+IrB8Df3drv7r3ng4ZtrZslVM0e4aTYLt0IjtwTLbBbRZC3owS7KTL5w8H
WYraQ2G15DcfQ3JnmDD3s+n3zisijgMWc3qssMFL5hm/fhEFgxFyqmf1no34uRxDSncm3SOkvrOX
GG7F5Px23qA10cK89z/gb4mZYC4KQPVRUI7m0Se+L8H8fa2+MBlaBsRWy9AJWsvvOp4lTEYbPBCM
dDkNWqTGxkLVfTpAqn5IOK2nLGWcGpazbAyo/m3BHUgcnipnpqtnId/09USMtHyGtuLVhLUnGgMI
/tvXcVZhBNmF/KG85gs2CfAgtH2+APhu9it2boKIuVyOpPuJ/DFvQ6fxZo/GgIcTVLpbXT+wdxfZ
K8Ij/u69qiBGDXC2R8ls2OENOt8ex3cB2viF/sy7bJWaa7z/QsMVrw5qQ5LLkvdzyn9iGihcAYpK
HM49WMmqlnMoQAyHMmhtsCANZSqHeV4R/krIslXnU+6dMYsDRRpaoDIineATCKZrO9iwzdSJsr5H
Pvg++7gDWbP2mSZmkBf5UZHEI2qSPSz8jLuZ8AD4BxiDzysHnxIpaShUeOqWq6VgiCJWJXeEjNYY
it76wjNpuuSHcyzxCu5oTOFmk5aRFkmzfkN8r6cA081H8KTRXBKcr9xdfeu74l+yDEO7+pYs2wrI
cBW7sk8MVlkqzj5b4EtwVNz7TEarXMYma1Ba1yRKgM++dsoUMRlBMWk18dJkpoPB5oNkKqecqk24
IrAt3ffQTiz7vaIpoJhlEnHqQ/cDEuocRn/6IaQk9gZ+HCmtTHuXKsFrpeH31nwFBOcYQnF8efJp
onVIkQJV2LR+RWehdT9Vuga1n+TuW3nsZjyHwekRERXFSIeWruKqphLX39qzEt6q2XICWKZi18Qh
1fLj+jhp3oXJR8sSva706NYfJpxvRv+/jHTZabZRZf8yqxhr//zT9nBkYRBTBsEr47kZDFip2HHK
YXz4UIOsOODUokoNv3Tfhl3OOVfIkKMCtQUTAyhUp6M8j6N5l4N2HPyZhS8ACuVhBc0wJv1piCUQ
TJkHvNM/kiR9QlixtG5LOyuMeysUtIpE9+pdBzAAh3YYWmG/1yLOXJA1Zy+5nJD2iJpfpntYH0gS
+dtKDU4zeN8CgIyJfFUdbanc6gSmByw2mEFqWk4w9btoO4+9xTrM5Yw5z7MZSegmFoVKXL9g3VD4
uc1lFzaUj8d5ZgRe715pm50oN1fsRdFQzzYv/cUPBWqeQbWN6Pynxacw/ytj6U3xV2vYcSw/A39p
bsWJE+iUqY7u8cIxWU39P2ZhbRwiVIMtDmt4TeZShOEs8PYJpt1Ra3/3s0dWgdbhWKj/UiC8nwzE
RjymsYcnOb9OZrde9BwSVSmXzGUe/N+2OgbMhOaTWiTnkXrzdP6M7iUlAgJ3niJC3TJJqKVOxfRc
piQEC2N6Vbk3nQI/I92MQQouDuMnMP0grAxZh/Cu/pgxIqntM3clxCn/ZsmpRfRzfiVqaOaz0+ho
BMAM9h7l5X68OZoHdGwL4PkniUUmHC4zQRb9Wi/aK54AShuhQwM4qFP3JIzYth8z4ytP6Q+LSoKf
YD3gmQy6HQGIYzj4PJkzB217BBpQsrGy83uqOIMsxOfgQix1XCYxsV7RjtEPU9/dHHGxfrYVciHM
yzyiHZAS5Ubgnjjh4K6l6gQqKmVRu28AkSRETIyVYZL2XJqz1EVjU5HdtTIaNu1marfbITY2fH+3
J5Q20yD49DxueXC0mXyoqlCQpanEOCKn8rO/JTjaA2wHJk/s72vhmrwgTI8o6XXZHNb3bUs1QdRu
sLa7gKR8nNUixUINaLfnFRZNCQMzeEEnRZU6VgJtHwASCTtQRPjx9DagaKfRyZF0RzXEm2Q7RgIX
v5/VDeBKG5XiaVhb0++qPkyDqvrqP8o5gVTvv8KVAobpE3CiSwRAqws5aLtlIFQtlPuuO4eKyDf3
3Ib+dNbBdxFyZHztFBhBuFtJ/4yI+na0DTL4VQizpUVi8iq0m/Bj7g/RrizKV+nmbw4wipU1HaSK
ZcPy+zvHxVq2UpzIzSTVtpYSSNSrC2iDrBBbAa92GqOxc+GimmvLkPAm1xYsAhK14w328yrAJs+C
Pq34j8d2qVxgEWRmsWLDW5jj4PNB9yurpoj8SGwcGpCB+JpJiNaqjOrwO56p43l9+qOoIrPWZdmL
n5WYvDp57HGk0KTFINZZsB2uTNHmAugsnNosm5PEjAXJPZ3XYkAejOOQcCv++U+BMqv3zEtde3wL
1kPm08+tSkdtkFOPIbOOBdZMhuBZle01PZM6jwF2kZiePd99gxK7TkhcXNAzZrTwIpvlGc/rBLIY
P6DOWZyNq3qmDViSvK5DVaKAgJw07OkKy7FRjkPTsCjL11ZJqEWwSYJabhtluHbvFivcsfxhY/tB
Ob7gN0red8fGlUaabgJpdqTGL3j78On9LEYmQs9X7gBAfEk1m6wTilEm7m4x4dnwNYZj5c/CvdYw
4q2pdqNFHeIe+krWLABfh6q/ujCq0GYsDkpKl4kK2IbFeqNCXgnOiI0NYL3D0Cmq/NHwirkQJr23
1Vpe+xDDTvP/DFbTi9GoWErXjWmTyX9vmScREuCxv3AUluEU01sa0964SPrnKR6cvKZDWdaolUHF
zvKY/Lu9eNda6GjYHmoo71HBNoQyiQMedZ/fR3TiacqmOnFCHeiFWEkWMMgQVvC1CMyozCXePC3g
hESHC8ILnY2pou7hVQ3Q3QpOBBYx/ov+1M0JP5zRzoeYcZlAmfn4c3wcao4rARCKqzrAtAgEw+vJ
FcgZoiE4U7lVB25taLOVWiEMUemP9WTVx4/80EtShD8MT31dN2BFSdi9JGgZZWB3EU9Gy4ErMasG
7nwEEG13daDZ0qvJpbQmglHc3Tc15SJTD+/yf0ZbqqTqhOUK+9TeEC3MRX5fujCFjn1yGfhybMY3
3mBg0Q+2bvewxa0R5PiqqZq95rcVv1wwcSoUPaebV6yxSwUvoy6GxzxalD3K/p038SkOacPEDCjk
Dpj5Uya5HmoTgLuI/UgtsdzKoOhAVYQRsGMlEduhZ5LdV7H0tcsFaHT5CkLehsQ1r41w+S+84r6Y
fmDOclAbkJPou3ubUyMkJ+Lz6utIekXdYCInK0d+fO3Wz6xyeonw6ZFDpyAHn9Yn2fPMIsMvpbqX
zY+Iry6Fcjd5Yu7cKfb1GIGBmFNUUGZgqT/ekf/dzrkvJ3dmwCuHO+zNZLd3it+PBRSGPrQG1PM4
pCuSL5oibf5wTEDbDXj2BkDMBC1pfkul28WIYcgxD8njrWPMiaoH0u+JrpXKpUU9yXhUuKh+aZO4
A1re1h2n0rXhIzkJczwaPKfzlXj8cwWrD8T18uOfKHzAPBgIDwpW3HFhKnH6IloTsLYkGBFar33C
BVBsf+TBy94IO1ZnYBhvwvdlGrc26EmqRIUzPihYdHrvdQ0sx104YRfnlhjr24S2Zb/dXumiWQrx
yVn5Or5SELBYTxZpHowVDmFtjkAqOfLYDvVxaFSWSoRRUaV2SjukQ+uLGcsEA8CkOyR/k06gJjfA
8vm0x6qVyq7zmFUOyo7cG/8PuPnzsCELZ9TV+vJhgmikvz1A7vHaM2KH/645vcdfZ64TOZfSTk1K
XhwPWLCCKxlqpyubc37j8lnopANxo9Xc0xsj00h3KUuU9ItPKR56+S9ZOVk5Wx2HKmMHq8NvTg33
Lk5EtrGIdSDYPNEO5Asrg7nMnKww1t6l6r0aJQ1qsfYX2HrhqE1whJZwm9DMBWg+QqSGNINQOpPr
Pj5asOzBzQpXSSTt0CB4UwpxAclDmsy2BPRbzsMp8a2G2mqxtdlcR2MJQ7WMbVteWXLHQ+ALG6xa
WelMyOw99iwhXQBP5g7C+YTwAJ0A1VM3upCIOBGsr3QeKs1HpJibdMXN5cDuupO6Vu5YT+uYwfdS
mnUHR+j3xkQGK1W9SfHsA8U6PaLMCzVyJxOJjvPP9n03rVfI0R2lAT6YbIWWu1X70okAbGMQaWt+
qcaqWnViFU1nxr+lx1kZ85Ij6H5W+edXtxOEsJkuGjuKy6MpQ5fFgzjXbnKdoUbEi6pCDPcfZJXR
I6ZhKfOKSQrB9PkoZIZCiEIksXXknKLV/UlHZxxQasqDPitPhXK4lV10I6IVoXfCFg1Xa2ZWTHhF
svC1/DF9RRLzTBfsTQi4hE7XEygSH/sOks9NrJhGxHHQrP/WBpRX3QlaXk//WfPTFTNxf+qet9no
JJkyGk2g4R3KiP2oX0w48Qms+o3WNWsk4+g/6bnCWGIHyNm2rs8W2/9dI0Tsya7hQ0kZCYpR5gbh
evMiA6JyPOW5qDOs7ectyKMaY04yw/NPMOWVJSreUPfsfkKGZwVr66fIV5XzeXQ6e1JXf7kDL9xY
iZMDiW9pmtF5CENm7LC8mcEGoZCqtn0EwXpIczf15AAfG8ZOf2h5JTzfmkx/SeK9iNHL395FMCdV
ehwv1PQqTCbaWU02C1TAvtBeCRN0lLSamuQIskyt4tvwT/AsA9t7yoNyHhonnDxbnhUsDgrYoler
b7LL3K6uE2uM9Bo3avlOI5CdpBK8gP38w86UQ82ZS6SgRv6vLYxxbxZh6sG9JmH2So9/hBEhZ3C4
5qMNyCchKI5tEo1NnWNx/+VPL44EEBy4WzdZzU/FodKAlW9lTRJmQO0zSMIoVNDC0E6GCZQjL54B
JQPuw2sBDBGk5mP1tMc48UMFQSN43/wdTVj/FVrq/Y9WlgBuavJsKJQaUcCEKOGhJveFNuXbHHFh
gUuOchYn+EZKHzS+7OMC1DOjiWvpfR6MvsHZqQ4Rk+kptoU2gdqGSfrnL5cYE4ciRBGUZh8Qzchw
GSoqpAH5jNx0Go5ErXfB4bP354vfodxgEWB6GqreVVQL0JOJJhWUvCQ1DzTBmTon96HdHApbLJm7
Bs0ABh38KEIIO3/uB0b86h67I9pEGCp2HLKcdO0SikXDwMSz7cDmft/NJq4jaJjnuHwyeHvQt4cP
ayjRyB1SeC+QW3tbC9AD0BOZEjd3ZoJpa4LBMrHtypoG+NLssNNiHSl18BUhrGPiPZp+bXl4qdkG
YvlAeaT8ix+lxBwygVT9QHrJaRZWKMsQpQRn3h9YIw+htk5MdGjgH0XS+HKqaVKL5bnSZhML6KY+
zhGdcQq7o2IeM6o35sJDsd8XefAv3lJzQze9PCTYXyhUCLk8bC+V1k57m6DFV560X2RBVBlWxyHp
ZweXH1tpnfwdPvh+UViItR58axIwSF+aGz3ZcmdF3ACpsUtl6c4iob3Km7gKq6/btwr17+qWI2vF
FzyZJUVgtp8WMzaw8plBp7asvjmnVsmTHDFZa3gZsDb420R15S1+YWUJvU9AU8Md1WRmm1uX9/F3
uRSWidbLULpRWSp8m1kfFuJSt+LT8kqZ61FM1o9pejaCehq5V0KMTGPl0mNj3lnqHBEMSIcr6nBw
Bz3d47ymTof90hKOb/Vq3l/bO1p1Tf1a7wPjoy6YQCJaZmilYa1kFMzAM+SB03DVzv4X+B9ZPHk2
KAT/FDVG5zk+k8GqvMSqugFjMaMovznXfskdG3lz6vUS2VC4TIlHc6udlvUrLAHWXlii0XcloZFO
ircZ4FfhgqfN82q8R83XWXjiOgtraiQF8Z5vGaNTsNXMb+FBgho8jRfnqSBZq6o5L6BqEnogoIVn
1hSTxpqM02d/2ql/+PbSl+hEfgThMnOHVrmNMrknDRiHnY0+cr/6NAvOZA9AnVw2wAks6ITVG3YV
CGYYVYUQSeXT1WOfCCDyV5rEw0B2W7CmkBbIboMaI7LKZ9b1RRf2dxyJqYfibzWj3d1gKuN1cZ2D
pkj3s8JzDC1H5AIUWImjq82jU3O487A7ir1rl7WlsIn/ylNZPAy5OX3SttJUWWSizZ6br0uMKP44
g4e//96GzTOo+6bZqsiDxmkjR2a/vggfUUlqTLi/dtrbkBTknDwjXjNpnR2Yq/EUux4phFBG6stH
Wr75768TH3fY9K5XPLem98mS81xWv3XuYoq45HRHilwFthSmdyV2B1bt/AOeS4HAAMcykQhQ9kXI
uogL8esoH1pW3bf/p4YauQzDReY3+BKA6yqQY9zCA/MelbNa0zQxvXLIU2a+1xAbz5fO58AEbMpb
D7jnbDU9uMCClK3RPYUpOojfLP3H45EzB1C3OCFWq4TrV9ZrSZsCgvpt3pWckWulv5Y/aude9uYa
40Ry6FpDSg9hPv0HjVojSm77d5dyPoy3xlxCv34HY2ILv8DzZF2Jhd1NTQ1DS2wkcCbBAzuU7Kdm
a6WNQ05fOSyL5Mv3qwj5oSGQeZ7aU5kP1974vxQh152d9xp4qqFGfPdfDQx0LoO3SpGz6NkMh8a0
jYAt97le9wmmJnI6+iTBpzdyTwd+hkKPXpXdZR6O621f6+9fG9xjywHygMbM9UEZtK5CFpSA0Zxo
/xo6KkchRnwBdiXWN9QHCxNPSy876zhlOJwcqNyhC/yQByF4Mqw2VFdyOOtfEsYOp2MIEts1nmI1
Jgf5NFutmpWH6VsY+W+12AGUrBwipcitmYn3ESk9lpBxbcn6+hUhziIaG3q+HE3JoMSnGQOG3mH+
p7fgNLpMMG/Rrcwxmui7rzFTZz9r48s1bXLuanfWfcRERu82M1GksKZWcvzGsr7yN5CkPT5jVTzD
gUCaAKbqoj7Lk1gAFDUsA8PLw6lxiBpPZiaUsz+7k4JLniLaxyqZOvmWDkWnLxxhIzcDQjf4bF9f
UyMdeSQvkU0rJfPt3VaiTdXxgWvBs2SZjkQL80c0NteaFblEiPS2MwoXbMqkxGgj9i858+qboaeQ
H4/8340H0EwRDMiryzuOAZp2B52HFZgNXns9GdLPyCXmGX04ObdrPp7tJtMk+JRSINF0uq5mzTN4
4wOuF5TPzgUKUjWHYFttyq10M3PQ/siLWcz7X5O/mpZ6nR8UjGiTREToNvCRB3JRGX8dgSj8S5yP
S+nCsgyIxKdgihzxJk8cHjMOGpbpY2Ha5l1+cvoWclH1T90DZ/+fJMkvaddxeNe6TwnLXT93knHj
bt6ueHUCTSApfXs0thYjTYBtubiHzSVYh0FdN+unRA4hHutcqiz7q0ux0hp8vFApqFgfQe+BJ3ax
8aDOyRUgLNekULnmegJR4IO1hSyylvbboVI7ZOzwKIPJug215CNyZmbxfIu+S/CJB5iiEF9m/zMF
HFemi2XL8Mbg7wPcp4K3kCEUgw821XeEgqcGio7oAUl+orDYugen3QsZXDVRfFP/ViKGRntmQE9o
qlMv3EQ2l5CrQPQhbDg7AVixQLOnkuZEiH/VzsbnyX8TGjbHfUK7nK+uEfyLrbRjnsTMrroDsMsl
4PC0gAnwuyBX0eBq+vVwds9ta8VRDIYIGawWd+yL97oeMC/GOCvGmRYFwg4y/iSmBzAXtSiLn8hX
OttJJ7MyzJaRN+aG0p/xhfHmewv53caHin+/UZaiGgv/ZiYfGvXkxZp8qgolK6Qkn2Wzo0l6RiH4
NeT7VwvHqc9rCeBt0uFoZXSqZM1ShTnLlbmt/5FdC76POd5CnMzW0LljMDU1GNwgw4efkLzawcIs
dQV9M5L5MBRuQFMN5DwAVa94WbnUdVesvY2TNNQUzZZ93vUoXHb/GTfrhp3TxYYgFvqn+S4loZIu
frzJDWlq3dDcjO5l4/V2+tP1XJdi4ghUsn8gOP88bKW+bn+C3VtsV04KYBgCooGLxLUKUnwigILS
l4Ix8/PIEqbbdIJUSjTiew5rcPd3X2xMlxOxaRC5VsZxgzUbCc/0ocUxNRKzWGQLPPd58eU5UHMt
V1csEj+AE0uoUTX1ZzsJkrtyHSfzodWygpdO5Nb+DGhAwlON16xJzavMR1/6MXdGisy+13AQElpH
LNxGv4KDda9FCiHWcRtNIM7+3Q7Aj9FgFHgSkZLjXEmnS5f3WDLXjT+CvWry2/IBS1YriCdNnCKo
EruBI0smxQ5eqSTdDRChIrUqZG8JjOoQrPyR1Qh8GsVgienXulooENEuA8LzHLj+Vrc3m34mhTaj
JA83yqe4NJFiw9Bx0bxNgjoT+o9vkEORpbhxB3+qpT3zzu1TXJmGV63lHSzfwfwQ+ZkoYmnqgglo
nLxgq8mKP39NtO1xm5M0jcFec9aac3ced2vSlH99ohjmtB8EBjrRPMuAu515jMOKUTTjprJXl/ky
BYVG08rnwl3RIkR3JjZE16GNY7rdsnXT9OipLdrLKHVgsMkRgw+CyBqipGe5jEVkiwgupNMGjG/8
pXZ2ExqLMORnHSS6sEF7A8as3VHoILm6VFB55Oxjrwi8Sgz7vT1wojYiSslB6C6qXiY+SdruCS5C
hQxBrZJDwrvw3jWp3Yk0CKt3kZFhJKb6jCArH+vshNEA9uo0haiRVFGW10o1Pq8wnZogttqq1w3/
B9cRa2ZvHs5d2v1oWdWWmRgvl5N24doRlu5fOL3/3ytNraGppHqlOdqgwhFheXQV0uFVH6U6biPC
FEkLT58Yva5SdDWsBZ4Be/PqmF9Aw7GArd91uR3hTMLVcm441Mux1Nwg/aln/iHZEe+m+MvoUCqJ
3uhDei5xtDbJvLUVEUZp1HzwydZfQ8E06FZyjiMqYSP1e0wr4fn+uj/evLZ6FsCNFpgSh/0LrwEK
y57KWX4cSTPfQ/yiX61qfa9+u87woVHBqtbc8lwjWyFH3wnv/cYszg8ej9UY6WUtP1RTD14EnLgN
InW0u40FdWP2rA5X8/AXwuwAfnZHqYMtOIhbYUZdOwaxGterzbId/PTSDHtBG4ug9kd3lT8FbtOQ
yx1/iO05iVV2chsbNlA7QisMsnGuVHi1J65mvdQEzJr0VUqQeK3L6esLvJqbOXCkAdYvnVLrlT1o
UHPHXrQ94hQs6MYall6v4+o6Q7MOdD1IeIhlPNd+3oZx7L6g11NzjefEG3g2qtWEWLwf4xyNvubv
AxTl7XAK4UuMqsmQ4WIfIW30bx6o3tALbpo87oNSaPaZR+0cKZpXsgyrN8Dyz8eL8iV/hM7MwCFH
RHHqpNMrj/Jijj3HMcNgNBN9Y96Rs2PKoaD+2IX3Jz7/elzQVvlUsRU3eDDVS/Pxq8RZ8G8Q4ONo
iqcywJJOZcG4OUs0seZ0lo+J/9O9Q2/uW0r9Jogez1ZmXZ2HkSUaqAw9vucl8clm86xSapQyrG+O
EvvvlpWtV0OZKRuDiz77zOtldBIdvjG7bKVkFaRKZgCKAI9A8kh3eM0vu2psyIJ6Ef3YCNaOqAwy
hl03umuRmys8CWqV6ExUw/3lvjIjXhMTjT8ZlvtvKjnhbUzDwDHO1BhBBku2D3UWU7vRxZXSQwdS
Z6foewgtLCzq9pV4hg826xAeYENqIvEBtk3PMlpRB9lWQbQqcU3oemGNQtlnXGZxNNbWmHEbcaVz
+Tk2n4MpAYnATpmOUpivTDxAsfEpxoU7SWPpTKecJhz9iN/kCYB+HJklEVleGjQlo+h3GNkHrWgn
n99H7821KtzazCg5yjxXo+72QaxeJLSVnEf1RWnM8yJWHWUPMIXa6Iv/QjTVgnXX+8XMX3g59Vkr
C0QzeQWUQ1AFANUAHvybjISDChs8e/LnTzHuC5hA+RmNRpbwyBAElLVs55T24Ax6i74JmeinY8cO
55Nl/y3mZX34o028t0IrOhfJmOidxv29XVCf9nc3Pz5g+ysmpRT2NBuW/OjAlQHe9WjRm9XMO6cI
kde7Ei9kM0kW3zZgAJnrvRJR9kg99hObr1YDA2K7Fnkwp9/8pM7CZUxx0lgaJ5Lxwm02/n15reY7
zjL+A4ZpKS2+G6CGa/+PSpz86UsWXhdWEz7uTlLdwMEc1d4Yp3hGgJrfga3YgZPHrByEz9Jr9dEe
3IxP7PNVi8Yn5NjvsHk5eB0T5Do/V6pwVTG93R9TlnocclXHri4aVk2QXd1x5laKODlWexPEN67E
wUyf+rlTZXn3PQTIEN4p8IKVIMeKxxQSl7Bi/xJEPPgagdp/fvGOg1eMvR5WmiENIVsmqDTGp/XO
x73t7lHIbPTuVPAGpZyu+M0Z5XHq9dNDv2KEou1bKKDmOVU3zF+TiP+uIR/34rSZtiaht2KRCr8E
Np6yYglUD8lVzSlLKTWe04ANuiPo+JfplNsdE65aQSPXd6gx8dFBh6J0uXqPuvvO9/o3gxQS6YOq
GExa50RkrrzeEqVbyEBkV/AbVmJSLcQY9DgmuAqtj0FBJ2p7VVaKAqAwI5Y6ak1hI1aTLvxqiaND
ApK4hNSQAjr4GoOnqGM3kszZVc4cM1+JoecZ/DYaXQ10EFiaAhSHcB2QM2FztVDYHcBJ5nxEw8a9
MFdCdq1sQKjCtJL3TsAYo6FC2o3ZmGmMO1ML57K9px1jFQmpzfomQBAFvSCtnFjIMHdYABvoAsdq
9VdbA3Rwg/iJrg0JkGLfOmzWnn3/FC1kxl0HmSgZ4HYSjrGoGYkBryRUn243KN2t7VsiJTxVcnic
EPBZ2wnMjLUrb/V6TapuC8TfMiEcAgA5n2mqdL3Xl3AnuKjunbc+esifegVOBB+KeX0VCsU3Q9FQ
Br0Kbs8LQo1AZitqwV3G6tst43qLuFOZd6mmqoiWQNbX0qKvpLe1nssezy7+rI5k2KsL4AwLm+li
MYH2kTl8nZDAC8axirx1Vygt79OOum2nkdhvZnauGcaQXixPiH8gF0o8Yf+gjDSEdL3EIFyGUTwD
vTYu1qFOzEzSdW8vbyGt8P1+Dfd4x6VGDbxc4aQ+peGPQGuUxz0eNXKJrG4Go3sLvsXerNjJeg71
OMZBxP6CAwWDtsqwM8rS/RRPeXRM1CwVr7OeoeUp8toZicpJCbw+dwy+PnCyMKfLea9YiY0XJi6h
B9Vv1WPfKvk1NNCDj8V5gE9vmzgcQSO5hRDQi41LbP6S3os713AEAdmD4tqlxgcL62uB+6r0PKPS
hLk+b+RCOar3nUt8yfpFwpFoDVmu7XTl3RDF/9zsKQHJ0RfDELxnITT+fJLMI+H6jhPobBhIUV7l
TJ7r5xjmYwA4jXbdTH51kU4G38Ztq8Z16XpHuu5FrtPqX2mFMYrtc4B1rRXo0t7QtJJ8Kdgo/i0Q
Vl0k3v6j9Bz8ormYwxX8eZHuwVWUGBvMFWycT6q49f3cuXELkAgTo883WwEDdB0mnoYYDagxif1m
P1eW6eszokueoSzJ3WXL6Aq2OeVbSw+NwpSseXDh4W00UEAqgbUgHn+iVx59+jI+W61Ow6ACoRQz
hl3qbdMCHxmvut7xqnG19miKHEuZNYH1nHUWoNruYDSlFexT9EXaGpZ2WMlbrT8V/ppd6TdSyHuL
NBp53phCiC0ToNDFZ58XbkDiUVXUA4sVw15AgtEsvgnZy78p20t4GzFirHj8HvBbc3Zio6lCSsED
Hjl5qFL82AD/EYmGWrbKJtfZ2+hMaNPUQ2LW4Pz+GL6RXFv7g/yAv5aWaEj9FqaoYp75YyZT7cat
SGWVNy4niDJ3OTMIpoGVEGBFJRA3g+jpoIANDGUftilg5KELdDoEtXUkyO4FM8OBeR/Zygf2UnFZ
tmN2ni71+YqEa9OOclVCEEei6wIwbSaQvs2/SMmu7vUryr4CZhCQHVuR3Qd4UhEaTQTFjeP/f6Oa
kTDDhzchRC8+U+S9JeYyQvMTql42Y8bbuR3izWvAiF6LuNOOvXJ9B+bt7sLV5XYOAtW+9G3dNicX
vU/PzaTQp4Hx3pcbIzD/B+9294s+3UlaP2UQg7AEMnhiPkHdgLh7betDza6gm1ostsNNkRJVXCg0
C8upZwoW3NbevRRPDa0hj6v+FTMRWeHf4Tp7eXsY23ItdUh32Ylv4n2smvbn5BuiV64IGXPAj7kB
dBP3WXhV0Ht7qWyEhUWh2GCdMScnpiGd0ZKs+bJznYlIo0WsXTIKyc93XsL85U7NDHvZpCnWZuZm
G9/0DV4RZj/lyEuApU1EtqvemhL82dxcVTiBio/o2hrIuyJog4KD9dJI9i0BHhjcNNyMIv3P7T1f
5NlB2A3f7IcbyqmwuirNyQ7lANJmJb06IdH7+pm8lxq/c3yCsEy+2EqFkExsgftpZLhLGzRBK0Zp
eEJsKZMJSRA+C64FYPIHVbwL/UcPWPPwB8yLNu7N1N5NURSKJXsVA1S7pLodUv2oO4srlUoHV48x
uFqOvpw33yBrTBEmIqlMIY/BP5ktm6vQmDtNKaf1lOKfFxiCmeZuQmEFzwTOzAfrRcCwsSLEkJzx
FzxMG+Is3KYai3z7OjbdmVlhi2+6erPZCxYvQuH+dOr5Opn5CAT8g/ZHjmqehaQxK01hmQ6H8ipM
ReMmYJhk3FoH391StPyen/87I0k9hRw/jE93+bZ5t/GfkAlX79yTS1aQbh++BA1QhcxE2sFHxuOZ
iZgVAUnp8PzDgPvzjkY4jh43aNgBaYwKroH4P7+fnKuPx+iB8rZl+dKI7zpgLqsui9K1Of1byCTw
HO0R1tLDZ0a45Wa8sLeBOJFaUNyUa3ndYC13lqAJae5pVHOyBq56wpUI9wgAMYQvwLl2Zotd3kCG
3lZlWy6qM4bunVXGE6qj+zgbQGuZ2pod4Yr08R6jcBqEYw7H+DKlJuzP1pVZpZ3lPHqso+TWmWge
pTLeKXK1RwRACp9IiWmCRHKvR7r7Lbkt4Yj+++1KoMEaWrTjwGvYgEdxW5noAmlfHEVskjEmMDef
oQX93Wyqd1JemhMAlIBfpcKBjBhr07b7DmOH1eTrFD85Wx5TBas2FF+l3bbP3KgZnVog4JH5oZdn
CoZrheVAD7KHLDGa621a0ZiLSHArqPXusC6/6BjkSktm5BJ4Mo6o6ZXGEF3gyj6bEWdqDRnExtGH
n8OxSIcM3CUyJX5orA51Dqi1Nz2wXUHgewTR3AUGPliYbkHY1n6Gg5ktIjK/9KA93AWC4GcZEjNt
9HbwwLQAKftjtrnC76qTTn1Z+VYll8C1yTVEfFJLEJEfdAfycNGJ2ai9H/TltK3HVXFPBxf3QfvY
JWaGIxdJE5TDOU0BmmoV2NSile9G/FyqlwSajauEZKTzH2Wlu6KWSdB9oO1nQOf0l0+wX79zH5qc
0fbJcE/6BknJ+6ditxFM9xlEvJe5kqkYTbVhM60f7BmzMf1g/pZUNUn2lJSP1jwbPEaL37BKgGvB
+wzxLyCqMe0XI2GZavn9idsj3VINgUK6Dt348w9i1v02fibbKqlD0ByQqgdTWxP/7AFxtDTWLvNE
IxgxpqCcTA/De6z5Qy46FdDhLECB8VYgg5WRzfL/Gi5VLIieMO5eKlPCAOi98ruvdvh5vY8TLPVV
lZpGNIOah7ebNZrmNEWMWoZLKrThu0kYTVB0gC1g1MCfohME3DkKRFNCvXjpNV17hasqe/bLc16a
37NMgP6qprq1cRkGGxbx3YWJjwm+Hx5u9+kAUw9JfnpIqeYNk8tLRSPpPghdvEkU5Rplj5iz66jW
5pL1wik2WDL3ocazAgCuf04V6IYPCzKT6xyUsb8wya7QdkDhf+4ZriAog+nskMsQsM9FnDVVM0FX
AtlYiWu9lfJsc3cuDGE12QWc7ZvOh4Evy5HDCzxZhVBZbnQmkDiH8xIQdhR6CwzyLXfK8exOnWA+
Uy9aBjxl3OS/643dCqE04AWcs+cVH8KQunuzl/Bow14iKFht9iHSLvH5Kat/odK8gKa0UN/7hU9v
SpmqjoarYMh1n45v0rqvUsakWX/yjo37iSChqFQ7j0mWUMK9U3vGPhnjA3bj/dearDLRdpjy4CC1
oZr73i3YAr9p6cAMZUlhvfK3ix0J9Zu3Skq0JAYMVc7u1AbUJrI3icuZvHo/FIw4CfZm2ipSju0A
0JJuZCq42wECvQujCktI19fWTdFfwjQQGKG/WLisXes+3nnEh8enWLTZp254Wwg0rclxANlerOET
YM9RQb+vz6VyOCiacqOVHXT24UMoPVzSatCaWv7RGlJGam/oQep4fGmh+YQc8fWj2etT4SzClJqG
sfUPvguezZ52oRsrZvJzTI84mYoPLLnfvA6DK8mfZ8ssuWROI8+ckTOl0gc0mQ1toRJUvQ/UJ1p8
h1eUREeLvlVpUTpx8xMi47jWm5fBhx5vN1mGVsq/T0ydrADdS15y0L54yEgDfUW0b00+rgsdh5nb
RWjcj338N1VxFQ6K6dnEcftCyCfMwSLO947YdHev6OibF8pZqwW5yPjsfcQ1T7y5HtMkXFYrnj87
7v+zbFlinxB/vbVspFUhC/NHB1BBfoYsOzZvwlPO2fv8HX1pOC2oq+nGlIHJQCCdVP7tChAhYTSv
aW8jAxE+0icG241LD1+ed3wZ3dVHQQGowaPYV71Cwh0Tqapcu9acCsKKZ9BQy8KzZFKcPE0xf2eL
gitySHZYdZ5Rn4tnWTZZNU6wmWkWJ4juqsxFeiAAGhXw1w04aQKFbQ00lSyN359grKaaugc0yRJf
azpKNJt0lehoUzco1Va55OZDPlGVQSbfLKF6VIRwAPvwEEmAnX9j7cqEjzqrhoJCcty12I5YR95D
68hJBDuYhM84MS5QhSg6oJMvc6CZ3OlGFEXZg2ChwmfSAVF+nNLm5cWFHxXut/6jtHlRbC/JuhMv
P6FSHUubR2sH+Y56kNYgqn326yaVXXJ41ghJZ/q2aZvfMkIelfjGumCflk63XGrN+rW53Ri6HmBV
JKKleSOwWNRiGGSkZu2KE/CQdAcGowTd9wiRGdPG+O8OnxBA2fNKkZgFl8XYAfVLg2pYNaOufwnx
eDa005mPWqj/LWg5Rtingt53OP07cmbW0cfS5eb9Jxit6CS/6hb3K9K4+FXhG7zH2it0MJIivWn9
qejjZQTVrn7MLPlezOPzON6i+QNTTcgqsorVZD2cIWrqn9hB6k9guIGZd/1HndAwdXniOLIJ4klP
5xkJFAH4pOQrL5fnkmL0Dftwh8Upi2axktePJdo7/OudivJ51WE3Kevaf5nxMWuhu7zTzQqjCFkA
yqZQWYSID7nElcNcXjsCf92kU+FKiAJm+EKg8koN56hHFj9MC4gX9jHmB+Ybz54tL2pW+5GxBWu8
KsDqOu3SsYnn/8uxNQfbtyH2TTEN+RYcluioJuBD7s1SBprD0967OTVfacSG2ByCsP9W5dbEEj+B
Du/byn+wZJufm4n1JkSvhMU/RqwmJ85IuYfSqAUuTrlRUdjN8YBg6U2iswlxBVUioEn6SD2bN0Mf
6FU18HKblvB1BuYqkFx0MvyN+c0noybDoow4GS1PW95ycU6UT8Bd3SMBfanaIoBnsRo7NVBQgQNG
V2B0PjvZMlByGKE0ljXAArgjFbcJnpkOinezCLTvom7rsOYmiFejWeoYex4UCnyptCQPIzxFM+rK
MZKtrxcNH6njd6ZTtNAlEz23fp937hGBsAa8u4blxcUA9HtC5XF3qWhF29PzsXd/9Pbc4cUIbZd6
r/Ys+EeYbv2kdotbfsLe/UHwaOfZAQGFSZTw8CjSZm0vpQpf1jUpblvexTfpDbtu2/XN9InH9w3r
Zav9kYaJYMzOAaa7D3EnruAVjsv+14Yzw6D92PdScsb/oZJk09DN+Mi5NPmssX9pl11vFVkvnIJg
NvkpcGWYa0A+tDVk3cm9QcaXogsL3hAhVMW9KQs21WoJf97DcMa9GrMN5XUtXr+UBVtHoNEIrXYd
vbrgmTRmZ744tXkkj3It62IXNF8DxONFBuDG0RKC4hKWy+OXSAP5SEHygCMC8XI8Gzq4K8yA7XeV
6DhoCjP3J8JGRrGLVl5qzZx6pbOop1eKO69fSozYYydbju4MK6jOOZFJ+9XxFod/ZU4wXQBT5WNS
/cOWp+HyyMtkkpFUJAevDhNzIXH+idvBogmZlbnHz0yqGJM4Ffk9VZCekjnmC42AWzQqZcQPmmrE
GPGxl6+WLPi4EqCpdvnGbyWQiqXPdKa0dFizwyatun70xqzINyHMNweW6KZTouaQLIv8cy8svVXT
vin8ib+2N+2/keY+uevEwCAAkpGjNw/vZ5gBY1ZKqWXuG0c4XUNZxq1lDKepCGuPtDH34LtEXDNU
HumLVqLhEl3CYKBtet1iGoaeJAzMyyLdeRp9l736iqrUSXDAvoFFKoLTnrOqccIZMTe8hLHqF25l
bbv87F6n/bpFT+3eLrplAWcI7WUKRagEKRLxMnf9T35a7OkuynlOKvooDjAO43X1nkkcvGbXuUnI
O/8WSDJpb802nthXrKVggosHhCItxwni2ZeVk7N9s6vDiMR6EtzEDDZYSLgwvE/018G56QHBIOUx
EXSNkAwNJCa7xyo2/nQfxUWUp50hZk9PYUXhSopBZM83KiA1dyPFnL06PXWUPY6S2PM78x8/myXU
4i8oblYTfXirrdgeTP9Vw6PO5tooXno7c3R6Tuj3DlQKLVm2+6GW8QUECZQf0YI0G9e/iQd8vja5
2I6SyoNzWplnt+L91WFbNx7aUk3z4d6KJXG3OUbtW/QecwyUrDgcyupwLuuwNKzRKbGZJUGqMjV+
9D7jgrO9kurYfcYWLlFKA6LBH6Kzm4vKXUXKDlOBjKmvRmsYNdC/9k/+IvcNKKvHZCtWGclP1ldW
MjKMxSxfzU89iadvfoz6mBtl1saWWorY9pbQOjgcFUle9xmn7OvaAFmZwdg1kRi5u/Uu+CxrBRUJ
xXyrLNdgGDh3xOk/WJWdcPHnQJat2EKGi9LAY3G6ri2UrSnMa0k4pouYnUoiv9wlwEMMM4+YvqBF
v1Fl58iGaFTVZo2gZp6qGKFplHrk+oQaVOY6WQ8nBwziM5DyAI7/9YsPpB27Iy34p0/0hrjIDtPx
+QDjRsqK1CeHz5+avBg113+9oYaVTuAumDO31Tyk6uVnSLPvIpkMPRitnEP+0mlGaJDv0xet5Ywh
kZn/iNXCjH9z0B/Z2XzNUxAMFTs+DOOiI/q0ga9nWfO7f1cC4zW9++K6Lv9brbL2kIRLtz39Oekx
SConjW0x5CTMGkh5178vfnaKlrl36o4xcX2m6TO4rbJuuAQoDaTcWXTUo+KdQlPN+vU9sQXcPadg
F3pBHDNTwEaiX4temv+LCT38VoENWUW7XT4uh3ELEpiS9NMDKWM08P5NUl7oyfEhCY5TghpCj48i
KpfduCLpqEjpb8OWlkncR8B7ieliyb5TgcCauRj9TE4mfp9n34SW6NPH4lkZ+sBlfcXCRPyJF/8p
KdYwcvg0Ml7XQKRPyb4QBHngQrQFM+BC/7EppDwOtEmUT8bIamYPiELx1zlvhWOUs8ddz5A/dhco
7hm74FZt3bn+6C8nP53Q8JqdVZbvtoo2FfM3z274Y10I766kjTVOk1YSuRYxWnbPcY9iqYAXRvpw
ZyMZ21a+U2L4UCY2BxXJA9at5zBlERIgTm0BtGY3sChxF9a0+0DkWyMZyHkjzaaiHCvke4IeHn87
MDZwOhU1m8kPL2pstv1hFsKXtG94EEZrZf5VgSFYM2hPRiYOVkjtXQrNkNBIp3uracNst6H75JeM
yHc30opP2O2/dvLzA69+Gpyr8A0UgVbeNApicBUSWZRs9yds6LjsvosLItpyBI7hf4+GNq0pLs9v
SWHPvH+D1dPOSRGfqeA64CsGLhQ3/GQvoD3FTwCyzEAQ/SlXhAGpiQJy2T22kjOeXjQ50jyoCoPC
6lW+6tFqQfJzmUjm+34LamaAHsM+ZHg9d8ARGhJNYdZ6X3H63zxm6DZXrG057qvQscYA87C0HltQ
AjawfL6kwdoPbEZyeo/dAc5KGsDe3pQ/6xGwjvnmDrwDNOelcn+TsSkIkVDdhZDkR+OpAdRiJnNq
ErYN21KHsRVJkLqXkMZ1JCkcPz8oVVB5kLI2nsBRL1IW2SZhqm6q/RtexBia5HopEpcyuSiZTEqW
c918uo16lGvj5b1Z8fsvNKf1TAcuEqMfBxmPtb8NNkUb2j4B8IEZmwRXQC118E94epJo99LFaso/
Wr0qDqE9UZ3lxOMuYntUtYTrZfwCRF/ySXcMhRxv+Fi6zLkd9o3qNqpdnYmzSD2sxMEtuoYjDMXB
aOX648KSxHx2CzQgKFc8Ue5XfrfLloivgLIlnqCf3avzMpUjn1aYwFvsNBH3zrasarjIlFtHC1nn
VEvSUDdMxjphFVOK+VIRbjgOA15g25xTVU2+unNAZJS+4eKvpU/DWfQgDq9IpYm9T8//BLuNkQSA
UGMIGwjKimfNa9wfl4H9PTsxA+TYF/xwDXDUFT3/WfvkbNWpAOfNpIDfXt+Px9pxuVTk4nUPPbqK
IrASjACREm1QHh1jsY30EiXCqjntseDeShw9nROk9i3qhUxNx3pl9yexycG5N7AAY2pKJ899PSqZ
ZrTM0TvZMJHBAJe+6AvLyU90hobHO2sD3QLsJZy7zIzqgGobGgusEbOvcw0ncYymgKX50H9hCFVL
dNBJUr5Z4JObN9O5rMOJ7hTTq98bbJ8yLBXzApiT14VFkuS06pVkKK3nTGqgnbhnMsX45ZcFLxmA
JudbBolxJA+aULoeYSbo6+7eT8+hnA/T1l78ycSGpuzIUqFDXS//ML0hffXEzkm3ycdZmwifHBl1
BoSxuJVn75greXEjq2KNIpo2KXlTUsqGrwsaozdA8fYtoKgfJreTpgNdInOrMc+I6/Oaa4GzLzEI
nQYR3pBwkLSLu80xRcohJoPIGcQ/3qy0gRogROOVgwA2xy04poMUS8OYBhuBQyaO2UM4AFRPyzTq
CMEmrv2ZcuyYWID5lGUnTKzUeE/bVsb/mpHiS8bkRwS+UNxl7tLZLXDRUMhlujcQysTEZRzsNKy4
vmGRUmJxk+SmaJtkXd1q6hjazHrDztn8t5nWCnOiN2SqYCjF35YUFXnfhqViYgtKI9V8eioFhvSX
/9Qf5fQWORySYy1MPsMEE0ZGxnLmtfQRf2hBmofUPcjN+ITx5brZaa104O34UiENxFMarnfstg2Y
bx0XOrmNCQT/fa98uGLJOBVnejKwVKL/E0tNGjg6DJR9fSkt+LlWzTLzFMnxfsnZedKFkd8z5qOb
9Gtwk2Gi6e2NSTFF1Adhd0Lf9q1BJCFfalhEkUk6BtdJmmWHrFSkcZHSXyLeCRDndJakLs37GCFT
UNgj7JW6Fn9yfe47lekTQT3l/FlOR3H+gF2Vkfg24bXBlfuUePAgNOzva7o62jlLjMgTey+5arwi
HwaNCFNauO8OghwtIF4VUJ0TSO2Fq8OC8LhB7SUga0u2QTHQV5X0+BfYVN7GCfkpgMbSh+L3P3pB
G4zHB/kFfKX8fV4pxf6u+tW25LYurHrcx+gIx2Ioei8NPEQeQPDTma6IvjWwR/TQRPUKZuio2Da8
qgvWMdBDFcKVNzmGiDywq5sYYQPST1Xr7WJ9bH6i9OnWoLgbkOPqvYfMBothrNwk0o9MnoewoVjP
g76QWu6C2o3YeApYShIOZ8XZgDNGbkpmiasDTPriRwLqcMEHAUjDk9V5Ye9PgVdk+xfzZiezAlNE
jbKRBtHpKCPgiw4+mv1uhBY3rOJaY75hItDChNUUcIqQuxSt62GMxjmGmbJGMN+zsvYv1ISdJNb+
/uborlj3IvFd8VCu+hibByb5K79ei96VGdJ9CodsJzPhEwA2RbR5R1+1Gd42jrnUfKSAJ3aK5b+L
swd9/sTdN1GJzYDkfLC6BMMKv26eyrllQljxrMWCk1pWO6GxMCspORKIQXFFjnqXFw3a92u38zDt
J/hK7daI+OFuS5baPTJkiXHOcVfx9kkeNoHqZ20Mo0IuNIT1UKuth9Ry+iDbL2X8HCd8Qce+cBB8
NpQUp4DLdXtAC3HVHw6tNNkGz4wVOUpkDimAy+YgQPYN2wVWT1qPoi5zI/+j1QztTsTBJeLLCaI8
bIRu6NSBh7ekmZIoko6FW/eo2YScA/VFI8NQcrceyFpBCeDkMDWaWoTyk0qzQFw5VUmu3zCLgxT6
oIs7em8oMLIUYAvs+VK3ojj7f4gH+tnN3WJ0gkkp6pmwh1wA78hfIsrNm0hWpBJ9sZONEREkRI8O
GNF6Q9SoNyS+U+Ses2AZS/sW1IR9nuR2S8CoqEeJ9oM/A5IHbBiZA2dUcA9hAWwaXihlu3yzXt+s
iUy+uCp1UlFHjsoIyBiJ9ATj7Fj0WnlwVBSaRsKyhWA8b8YrwRpM5gjL8HFpUISIB19ePpat5u/5
CZ3VlzpoAyBcTyIG0wiwaO1mt59TC7EuvbqyJwklO5isEXFvTYXrvyUt/HkIkUOSnOgKjahAuRke
jwONGz/2hIy3qLAg6fKDgC+BdlC84w/jmIwsCr8sY3NWWYe+vLj6yFnNpcgzdqyz4LVKQD7On7wz
MTnqonXpECPkPRlnSMVh8Stx5ba5ZRh0VRhDhWFQ7YyA9SEcv+ZcE0eN750JV/pX0RnCm+S+8EBv
YiKBJkSnoesM1hHzpEcRvIiI3811ycywMsJ5O96476LQ5Idp3om1CKuzOuk+QG6bu3zruCkxhA0x
AWr+amBv70kWbWjjV0dXyUr9I9+bxw/upmxX7NlMih/gbSwjMi4MNF2Ah/wNfpSu3+Uy5OkrmHGU
k4QXkMrIX/TWV0091rrlMQmo4XxLbE07UjeEoVxssTRYDVsOiaKu37ZPAbIYQhVYEuP4mvrZ7SZG
Tqc0YmeLbivMpLIwtBDomrNc/f12VvuC/veOJFHXPDMN0Qjmek7JV7tLcsXqvuO3rr6Y9vkIeUmi
rq7GfYP8L6jYlfAu5UwgSfDqU7aErPiutDhB9mT0XmVCTgUw4W2ydoXj+uCAHmYHU64xyXS5OwJO
0zGIRJTaG/FPAA7tMoH/b5JjhQjJSvhdfuGKX+jdEFfm9Q0IcAEwaW/hpG7Ee+kJjQXe8LsjOe+1
nU0QG7Eh+MsdTvz7ArzTCcn/wVjvF5LjGSrQvbWjB3jSXwvrRRzHlIyJ4B/Lxh6kk3SrZzUIeRR1
bW9TDBVQzk2Mmru4XsQA8Ph9o8C+k9FOv2AUUS76HJFa7XdsCeXJsRl1fd4FeEmlG7Dl7sPVqH6s
DeFTaHD4Lj7rTMciGhsbKcerNe3OvnxOeniTMitU1rnCVvgK9OUeT99nh2X6BkWrG1FZd6rqcg4L
bOcNQ71ipOzTUdxyWeZBoWssOjOwqaGEwgsSFZrBxdFlepFG7o/0RfpXrZR2/SKQrAQaZX0wyqU6
6ENzxG5YzV39s04Wqt2s3nMQ4sD542iC6rlGF3bAWF+oymY4PCo31PT+d+ujwk41mEwFmZPiMkfz
ZFx99EOJ4l8+8RKp0kBiaZOMqCMVA1lSBTA1zh3/oKPmKiYDN42X8HXTO0KajWTL1LpAVnrurWfg
KnNPEuuAabAioEvOrGjgEJTsyxrW2Jp5FNBBHztH9hf2ESkM4D8yJ0kJpYMucrZrD3gOEadj+to1
wX7tV8HOmymPbC5AaPPusl64thBhM5zxRlpF+HJQiYlMrrxFtGVpO/8SYmNV1kg61N4iJ2PpsofH
X3kdYb1nkOe4bYmtbSp9ejBB5JqFFrDgICLwclhh+81B6tFf7nGRodODwy2Bmzg72rlVkJTQIqf6
U4Z0havst6LfBlvut4q2UtqjHu5sQpRVDwoyGLqNLtF+fRjzn1gV+gBBgyvGpTLaq/zve9/7cMea
HauQJE03SRV6YmnTx7b1f+SGs4RB02yMuEW7R3Lg+OCvXBtoypk8FTenB8UHcUk6nLBAtuX3zMDm
ZffIZpNTY2JwSd+V7xyDeQWnkz7yMWsP8/2SKnje2yrpBmFgbavFd7cssgZvVoht9XzFXKCRXre5
OhfMn717boE9UrcptxW9qgc8/2P4WIysKsc9L7XqY38/0mP05sTXWqAGAuzCmtq2A046ifV2m8Oj
Qi9maLLHh+cEDpro6gFvdhASsT1znjmTd+BH3OpmjkyyfhPMMErB9mLRF9YfXTW5aDLi06bGSohD
Cqf3sTZ7Qd7Oj7lgy6quvlIpHrCheoXAh50iMsp1eLF5dtuvAz3eLzWrrO8ivKwwr9bSw0gvPSsX
cApBleDGtKX7q512E40rChYjAF87BshHEraPQA7GDCEKpK56+PrI4Dco9aiktF1J6xhNuxmYeTXp
ayX6wAYpbFGNIr22ci16sPWlRFMb1fNEq564DY0eLnyOHt2//voPXoAHyJW/73L3USIA0FMaatlE
SmsDavLC0QVB2g0O/hsTpk/ezJwkQDP20X7J2Yb8BMAKazzxWFVqEownEhFWl/iRNwmMajEuGozD
NaYnWcl2urTK322gR3BzUF87tnHL/JMFRUDEcFtbvz+bVle1jpOnaMkfmlppvJxSOlKCx3H1aRs1
UM8/1/wncq2VhFdlUnRitwzsp2J+EUY6Qj1hv8QmoVNpq/Fr9dgEjCI+VxqpfEdu3sE3wkIa8A7I
TR+AX5Y3TWTw6+9WXdK/u9Nrl+Geg6YkKcT68xKd3o0OmizjqS40iiLp7ZqUcNHsFN1nuXR1J67x
IMi+F1aP7LRyoTb7adF/LA51ubAmB+9K+s0oMIcglecN69awz+PmvTRxaAG2zOHZLOVI2PxiTmEc
r7/Nlu7fMwJVZION+1McBZS5ZzsszOmvJKG2lCimLrxpzMDPLeWynwZ4ey8RHHNhYEg30+xDS8Ip
QVLvFpgTQ7hsbokx8VXjUFPbCmuD0rhtvzD+f6PnxknYZdZtv+PH+/qEkTQG+CtA+dMTyey1PUnB
9eqxzsDFPsR40YsjyIkHjzhbz0grykZSrybolLYW+XK3Qa0apWxjnqVCcWdwdspc8v0a4rVUWtks
hJHX7l3dPJiv6UgDpJIEqVvX0yqLnDnggkmk2HStu0iH6aQnBDS0ZiqmiHzSpXEtgpjc7n+Ho58K
0+JQQXbUe4QS4CcFxlVngnRQsQPsp2wJrdIQ1KtcbyYIZs/gWL8ITjpe089o2wau5QKR43nw7Q8k
Qd6jGWJ4xhULCMWwkY4aQJlSo3ROKaVFc/L5GIxl0ejtiWsx440RWTmcdMcUNdt5yY8aMoJVW7xb
Xi9TFgc5EpESqNNE0whNV06F2F15FqOJWh2YYQkhT16evsCzA4WhNb3srAoYu3qu8o5nmFtdg6fp
VMoHHvYZUfSh9A4k1b0vl5XRdmRuI+wAICDTSIqNfOwKYrTEHbAVQUJOweU16rdalCQBhVSSVHjE
LcDZbhJnDjS5/P2HP/XvfEuQVgEz+7k3se7tzWuBvBND1I3AzQwv5lYPJgMNu7pUjfVoMen/KSFR
OT6IEilMkpkWThFxFZqMB5EN1PT+hdGtEfpgc3fgpYcuJ1Imn+nbbfsn1LpCqaHb3XXLGOkUNgmA
zr3shKWMDwxv8GKPgjVA6gByp3nh6DaJ9ZfbvgoK2PL6bltaMtVUjFj2xDl6r0UFOOI3iyf1Tun8
vGczrnZ0U/sA17haWHxzP5UKWE+jY4bbX18iWYHKiaU7fZb9sA4MQJuYoCFS0CZ67m66VSdYF3kC
Qx6TSj+1voSpCCPcrJwUWT+X6v5bn7JeB0BeHuB/m+TvUU1mjQJiq3YVsNcycM5pFULit7ekrsZw
hwVmYAp092oo6mjdYZG1MLskMtFO/ixnyUgcDShHW5P2ru7Hpesi/m+BRygHb3ojCs8wI7uso6xm
alZyR1gfN4MPSey+2NjxYANzJU86iQWWwRrTtU/6ShcX+4beXWsaF/jsSPzJEbkWlhOj0k+jph5o
lvcYbXQZmqlgxu/7iao7jSnhub3zEMscZTvlTd3jx+yz2c1EiPMQaRLg/N5sinJrvRzcy+vpflG5
qEDGbUGt3tKOD+w/9EKzlH/cMX8IQyqM236ETuQrtUAmG+xsUJqwjB6rocCdtTgc0x7J1Np/F+7G
8MeAgDyrHrE6TcHT3a9Xl3gsRmcK9SHE7mPYh8ZZx6wMu3Z7DR4n17rj3cAMPEt91qZhqWKx/BJ1
P3tT3bPA8TldBhqyyE8jhZPnfGGSi2nTWl7yoWO1XXDkr5lae9JrVPXHhmyjKX4SYNpvbOusbfRL
3EgAoZU6S8e3fiNlJ0p1w6auR9MZtfZNkT78t4fTgij3OMJ8Wkszup80ElJlJK1nh13ZjpHZtmU6
eZbYVZtxZiQdq8Sv54VYpFcE8jdP5VvxtRIIsDIOOxpEvioZIUwfVo3SXPvHsSs+NBGtUCrpCKyc
odjGhaNjE4sx416LgNURN0YIJe/+Egfmh8enKys40hScvUt/nyl0s5GcOrIt0VlKyYlWGzvs7gBH
yGKkGocwh3bOFlfIZbM2D59V4KNCfLEaX3dLVm7aS451gOoTlZ+EHhsTr3bx9QNBYqCsNcW/0lru
Skr/BhMcXYuqCtpddFrO7W4UYe17DTa78q+rLc3gIlSTYdFNdHVg/QEu6sSyXHSeZd3N+U7cmxc/
555KYopfCNzVssXX22woMcfGKLfmvpjGkkPB3VDaI1o5C6dmcDcT2sompzdvu/qYq253RK2FvpYX
5nbUQZEbRPeniqX7W6bX6sAgqjMIpE9lf7JF3+LguftCFmcodWgDwhBRRI8ZijJ5Y4pjDR93UyG8
EVJK4jRv8zSy4v1Ayuo8HgtZUyo5R4oI4bKWkaWhU9W8qhfQy+OKJFAM5zrc65sRSSbYkcGOzX+q
v4/YGVc+B/C2zFGf2eup0TIeMW+UP39DCAKSATDJXfybNjNVsWOpTjsZ7BaE+0VVQf4IIdZLlU7Q
bE6Kvc1omy7xa4+g4y7p+xbnDIzrR1bEaIL3LepuIyeeTFKAkT58nLdqhUiJZFT0tfrxmlFxnkkC
3jAhu/kx7cV4aNnR8bt37lz8NERpnMRvuUQu8udye10g7yTkSRPz8eoC5So1TzQvq3SIk80F0zqK
eLkP9BjCgdMUzFKKtegDXZcX3TC0VbEt4SDVnlmPpVpOchXgklN4T3z/6hM7y+WJC6IN0qgpNoOe
1VuG3WEdprHtE1ek2YxW2oynHB02KV+mpzfDz8RPPR6SqePpt8TJjrUn5XChRJrJx9ad3xatGc3x
u/OmEubajVMBxPnm/9ZfPGiof5OiDkF4n20M2kd79PkplMha4diT4Bgqs6v3/FZLopecPaUTOxJn
61A7F25fpN6gbAhbaoZMGJwnB2n0xs+ejF9hWgUMmiFJzxlKDRq7lBGfHmOUN+Pq+GtVFYuOh0bz
y8Re1remURoOebAkSzoi3VsKe8u70wKnjNYdT8Nc5kH33DGNKDsNs2vv8MOZIvwxYhokQ8PgJ0vH
EYcFEcvNl5qMbVMnp7KrvwWhrYOl0oEwFryl9OmuejrieL56Jgs0tJRNgm6lNkc+CnvPC6Gbn1MZ
WXHGbyvGk37K5FLSj3dK/xmdQZdBJwdiztIQVo30AmlTvev0vbUc5DvVR9WC9LHuVzIS3IhQ/9Jw
wwHkGVpsLO8AdL+wZhaVMBUFfUv6dk0a+xTOmJ5CAOdK/xAWBvGyQIef2+tsPxpPIgYc+dodRyFj
koRXnIEjhvBKhzGBFwX+6omGgFJgG2qftNArmPO9m2S4nyvbSvZ/C6LZDQS217wtZCLMhnFti1fN
L9e86Obxtvvn76NYwXDPJ2fMoGNJDTwAfm6wslFRznw4vD/bT5GsQFFeQTn7d5HYWBtks+inPyrO
19lsikRI7Yp3bCjG585FwJIzaDwmt6+qJ6sE07mU/13ovba0a8whprb6GAEnY0AjXrhipOxwZBaL
pjitaDOiLWpbDEe/bOHuo+lSU3J1DdNX6WoPxwEbp16K8hfxtDaSkIu1qeMAhe0SRZwpbuj9QHDx
MEUwa/nDE5V7b85mEZotrwvenUbyrb8FGcMFdPCCqQB3Z+d1OJffyexJKDjGA7J0LP3HKiP5a1UZ
YWn+8cNa3Q51MC8cTPY098atowk6fVtafbbuKZHN+IMqDo0sKDWaP8qOoC2d7cA45usqm8d1wvev
54T5amYh5NdwIklIzrjxbYZeq2CnHBm/VnLxNKrA59+4KkEZyPwLLAPFv445+3fjak4FNRzOuT/t
JZJid9RZ0hwGXeaaP/vVzYG3hPZgewVGLg2jPZkUAOhHFRHcGsWDQgnDPpdj27Fh5UDwero27E3B
tzF+f5jZRKM+fAarOwHpjmSQrEsEikHpy9w0WyTBoRHI7a9ip6y1Ixaar7t/lFbW0Oxm2ekApyfJ
AUxv21SixsbDZdl0Qoiwsx32NlTslJl5wfMQOk8sRdUTqdnF5J/xwIP6SaPViK90+wbUmoHV4LRQ
Csg920Se9s8t3g5T6VhpsEExp+CGUd7tGfOSXUg/OBGdgojOahqTzs4nywl1ThTQbBUBPqrjTXu9
I0uqD4qWdoUi3BqC9cstGODsyVmr25n5Pt/oXgQGCViuhwEa/mqvhsBKSareyDhFiGDmBRda6I8y
e/gY7QcWDs6NUbgKSTKKx+PJnwqfXgEmP5lxlflSKRpVsRCtEYEf0o/4xues5RIRSncZvJ8VkeFt
wEUh5a1Ce9mhnnGAYMPutFu6KaZ+KOzwSksLKej2OyfGrnA7DWXFlniGso1QDRNM+I9CI8p/xl04
lVQqarFylMFS6Qz380zNbY1dLOjaVSoD14Y7qQoxZzvCdyhQMuii3Zb0eRmCPDkchxKgHFo+qDHh
DTcG/AP2At4RsegJgrCqtbx7FSK9BSHu5aybDzYiFhv2PUEldL9vjJMIVXaXKHdnh+e0ZJ2t2b0V
rvR7KNib1q8sDkAdlYcPxTl1jg2PD3jJ7a/e3A5EGTKvmyLqIDmYNgss3jPc0KEpP/8020HMgs0j
svYQ0eNcCGQ6/kCUcFOX6l5r8YO02LlqQkq7/gB//TKXaHmUau38DK7ei+BkeO9NfcmZX8NBWm2z
oM0SebKD77bdqM36skRfPiol/gjWQULVz8Q1s+KQnq3Rwlwl0Pc3Paj7XWO94sxndXkYCFpC7DWm
fHwjY0OjKi/Td4GVjPZUxaMBURnX4mvleMNtlMdWaInN2Dn08kce9BaDHxGpCm3BhrhQBWJQmSav
ePlhfskwrcpkVSaHaxYFhNaCh6rexFDgNWUKQs6ww1PgZjkiAQg60G8+lOfsMHtxG4rFaFSZQxfM
IYmWq8ICN/edRZXn+qNjYcaXSZVAPvXEqJjgNuaSuq0kxiX36s8OletdGGh8MW0UGY/TvzRJBe7x
BKBBZYfm9PMHmk51zgxg0gXKVIoei6iFf4gfiuriJnecAnpgBHHnSI+4PUgEI7CxeNC8JN4vgCWW
WldKDvTK8tplohHmjyM52dLg8Zv8aKvrs0lLVDdkNieAV116fZJKpgUNqqh+kJZ437KzxiMH65pp
M1tymXaHnm2BubFjYg6cuv/CeMedxKU5Lsc5Vi67opy3+v+X0FcgQM8v3UuHcAD7l3o3U6LW1fbv
+Kyl4FlasOY9bNdjXvSgi6Z800+wqa5rDVsGsNRaqT+c372YkLCg7tNlnCEDjIN0AE5dH36QXm6v
YFZv9H5DRDRhhBGpeyQ9uBUB9XcXHZGFhYDg8EV6kPW0I8q6SZ5b+HL5XmeBaVuAcYLXsJHLzzob
MaQwOl6cnStvyYLFxFvMaOKpmncOFwL5IxgUI3PkBfO3asBGD9zErHhrknHkzRrC8DTchlT+rbYH
JF3/28jUjWGtNslT2hU0m97uiVXMhTP5ao+gcWHJcW2ChyrRNnaMmsb85DFvva7Vh2ARPxXXFjUC
zNe8XMFlIs3tgs/xUKITcBK+neASJ2DXGf0mxJd4VHOWSjMDoaWYSYpZoN04NRcdWZYBy5Q/nCwd
SW4U9qt6q4zT4R6rr080ZnX9AotOW506hmtn/g6QBr6kPbyDjlSh2KvXt+4z8wWsmHkek0021mB7
XshmPk5LE7Cqtk42tax33hxtWYMnn0JSrMyG0GwD5jqouiuS91CoQsBcQCgpt6Xp2K2ScQiWsZDk
jReJWs9EHhykWHm4GSxKD5nm/bSrgJKbgUyMwN//SGqI1QKSANusC1kcHgp/lkDS1SZ1vztQvTb8
0v47HugNstG0yrRJ86kbYKyk0jD3/HkvsQ/o5MtSGb/aG8c8zR6gF3zhm2PtEX+vw4kvVHDpi0iX
z2G8SLUzZVNpnAC9MMw3H816sivJW6AZmEJJMTCD35F7gCg7gY/+8EAgJ3KSvqk/9VhiMDNxzr3D
HRoA5gaS8jCUWPNsiHa2hLynLbiQM1qQitlBJir4TLoXxN5PmeRkRbro1u7lJYuySRw1ke3Xrr9o
32YaFzO/BKA/MOq5TJIwlv4eF8JbvvqNsOavWfY6pZ1naiW3KEC8jVuVOfExvzdbvjCDZ/6gZ6sN
Vdupk5dvZmONPIGAS/9+kLVnUcBofmwa47dQ5jUkeLqG5j1eB2Km67iXQf8N/dTifVvCYdMGqi6W
Oo0p+8hN+t202ObsZdxCT9N96Lm5IOz/WZHIYyzL4mwhHfa7xvEruzaNFutXqmD0fnCIp7+xjHpz
XU6przShvuV2qfq9XSc/I5RP9pAsVoq5udHJIjAsWaQBdfZwiLb6y9dKIgZf1dbxBsI5dFpw0kYu
neQY1PHzmfcLD88C9K1QjJcjtobnUM3ZYLWO9jIEwgUswOmMVlA73956StXhsZzcsS8IbMOpFE/d
tH4FBT2FuRZkYANTgCGkgz2WLiVxSVEpGmNTS27dzVMRLPilhkE/deJeV8nI9iAInvMHejIlcWqK
3mCg0J8ZlcGHrYZ+A29X80pY4oAW+3z4Tqng/3Bn/JiHxjRWZKCIqgNBw82gTAIA0/Lq5pxpyxqy
wL7ufNSlmHhkGoDEELo0w+RDkA5hQ2NQR0RPCsCtx/KA6j4eYS6qzN7bP8NyjZeihD/80caXELeu
z6jkZ/u7erciRkFbGln5fdgqNgjpPxD1Mz6+wy8LhQH4hiROwrj7yhcPhuA1EnkSZHdM/4gl6tmb
EVGQsejXyxvgUP1SK1panhKvrXjFPP+HT/9MzNHseR6Sg7K6FYW1A+uvo9nDmNHnvhHU21NrIsxp
vXvCR3zPeaEKCK53X9Kgv5/vj1MqOm62moBM3/rmPgTTrvM7CbKitTKQbGHc8kUn7FNdhDdOR+Ls
A7wqsKx2xbxa2hTDlcvt5ZvDboHWQ1gZiiYkAkt4zCPLF/yOdpxI35/wnR9Isp3D8gmLbZdj58Ja
cyMwHeOPJS5f4Is3C2amj47TCZGR4AN+d2rTCkWnJM/ho+nP5GfJ1LZJ715wiS1jAAtNcjodP+uU
/PxyaqbNyQFt2p+fYfir/YIM6jbxuM7aSSCJ1yioBkn9Qnb6t2rUQx59/k4J6uI+AzGx9ZAPBof9
LFdBFETMsoSeoMwFDf748zFIWOujW/x8fnTUmRdsFEfqZyMxtN/A+lwPlRHc/oIrezxwTBuvPTW8
NBhv8eaMVG/IUWC0CbmCZZ4dEmaiyB/mokrLn5U68VqZ337O9VPSTmD1EPCuRNIaN0FLYv1vwKq0
sbPdxnsNiJzq8AdTp9k8tUdciqT5g1+a8nkdoP817fXyZirYGSPVMJLcDLsimMTUZLv+mAf/zun1
QtGcLzh9hUDAsTndftGto/7zo2HEgc9l3H10HWJ8eyZk458kozVfq3uw8af4z6d52mvFvYTPwSYd
38/EIjaPcLpvouzqtWbdoZ7/wRPn95yuX62ZeZvZ3k5hTx9BIVKFMMy1GmHlGS4Z4vZ/LKwZJmEJ
0lAK/kpI/ouJxzmalS5QIiHp+R327A605zl7Qhue+8taI/5Mj0hYOPInMRU0h9XwFgcQiNKKBUHv
rDMo8Zsan1vOF7CsW8qzTLB7HObiZD59+efcsrdIf5h8usBVRoJcSt/4vY8FYn5R9JU/F/s4kLdD
2ICFJeGLd1zi8h/3Ft1USAYcadTe7lTyOx9jp2LBRqHFsl2LHhW5EORtw7Y9fcHXRQic/dH65ouM
LbCRCtwqj7NDuVFuLVPl2DZI0IJaaj34WPiWjDw5Yv9fZV6wyGNLx3w8N5swVYgVCqcX4H7WuWXY
/MQ3F6fZv7TU/7luVQYLmVHdpnjwAU426EIc6MGTuSPiA2hCk3Z7bNiSYYZyxiyEkd2jnZnqYDru
QOphyULO2qL9yewgtTngI1oBtXAtKvKOh2OrOWSkY2l8OFUD/931hVPh+ufkNjq16j5HWm1FCN53
6kA/LPpm+TfJNpWNHYd8fHQHMrwq8VPoUBLfSjfMD/Gyx1V/V2SEk6p7zG2htcSxQCvrjAcSO7Lh
HWKTUs3nK5B/4a2VcvOwM6Z01s9YkdhD7KRweOEIsuS9bsjxzXryHLnNkButP5LAtLpag5K0aT7T
S5o2Ay7BaFCyyxlXu0RLTtVVdK/q8WYgiq+cxSAKn4mOPWSOLT6Z8IqYbQDO/+sPHrtvp9y94aV1
VB/krLeQjj9JaDvfQpx6urWE2ya6QLyDBtIidaK8/WFj/mNMO8Y/pxg5fZoN2ycz36Xrz9vP7RIo
9Bqoqg4922aIiTdzJyCvj8rrZaI749thJVdbnU+Ud1M1OPV9DhEq8V0EL1ogBJyDfV/cCHGLtF2+
E+yPGKI0Np+0MJY+6bk5xhk33P/h4AeQQyOVNpJI+0iUe854wlgMocdeIvFpQWdTBsxUZMtzY8QW
qapqIfj/SdNKtJe1h4p3YiClCMKDxdLCWi9zi/RaeeZHMsHKYBk7pxz0REYSh8BEozhZyPHrQuGw
LngUA8jyvlmhqWduUE0gb/ksaRSlW3Y+aACJG9KkYEaLQcaRa0WSMtwg0XfJjD7xpXDd/Fg8z8v/
KmBiuM+Nd9USn7eDTnXNEhOIlHljPEhx6NHpgE79536LDdANbpJS5gbH0xWIqAj5GLT2TJLXEnsI
4C4gF8OuvQuq7o1SZLfKBENxXGorXFYiaALnhstXCALXfp88MnveoK6+L0JTSHjvhYgOyQjcpxev
SzPgQar6U4jN+e7dbu5Ei8nYBA6ygC/BjWzc6s65uOHsVdaCnivJZl8frNWuWDNRK7IUxCQQHEtj
TR1DhRRBXVhpFKOWKbpt7TIpmWEt6t8B8vwKTn4qmZFnowXzyVyEbdTqKEml2E/GlBGUQCpl0yRM
jG1ltkVI3vURwOdZcTUwW97r3uqpmA/T0gmR5asYn3so7jEQgHOLOKo6MewB4P6qcEcZ0yOexAa4
iWc00e87C2339Xmojmneg1hAgVcMq1aRX2BtDNDTINCXBrMoHWRph1fqK+kLf/83QD33Ty2Ausar
Xuyi1qROF7J5QYk7kU+ZRs/GTjWisXAyTrHyYfaxGrex1w5IDfbmxuKk/5faQjlDjyWeV3P+8zyo
/GvJsSkP1YIjI0IOV/7ruMl8bV96v+FE5wOUlBFtqGS/+WlMCGofOBWgeDyKAwNI/ylxhueXAPVi
M49yid1vJx7g9BURJyHUyE8on3KKeEJSi/xBq4nJOMOH5lm5ZlSjrkEyi/19nKyQgBQ+gpV2ZC+m
dAGSq9odExHn80NxEEnkWWyHGLBX2uBxP3jT+CBkuFWsES7F+360sfXJAVX6dxAjYdHnFRjHC5QQ
kkEIUUdkt/hZDisqik59A+nOuWZSryg+lLvo7s1zk1UYueVZZ6popCKeS6+LLQyZKQ8Re8r0W0Vq
UVtwu4TJ5HNrxKblk2EVvIkn8OnO6Kz1vprHrkFaz6clW/q6zyd4uRPMrIHEBPRY7SySIdv7YSpw
/xlhRMDHtw5X4CvJW1cM7NtoYzth+Hu1/44lVLkdpQ4niqQenV5qdGalIdMjgSrDXkiNYPjzyPNn
TapCOQrLDaCBM7v20SG8NddQNyyjlg4EwNujxyapGoVs+AuBf5NW0zd96DF02I0bDbA1crFD3LUZ
Qk8CHyu9KR9aokvg823KR7zD83dmviiE4Ny6E4IRvpo/wWEzLyjSdBUsx/9SZTwjMKgONZYKS5iG
OZ+43D7YzoCXxsHTgL3RrjcNXQTGxK4NQMkeKhg1YWSMYrNa6UHhtJquqoT15dvLp9fBRoUa7++T
sadQu4hhty7BkSiHo9S77HTC8tp+1c+HrZo/fVxjwzTEMEmfNk84jkZc6nYWki8WLBQg4O1re+oA
yGQqqjAjANuwxnz1clNYMFKvCqRAxeFVfZ6fUOWXlAP0HiGrsm/NgWAzUVovtUHnjQI5tnnCR6DT
bf1JnCyhKLLLcmha4PNr7XQ+pbzquS5qttb7JoKQAEA32a1VRovSl7Cm3dwstq4/y0qu5tkdjMDV
0PUrECIZpi2DgSKRWfF4WGYolGt0ciLn3MIYayyBJvPcYMaxubkobuczQxWmeOYamkPy/podkMdA
VJyuesm2DjzgHWXm1iFz5J/RKeaySVzhwaC3aLK15y5RG7AGaUu/xz65dcZCRd/UaSKA9MUNqF0p
g966RWvRx4kSuBkt4sf0hRni+IIgA9siH7/wIIzFyoHqmzgbIKyo/X/WPqfXEm7LYmZtOj8TSls2
SKsuXNoVAkRaVDFp9+pCeCU7hFOUlGQkR9cImpjXKrfaUS5n92/D7pZqqihi0H96dQuBjLOi9val
vcndLknYD83eahFQyBWdRrafXLe7ipCoqvP15VG2gxzH3fXB6ls8Dxr9j/ZGU9oKY6KiGkaSiVs4
GqDT79daIY87rhgN/6MTGjtIlomgdqwrW9iQkRnSqlUno8LBCz6yMaU33sX5Pue68YzaXDIxxlA0
QykNqxlMnh6kzhLS3xq9Jo2IziJFt1PjuFIG+eyesz1YFCUGQqbus11+1gdHHnBsBGeDPNSR8XrZ
eY4BQK2DcchAif16AM4BTv6caUJiB80uYhNxMTXtimMd7ven4xILMIm8mpu94D625zRVBjC3Sp57
+vcTCuvitV9lmQuvU2uu1B9qZFjrhpjyl3CJil4TPiEiRZ87NGu+qOFIbSdhSaei03xRcw7iL7T2
7H4C+L7q/sBRdGnN4FgeE01JRsonDvUxXMeUmzSI26HPhdbfvrqxowP0+X74FxRnsWEXQISW62Wn
nFle/hrfmQwBeLxxBhNLQURGpLYKETrN4felR1w78IkUCCfdX+bEC1yjACmDBw1gCLFyYpB8/t00
IK589DjQh0lAK5zuUItyPSemZg8Uh0dzsWCQR+wpqi1C0+ArxtQAXwleTwOw/b2nzIS1rcraggwF
GgGc654p2Rey5UbEz0nE6cUkc9QMWoKf1BwWzwxH3tdFUBJVszoT0JMbyKws2upJghHd3II/h8Kw
iObSWuETq30ZDjX2SnxeoE21WOd2axy64Wc0Va6SRnSh1oUKLMND7mCr/zxBIabzzBfvBmzpXpNI
T/b2j9NUokxE5VQQszfSVwhVZqBW3Sxddotk22xhfJBh/N6OAf33rTzAPVH7cLhuDjGx17x5WIlu
DZ0GF+PtA7necNpVQNM8rpN/z8xmDCIkS2iKiX0c8fpFMiDE3gL1ejocE4NRiXEwDzrcCSiLKrf8
caxYSUPLdPD3K2rvJomLRKbVxDKtsdb2OxJeDQGtK1jzMP1ObYuZ5AP4la0+PsoC0PxGbQZXlmWp
GR5Y/RD2hs6VEunNhNiZVmc5H5sFMXUoYIDDsUpdDTmIrJvu4k1HLFCPK8RrEVwjL3AqTuD+pstb
YqB9Q48gi6/apfT9PLukdT2BvSQG3b2TWcHVk9J7aW8eR5grEGcdDNIcfrJomUrBZmoxhHpCQG4L
b4aSd9PWMTJAOWXziYEKccRjylsdO3rxp5bIUreOhtQqXg3SenwtMJ0wA9oieq9EVvTRFTo6imB0
RT1Tq+iQi4vHT0obLe8v58jTpswXtO63frmb5nLB1YtdMY0RRjpbDsIxovZWkU0FpjDAulGVEsZ3
t26i98/cPSXavNBpcydapz4XD+o4we8Zgz6prIxjYhBdLagcoDWRWyqxrRPZcsmAd5Jpj/gv2y0c
owUW6zqVf9J8kzTllYiPnLowTl+tRYsgTbG1tZWF7fnbyeUBZES97Cd+R6PQai23f+lkXHCoFzVe
9ygYQhUP5HDWZ88sQpBCwWR07lOP/BEYawHdRhZQUinBBY0cqe1Z8VCl78tr54L6MYWOoVIfJ/Zk
r52Zui6OZNVzbaTPWYSbc0OzNqp4AypAZSbiyaU22Hz99uUvyn5M34pYyeu/TEqKDzBTkoPHQtBh
vyd0nv3anBzqF5Z4wpQcZ7afRSeC8d0iXxCwz3GxTh86sf3b9k5ZlOKJEZKBQzeWYm2hPnfw2EH1
pwN253BLtcyIqUz1NlqF2UcxLEWciisdyp89Tzp6jGwaaLMVV0FXt90pwhirHl6sMDdUoUGCeoQv
hgqNlEscnoFmVxyMxU0V09w9TBoTIXRAGZcfRyCmuShocnRYvv+bz1Z0wTdtA5safjSQdP20yMic
Bpox7nDTGGqG12jNz7lUZ3qR+xhn2JpsG0g9aqJsZkcWZIpui81PYM/lTKzGHUvi09kNC4Dlsjuh
o9yNvWBqjqa2EV8ZojnN9V2lYcP5neahUKb3uRFHr7LZXZHl0S9bLfkbxzYaEBRFUqL2MV3M965J
UbeSmoOZ89LbI45owfa8QAFsqO2TGgwKJ355RqCJKlIy+z9ANCRXRvIRBtoDsE04f+aSNs6abj2i
aDhN69LQw1tknvPxugKNVXduRdqAy1EaCiaLEDUztrGuH2M6Kx61NGcbBJgeYHcoz5XW1KwVcxqu
rkzPoCdt04ZjyJH3vCm9ISQFCSiS8nW41IQ/pfoV6uTneIT83zLtuDWWlHZoL1P3tLQa5J5yHIPs
vw7L/5LUrxtadlVGL+6e8ozahDYxz4Ls/AD4llPN76XlUk4BMN4kPkETRt7owt+aXZ8ksOLh4b77
f1GxNuAW+gFLphqU9f9eQPYhqYjBJRK+qqYjq/NnW+L6bDsx0vdfCQ4nI/5E5MEC4aMAjbzUyRyC
jFDgo1vfgni6Gjr4c9PsiB9GsUZ0PUs9Vpu7L2heLVTwbg5oJvvSYNwqLz+pQfgHQRYXz5JKceVx
/aePQ5ywuP7buqetxn25o6+IFkZB0oWV7JM4IrmSQYGJ8DuqJiiAuYy3ojsXfHPXnTOKkZhWi4eU
vT+la+yybi1hNi2KtUtHck2Nyd4R5hBcka1mHLUoDDNVyR97hSnTXFnA4LHwIMMuKJhGfDQ+eN5h
22gaCrJmULmEngekblMSyHbmJaC5KKzOmFqbKCe/ThCUvb2WxKGwxcDHPPxxTkOvcyoYsJ+ig1y2
AigC6FDjcSqkZCLAirkni60cqEwxv34khbjv2z4IrFjoY8KFn73bHH/2aOW7s8LaIuQ6d6atan36
cFp8DHsrnPrzbfnIa0a1BTOOCofO5f9PUvXDC8w6WShOWMDuXyc+IIC2QYzY/uW+G9lEnYa8Fehd
EOM/LMtx7Fg8oin2Yt22dZ6nMYqcjHz2bJGAukQ1wMpXpz0Rg/4TIkh9WQlfaV3eXrYrYqfbXn6C
hNYUAywlQ+XEWGUPLBjTM9tb1JfIWZtWSAd3P59NGZicZCQfs6L20Jas9qvBzMP16XY3v1j+UtbP
N23sHRob5LHcbrS/WtgUyoHkzG+EYdU/u9niTUf/3/TqzGHkogpsvN+/zfvRBDC4ZNyTKgc+5QR6
mvWA5z48f57gewKfuy0i+/koVhtCuE5HMF3re51MtXoUaPsLqZUHyErFuRUJCZVB2SPQc+YfGvjo
V4tpZTkCbv/6LyXeNpHtrE295T+l/iIzkjQYAo4bQ1/aYPf9ofee5Vr8v8S8p/fNauPj3NmApAVF
wA7YnktNIVY0NaFfZDz46JA104TfsNxo/pQyVmlpKH72Ir30mNfxm7AYWsW9qdQoiMyvHImcG7XC
UljuDbdjhNfMwgZWxJ5tLYTaSzNzP/sPRzT+2OkpL21JYgOdaQ6Ae6bl+y84pYPkDLcpIGp59fHO
maO/Sh+R5u0NCRJvgcecIzh5MDdCe9kbNhKZvLrEcimH+5hkLIShQQ5WR5ZRlm/ZcwmMj2VOhD7f
KElSp/kmWsgeDZBN+8ohiLh2IJ3IhXbgM0pfWAIEvdUP2L/Hsyjs4wG+dCHgAH0fT+/H+JAJ/lgY
BxEQW30wB+vxelB3trw0VZzdYT31Qiy999LqN5SWiXb41Ib4dHyMoRDIQDbir+3xEMaCF8OugjDQ
TLRKb6t/gfgh3+FbkEAqCsaLEISF5Q9BHx01NmOxaLO6qeGAAXHIqfcf4Pr4S+a3omT/ZrNa06wD
Yc3FSbHU4HyfPBAzYOmOTH/Mu7vGCQdGuaUokq0tE5DEdctxg5V5BU4QXLm4ylPT+pBoxgFYHRs+
ed2Z6o9bsnPFaZUWhK/1ud0cXB/L0LdkFoCsnW/wRplGLvsScArEsbie4lNX8GbOzYSR6gHr4Bqw
2Rtx+24Auh5rJM/vtLKjgnz0MyjxByzt5GAbsqvQzZWMsDLQaqRhF0LC2cEpDCFvLvISi/fMC0b8
EVRWBE73EtpSy4O/xHeKVJpcEnqvtRPnywTUxOI/ufEQRn0senKgSdvrgd9qn5gvXxP+G10LqHOL
aBsQC/dG8KCa7Y2HDWkl8yGQTK9g024k1lpjPlmtAB00DJtA05Wn0FqZ57AELf8afbkcqNPnXwMY
w+bo4GgerJKxyNlayw8bQRnaIQPzs1bDn9+35pmP4PEYUgqOOuSmBWk0ctkWAUbYUy0adrrkEm6e
5VephPYKelxbOGDWiToe9VeJqIdG1VbuUz7n1JkUeu9LI17/9mE/FsTArowgNFLjFPF/tNG+Ps4V
iyfdFNCfTcvyR/RslUCL0z4JGygN+AgcKHsOqUJak3YPO5zGkUqqKW5SNxxOX5DNWN2Hz+az0CSO
GbXVEGF/Fqet+j3QBSs3ty89LfvSBtBu65yi0UJC6gygtepOhbk8yovoGfrOmp9F68R8V2KEsthx
ZktdVUYaxZpe2+4cv3Ncm6xDgZvuBnYAJObES4YrY++uhIMyV1rlkc0184JZgD3cwdvE9OF9igAt
xWohZfMdrGHPMdgmDKN/EkHubUFHwz8b8KIqlBmibbg4m0SeTwpcBjyQijXA1epjaDfi2IB1h4kq
d2Q3jsKy2RTJMo7tsPgbn8HXs3t81url6GXe8WHbnNO9Vzw+2CZDMjC9c8HvsmzhJPRCuVo8gwbc
S+SauMlT9IEj9zUj78i5mzFolup9keEM2d8WJIxdz71QBBxkLaYlC/FkdnftBLmM74JIGo8BWUOe
U7Jz0xFbhP1183mQZHKLXBl+CWIKJINt/SF0f5ZVhPIud+aDhW2diHrP7Y/Rli3CvAOBid3e85em
9Jb6uMsIbm7c+8ZjQVAEsksuKi65+vvOF6RNUeNB4Cakw13tpepBxrm/OuBkypi0Snuu5bqwL/k2
BUZCV6lEut58f83IU67xlDfSe7vHe7XYRRNTvg+oRkEIpXWspIZR4TKT7q5FnjgGKi/g2rtZ0ttc
xr+gnJv/OnO/cklFwBtenwt6z8Q+nXEWiCUdP1STlETt/eAhKX6PYj76R2UcKzhgM9jCLDPH84M7
7idIMot802Amxd1guSXMIuH0yxRAXvxog4j0q19p+ftpX947tO4ZH7xPjUmoFQG2NVAeE01tla7M
LI7p4nSCMpgpm0Xg36NK66OO6WnKIfs89hJJCfWWz29zJsIbune4ULTLQT5IQt+l9OfnMQKdivvr
KARgj6rGNAlRSA6d5gZzh2XqZT42H1aotNiZkL+eRofYOBXXe5/kOMh50HeBurIBUjIgfiOqQIU3
jx/z6o72AKL9GKwffuOfa9MXwHdoXeAZ7k+opzvZE4AGp4c+pN9lFab6vAWNnuinTOvHG+1bgIls
oRDyYY7+M01YKOjvOPRMDpq2evmFTCHLALSrZlKkTZcCXUtcQvEp3aS4nH9J8zFgycgZZIw+gTJQ
IwdxemlV7RN/LSZfLSq25uNBSR5vGjGgcgUfzrDFb8JuQ5VyHRJobV/xDOri2hrW0XHJ/bzPhR6j
Vi8EuXuXqClkqzzJbB0eD1jjZelkVfBx/OTePZWcU8wt9M+DdEckA1Bc5WuiikVWs16iNXAE8zWt
Wx9XdnXbw4neub7A9wWFkFpaSdtT8iw1GB8Ew4KRlR80ozxFf1hj7iS652U3RXVhyJ9c9U5zKNqC
tw2lmXbokcZA22gW/M6nyl+g8qjNVEPeM6i+ESfRIEW9qL7tZU/Q3TDqIw3M2zHKeFUExDGAI6gX
K51g6w3ZbXoLHaeTcWPe3b4Ncavt4Vsr5ozu583mYmTE3Jybh+ldCX4B1AFqccUVtAOKFN9DFgko
HzZCgXzjjVSKTO2uO+LZKeKH5DSiJxfBcfjmbFv2/lvBJmDXSgSS2wKXfzhFVWLTF1tp89UifOlY
I3+o3xsRC4JqhwywjASpDL4bjVwDNaeV3vRizJi758omMsaMSPCXCIkLIo4ic507LbVrv1qRMIeo
AA05WxymjsnliuJ0B4mWQOWtcvskQ1crhvJshtEkMNB6oAy5kzC8Sb1UxQ6vZ8kW+xBYRJ9HZDfw
UyRzN8ZlzPFF3MIfVTTzhFSpxcOxn1l60YgmYNXBxBSOSJaqSjOtor9ffMZHvOhgEYS5mWZcIiUd
tZPjIiG/VbcjYHeAtE1dKKKo7W75u0g4bvGh59FS9Ho43w1O+j1raf4X/wsh14GYXSYjr8239Zl4
7FM3K1KsOMBQSf8VIwzfxyQZhTKeusv5MYIXi5gctmg9MNpy4I3Oczh6yjJ7cUR0Xeoby1uB6uPe
/ukeb50dYMr8BtU3eAP7JnrywVxGLEzJNmo4BL++HtnhYygP95SiV8hTbe3mSbG7fFgNQFYSbSst
Hgf6RgcXA/y3NA3PNybEzjNW6oOXae+QnVdd807gEeu4WO4zsXYxjglvRDZjVMZScve+LK2TAPET
QAINTCWd/51FPycMFkKb/JhvZIx2AXge4/RE4zTpA9eF38YPm60vGbqjxZ5jEfxJY/KE06sfd4Rq
4bAPSuVTyFTigjACtxvVdUfAFiHveL4ss4m3iS0on8Q5cc+D84Q3KQP8qsBaB8W780W5mDUABnsS
lVHuynvGGOHsr/IN5SsRk8ippO6RuS991C743XlbW+6Jl6XWl7hJLo7iV8/dSoGCcIG8kfi58rvY
M6N6hvOMmYljYAIBgiwVKef6YpX/EaV1eiLAs3sS53muyMJdpKE/w0YK0wn4+JCAf9lD1CVa0qZ/
7GlbVetC9tn59/1dR6JCXsxDt9rlqUtkazSk8K9/p22+zellJC6ZHc24x3T3UKTzl9cenWgfhCKo
XP8eg15xprJC1EpHhz+StmeELVSlEVzXndvhKzMko65da/ltfZBbOm6DV6SKX9BXdW3pakzlgVFS
7+Vs1BJbaIo+8nhraKVpa+60xCu5pTnoxKaXN6o42PJZlRWwx2EsoayIcibHKeCjRHLB0tKR84rA
f3vrMBmbC2vEO0pNw3ZJ4u3UoSJV0FuD7S3hBrzG0OmD1kNG90L+msPJAjWO2sIyHvcMoh+MYxcw
8TZHVz3W2qYbFcq/ZgR+icJAHlNmeHMy07D0qz2++UmW1Oc65yN+T7awchMN8kJH2MidS1TjFgiU
IpaS8QVgWkc0KGLyMMH2v0++SMGJbLUxiTlQb0/LKAaMTgGalEhEFz+vIM1iA7iriKzb+pmVfL1I
X0oBsFJv10Nsx9dEFTIdPn2YLwnNDDgLBOEeps4A3GaEyFlqMvff2JHYlTYLqju4N4AJQgFQKLHv
ThVIJzFzlgv/YYoNqpehLdeRhSh/HfYIKz104UneD5LQH+nGkbpauFqev1/D2QcB6OvXb6IR+4I6
2h++x3aFGdKsadEshEMynqV8eyT4tDXM888Z+e9axvrMy+r0mNHnjR9cGnPhMfxZet2yreywd5z3
Uc/1kJ2gPHR5Z5bOQ/OZ8pvKTpnUIqMHQfA8pNs4rJDBbVc4wSWoZsLor/u1I6p/ZWS+4Z0tsSal
hp7XsGDNsTkVkpTs4bzTSewqtRN46yoKw1iFhhNZkS+x4pSRSOMzSQEa/xdpbG1KpKrskROmlPD3
/tJpBugu4gb/rmF+uFhf60w0bqn5dU9+feccjVxHBslxjDA/u+LOL2y4OSMzs+Rs+QmoYH5L0Pf9
YugYUwW9ujc4+S2Xsu3T5MtVfAJkZXKQ7c6X8FYv/Pw4CKii4CltCUv1LE+DWl60r2h05yHLxDo5
XBfe7nfWqDHkgcOc479HYi+/A7Cpuf5Z9OBFAtsRu6AgPZTYSfHtZn3FQ22vEXkvIAe2sts2zTpe
ytbltr5XPJknV6SzS1AO1j89IjUPl11SnTWpOOmhWjgT7V0p6RnAdIoZI+/DqrZhlqk3Ba69Hf5/
UqnYqOtaq4bjqO4e1B3Tw0ba7xXScJUInsFkIIEmEcm6CXmnIEC8oiBeXf9Xd3algMwPlyQd6Y1g
N5nqpT/FtYQLYk/huednBQHs/dwZdefXUlxb5DVkknQWuB9xE4tuEJAvPqHwQACo8GILKckYm0aV
8ZUl09KsXe0p04jcB09T0toSaoeF4or7fUCQnPGq1s5sWsgqncJ4BiJIG4fF53XR4nJIHzQXaz+n
2izY6QxQJi36q33mehclwq8TODw52ff6CAv1TLt3a721jx2D75f7DFTjSQ3cGQh+BOWZr8zIxcYS
XkNI6Cg7tvM8eCNXCQT1KSR8JRf063ULw3nNjnePZBFBRTIbM0F/grt0gYNNXidHC8KiuKp1YsCF
jCpl65S13RLETNchems8pIw3C6fPLqCa0AWB4//SiSyu3mox8wqq8rIDV6pv5O2OJ4VG43No77Ff
xktzuhBwoF4WDaQSNPVHI/ede/vgaXPJmPQyy0HgEXBgkG/9uFS/l9TKISyj37sT1WIfi29YgOfE
osZtMBWcixBrXBSaN1+JstZ48wXJbnEGOj3RRzyRjnrIV1OZhFcO2WpeyD0HYcg3/oaNMhP43ORf
WlC2hzYBgxk2X7XCThKrrYpH55jef/cyxP/9LNLHPsjcxJ1Ug+UE0JBJ0zJlDH6y3xDe8mUwRnkX
mRZlBO0ghn9xDNfuEdQPwG6pt35f4b9dnS9Jc1R5tMZcVto77Of73AZ07yk7pHODDNU6FQssa/iP
tJQ0KbK+Ts2GUngwI/nOsfMpIiCcy7oP9cfedjKESZI4iee6VmeLO3uktXOOI+elNXbMpxEiovA8
oQa3F0+PkoTvKtwAiXK1w99xM2Eu8BftJrqpKvox6GRawexRteim15P87sDo5ukWCHmjRQpOOBMT
d0MlKj1T3n1YJpqR4TD5nd7NlVI+/pErThyPX1pKjK4MwTbBjD8MBDGst0I3/LGi9dDIj2PqPoCp
KAFD1b+zeTevGEK4MyNYB2/JoblRCg3SukBj+zlckBzIpXrkqCnyCsg/ot7boT3wNCy41QfRx9SD
h+oQab22Npmq4qOJAe/iuOMHZ26wb1i/9EFSZ5TmxoEPoQO5D50whdKaq5aXQS1+dJhZ4zZPqAFU
3iYcomH58pbv77d/pi20qYG5xua8VOWWH0helWqUc2YrRqD0WDeiQEerYQYHw24HWCDE0ANkIo4o
rUBz5xFxYBy5DJr3jgBB0MEger5AmPUSnX5nzWsoYARUsUV0DS41ED2xHSkM8o2fJJJWw+j6pHhn
UK4LeHNANj7kYv+TijuqodbUw2ad5HivjqiUwuQ486mzNHqBTwUfEwjqeGNgC8VEGkeO/YlyMf5P
whRulW1JCQRUrpH6jufYnflOkuKa22nBQ9PH+flY/sOpzNzv6KQzzK5kcSQ6q+AJk1/9Fsrk1xXu
EjyBMLKJCeYeMarTGLpos4qu6CqYWQL8qh8khN9ZBEgGB2w73SQ8fb3d5DnwZpe7bIpui9IuNYnK
Yy7kyy9xy72OhV7GEeylLRp+qM3STCK+mTQdlpNvfS01FF1VZzJSWrEOhsL+v7n5YwWgZN4cwTQP
+epEyEHBvdtnVwFzIoCQWNR14cx6bdYHLcHxhzJp85TS37fVEE1wl/jU85GKlcJY1Vm2yhXrfA/0
LHx/lWBLCzlTjXGkEfi4q9sqks9Ttxfy992dhCkwxzZKsITyHyyb9iuSQ9Le3Yv0HvPYEnm7Cn55
t1Gnjz25+d6Nz01zaUpYz9JcmAg+NrBOiyVjjB7btuB4+m/DD7MxJwrYx6IrX2NGt0oEhkjmmED/
N7AoXNEltBqZxrSg7QukjPnZ7Kg61e+d9YWUTqWMrsPAGIkrYMLZPcgwmZ0SP1k3utKUqp9Cw6W8
lwjddLUpLjRokFoq4kOcKc6ZBO6VPTgVr5ZfnsTIo8V7+IqIIFmLVV18o3i/r/BVu9CgzE7ETc9A
skW1J+OdMChRqm2yFYjzhPrmdai1Ctkc04YJP81pu7PBAJKQ59cZOfS7Sr1fJwbPbppiw/K00/dg
xH1CkFQPELFUdc/MWJuHDf4CxXKa+gOCRhoy14HRmPCsCDFB9SURa7V/huMEqNuNuxnVoKbN877+
cwLUwBE05/qJgzs/tQgfrqgPMmq2n8cgN/DNXohU8M0cgmh7QeDLEBVepM9AY/YWtePBwDSdTh+9
8HYi9IhbRXDGR5SDeesQCFCCr4B7ONqkB4DqI4rv536J9Tkjxpv5ck6zgZ4+zxyN4cHJCfpPe533
Iws069SJue+fMQD7Ui9tuIqS4wZI4irX/kvZfUyVQSbcJtGhiCWFPdKRWKa+HLLrXYk4/KO/0vw2
C5O8EAW2J9ruj6O7ji0vVNUu+ju7KLdn+d/2mnpods/1aH30UsNA+TyTfXs/YWRlkDTo519My5FN
70pkegMNIDhoRr/la1JSU3rHdrIfCcSyX7WU9YaH153Brd7zuZeBCCL8+ZEET3aiZO63ji2wLkjf
tgQZIUMyeN1nyvecqS1CnG97YACI6UymEVCbRmXRC5SLD9cn9GWF3fMSPBJ0wnGSInBYY9Xhcr1Q
NSBoG4XU5ZV7wTRvWyTR6YCL+/edp7VU3zo8rPdC7xjVvwCZUQMfuH0rWSvjuehvKL9LUFQoMhny
A9WAX6PlKon4IKqU8MqUmZoerIpYuEUWJj408ERXVN0DGMd6yFZ8GSevYypadPdo7smI6281OCqQ
QaTjXEd3OyC1KgWdr8ssxhO6dxgJPalOonTandde4E6Umm5ZqO8wXWYR5S8mKh145FpG3bT7Cb41
6rPVAMLJLZ1KcElNRih7gX24C7DBmAIpto/YcPAlBecMOJY1Fkr9y8CAgGDO60LD3tPU/W120+t3
3IUH/0ggSw8ObvEOi136cXba9S1OFxXeiiX3EgiyEL+kNotBufIewBrwU38Bbql0FpDuIioX/gDF
3cA+9+tNGdb478CTYG3MYCzUaIwnbfQd1m0GrC2jIHLGyC/lB/JtbanciMUlolzTGs3BWpKqQQP0
x6LLE95F224Y1xS4VtHFdmGGdBJT10GpUo4zp9KTEu01GfjAa3n3s7dJTzhyNji5O2Pa8ianotEc
ZDO3lMGfwq5HtBtZyhzNlQqVRhzHGn9U+d7b5T2V36cigatGaN7yXGV3X3B+E8yMs0C4htma6irU
vY0y6LFbLF/OtGqcrQN16LVVftiB62zJ9XDJDMlxnmYuEFb1d5qiSG6DMCmvqzqTAiqmuWlUO8nQ
8AM79HwADNZOsfQe4maRAxZcQ+cdB9rX1qpztxBpb4L4m4dpDnbdifuo/SNChKjg1nd4ee7zw8S/
bKNcKejRKGvWVKVeBxt0mliYbuusXZ7kuH/Iq8kUEjO9Tl2MPFOrNZZUKgq23rKm0yaVZ4kGSc8h
YmJ30LLtCesggTvNPDEcOgfHm7HfxbhY44dGu6AvVwwKjExlinbe0Ho0lKRypItmbaQnsrWAWmr+
XcPCw4N06wf8/oNCFVT4HzTuMQN8CVCdRnD/zX003AFg/T4fe1jdMJLDqB2ZqULLzxYxJfgXQFpM
n6inUPDWnp16MgR2hPZji6T+OOduZd6Z/avaS71Q1a3mjw2awFWGPi6xIjeuwbCOEpHF37hLwrPN
deSRdEsGkp4Vaopj/QlYecAG2xeagXrviNHiJog6JXm2O8x1w91gGsxkTkiXZQp8QolPHX/jDIFA
KzriDUbgQcm2eZdguVUEax5fqLhbz4FUDplgJg3gBUaDkKaHNJxzrLA4ry1+EsVmOW+ZC7r/M748
8eFXay2cwBz8WbSDtHTunBB0EgD32XjhAUeQ1kHkNaW5TUPc/7vYPA9clxLnMd0qBBazTmGGlaPp
ESVz+65hoYc1Q8KGK9prkPNX2IOYLvo7JFS91F+hNW2WsaDbIRddyi0z/sQihIPBTFk3QPJEe9x2
nV/xd6jxqpTDQK8OP+745pJjqR9Z/HDwzMMXAu/eRACBgslKDapucwJWyfWoAwTFpX9lbN/u6Ixa
ObBpOanJd9ffKfpRW/9EaU+9tVVMAyO4x0qcYe1JTpYhDHXQeFOiDaCBCOLEvGQOw9OMJgYcW+dp
DlwJilL87SwLiy9++ucRer80CoRzxLYSYWmbeHnV/X3puZdWXfqMgXlxSXxVQcoNCZqRqCNb+0X5
Yh/UhEeqsJJ5zZ8NxUqQeq5QAbJkWbKNh3peUcE4s/dC+Ko7WfPgwke9MNlA1EbGEwOUzrvTAh4Z
E7kXHMWpW38ZuECae4xtK8m+LAEWUOBBsLTcja/2nwBpF572r8VzXhRYQMiJtaCdMotliEDaqpy9
KziD/+coTglJIFYwSaN0XtGDhz3+5oYK+iwUM5r3Z/aC+hgp5KDCMB6zk23Qxz9fmOlvBCBGNp17
Jf7IVjSTgpMsXmj2zUDmoYjt3QF2f7VK9cQt6lBQ3kMWiSMYVbeMxLNjNa3cDTkAhmxyKhaJj3wl
vhWc4Xsdz93cjkxowf4kjxemw70U7J0DAlxIZHCYsJSKVg5gHeSprO47zJ1Q6kwX5HPQgxHC/5DX
lDD1jTGi3zx0kulmY+KEApribze7JjtYwvo3u+CNk1uDz95CtQy8RUaIacIv44Ym4RpMmWWepYUn
rewaI1SIP0/ySfliEQ69JA6kpC6MaZQgdfxQRfj7uxgdKN32WeAlosttJPD3K9VFXRs+d2VY+ufK
zQ4+T8DlL0g+HkNSl/NTtVXtPCUt7o2qzXNu5VkSl94WLIYY/SgReXNROaNElegYcv2SNwCuJTQr
o5zh1b6wozNkBs5PcJuNzsgprtMlu/dINgaAlXsTvdhjTsHGY0IWPcsgNaJUcyct6CAxFxOuSpOQ
cPHdSSsIqMsxzYjNI7u4p4OjUrGaeMSmtmpEgA2zfTfRQqWWqoj3ZpLAMO/SOBY7CSd0gDCxRNS+
9uX38bfOBiKGTl39HWUfiuGSsUTqHMvGtzBTjqlk00L64RXDIeuKw3EUEJbjB0EWWi4Vtx3ZUJuV
jefZikIY78HKWW1bYkG7+pgr/OJexZbHOYP4KFIf/CQ6d6V9qCiSqpZ6xlatBnAqWEM0d+GdsXi9
1DFTkrfvvuISkDkTUIKnapwxIXCy5zO+Wok9yI1xR82y3pmiHMTEgszhbIZvJw8SJJplhDOEpeyJ
fuCxtz1vgi8MSEws3/tjPXx57c5yACYslemimShYdaSo0pOkcludjTzT5rhjdXH0SvpBzl0eKdMw
IbRjpY4sJoqNzm86y+M3IQ5GoYAc7N5UoDK7ZIO7YQlNF4YYfGH+y4VI2Sk3h3doS/8w30U6DcRp
355MyA0cnxdiq40fpT3gJBDJRcQ8SHWI9Pgz9iwa/QzvMHC3FlyWhLBE9PQQavSv/z94b5iIWZWv
1eX2LBA6fHfQpHt/NqJVjedI75ykhniNc/0Mw7OIrFdme8df+alyi00yRN9/4Rp/YVJHSCAmiMKd
R2LLuBhGzlAq5EKVu9SY/JdBj8ypUvt4kRQuWIwsY58MFjcIBczlFDk0X+DUv4CftRmc2GjcijYr
DCIi0CdKGNA60BFOnJe8oPhPuP+zVN+BESmQM8qmHoNFeJIf6Xgu2ksexEPVb+SlXsLwoCunY5EQ
4P4zy+243BQ2KgHTEfUGgQBszLg1Uj/FedSooBnOau9ioX3AboXkjq9Fg9Wv0JWmOtkalzRO+Hiv
Ewz06E1wuZJ7fASVAHUj8334bvvHXr8MdPTGlmAorGWLGKo5gygEvm62Fb+CHu85okLA+VYZ4c6K
iiAKFIXcZ++YGDK5C+Ct3u+RlvT2ToHwG0cdB77hg2Kd67unfTKbQL5Xi9TrW/7vJ76iXeI5oxsz
cF6v5UCmBtnSvRvO4Z9qo4K5D3XKqexMgPXXNajryp6buAxqzQefIOqBVoRR5aowvxPdjmuuWtm2
lrY+ty5FaAUaHGSJJGBS4SJYx3drEwBlRMBTnt4y5ImrjQBfWBRhnXa/UM8vy4ng8Tv/12BENM0i
yleJPe3NeCT2vCeP8L+GyH4vLdhAfgKGaXGAWOwfvHyf4FF+2K++kA5KxwvTUPDqA2+w8gROwQud
aQzqX8BEDDBfIQs/RFT50PBMH3WNyguENhJ2+y18uO7yWIhMtpPy7LA5y4eTTEprfKjct4Xgs56o
RiWRpq2dDC1rFd+7o/hufr2GTfRNDHndBbyxHTYLVb6IZH89oU0Au25idznYHupORZXXupotawLa
GnSLGSHFs1AyJ/SNQSzekkv2Er/beajqxMvDHIPVmhQOSbkndTcruas4TvHqyPiAXOQiNM7AYKNz
4X2Q0aIp37UqjJvlE3fkEdULJ45fm9wbaV7KJG2KhsG04mTveMvm1We6aeEXjrDPOmv7LhWDr8oi
D5Ey/6VP+fxkvFEXVw7GL3BvgbrV9EBVzwfkbDTQJ0glVSqnmvzb/17K2ch+2KYcvrGaokU87q4/
AhtvMY7x0UUOU+r75I8f1MsN4gyfrRU3DewTsA8UQ0Z6xG2WqHihJGu94vAq8r2AivNq1ZQNZIrh
6qNLJABljiN6UHI63RNsGu6ECAAKAml1d6UXOxyC6Sz27yMFkOS1L1G671iVD97ZjuErHe0Q2Bm2
830WpjSLETPPRZY5mJyw2FFxw+K81uBe191ATuVScTkTPEK7AjN5IWDyETN2F1gcG4xdD3k9rFA7
JjYQdGv+NYGJVTRjWl0eHzTvMLS7OLGSyKTRj/bC+r+puPUWydcsZuOGfCcKvB0HcKfO2nVZivgb
HaZGf09zNqcYtls3lMcJH9cqE+0dDMv8IxEHKjh/SVXeIG68pj35ivjjSPtqSX1cF0tCp70ql0N6
XeUu3KdbV3tOijfhZ/NdEqEcM1cUHpgBHSMR0wE76PmH8BkZSRZsvoG9/GKD9WZ7lOG4Dk1yMAZr
yWrAJIo13rw4ZwGBuWVJjw1faqqKZI5d1rVn26NzC/AHhqIdyqGeHlQHOhNjiT3+M5/fUS2WYw54
o3Rm0YA9w82wHrXQFdJ4ANSr5QvZ/sAW5sxfGK+PN8+xyKMLODlKW5BbXT7XwLPRlA/b38UwowI1
4QkdOP9/cdgi2mWwuyIra4U3++0290pETJmTcNMPIMZNgbwDHy42IpeFy+ZcFlV6REB6frV5hCxW
eM2k5HWlk4knt7BRv14zKhWiNr8bvHBOm9Q/H/xqyyF22Gw6iZGLlVyDRV4x75AWo89NaBQV9/OA
YyEBsZZuCW4a1vymoM81iXKlpjydL9kqFTqtZvDYcL6wK6Kk7wtBp8rXqd4UWtt83dLDuqPdHy4Y
W9rFlMULyDtJ0poEk/u5IZj4laklDGJG+kJ9LI+FqG3t8709uSz0lcjOmcB8ewaPgyOvpeJJyCcw
20Y3+dZ0UcyjMgoJITLp430EJQvPfY3Hprg89LNZbd1mizN61LCH3ay/FCESZ0ZlElgeZjNYKXsi
P3kxpfdmvXxTfEV5lR04Q2Ye7fyj+8oOgtLfa0SFmrEnmNUHdaewn2TabdKzqnw667eDp/51MCvE
MM0WMhPpfUI38PI7+lQ6+GYsIZb9rg7nVrT/L12LJ5AcyLG7gpbSTf4Dl7wXsuypCSZdwIZ7X5zp
vBIRKSoX8S/zZeB0GnpqDhIyHntiLR0i8QffKNWqdFJIZA/HPW+t44jJ8dXEDX7/uEVGHK0b4d5S
KYtvgcHdtFNMDwS7W3XfSrFGCnrPB9VTKpmuwOSdbZouHornjHaRvFrH6jAFFok5PrrMYrXboaFb
zJERpaCBSO1wWA3uRu6j8LTY7HNZDArH1LCCkm/BiGlp9pw1GyrOBlK/bxDUFEd4ZVyXPLziMYLA
GY5Yegn1iBemYQT9xsjitrzi77sy2ASFV0EO4toZKaWpDEuUUCjLFWrFcDrKKnF9RFcsQqenO4hE
GWxA/0Hbw7Gn676kgBCxB+xh3iaLYj/gVAWPapvAU+4xqM91xkP91NGciBeavs4jw18ijs23Rdc4
sNKcarOMlpYqRR3PdFQjqfbc6PXZ/tOSczKjMsKwxCiLaatuKLYYqyREbLhe146BBXePuUh/MVGA
a47eINghp4CgDqESWVFFTWb1Ep2QfybdGfjBBpcVgnDoPNOWPcfITAoPuIqvfZvLxg8Dj+3WQL3k
eIeQPqTvhawuO+dSudAZf6U7D6HfQvqW9WqGUIPv0lSckxT+Zbt2oj8Qcn+5smB+qUftiiCgQOVH
72M3ixI+bmrxPbLpmuytcu6NFD7Vsm4O5PSYOWr/sB9SeOBOlKQjDDvzjEkO2CR92L7DhJbD5F3r
JPhUozjzLg1mQvpPpu/2hrWG0iidjdOHy/+9YkhntwpyTxCTs0f7nu9Mhy4KxLztXtOm6tvp+yDQ
o0dZPM/TCH2n56NQFlyh1sjPiSRdDv8pATBXNfC3x5ihc3dCPChFnmNLcz+q39jmwMtX1XfFkP/L
hzBQWkfXancZrfUlkEKHnZnbzgLK4lebKzi5L+hObKBQ4gGnyTKkgdW/5uyYCAC4palhEA/f2nqd
gUH+O67K8zL2tMNgULkvc8v6OcdAnnhdoBP4jrPDxrZxIS6HPmQM4KdTjC0Sjk/Bi5jTapF5fv0Z
glWItInqZ3JbDoRXkCOhk0LktGsIUMIQOidaEGnqbWAjp1fKU5zt6IhWkFRi4QFly8cihgngYCWm
VfcjBuyp9aMOSifnA5nwkA5lZKwKmVloNPNKqj1lFKYPPMSMSkqEpqeTPc5itRKE0Cz0GbzlRV+r
r9iZltzKABKjWbpxNOIP7DNaM4kVHyamEzRB9Xofw6L2W78pUUTc5nXMgSvFfrtt5t+g1BJgCaLW
AZjLgw6WT2fwizlpgM3C3bBQcCyqi9Ob9AAYNlQT7V/U0o+NsdDsGCp5YBJOr4ds7zYOLJ6aIViZ
OaGro4dHbHZx6WIg7J7YRuu72z50Sox9fgeNgBIEeCxbTWdkIs12idWQ9npU8sBjLN+jZPrPkppm
eGExCKWNsvtNKyMjqR2GvAG4pE2k0nZyiKCApJUMMuxd3x4pX//4Xelh+rfcJdn/9YSJXKOZ6t4J
FXmCBSPLnleSLoEom5l4lkAvLgZT5GqfmGMG93+EuIuvRyjoBRuy9wW088DBil/j/madJwDu7Qx+
S1b4fXOTGZKxlCbpnsca4S+1mYXuRpBc2IbtBuLLA5nEyeSTj8MsBuaoCLxknVa/TX7jVyoG+HmL
39rp0d7EjvDcQHLDNcwGrGblYsMYRfauZJ56YbX66MdAU0yl5Bozact5Z6Pr8i7jJv8g+mXQJkfF
JBJ3htv4nlDMGJCJQieuIy5/EwVCuaIkNERVLgYNftlhg4Z9GEKaz+aGnTjysMxNAJ4d6CNTDA0F
FzJj0ptfydB82kgJMsmobsMY6l+Kp2EVsWCKV7NuAXn+2TLt7MIwXKT6IipXGbpgKiWO1YhBDYRs
6NAJA+InJrRJNNVVON8o9ic1oK+4Lrb9+t23XUjK8TXTocMT7Hcn/KB8RX5cjFGm6JQDu9v4vC/s
7gaD60/R/7nklo5SYvMtvzxsCq24uz5dCTD0eJw40HgX4wZ9hd1vR0VPRiHmolxwbCZPk9Zv0b9h
5GMR7kt2QeSl+BEDflYLgreVWH2bCPk0H3VywS/MhTBMF3mtAsvgqdGaOpTs7QSmGQB2tW4VfI9j
IZcnd/PXmvefKWzXosGTlJ1JqvHR+9rLo2cCXF1GF1KXbx4DX4DGQHPyo9KlzL0KYUh97zkw72Rn
Nbzn3PCF4+7T+q6SkhgiV8wNA8nfo7aSTXOU641FWGaQhYVp9buyCN1g+oSjnjFE4He6MctFbxCw
8gp39I3raVNGNSi+WMtIOEjO76x5cq820vsywFiQuV2mtEhH9otga7E5vIOq+qoZjgucqxRUIqxw
dOPDTJAiqtlkkaaxo8UgashThVv8yyllR3pJjVsb+iEHll5f3CRJ65k6buNtnmnVlaMcYb5UxNRS
OhgEdEsuxpDpI32/0Pdy0NzLboqNg05I3NCwP8Go3uLOQREwfr7xGJ2OpK+pn0BJHjiR4Qp0z9lJ
WPHJI4WdohvOiNl9U7kEjKAsZSQ1NoWsjgqBnCCyqSv8jg0mXVaCXTzTvFpDHOnin0RSpxBpdLSk
cjaxcFRKysbT5eKu0/Z3Pd8A8a3dhmFQSmDP7Q37Ny1+ujPV9QTVBwzvQ3zC11Oct9Fe2vRzdQ40
rG50zylnL/iJO36arMNitgDtprnRWps3TdoQd7JiO3P/3893Uf4HlwKtroWqFRaSp7st50/vYk7t
Qxekr2Hy5lwqU54D141Dnw/ulN8JOKnBQJPuDAJ5IhlVr6eP9QcBO4JE3CcADujzVZwPqYGVQyKq
e3+moauf0fV0sNcWuMVO2kqps7MnqjAEBg9Ou0j2IKEX3baeeQIYup/JVqS95/J/RjaChWc9yiN0
Ya+1uYg+E9egA4ABps6YxaEbSc3NN5IWNnI0bxCd2ktaq/VOnoHLfQjtuszFmSbtDU11qx7/v0Re
7YphOtUdbtlbawjFaU96nKBhtXs+P88uklSwScTOywRaEUqHGoostD3tMKu6Sr6lxaHDyKpGNU/G
WPX+++Jv0UjjuMlB3G7dzMjPFV09o/j6KUUsK08TyTmbeaM2OtjAoz+mXM279YhH3q342Nm7WvYQ
yvxDWYRMw36WkzJkCzsSJ61fjr+avacK+qifwJLUPr7z75/2O2977/bwYkyuwFe0GTtGO6DnurCB
y3OF8//8LB6AQ/6O6b4WFuod80iU5XpWJ3YGPK+qObaVJhqyQFL5jGonJFn/7+32VFFjI2xy4vVF
e8jCuY2XOR4yGov7snN5PPpf99qaSrtKuxWs8djvItxv811MQKFu80d7dc7TxF+DhHejw8P4FQRQ
kHvYvRFx3bQr21d6lEb5j3pPA1cJ4EgLt37BQu278Mk/gowd78uKuijAv8bFgX1ITeIaMFOlc4bF
zX9Us5dKVQvqHYCPhAouXdXOzmPLiNnS2ern7PhBosqc2T1w9u4uwEiCJjQFMyjbIKGY60WDyXaV
BFPAB4wZg3rQg7UGyCO7e9d0sEKk0FvmgZdB5sHSTxKGHIgSXTU08OCxTWVRnLSk70+lu7xXdHD1
+rHLvBpH/2xUjiPEmORg5WqkZfjMaMICKooJQWlGmpWUk6/Me9ehQySFqOlc9wFXSzxTIbtMhn32
5ujPz3fPoj2sepVDPEZLGmySOK+ugKoEStoyNpVCflgZEWfV15RDLKyhJ9CbmEM3DFJEvwwCnKmP
/THUqz8CfArPXyTEgS4/bRvc8KS4rDBp3h7Wo66vOH6J2n5Bsg9Q7VFHNBrDMsYbW7K1sQ8Or0fE
6re2RFjNuu6Rtpu/GJlUJHM+bufjwW2oQpl6ozeSp5bao3KXb5ZpvK3y7gAexUUn4mw894zqjKlT
+D63saDaCPRhK6qtoRlwrnTM7q0TUmGVIXQ1QeIpE2Iq8lFchR+7eqvNO0ZPtCxJ5ZxQu/lbSU3d
z+Z9xfPFoF8RQ3Qb5KhYdJLqA2feTlouE/UNIDAAJeSkLDp7QJQ7LfyUnczNiGbhmq2sW9VDKRx6
3Du+xjHkmFFLdcYK4IFwf7uM8I4GHmJzn36ZLmqlZfx41Kd+cvUvyGUP1YlJP9dfD3V7So4jWNaW
0Hl0ag8GrC4kFVj0lCE8mWBk2sWPrzVp6l/EFXFK3dzLCX57/6a9Q6Xi9gBFqgfd2of1VYYrw83P
1jTN/xqarO3brT2BOOA7bg5C9WlRcg71fkB/sYTUBYMorMc6O+Ux2ypzUQM4VOUZv1NMwFWBwann
whZ9m40h0cyJT6x95sSfy2cJBYz6Jfl70OsgF5GlgXAd6aDZYgn4Hw0AaEKB906AzA6aE2n6TqTl
ihTqrhrdigODunTJcAS80fWag5inDcz1rJpByPFq/T5uoUwReu+J6Cy1x2GHmq6IYjVbAAtfy879
JTczEj8nXYFh71zBGFdwHeA74+1nsx3/4KM5dJNr6KuRmmcyx0yOZSB+YI5zcrj7fZEq6jEm6Aud
3GZPmFLIAHks03AiUmF+PkzoszfLWFEooBXCb4/8TZe0JLNCXE59D6xwaCQEh1UTZAIRd4znDpBX
8qY0csYKzvXjipbr66xFek5/5mkfD6Pr83apQwRZGPCudG5APg7S1HCbYGqG5G6244fYhCU686gP
kB9LIpxSVj1aEZVMRXi2QV/57xxKETUoRBlCOqYaEfrW12UBePbgfK8CxWvWjGSpUGMo660QpGYm
YIVVnYn44VUAWM0NLRvn8tdOcbFpS0bHHfU5OdEj8vBDfPYY6bOAGYU5dfznu+7g9q/kUoK88dLf
C/+AJHMUcHGYCrZBvkTrRmk+cguhK/t7OVTmrlNjZDynnt5xumD286gzLvaVRfRNwIQ7Sy62NhGc
0uYKoV9PMqeftkaldZyA8nHZsByoFOZNF3VAss7uLqaRkqOAXA2x8dQieh+eVBBSAnYkhLg3aMg6
pN11ulAlIyu7PzaJePEkXVMBM7cUhZCd1j/h0Bz2DhMzyDtzpbgT5lSn+sQPpHVuQEPweApQ/O6M
xYpLcye+0J9Wnv+h4MW4BSB5PSArssWpJFbNZoK3y7kDnQ1ojfdX25TevjpRux1y+2dKyTGOYg4e
YWyGPQSPrI4N9Raf6Q5sviFCwbz7lmwhjEwmNlV9NkVAtyKLiquxtxmPQRUjSm5TUeX0BUcw0nd0
YHvGq/Gh0XgCKEvaFf9CyfeZkWxLJFCo7x0A6gN4gt+F9bsAySZ9vT95xCj9V3m61TFhA7LbxpHK
jrFZ2B7OywwgqoOHLWtj5Oq3FfVoB//Ea1EF0GXtxisigHr1FC2ejPsIssVygohHY2FFhVgV3DFK
z23N6Mzk5ljbcIi+rEj2JuitOn8szlw8AhjXMz0jarDrHa+rcuIl0tXdqaGHvGDnpGmm4gpryxYP
39MEz63vdIr+T3KX/GXQ+1FrqTZEOtKMrFO0yrS/015agOJihu25myII6tbqkZL2aX9kiAHN9MrO
f6oWEYjdQmVBG9iU719s5dMS5umQx7gxyURlPg71otnBbQFHwFsFrfsRDSch/XJAQPkXhLfqi8+S
F5W5jHyOLZpuaFCmDpybyI1+9HrEB0YZ6wvhz1CkAbsDVeZe3Erc5H7tgdfnuhSV6t/Z2Xxroqx1
qi+VzpS9IcqSx+UUMIC2Ml3KCy5R01Px4BrcDhHzceJL5e15b/meGObQ0gnA6yr1UJ+5u43cMHrq
jdW4b74mVQLZXa8rPJEnv9SNijeUS1PAPDnum6f9rmwiahPsBfsQgfwiKGln79LjgvXebjaNCFxS
P89dS/S+469rp6uN5oo3njMaID8KbFyguRty6FKTR9lp3O1GSgNoBDWGhT6TgfTeelV5b97uGpYz
AZ60QPh+FpX3xZlKGnyYUViYFse3D/YsTzk2nnKK4JYycjgEYjsyz+JxrG+u7Rwr6pDppMGbzEQO
gNcM+kBlGcHJuTSzzUQcNB3QYF4uVgHexhnKWxQAg6nR/4sBOqSTiwtlrKJpshHxZ1qPACcvU09L
6lP06OQ4je0c/fVcfA5gmxR4KKpvOZ1O0FxcsM7j8KFe6DYWD60L8n/0BPTZwJcyCy6Ge2HPUqhF
Ep8MSBFpSozcAcrVkbXLFkOpQYh/VVBrGG127IrmEJzDYwtnDCeCBPauFSS5IJbbPO+y2u2B5AJZ
V5FmnEk+BZkdH2NTLwmP5ZL4k7L6ASPKkKCZKJaK/35TYkaUzpQ6b17b/88nmOXCunB7ZodGCLcp
v9RbwoZcDwQYsutpqxlhwR1gVYzPFzGvlzUtydJLypw4/Gzha/BrFzvY01/z1Kgb8d6nY1TxWCMO
Ovj+d5UUJN/x2ZdS0a/tLh8XgsssNiSPZY3wxZabhMMR+yn72d+cl75myXt/kZTi6YE9L62IwieJ
pelXaGoYsmRGiVQfMQV1d5yhIV2mOSRbiRtMV1Q3Vq2uyZ0++irMzuU2aY8sToi1dN3VFpWozZGy
rOhVZh+vyCDXPVLyKH0Xw7QgGdbtN6T0ZNpJ/Hd/ScRQCGM4vegwrXKym6QWT+C1Syw45OHATNMX
KWT+3zljiHDBspfUzMLMOB7Xebrp/xXp4/+VLk44Z6ozYeuxo7ESLXVyXNPwSNiGlo/lD6KOpaJc
Fo+pcLQkdR/UQd9uOGRnR2uf+FzZxU1D+xZH2Xp4mu3IY/yZ6QwD65Hyo3J76iDDcBF0EcaTGqZ1
6YyQEiIUgYFshR7zvYPFJ0MJrGQFwJo9hRbAMZucE1AYROP47uEX5CF5ycMZgL9HemTCsdaKeWkY
xZD+V+H1IeK8QGMsskBAYMyQ1U92hqxQQ4rv2xu+dK65ggJ190rum7WFrIM4xysA3A+5mYF0J1PQ
mEgNDA8NCT0HHRVame24ckM2RlfpREmTUr+HILdPO3PWI1LVkxH5ewZVPrkrwcyjwVe6TKYTcJl4
l+iSI6smOPdifcET7MJLgtEIPzF4vw0yrQruT1G/wBjeyXlCxD/APVRieJwFVp0aPMS34H/q8kSZ
vzY6trpPM9UpzZ1gBr5umQ7ZeECM25IkLF9O91vdl9sl8HmObNDJE2RZ+eL2Ocss/rWhTGZmyS9n
noBX4fZ05PkJYMZkgA9Z17h0+Ljxfuje0zU0uAeKmQmqBopwea3/uKRlN8Lfj8h7g9y9KYM7U9XT
Mq6Ftp4Pb7n8ahZ6W4XnAROryqQIFokvrvuaQXWRwY4FbJMcOd/n+JHNgcOeM3ERYD1Shm5N5did
Or0lblG6Nq2bOEN5Lv5RREmg4Vt4JLkeU7thTrSeSyUnuAxVRvE5BUkXJmAaE+oH1zrfYYj8SKM4
0o2NATzOCwIM9CYN9jy7xd8eqvWeKrn6rB29C7ds135wFVWkn6cvEbv5vGbGAqTWYCfNiOgqNSzO
DQl7jiL4k9poh+ZYZj+rSGld/51FPY92yEzCU2I/Wz0pxFAPy7iK2M1AYsnxGNNt6NXzppOUON3+
Mem08nEhgmDK8rLwfzj8aQX8ulAJdQmvamNzQdvOB+C/xpvH1ESCFyC+gHiwQGNYAflCYueIBoIi
Js+QbTQ8gh+nsZ/1YG7OHoT9C36xqeaCMeGMFTknzDBVYWLAH9rx12NM3g9+Ean3KAParkMrB8R7
pGFUwpavWRzTQelgm4J9SFLhcaPSFbevNhiaKiyhhcGqj7jQLIcqAjU4X9xJiNhH4BLMvJjnjDjo
A5guUefpKj3DUQW16hRctHEqlZyOnbHO7ciz8nm6t0398L+BxOeOm61ww04YPsM2boaQkgpqHLxo
FlDxJbbCEEVF50+mrrHAhHX4Vd4lDhHRBFFM9a6rTCibS1TmLs7rkvSI+WEGl+PdWFqlfrp2Vw4N
n+tm2Z/LA+t0tKONFpQUlDhW1ELnZHpsXRtTz23mn1Q5p3YJxGzdbESPLoSqAo1UWnc2Qc67anQD
OV+kVHKk0c/1T+XWpVc0IlO7kh6vAMwHNSBcAWZLJ0P4D5cT5FT14fkw0yXJO6C1CV+bY9+Ht7Cc
9Ki5MI/Z3i+Vcg4346OiJZHQq7DkajY5qX4qY4IvkGURNgY1vVEfgdoTEHpciAwr7rtj9RwFKnEW
Y1IOkTt7RqAVViljaaml+o9kmCcdMRejtMmziLTUfM/zvV7m39FKFDNPIOHpNE88H8HiHkhJLPIv
cuKKal21JGTxlqSEJknhX0BYdU1bL646kXn6OFvzBSLozJ8p9tNH0LLSXYYmCC/YNXCPlGtlMl9y
HnliWT9vTpSVlfKH7eIaWDf4iB5SEUVyGmyR7MraJNHvUvUERNlG+tAJO6fPVqN2OwUWDYhNzE5c
4mz6fN/HezvtJgfeRTeChX2zP173KZ1NQExgQIjmZyz4SJ07qt+Zf9LLZM57skXcaDpDw7JVE+cN
M+3MPA4s1r1QZvP7+3+Ct/xfvteLR1Lx+sRftrbcPYP6CsxbuvPpAxj5OejyzedLbKpSx0RaYY8H
AkfqlE/Z2qcAmVFk/g5sAYKuG+MtIFVNRqOS6AKVhAjvgLvNw1bU43iEUdTSWI9YKrOkorjKmoty
WonQnmnqhWDsug1Uhg2wTKLz1lpJhihy4s122pwS6aL2wvEt+F7XK1FnU3x++LCXlYmyNgs1RZvC
zgTTapvX7h9UajhKnDLCIfFQy0rrr+CBLRXza06mKBsrX8FGhYtlm0VABNTqHc8QbxNIUGfIMfrj
BVE3jWckAilxEx0qReRLZ5XjO40BcEh5ktiZxd1TehwcYuRHryqUZ/tuoaiLSFZhUAkkhQhngC0F
k5CxsYNWZkk3K2x1FI+mYDs7+EBPG2btvw86+C0wWq454FfJoRUtULR3Z3CtRc05M4d9c9x4YbN4
+7S6agr1kscNhoo2D5Cghie7r6VCk5gOqSZlYrR0my9ixnOZre1kUhNCbZJmfuEtKOL1iS1fHhxL
Pd0j3EIfJ4s+HXAvfFl9AjjgCHi9pbxASxayptDzVqSQ//vz6y93oUwIbbU2GtEJm9i549sShpjY
OP+iDFu5j+gs9WnFP3dfFK4gARXHq72eEMejLbe6Qg651SpNn8eAmWn5RYXr38lysaEJthEtm/ic
tBkev8fiUmFf//UdwFC4i0yaQKMkM00Z23HzyjiJK1zKY6ciUDdAg1ioZm73r84eC4mCXxpUUyCm
Rg7Kd/Xt8L7V3FM39mtaT96nEDNE4kAq3NCGX79TAGNDLZWIYbzGB0dljmq7fCLjMo2C6roTk6ls
Ma/L/3LgggEDBi7r3DYeujsRPreVdDyTGD3lpHO4s+P+tWekVkVC7SQcYvHaa57p2aj7KUYE3oZU
kmH4nyXj3s4WbGpVGGO4o6aVMa2lBU4og5gsTKkFEmdcRGeQgOzezdRpkt3TsLsD3HqlSniEcfOp
8hVk+jFY1NQTGG3caMygM1qcKJIBtgoErxXM9ZNUn5+O8mVuQP+T0XqKj3gM2Fv+rvmpcqkLUy5b
jYI2tUGbYK4BfWqZbNxyQYOInKPxOqbyxf8OePqYlPC7QKqN/T6KVuWkKinV7nXOBN1gB5PnZeYd
69oJnT7I3U1ZrPiRFhXOWR6GjvY0dqgHvoR/r5Q5hGOUyGNMR3xyL0oLK7PqjrT2slLEdgYIOAYt
w+Jq5n0rusMC41UJxtMXdiWLFQzO2FBxvymBYkj9XEkLX/wRVtgh4AhwRAS0Y90Jdr405c1aOUHW
6oVhXSDLhxqFsMNAL8FddMOsIBQbd0a+MqLeZ7k2oHo35A5iESUdNTdmWwXN6HuToHdYeAo9EoGL
Cw9AzDycXZPU1a6pw4Cr9pCsJJ4rMdiJhWuU9XfVcbwlT7hpn3YkO7tvEuFxQtn26QXMGSPcue9p
xqg8Ztg4TVlfZieXM2yP1HbZteIRJwE2QEPJHtnZiHHPZ3/0u79TNOLytesFwOiqFgIGM23BqUON
5iacFe8Ett2PsxnsocTdbWnIq1PQ/eC1hkKP3KGzYagzXBC9tDpQB3xwYxBmuzmlF2+v1rZDRPlD
F7exPKqiSoFBLohqchYQ/xG7+mPs9AemRmups1gi5X5pVEOo5ZmdROWwxMfVKfbZhLYv2Ib7vT7f
oI0kP5QeFNvK5634IlrRHY504R+XAZigLbwuk1CabhMiXrz1LjgtO/oVyKSbTLpn+imGA1lh8Akc
ogtGca44CFtdmhrpjpvz6GkUcMGdNFPHjrS/50CFkgEr8Wlrj6vBdKCW4m518EDDgM8WFmdZILV/
G2Tqdt4skgTgcjRBBcntig8ZchxC7JUrb7RXuvmkAJQ0th/etXoeuHqI2cLFcAx6BPh5zX5vOWJ8
ltXZdisy2s5cW5na/QvfH0X1JAFu9eOJql5Qd9INdVHlbVlrY2WWartHKNeNhqcz6eVZjxPBbUqt
Gar4oaQoLlS581W0xIBIuOQDi1x3G1ahawMlsmHonoRfHDv7P6e4E5nRj5Gcmes5K3KHh1+qTktR
iMMcpCwM42o9wCd/nD1rON4b0tWp9m/d6nhHEvml06hL+JHb4u2BTOYdERigoFkqaWY3mfA1eelH
MpzsKbKMl2CWcPyQWeHLraa/62kO1D8PNOceC5Y2zskAH1btievprsp2KwE6xpy7ykNbrS5poOm5
rRvg5uB6NthGkKZMkgDPvfmbu2bJIXiyg6QXFL84hSOmPdEGhiLS/Yb6TeQVjzDA81t8AenkvJZE
NPKBPlTboijFOJ8FxdjG23kPVXqDvC9Hm9SL2ZR/OputaTEd2o86uEcMWra0Tr87+K0ireW6j4n6
bN3iWfDNGk8CA+slntG6ALIcEjqBOHoXDbJ0ZUj4ZJj47v58fP7zEDZhIk6qtFLdQ23KBxPXj50M
oaeeq9ZyHwgzz4wfN0fRN2VbmVwXJmlPamb1ReVn3HRlN98PDLyP9sMRmraDMSjjaWf4J/vJ5tKD
mfVvSnRfldA5yvjDKrjK5g/HHC69yTkD6priiHRTtHi8BJgyJVX2JwI94Eux67mGfCb0L0+ZFZ01
d6v4xJf9M0RlGr9ZHKxuyl/GiLpX5pepTn+ee6sNhHRQADhMdwzwJ2CAxgup991ONJGmXuZSCbaQ
F4f14u+g3xOiyH0CtcWHz4cFhd/pB7wrCrFLx8USPsv3Ug2PUMf1iqQpaqbpW9YzaGAHD+j+6YYK
pdE6JvPA9TidrGpxUnJf/devA4qUIbGdV5qnTzTe589FU7h4hFKEmHO4KSpDkGMVUvvTi1x08WGi
gnsoczmAnp++bN3RdsiPsJ6fsfe8BkjiKYqn3QRd4+5Rt9O0CwS2XANqPDI2OU1BbhryJP/yzSRE
gXhbGMIFDLH5Ks1gV8RgK1IMeO2gpBoDTLvSm75jP9pH90Omnqs1eG9bSBgoi48q7Rffx3JEnbAi
QnQrP0QMBm28nn2UWycswbEwiuuRn6beKmQmYfa9KT8A/egja4xLR1mT2s4PZ1E9uZN8w2T/9pfR
dHNb7QZayFxXnuuyy+fnIuT7BhO7nQGEiE39K8SHWXm0bVnmRl28eRSHPGY8onNUG9xMm6sSXsW1
YsraOv82x9EOdRBLdKQLQgEADj2DnJMmWvuhaMP9eCZTUKNv3SVDER/zwnBadJxRbVFTSYcn23On
LvFY3TU3Xn6l4nT04P7Q0WmYf3dltdnLMG0LzNgAhEtGitSBLTJlna6lPoE9xe4JfAp8LkSpXvNp
GGdyMAvINpj9BKlHD7yYyui3rYi8rE9Yc/tEVymh46+KFUN6H7GbzwUl9oLZCo0LjQAvoRK9EYjL
AyxUZFpb1SpbNW7YZSmfLmBPHVitEW4d8FACF4y+mrCmYlfmllERYSBVlKzgh4b1e9vfEa+pb0S1
NNxfgskc4Ryacs6BZf9M3TVRq0lIqtFIrcb0t7b+A1vhH659jA1S/tEt1DWojjvABr5UHyyZg1ry
zSZbex9pinxx5qH8vAHoKha/bKxO46YCRJeZkoqud+cP5lCsW+CZoUiKdQSZBhFIhHUkGp/hqlDJ
bgi34WUA82wvcHlM9U+ngjd+iezW8ozBB/yb0SuXVo33E+rp1RHs7f+wmgzAuJ8vExKs52oH84tI
3MkcXF38DCH09VZsaLt3pT9dOKT/WOFLzp12xaey2+r5ptyifPZgDuy+NBonsvmxu5bW54Uzg0Fd
SCDFG2FVsT7+kAXlgnvWFSvvZrtYZlphCc9MWOlnghX/p2KJgzVo78KcTqDNbk/upiyOYFeDnr6O
QIfyY58eeWFqbXSgFej6WwGX9KBACmUAXDYAqqG0mJxLhIWw4ykRKIfqJfjqsSyAlaY/TkmGhvN8
N1Xbsh+fMuj28ckDfwL3hCbAMcVM6YsJ/cHe8mA9wJVOac3T0XArR7BxUQjRPXLpYoW0edjlDxYz
HcVcsBxD2I0RfpWrpy/rHz/SibvwKDOcBgjNXBsz7FQWkDe9cc+DefBQaIsQzENv66gyGMP2rupO
mc7XoNWOT1iAveEQJzD2wH2Ffq+i0mwF8Ez3rt8FZ+O52Q6wDkNBlQN25I059zhCCNAipghsy6jB
2M7+E4hhTw2ptY3u+l/AyJXLNUU9LauzYXwciUFvFXNaM0Yy0xpDcjm7SSj3JGYI/70+6rL9zJqC
5pLVRqOHm8P5s1NGnvJQRIkkAV+V0xSYIBZTdWoimExj1jkkeNL9MjXmW31XyQPRxExd38VarUqI
CIJc8tHfXDxTqTuzsgLJU5weVLy2poJzFs6GRAvoAjHubfy27l4yEbBOo3GzCIDRwW9M+9ckkiWQ
h8ywZJeZVUEMDTT5/PxIrY1TvehWT/W75R0Yowyvkl/nBLcPxDlwLUBSevkIktPsSroXITvL00me
2roipsssxJYMJwdeX7BpBDgUxAuIyH09id8O/qUIarLqqXw9CiJBTtxFH3aD6b4sJelhluSz9QWJ
wdSHIdn001VEBmGwszU95mZk7dPS6SYDxsUSPpZlFJ8lBfU2dELg6rF/7tKtztfl5A3RzdDCE/cZ
z0hokFjGg2eHfSIySOkc4d2Jw0Ax5V0f5yyBoefyj5UGd6yaBePvPz2O37kuahowZd/nrg39vyJ/
IryeUerIYr151NRr7RH+deIpPvJUweQU4d0iFDGjdv+0YwboL12eeX0E/yO5bmRvZBdC8DPr40Lv
k+jquwLUo4EmxNEgRI16rcVnzJZ6DjQ5/v9NLtpOee93nQoX79X0QSdYV++AELMiQbIC5U+iGqvb
2mXy1DEy9l/rR+0BWJ23DkQjqbXAGbOfHzG9zWm/RRKQ1swfZMBdGtXrNzIvx2lVoN5Cow+jWDf3
lDzHdlagd/8KgW0IBC/cYC1MtAJR/B3fdmyOBa00URMF+jBot1qCsGhOWPQlYY9zgmdgZnvJk3gQ
Lhclo/Rv6gF2xG93tnOxd04Tls6psa9myUouGrle6+uwB/YCVOxexIaIQpiCcD8h+Jdt210Awgqo
FSGOcTLW+JnF8ekbCnwH3NGqUGamJ8nKx0utAE5Oo6sUCa2+pwaDUcgMr2UHfTIJlojD5RBjECfd
rOZqiKceq9y/cgpgWUYUCBeNDqlDUCD7F0ceK4vTUvUo90Sa9lXkbe1wTE+M2VPkuvjKI0bQRQrj
JiMUvU8kxRCdiIoGwCZcPXFajy+WonN8YK1yl3pZhpcF0FT1wVXj+h7Ae8twS/0eUQSR1etSNqie
r8CB4/fNgsbttsP8OT/GaHartTc3AFB1DMyDzfPOKcSruatLTKSwhq1nD2dxzbwMmrJSYT32j+AG
/ScZYxEm2S9Nqi9CBVHHgXpbg89gNgbHScS15V0gMd8UFbtEUOk7yJ/Vi55hlVaqECgZWk1gUdPI
7qrkldhSctm0Wtp2U2UtCLnrIxj4lHDhJs6TZQ9jyji0lvkeE3gOJqFczXCYquPkggE4KW6K9dtW
oObXA5d5mMGHtjvW6oNVg2RT0Rb6UuoeMkpZstMXyzLJfMTzdCFbEnmTsTCwYXKuQUvpkz1FdzR8
wcz6ZUErYsgR9Xs1O8mgwAT3vcV9C/AxmcnBBr/BLIWgxKZlgt+35+Qo0T8CQ9x7HTxfoDtd6LwY
CyKEa+ne/04zWHIyBKIGsKg8336Us7oUzMbpWiT7+4anHBm1r30xki5It0R2yXjJ9cg4sVTKDgxC
p3GoceFRbmAR9/5UaKBaeZQ7wAi4qQvzaMt4v/+J1MIjcShyjJEshEk5V3CvT1PQrPCE3lMe/pIb
HzVgOymfsqgRDj/Cstf/UwOhsVYc4PjcboHYtZNb87ZVtyaooW4BEolR5W9t6lqOAwHi2DGr0OBV
5D/FtRWRlTfvxz5kPzCZQ2bk+/2x0J6oUItp0ZyGHcdufYug53J/hrTW1C+nncIjQsNvGP8vWI5L
FSORZezjDW4tbyowLp697PK/BjGaTKuBbV7aYtZ3PJx0wc1+355Oq3cHfSILasCAh/yT3OvsojsV
tKMFM8BlCYHMKCEL8HOLvfZVaAkDKn2xFwmnh/ALLstbBIpiVGYhJ3GAEkTdqrbjJppq9X5VEtwQ
1opavYKWOQxUUo3D8hESzcjiezjiZjNuI8pJw2qEqgg4DzqylQEm1IK/KyQFQ/GWrr+UQMxwRWUo
DHwMPeNRmLcOBD0BpxzT856oMqq24SxCC9J/7HEtPA7s/hrXkaaYvTVGuPTimrb79bgYaBmozPQ6
/qRZrRl7ULtbUmD+xDo6wXomp2+Tuhb2IUy8mjOEfx59P8jnybAx8S7az9TSaCxiqirvB+CV6f/R
pzWGYeNTm6suBj0OjlIBfXLW2/qm1cbmtEifp7tB4D46bHPVjq8WkfW44mZqk1bDJ1dOEP0JczQc
Kib4uBLd9c5XpzELN1JSe3TVxjHiESPDmUOqnJowNC7vi0r6xMUzeU8ZMyv+mA6/MvKuBSiaMOdA
0tl37XegIRF7fWmvgD3AocbXGXbHKJcYt9gtkOhtF+ITwv5UDu82DdVQzSiz8/jXVOc6LFG4ydMf
nq1++QdZJOvBmEsyFEYWRSB16wpTARqK1z22JARCkrYIG2eenHVivENqpuLfZ8j2ZfQYARGwxgxk
GCsQMlOaN4Uzc1qK8PEuy5PdfmMsj/YxXtTuqPZ9EJSxzkaKsUPX9wEmpBfNkJbIxnAjxPR02Ad1
7xh8LyJvWTFUQAKt3HwopSJhLwYKg1Mvb/Xn5Shyb+Hs7mDEqzb4zHxTKAAOcYK5G//JoB7Kt4gC
nWJXeqysvJKKy8Uad7wiDKlUMYVPfjtPsugl9Idj9CTZD+7FRS7VE+GOzBWIhXce+a+NjpcssBa7
8StHM7pcJqKuM+gx8c/GAihr1rv6MfvCrMzVaR6MoDdvYXXRo/EIj0axpy8vKQLI5WJBhi1+1vU1
B4OGp5hV8SmqFFG1e6YcPwE0ZH4ts7lBjlsdQ4OSWXokEkpTf+3wLs+AIQ2fReisph5n5d3wy4LD
GOOlcBZFj8M2rYz/DeGCH+pWwcxKrXp2x28OJtBDS3VN1z0SLwXXp8imT+c27Si+VzDaLjCggOtQ
zmDxoUjn10WcLj+QF3tzX+tgdn7bXoG7/N2IXzeFkrY43taON2vcHOpTgtWrh/RkHX8JhRZh0Ms7
xvFJQhgaCCZ0STa2n0H9l/G/t09brF4Rnr8cPJ9r4fzL1xN8nDf2eY0imRih8YZntqjVB/jbYoqM
uhwvMeiXCqM1JuxKinOD+MBaQTIQ4CQYK5bQ3OKS5R2pYJ/9exy1nivGQdPeCEdCiRDmCYU2/64u
5G3fBMFGqVPE6Aj7itOKVo0XafX4zu1eWaudu8PpELBuP+tjD7fAkg5zp4o6M4Ls2PfziAgXBpCY
QJuiaDbW26TM/BY475IK1Rktrf3+LvS4Fy9Mt4wkQPBzPf0arxWpY6FpRJMBSV8rg0OeZpWPW0WS
jByvdwbbv+z0iqBGO+ar/OcJxDEM0FhKJZhLIM/bwxLvpdDr4EYjUj/VCfb0tlLR5zFG4Ut9xCGz
oGgKZsE5MVj9js3x15YWLwti7qJeNf7qr7y5kFtgjAAr5wPx+4969bFGYrkDdDT1EnjkkkCXvO7k
VXaXpmr48xhfxQr+P1TMwJQ/RrPYXj/2tkvHmHkJDZiw/4Q6Q4PtdjgU49NXesuZgv1Krz3Y/guB
vnwDuO+9wdEO9Vl6cjSazJnoPARX0wcov0hdgwgLKj2ZbemThrLhFgXbVFzKhYq59evCGvzoWppf
kFV4su1T2uxSeCg+5OfgD7Pj7Sn72ZHZ6PUM373IsxIAgm1Ld3V081WiYke/aX1zmSYZuZwsI6Mx
4N4GefpFm/9RbIw/IhyiRRZkXww9VhMuqPPzwc6mQ/xuXtqPIV3xjBII7lvqXNo64bxtfjr180W2
yb38jXQlZmjZQVBkyGXb1MMFT68fXZp07hEDLD80RfK8p5oxGKCctCB2nP906EgG9+VxxNMTFi/4
23BLjLL7MtSkXn0kQZTQcG0pNTJ2VxbA8wIS+wNXWm85GcEEIfCyGTG6ZJAL9BqKX61sl0jMzvTc
AAfj22tPGBlKqtMQ7lrV9E5FUQgc0drfdoKQvVs2Lg1ZZdF6RNbTLmbCkMBodTeBM+fuqYInz4uD
eKHWNB+moJnPEofyvtp0aAuWmyNDUz9MS5AXTq9C0LJ2sEGejCNUUprR71pFjxfMCmpO957nUqQ7
juxf2lLt5G/GC/bpsvFUTTgJtuTHrTp9hG+NzuCwhzfnIk50vqTz/443z9lqXvIGj+a92bPN119D
LAIKpdY/b/E9JLAmQzHq4zmL5Vt5Sh7i8vnbU2Wywpo4YoA/tjmebQDOEggvR/f6vro2u3zzr64o
hj7s3bQMsuTJj83i+kLX2kb+u1oCKzdXGLCcQy5kKv4dPF+TzDmsfyG4y/PxXlBddbC/CfLhWlJm
NUv+giGd40eLzXQNnRdsz3ewElQYBuzIZppOZbwtXXWzCYiDhCIlCyRMvVZe5yIEatiyOSWcjjbb
lPJFhEm9wg12WvFOt2ii1ZYIfUMWm7nCArlNyG0VzyhdSNJdxrI94WuuVp9FGSniHewpwcMfBd5q
wgEyJkXZ/m9efLAzTeSpWqhoT1UQLuvHGfIBNgVvFWRyaV+uEpX5B4CrhIpa4sy9Egwmg3vq6Kju
gGYetFKsKKvCpjJvp+H8PgIx4Q5YKZ3fVXKwDF5HOnXhsW5jZHQYwHmN2oEi5Bryl8egoEonY3eS
77odayUMP2OnKBvzSRVRst6SWcBDRJfGxRVlY97l0fz5mot6kU5YvEbSnmLocWtTHuVDFjh6/U0I
feCZerP2CZ/puWGWVQ1xDiOX1AS4tNAx20DdZ6+yAoihShtdBC30W9Sna8fpZAcAlzlLmFJFCOVO
JCkMlFlbNWVscECwNdE0Ed+Cy4i6JB+O0BY14P3FptaB4eIvJJdy3MIPdeu9XdvVG3TTTMDn/ZkT
PedEJN6Qjy6r8aKxEAZub+xr8p4YqwVl/NGjzC6M/Qk3QghybmtqvuU/jVn9WwuTd6cy9gjiq98f
Rs5U3Pf6LAjlImUsscGpBtdL6X8pOOqonsIANOhTegp/ZWt+A5IGYp7+TJrYDFdZmausium4qhyn
mIENBFMDqO0hbBKcFH6eBCacVVgyfwE5uZI0qdwPcqTh4nKZXlv53DpKPh/YWEfeV/nXDrwPkfRB
WAlubmC29QaFb2+h4orG2h3PKsyzdfcBPXLUx4ZBc4WqWa7iuWWnjr8dTiph9Dtqb0VCYSeA9ZO7
i894mBZQJJMdvAwv8WW3Zh4y4R/TbowQ6XwKtytJZZt3bRdR5iomAxORbQxaKYhQk0jMMbk4GBkk
xp+vsO74XE4sUY2kNSi8g19T5kZgXSei5d50IG2i8VtrNpXbRbEVcm0s1ZYIKddoMXn4kjdvBroj
tzMMCFko81tHAKXXeJe9UZJQ5bHX8pUNWy9HsTCPAf1ojD7CJ55OEVlkAiKKni1rk3WAoT6fIVWr
z9hwYPc1OHeOOejGO/o1xysymPZrMZMGd3jzeE/tiAZxswjMvwXuH8a8AwKG/gZbsvVzOgEyFyje
BoLUjhR6L8oZwScioFv3gar4kygyVpxoZKVDukXkxyLGW3fRa08mj07iFFvSxyBsPkR89uQq6jZP
nYoWrVT0Uxn+PlabhHddhJGjkU2HqyfxObWKyA3TtUViZB8aMKukNxB59lFj7WMmX63xpTAnL2y3
yboaDHvyGxRHmMnl0bpyXFvqop1g+pv4s/nKuGyiyouxozMTzl/AZoCNGzgbUiOU4y663iaCr1ys
qTY/tfkPpr8c5M24bKxCJUZgoX/pELJFZwLi1d5bXgAPFxQrG7XfAUy0/MyPcEwShsPUU/v902zL
QZmbjV5Yzsbiw4Y+HlgFNDFjS3YPreGkDF6WfaIhXTijaH1SngcgbQa/UhA+8mrETYqWX/2/8DIo
uTKGEYbxw8UrPbhGdB8/IqCeD2zvQLZGn33lZWT0juaWoYLilI59Wb+SkOPKAJsyU0cPIvoOQK31
5VuccdE4BatTzb1JgkA7bbz/HiQfBFqCqzqRlH5DeM6TaZmabXb01ndsLNcBdGsytYYcySGEeTNc
7rtd93zt3KAqpDtFy0CwB0AVWKMh4dsoJz7EMvGJLKYK8LoD4AYVo76yNfQssC4Xj+AohxkmikKG
wHpPxAj+XrzWzny/qtROgXcoejIG4XbXevkient5YPnXkSkPTfUXR+bszubZMr1IJpA+w3KYTjhb
lxuCWuyQsZosw+CfDhQboWIGObc/J00zuEz+gNWno46ZAJqtDAOiZYgb7j1RxWWEzHutxDajAMKF
FCfnH9BuDM3xdFaNcHO3OuqPVlyaxlFpRauHQkvULnG2BxrJEhBOjPw7rc0RRUR9uunrPfKTb9Lw
3eQ8DbUwqPrzGlD3axtLxOOisjMCCKHtuM4OZxYUd15k5x3M6n9Lq/lwylaiJlFiECMKombdrNMB
N9xMidBcjAOJSrpyOdG2QAxFoeSTq3AHpmqiSD2P79eRyU/j9MsmiS6hzxfu9MmIQsqOryCf09Tc
IM04TKjHkUq0Xr3bTvomd75UB1KotHzCGIRa24Zh9aSUqNDN1fcsxFTkl65T9nxTP1bzkcHUYUOp
3GAU1ZT3MGYwtZTc3blxzNGWlCAp/r2Nq2GiKOtIXEi9yAyYZ9YKc8qm/3nW3vnx3kyuUscN0AkF
Tjee0S0XFu+gk2CLBgRJDTX+bULH6jUEDm+IJNdIkTbnTcrL4lGg0nOPi+rKGYXdQ3E2iZNWS9l2
+2wUJCg+DVfysiyM8m1vHrOWZJ4VKp/wvKWYMNmXIwe/KBomssqma99n56RvlbrKb6NW2MFXhD2O
gF+adoFxaX67BCnq0LbXmrZT/t6udvzMxSnOsNai0iaCocr53U/myfUM4pvFkEr1XhelXn/2yN7i
oIgtC0NsnwmxXgkoOqmpLy4/BkAXWlb+eJ6uPY3wqbYJhYmy2FzG0BIYjtfuXKyz5y42RXk6KjfO
708bqGbNtVhaMBr56qeTlI8O1zC1jpLH5y7LN9PH3xlJam7uV57eREv5vO3bFQ/Glk+HB38rZ5RR
N0cF1gMusyqihmTfTGWgQgEtjTB4FN6GrPrhTeBJFAuVtOkaqxDlQt18vUlTd8CO+WcK0ONec2/M
0+P1ZGit3dCtlcYto/xZO/0EmHlrGzj8gsMlqdh7cAioHPTVAlGfLTYXfeAyOH2FbRVjDom/7wx8
PWZpAPDAlNUxunzFp5rm7S03uuY2xuKhCTeKydhp5SrzTZcg1VuA26pN40qcutqXw83gtGmXAXwt
XJb1jbZR3YOQo44Xn63oc4OKpNKiJObMaq/wJ9D8YB1Vtpa4o/ASbpVmq8H5uSLr/hSA0BzNINHO
KIDW38MV2PWaTQF8onYafQePmP+WaxuyQgCXmsuugchxDCEOuDc2q+z+y5b6k1fFMF9xBBkD2lL8
R4HkKItQpyAIpvH1/oBcSFH7fM9/ubW7n/zp1LiE1HuBVaADMOEdfQvnImOmSEVURe7VwSu66GqW
m5IPZbz6VA9l4KrbRrdhDMIccxJOxQQ6FahJWgLVWPJboFfsJ1EK3PXYbHmP+/72rllHHHRJwfYn
eGI/0rQ5LdeuQQCO+Q+S0XADqvaWw9BBf8jrXD4U8MDcPxFOU65gENgfVGdh71CHzJr2fWsD0npl
/0IaRIz3OmpAW6xbXnZ16OYDVtECvI/sftMNAXm3rdv50RNueFYfE90ETX20OPAdNaUiZ7RyQ1Xk
PsVhIY59FYkRaPcdMYz/eZ+O9MaGkxljoWQceDelq4hOfwq7gibqjjrtT283fhMJovzD77YC5f7k
d6AkXEQflgrd2aj9XlSvhTuphcfMYXwjC4BCvIjgAjNpuKuJQHdjAQibPmJ1koM7yLtUpFmlRPC9
fZOYKWcNZ81pgSxgKy7GsyZPt2Km+ShhB2Hl0N/xxQHXQJBNY49nzRyPuCx5Rfqmp84IL/T8JC7e
D4Ss3qLIkUs8Ee0oAK6OyOryzEQNNFuJHwAdASFq/V6x/FhyTqoaycNlFQPspAZeyOj24AiwttvY
sIzz9PRcdfXqrk+JeSqha2FArWg91VMZSx1y47rAw172xWTatCz7p4VQqJBww/dIFvwFpnoNerhk
zBDdYHoBo/emsaQpi9eoO95eaH3fRIVA3FXlKPrWTN1O6iA4VfiEAoc71jFVaYMLmq4A5yqpiGmT
Dw5A/iKh7ZtS3uhiQPPkVUCRFxN/DZnFSn4xG7EGjag6gH7uLB3bLhw2wsdezCtxtEILWfh0wO5/
fjZ5so4E9wMa4Si2fbVqulRb8cMR0ko1Lhln+N5UpR9czzsw/VAnERg5pAMTlPx4aTeUMORDTz0C
5WVqm/cnDpK7gbpZ4AaPLxTfr91OgT2dtUBSt/21QWu0fxXYaokwjv4SYeySlRj1xOks3WbBcKkz
Zn/4SYM7YboBcIeG3YJ09WRWPrV8UgiCfWbLzIQNLWdjAyJD3upsrH4BcteF2udZ+nSuB2iQCktS
OvMImP2CZej9/9JLC0aFfYqAgYQkYL9If2JAgqnBN/h5DC2wE9kByCSVNEAeakazXpU2RBjSrm1q
IQGo1JgExCV81GLxz+sIe5BxVEJX66pVBYTNSV+FZqkrI5YU0YrByOiBMgqeR5Hx8K9o8DItpbsZ
XOuqVSNnwKX6ml4PjOCUdyyTLhla+YZm2bODM7TdW62DsD4EJr/JmsyKWrffCEXwh3/9zFDXMM10
h4UHogEWhgQ1vfcErvoBarCoV+7VH1WXKL5JjxejSyxT53KLy3Z0XTosMDCYy01ous9xYerS/riO
Nvecq1HIlF14Fs/xEuZEfywm5AH4C3DHofEZjolbDQK1OaRlWuxmIP58t2hgttU7EAutCYjsw7a/
hWeSOudx8mnswYs372aUdM7C+CADX3t2MnzLXh+HDUUl/uKdYjxpUAhew6yUfBYWlMuylGe3xMxg
eOp3pCO0kTBSxXitnVlELuugX2GBiOHB7U9steG2yXjMkusPlDVull41pqItC+xEfGt101fyr2+6
3Yobl4ehpTPBLHxNRpYeJfrHBISaaq7yfLcXI4NGOLhYZcyq1K7qKqAGC2RKwo+QHtoZjLBDu56L
coMNIY4N8sy7uBB9qJLPktGPfXMtmid6x+/xXUrHx74KlryypAvr8pulX7a0UNtmkJTI8ZdL0dpx
Dtles4vJm17jnZGstkEkqdu2XPaT2+6nhkhyWc9LKxe6plEVwKhGPyF3+RSONAh/POb74abaVdLx
mz61rpoHmBfFPIzo3GJiL3ftXLd/TqGRR2h8T4lXFwvHcWEtl2KPn1hBo6H+Ur74EvSQWNGJarp1
BgJurfo8Jw//75/ZA6c3UkGor8OEY1s+ODOWI+zWSPnS+CwP0SKp74ak8ayY9S5dWkz++TwdA2GT
54hyunsGooLyxaUw0S8FqMjxfkLI3YkAoxqOr4xyGSTfGCLkA7FdmduKFTzjcizE0sJJDR2Psf0m
deftDH051kLdYrwRBUmI9GC2TzJSs3m2NybKrKUND5RpNGVw4St8NWOvBGpP92RD0xwXoLASLx8v
1tSKExhON4Rw75H/ed2MBdhhYUACOTSZVozId6Pjr7dI4rQIjx/R3BbvSJ/eKknXm9ZCWBVIwZl6
Jn6nWGb6jPugDYV72rMW9oNDifuCtflk0vaWlm2xM+EsK8Jv6murILRKT+8njfyUwzfPr26r68Sx
W8skZR5Kg21vGnvb5Vp9UHFLgjPF1X+OgL03udhdZgHUBPzYw5hVZQkdSddtglfW0LeUIdVJAe0D
zE51sK0bObRg/vCO2Y8CYaPJ7TVQAiKp2szUQ3OMzDHRzY0yZaVMDLCuq1Ih+a3iuxMg89mO0Zii
XdXiGbFYkVO4/vIGBjktGaPygT51cJQbqpH1QVxqq6OHTiom3lLVqrqwp7kRK0jjc7KMF/ezSt4J
0SODjWoyaGzyMOz1j8KpqTeMwxpr/I7bT6cdpqIY9aWCafwUDzUACJT1rQpQ7DDksrc8eDeYHyHW
QG0HIJaUj4NKSYi55VGTGQWOXdGdOT9yyW0mtEIn+vEwi3nOHuQ6C3zr92Rj4Z/QeyFDTeQdrj07
aXm59JwX72o9igFzchc+UFIkyCeueA6RzM/RW5Y9Eh7VCsNqE8PnXnfJ48ItG9YwGjq+BfAC233j
V5nh+wGQ9bqga0+w8+CmjZAHDOZ/qeGgPvx9IRn4E1D5B931fXRid4Oxo33C3UQSFRX9QndMgLlX
zhQ7aX1ZwSIsKFn7NKCO5j8BALFo28kXRjxNh9BFQ5oeq6NNmAnB4P+tgGY/PSKXX4TS4bqveQEv
zbkyqsbu4DVtw0b0nkJeeUnNGpVs2il3uh8kmhad9lSiZxPwSib5Mby4DXiPI6EO4aY69GAJsjDO
rLi/Iv1fMDZHsYrmFOti+k+V/34cZZd58ksT1AGa9ohYCw6VQ5IizmGKbAC1H3gJ/eneYjAuSWSd
P+6RG1Il4gh3lACJJvwITHToRLMl3d+Jvb/8zNfjew/N3yWurJNvJ/FKPlcWBtQSnm6MuKV0VBoX
dIvuo3icd3vsgH8bDKsO2SOsh/v9PbyDSciMALHUq7l/YjBTau7HJZVziL6ay/IMjHbQncdwXVs/
wfLJXloDaZVWXELB/W8vtUkAlcMx4tEUchn6IfFd82Zbo91bH8RjgwNO/fsB3td9WbtvgPFShje1
HtEGVtwTi+sdMJ9r6hAZx3TVePYk25zcgISLINY5Hj8pmLfVMam1HjqTxOb4EEsCVxfO3u7PfU/z
Fd+XPTGNC7KOmgYjZ75cwfsBDDoYRp71T+RBAuDTmIrvI7Irft2wJvf4uUA1W1AD78mY7RVoCfFl
UkanG+feydSKiPUNi6t42yfHvnJ9+jF7d9JX8AEcUWg1JguMeTbtrAigDX52R/l5WhbDNtB0FHT3
UStIkvjbrWiMsKG39oOIlTtiRgUPRCkd6reLQHC3QiJ/tlzpbO07VBdA/19rDAFv8Ll8lJYSq1zj
0lqIGP35G+ztEp646KdwWW90Jk5cZzX/xTPq9KJ05kyXoUfg13C3bmiK3jGMJYUkFNWOnMFkE6yo
zIgj4GEJSOXAIRYjXvFz44+eGdBPAXGb3H+aNsEHwVefob9DSWt0xd0yNYIa5P7sLLn8tncWqcyd
t2Cj4jDHBQAS8+WoNDXMr6P9L6qFlo34vDenmwUHU87VIiSMrHSdAlXrbHs/9gVlCVNkWdGx39cY
iL4JWBfrmf/sCioAoLeqjy2yuYhFnYaGMEucV+10ibvUXVMTTbUm3rwF1PrW7F6zSSsyakSW89Di
0xZ9rUxY1d2+zawnEpWxBZ9abYtdCH7Ui+WXRaBhJ3rPsKm4l/8H5hVFSE7Q0vsXM4zT+mHeYOFV
cMZcxjgBmmofHqPmg0hV4ss8cCqNiOWKdFc/EoAr2VDgXrtLZYUx3s8pxuF89q8gCsKnjtI5yF2G
1BLQW9Oly/3w7asPdp7To/ISX4hk9+iC388qGdSdUt1dZKoWmb38RTzdkIG2wLFvHzhX0V6pf1wk
YAS22DEE8GU3+zhFb4lvTGku5jH2fDIdPRDknpRFVzvwcNP5HgXkVAKkw08ZYWestF2RqMKp5jI9
0AxBe5O+ACcJXK1y6q1zqIfUy1d91LZPcQtNAx5gWuywVoxRv6XuOT6Oz7B104b/zd8IhxgkUgho
b5pyzHjrWvo6+O3t7+ccEH20BZZd8ChHcuaQKcoiwCUEq/tTUlw78RArRhrxkMRwkSqH4jhH7xZM
nkP9jNaKjyFiGeOF9GpgIaGBpVdcbFRnoe2jv8FcYlc1j2hVflOkn/mX2jA5rL5e40f2KLKZqi9L
90DDrtLk0UUbmul3+TlZ7/vt8FGpOuOJEwEFWBxQIjQJNVl6W7k9mP3cb9CaGDAFqF3JwvAUQtcB
dwX43zumPPeKjh98+P9UVN+YvpU9io+tuYlCdgyxct5dtKl1pfizHB0gEBKRPkdjW0jNjzF0cyH8
0feHHnhv4eT+BbLPN82Ci+G0Zkygpp50z6weEY7j/PvhUhW6A3/Ys5rJXrGUNgpKm4cvfeaRXRJz
XDiwnFpMRmX3dWUIyKaYmQay7p+Phwt9hnMO0AE7eGO4pKCIWcRJD1BPKcVufLQyPzPPxQXcXX0G
2spJ7bknU2LoTH1UxqfyXUd/O3RrpQLi4WbqcMt4XMUfRrLphW4ElzbjJZqdYB7hjT8VQzlJu67+
PqYk5wu8mDi4S6Y1vMt/9dUszElCOVZq8KltmVGaYBESyUboh9j63kHVpRQzBw/NDhdgaKnVsZJO
Mheymdwy8F5Thevi4KDrwNVNtuNs+xY9APsiimvOx3T5JP8L9e3JJrNDfr+4/K49DJdHrCYjMj96
OwX9W5fLm5eyZFby21lv48aEymErYJfUryP94yXsbfttHc6/qQlUU0vOgML/Ukoq3wg52tXblCkE
oZIz5qHU+Bj/FeYxokIfSJOccY6TzSYCM9KDcMPOCSHikmj/8b5At/R0GWjL/jDmu28+IxZshzs1
rSwwFjKgD8auiTt5VSYWN0X84j83SGScmwoTTXnuCUrefWaSsuuACE/iEPTnLQ+1ZFlr4RPkLkkm
FB7CzYVmvJsbgTt+jKikBEr/rb0prYjn900IoFvLYitwUCkS+zvhn9rHjgk8vKVsYCHfM+tbU0qV
K2iYg9fqQ3W3zyuofM4NUMdSxwSPPODQVvr5SH6iaxeO2XQGjYrS1p6xwFcsmos341PXKeCS8Ujf
vKCowMLG174bO9f3CYSmLu1E9D/gPtrRKXtUnaMmmsIhze2bsH5L7fAEt8QtdyfjU/tERh04QWPn
x2ZiEXXpLQU1+dQxXiO7VTJiDfjvHiezyQLpVgQG4zIR98dtQXyj9eX1LDi+F3cWDBem4xj4e3KC
YPGHm3Z+1usSCEBq1a5LME6Z4M/jlGqRFSoNQWj0WHPq/2NMiXqjnm8xi6ZDDiWqWDillzbwQVdQ
9Iara+QhZhl06+2SyEf7l8KO4oa10UV5h2snMP2AeTQdzbDme1dUhfjsQ5QMKhtRKZ9h1H+pjGyu
ZiBNkNj6k5WYUH6LfO9+68yVoQPgrVdZF5cAj0THa1rhzpFgryYd9hwixOIJ5wY0PyvPcsZXQtZO
BqsE1X21wiT6kSQxPPisCOzrWgwlyT595ltPykHhhOBzSrsFBxYHn6CG8nrSjmgIDaEIsOKlsn//
ctXKbFMuiBThQiw7/S7DNerZ40iKphrKpsasMyBBnI3lzNZrRq+H3IN2jKUF+l03dX34FeFPcCKV
TF6LKXewzA7+LkYu+TPzsv12tA8MC6RmNgjhmPYaYnlidLu3W36j1je9l0METs/sP5aChmLptEl3
88qX8X60c++DbEhokhSYZNoo5U5AxijXBSonGsOj954r2mHlcaPBOo+K5KD0Hst2y3e9sHEQw9XY
YX1MKzhWWmzbVUuNvog717Vrj1No3wBX4fsHsdVUWyYkylPgiTPP4yS0rDsOE+bQ4dSvyJerDbEn
hi3/lmJLXuP0uOL295+isnxO3gm5V8SLcyQVd1i2u+o/tD7Vg20BCru6q//1lN+B06YfA9NXOIWu
K9pSJnkjrIkxuQrNmEH0xyPrHi69DXmC9IWSp8MyXY3CztOMzpIvXOqmfN9sw8ytsMUU6mlNFgsE
syGwOv1QNNJK+EU6aPNXLaNLVRaYxLAgFb8SCad37XXiR7Hba83xar09LXT4iqB25WWVe/1Xzf/c
d3liVmzNQWwglPnu2U8HqmZrWSnZVIliUVYZdVgl7VuekN1JIoqdYQj/+4X2BJEP3oxFwo8iZ29v
ZrkDbsfLH+u6CwHE2eGQwL9gslmjYrfuBDJ5x8DhmEebFLHIF5NYQBRNqRtGK2Dkympu1GT6KxGL
d/YaP7mnJK44MleKy3Xh3E83VxeigFAMNGSlbSvSsKqD3cu+C3ubEFgP+2VtzVCJBQdyu24CehNV
4T+mgIa/epkExBVYT831wTRfNrpDQm5C7khIcYV5HoOJd2aZlmG2hKLYus85rNAkNi1fOm6qsnva
bM4/I6na5Tm3lSr5orzb7Wowcf+O8LFiBSjD5g5ps1sX6wZzl1WXQSUATAds9fj0+4R1Se22GNcz
5lDzUVi6INdkE5pAds72/iXCwUVgqZjpNcW5sXoWL+/5nDp6OdRKVXXNSr/JTu8tqImkVpESQHcV
R38Q1qpNbgiV7xS7nMMsf7k7L4/dKu1T510hNiXCgwGuWmwl83WUG3Cdk3cJmsV6psHZVB+N6IWN
0QuUWe9E2k8hyaqV1mbTV0qqbL9Qm/9zCO9J9j784l8xQvGF3s2mNIjLbcr365TGSy6vaWI1z18Z
3r2H/lSvq+b597WajdB88n4zMQqZHzlc4R8+cjhOmFlituKaHvlhSWBHbicnXnPD6P1+qlpAQFvw
C9Cq9UOQorH8lySzT7006457xTgoQd8C78JuTmb+TeiI4xwnOSjEbSJiHyPAlyN01cZaRgkI8jbc
WeSzWYpCxp8Bk5wxw/GlG6695AHB4mFnYitObB1NF0W+Hge+qV9E85a1njJd4nF+EDB0JkA5xHKz
Gd4MvkyDzoXlqxvW1s1hvMuMZLC/4b0XmehRH7+IwclRLSKFoN0MR6hxIIeVuDN3BRb/gSWk/2kX
I8HLIAOPDpUDOl+gZHPhO6J0sRSs7O8PQMBgkJ/pe48t/inRs3RPLhxavCeGcP5kSv3LVzOe0ucn
NKz0tPsRfrZ2oCaIvC3X2Hn1T5ZtSfBlvVnbx8r4ICyDksiK19o1B53F1gvKyfPAjg6aQtVOgXLg
E7/9YzuMqDwUrDYsS2ISAcxaTFE7xpNwQxCVbRNy+9JxyFjXkEpIwNEIVBqP7cyQcnreD9AQWH/j
UHDnEi0a8SmhypBEliYHh9pnirSImx8dYdTPennZnFU2biNvVzItW2fKkBiSVlOvZjis7vb4Gu4N
aUX5fFQVq+jd7CH7vfel3gA1Fv4utB2VC+xlGhCE7PgShME0ivtvnB7glYCGJ6lMeCbrC7pyo9K+
wE201QpmgnelHqAZ1Uj+bqYM8oSnhcz3eVgc3HrOuYyv2WHssDqxX9gyHGfAsWi5Rk5vTD66+Of5
0DtD9YT0dq8Rr5AlltzhZRQw+bvREsEuTGIDSvQnbu+6zG+bV8R4syOHrfmpzlST8r1YhUbopuY9
wlcZ6QyiXVlLLx00sAqJPz5INV297KgZv3ss+iFRT3uTelN0BTQCUP9+KdTDd/ySIJ5y2zvp3WCA
bT8ZS3hqL+18Vjw/juysNLuxOjF3fm+NZKbUg4Ah8VAU7HwdAUgUI8p6TCHL9mZIUJmvMjQUXwaw
IDcyUe9HS6K/k+KUCe3m1q7O1WB0KeQxmrTlD+6TkRZ1AyBYfnX1Oipk+MEIlapgcn2fh4zQKg6P
G68cY62xV/paFJSx/AuXq51+Ssf6AuF92u+/dwwL4luDItUyO3JHDs7fF2J5v+FnXTfsyDr1cagn
77KICDbSEopHtrR4K3VqM0rMNU4gJ94d929aXNTSSDcN6hf8auVSsMtv9NpxenbvcYU4eNeIeZLl
UE1oK2mNOcHa/HH6jXDeQT25kBY1pJaTosKL/l8z42WxJ4SmyyTj/YBmHDNdmqU7ZNCWyPPMvBln
Vhtvyw0iE2PiaIh5rv0gsTV+lm7U55n2bAIPquSIp3aW8LUq7S4f6D5gx50MzjXKIgUC5q/fPaFm
ELe6r9lGzS/7NTA+y9g7Qu15ZQIqTJO15IYAEV56OniUsk3fXszEZz+4K17BIgrdpXk4OnRlZpJ8
++qjYCBm+vYnpFirx8Fa9iwv/mstFzmEbakx3ADge7qhLITRasl7d0Jd4mubNfwdlb6yJyHMkWW7
XF2b5zpzFaZ2AOzKYhwqoPv1R7RP3WtDrq/qOj3jeKqmywRPxTQfjfuCscoH1GV3gD+aJK2uCQIg
vLYsPuOig66cHmQ01MJ4il0WS06XpobnWC6VVFoCRj49czH8GEyptqX5O3dcUcISj7dSMVYjqM4O
g+JnLn2T4rBsZpeNFH/g51qIFTCb6hEi2DTPz7hvFSnj8RQxpFvGggB0iqi1V5sixIjoA4U63W7J
fVrUnHiOLPpxgVFYHtAz2UkmR5XFus4u3JHu2DnN+ka4FU+kVgZ1Nd17CX6nlbWG9uYEYfuw7lUt
AoPhJttjfJQJew6T435fCgMpkwlKEWzp3SDCw9yOHy+fM0Q0niYYNJRV1Qa+4f9uRqS4HM/TY3Jf
xRAkSqnAnj2v7pKgCxxsE59FdBcEZzqOGOu/lxVlT+ZjmKPnFjnoaLHDNdgSvXsiLNdQ73Cxakf8
+HztyT43arqIq/OcsvIxVQ/XMaU8Vr/oX+2xtkyvgjUnmxDmy5jd9OjmtvvnNiGlmvPIcjs2NmWW
SkT8V1CvQ9phy4GFItDcMyWndP7Ok8sFcMa/Zy6x4Lr7lwOBxBEAn2ERLfrNUKKbHruSYQ4cQuYK
7ToHbSiqy0p7VLwAf8j7WA4ttvNWqNYiDGd0KUOFYJHgeWh/nNEAwg5ODTLWmqx1J4/DCI14LYr7
PvpeLMtvSwMYYyp70bNrEu4XPjoJkbUeth4mlzuUXM5EhXCzaEe+qYDYPT1jgktKRvsVnoJs3BbA
A+EJsnHaBt8pfk9S5KzLi9iWJq3dhPf+pWMWPXnKHnJZSASlAnWQJTKHJnBFIXIVNuG0liDS1Dh4
J0EmqEUr0tA4ocWAvHFkP0QnoTZ3CxOySK/zE1uLuodqDpWEX5sYmNzC2WmIQBUR5MPzTdXnaDSR
QlAFzZYFMoiw/DRZdSNAFn/mdGdrEraiad4Q7ruzRD6lHpq8E8FZAfJeaB9h3ntjBgqE33QYbFza
o2CE994K27iK8rPiajghKOfjyQPATEgXmQEIFztLcNp5QeTLWfqFj2aeViIbs3LSjK22D/YekTzd
pH9hiNSEuvFahOUVtgYX+mubEaus5GRCr48s8veHh4dTZgeLSaaesEBh9PKNH+9HW0TOExl1wbj/
p4Tat1S1Ot0IxJmbC8eyLbDNUchyC8bd1ecxVe2cOpyluj9+i/nfeHbRLzZU/wLun2Tw0Alxc02f
HMdhG8EtFZ+VMEjfZqPCZD3W1H56luNkbn2Gb6ksfKQuHGcndWHA7SKyAfyksRozUF0nHHEID1+5
9kacAb+COixIKOSghBkySIoLC2eAp2nbNt228RIzK8mCKPWZjfhJrMpK5qg/iTzNvtmX3edEFzt9
DQjcskjiUXJmj6ikr+mRmKOXdDBTyXoMkGxSvVgyifw16kTpMV0frgo7lFZzI0vFsbSf/LGECz+8
masJGcEvz34fJBMMpHWSICd5O34lRILXysOAxKSWdwSeW8pTrCH1dPslyW+f753vwiLYsnC89n2L
vP7I7V/okmQz+UQZyds2H/lWOwsWiCy5No/CtVJ/X6EG8lhmif4KsZrjnsPs+LzShhxrBUicFU6l
lVG5rMGQ7rZE9LUKXj541N7D64pQjAupc/Lhss3zpXbqywvyL7cFB70A9zu72x1Uvx9rG9UHX+Xe
qaUFW61ed9kLzcRQ/1UpyS0PTd7AJraxwRbDJ8IZlpvCspQBhDXwsxr4UWKQJlnd2QtwKuhPRXu2
0RCHL4hcnlqTXtCJt3KVD+H1w/P7CKo4JCGVMXSn95oOhP51ZZ6rdMzcyDHgqQtNR4iBFjdXHQH9
Af1O2mYfuJ22fxZEqClaWI2jeuy1Dg6lqbMnoFT352CgiNzs2OzwnAZA+8vZyjwQh2efURs8HI/S
2AU0NBk9lvpeIfuKcJbFYxd7hJSkDTbHBJ/kwuQLRu+mMTGz7GixApDBANsJIMTH5SQZX8plMV++
T7cCDqmfm72hgjgnGP5qtuBj/ak+s+vNa5aStgVw1e19OfWE+pfVeUbWNjpYtfuiuO9UqdjHf22F
fWDSZkywhTVDFOxbIP8TfZWDPoajv74YEU9H5HMUP0NDHa/tzO2LbMoStUEGUBzvzUFlL5uSuodN
PnHvG7/hWlB0KE/3LMe9930LUZmRgZB1BeZBmLtvehtaNVKBXJ0yEDA/UJM+efETvJCIFDkn0Ibt
KOVtSb6bi3u+OmmUEfv5Yta4Pik3WFQuT87qouCYI5nthHAPOB2NHaFMF9uzrmGcLRVTzRXOdtna
9mzXdOFzdbK93OAj7ADKBC1DJsZRn2N6QHYQEP+tWZmDTCkga6qygKPlJFoxZlppG2XnlE3XqITm
g9NEKGUCnFAr7MYzh1Tq9MIj6s91EeZd9krun3DtEJa4gNQSuUyJn8E4exqf1MZNJefcQroJuFTb
QOMqb40kjQDwrqUoU14u3PKrdeQH8+sjHo/X/4mEAXOS6o9H68JGZn6cpQwkJvTiSZaY4rrOkHHg
PguB3j1GYTbh+5hLhIZ/81oUdLP/5lO6svEojVYFF+pdViFeHkQGS/+uEKmV+ISHBpWDXv44Hl2M
TROvT9wSoUxb8lQ2V7JMYvt/q9ucWVCncw3Sje17T89iL77QJVgVxhBVvEznrFzYI4gEzlL9CXdZ
NIgu9T/mNyBq+3iO3jAij1k96/ZAZytI6ABN8jfjruFv4GzBE1sKWHmEvns9lG+ltKMS/c7/IJAF
scyXPhR4gcL4uKb/sPA9AryJ8Wi+v0Kzt4w7Mwf4jDerVjZghT4rN+Nn/ajoY1LwkDXYhyjncyRh
1C6J7iB5ffZEoB4ghe7xKOB7Dxa7Z4SHmn5emIgRtw5LiwZuqTBy6XQsos1fKp6PnoAg+FAhSYJZ
4fSC92sPOGZfaFji5C2SfNeml+od2WKXNjepXQWmZ5jrvwnUjV1elgsyjIFopjya5La2LnJqIP1N
Gh7XU3WdERFCxybEx5nEOkvpCPWHcvRMpwSOuWN2tyAnaZmoLZlu9gk+pNNtb303I9WSEI8BnJr2
9CNskOl77KB7c+/gVpGeZeYAlThB7VNtj0HZTQf8KNl8qbjL45lgSPEEGknSJLF8Vi+0RMDGVQn7
yMdnoQw1GjCZg5CEbiVMHqCDtqYvGN3vka7EQqn3hohZ/xGHfCj8r0qcSjQmKc6vHhFmtukK4jvi
btkd+BS4kiRSD3/2M3wntxe5p3x66NbR/6TmcmVH4vrpFppSe2PZA7j2gsO9VNH0iRYNhwshfRi+
5FJ+wfJDGjc0JjmwxUURjv6GAn0vfnEuZikNqmRgEepzCLevDJO5nd8lgSeSfR+aBhhchIQwuzQN
/ByxCDjQ+jUpzh/X5Yars3JGIpmN/XCC8jCxWYcMq+2MANhCleZL1GGDr9Ayo1UI9CoX31f1gtaC
ZbfoDQCcoUDcUg4El65aAG5N6H/SmXSD2VIt+DnTGvEWnvsyxaCWlZh3skLOSLpTzKl/CbFeQpiH
0RqW1mRFEu3z8C3g1h1SKZT0QE9vWFOD3NjvQbZa9pfdGODa2njexQDOpboC0fZQ89eWI9p74LZV
OUt1UZ6sUrw9BRZIrUayHXq8U8J1yzY9L63czimphI5CXGPRVdpTJV55yIScIUb6An03VRb7kiDQ
Mek2FAr0tCY4I3Wq43aGLRiiarF22vI/qZwTxnNMeX5Vav0cmIelRVnZ0RGuVVA8MCvb05WZNp2/
yYnHwscbPdsxIX2vlqm6zX7f0ekBGRVaYQqdf8guj5CwSDtUotyri7yHQE0z9XuicF52W3D8uNQH
t/ODsdumaJWNFfleXZlNLcxFCXyYZQ3cf/TT7TaGy9s+L5ZOpt2julOQC8/VCkXFZHf1B4OR6t07
Q9hZCmZfQQY/ICIJ1iJIy+8z4PvofRrZ4zPwIZ2hSeyxDnqRHcN1DikBMF96+uQqCkk+t4kFmp7Z
qxN9yPEvtna/JRHX3roqeoM45ytwR1kzRBHDrvljmZOCSMGJbcM39tDo5/55GrKkdPAnUSU3f0L9
sZ3QCLduikKnQ2YQ9hrPhuWLlbDRlMVnieoV8OdXN7oxk7quO/Rr36oMN5dxvJyn4f8imS3iKE3x
qwUSaguKosTR9QO36OZyaMKqxFVZfPZT9F+44gMtMPy/FaFLEeYLDXumhappPNwJJ/9mctkkyn0Y
RetccZ0GctcZqLtIzVNzJqcZA2NMbFUzhaKEuurq02PmVUT5qfXHEIa6KA7KhCtN5XbmgFkCJ83E
YZ2Pn8j6rD7U7ENafoYSx5zBApeyqJXMOm+eiOHyMa1uR1DLSJMF2AqzRnjnzKOyAGqRkoaQFkSI
xbF/lr60nYUdilLBd8GJQSTc2EMb0BbwNE5ymXfLLRiS/tmDMYhePmdP/bwAb1qx+G6eUCLxig+1
6kBh1zAu2ZL4V+bXblAiDG8W6+gdPNvK9B+S6o0Z7WBsghQJcd9yI6Ku+ebNQtCWXjcUEIXGQ5lb
IGEVn/7fXbFEoXHCddbirp/TBO8Kv1+hOjCw2MEg4RhYGrnQSjHnl+6Q+KYvDYSVRz18M6fkofn/
yh61CFseF0lwk/gNvRLVwSmADA5GuUVAFib64DYQyx6mazM6QHtpOUoT4+cgCtZEGHR9zzNKRf7y
hwUQagYd784OXZ2to8MifrB00uMlg/Jb+3CpndpWNEOVKyUHhA/eMkJTpxJPD49dHTsEv9ZYz06b
mIiGtfXOwDz/YZIySScZxVZVsD22C1aNJrS5fT0X3mZg3msVnrfXUETiQqHLjhu6mLOQFPCoC3gP
I7sFdQe5lDoo7wwQPnZkgZzrmrKLpDMUJExDlfyn7wtA1Lkg/lOkXEckLy0BKEXgI9Ws6KIZ4ldX
g8aIqyP+Uljy30tDos5y/tl8o9B60HjHc82gkF0EILGImQKWp0XySGL1CdzMAXw7AvEuFb1oH+Gx
ao/Mf9V6hGTa796yqkCg23iWN1glz+Rqnzj93sXbrhh0ITHV3B4Qb1Zdcfve69h67jRvwr/L4VPi
ai5JzAzgaqQih0q99fH/viy1UFDoxAS1fA0kixFOpvBAkhxNK00I4AiaMiMFrd9OK2Cs7TkQCpD8
97zpMwVTH1tFMvyxuuaZQq7x4ySsW/b8hhij4BQa40WtV4GW58lE+KUYiYkF6WQ5FcSI18O4RI3U
jIB7GWUMHe71QKPqPeaCBeWxnZ/CBBqK+oTAxZFh8/tjdJ11W9AyO29Fsa98Fl92SgRzLZwqucPE
D2bcMgvyxPATJGiIldC5uMRIh5twzeRTN7wakfEDy/NhdugpVPnAL2L5NzRK8L+FnEFApwF3U5a3
Zp77DdstP3pzW3LHmndiZe9LuaKvx9Z4OlQNQSDhpC/5BVaPEJpQIvJpRcCBPy6kDikuOu+DO5sU
P0fZsaEhrEHXyTr0YjTosIZ2cmH8hg1NBgiF0TMcFt9wziS9QlLRuOYtr3Tz4h9mdENOMRpqKgOm
kKO98s8ThPZzDD+Nod0OUTZiyqe4r/mtIw/eGscDJUm/V4EUoTVYH6aTP1HKGza+l4EpSyapI3hF
qNd3BwD6VuFR1M/VpyTODv2XEde5i0/iz4ySTcXPxp/9kEGBSyyb/zgriicCSpz2bCAYgmZOjlwm
8G+px0lG6sR2UZJ5/dE0IoyoP0DqWT54O9VA6vaXaEMIUBnA3mTGBGQN159n6wbHnsmHbjbgySCe
/9Vi5xqfmE3NgN6UgWgD3jigp5ElIGdYib63o2EZ8hiK2E/KpXzFUNbTDeMdJhjcEj/m3jxAy0qT
lTPbJx/RlAfC+EIVitoQDURjo+jfdmmIVrwDaq9r80IpLHNX9cPJGKBKTiFwjsET7QyEeE7S7QpF
h/KiQyNPrrZcRDgOwxagwCT3kAY2NXxS6nVaMf5IOfyrIwr6En4VZj+0n/FejKTLBS1+76GiNzf3
8lEHRBE7AQyqrKF95aeN6dkSYOdiNlr8bBlndTougtwZb0FeWUyy+wHjMTd65HiqMKmRwSITgTXM
jXuhtCbnkyZG0pJlVByE8YN+mYr7LHva15KGLAbsLqm6P3zql/T+qf8ZKx8y/BqVwErRXz7/vGK2
RiiuwrPTsJOd4pDh2WFe8xB2gPiBOmYMvVZAAZjP7qopc8EWaBMaY6m2UTXDdqESpk6SiGKr2xvK
Ny6tNuB9by3R1NThf4QZNXZeZ2Zp2Mf9JpmPBjwG88hPdKyu/7ybOIczK1yAl0fLCS1sGMaVwbew
EguruXW94vzHOXonw0qhEHfVTmKxFIAAbLJY2vJTxyS8unjbyZJwrwl8rOU7rlRHBthOsZaVuZle
x1lvixmk+tV2H1DAduEX/AQ4Alv9pTkqMPkol1X88yxIV+pWVISHPpvApXvCa9d3Ygxj/oJtkVT0
sieVFpIUCEVCe1naSwdq84xAw+Ebwes2AKVG3OGhzysksdgYXPVQskfTXK6M81BDP8EJ+80a/vsk
Od+bfISHyc/SvJtVMhNtJg5yxkBFzty1eE8cr/sx7s2b3fbpZytSdkc4y2e34PVrce3pV2NzbJav
UJyS2E4A/SfADZR4sIIPiQNx+RYLTBlEy/n1XwL+40q/I/Sb4l2HpPqiGVzbzA4Qm2wxm36f5Et4
/YQWaknIt1KDTIqbMo5SYjuYZuBn/Bn2G+6RS0pGGSr/WOICoh36dAJb7FTfuA2bPVWlzvG7TkxU
p+Brdwlq3gkp9JNbdYudylLzMU/VJosYY+yVwmE9yVYE+r+KEsC1B6Y191h9Zz2o37UxOVFkyr6V
aLoe/TIdNmbbpFSoGqDZNiGo98vjuMSY5ympsMc5ZqdAnxuJG4ZGgjbuHd5mo209IPaJWlqCFQwY
4DIcxiUf520ysqvJh7c1nBBnws2TE/ksT7VamzAJ1XlUHZQuJmKZsuBzySdqEktV98J4c83IX2w9
s4wm87t4G0CYXLlFyL7vyBKqBAcgMG9Xtyob2mysfE8TZUskhAdwu0pksJjFH0XRr4hAteANMXcL
U4cimJJghrWp6QBK6tpA5UbIox5rwTM9XTVTbxReaz84JmFwsVb6GoZ2H72OldmDT6Lr/vlVJtfi
TjYPe1ZmuT6JVPv0aoqfHAet+9YisMCYU8HqKhDtn69v1R2a6K10eQ9LujiB56yWIQsxVt/VT55o
Y0A2iAgh5Lp6YY5CKFZD3DPkYwXVWEjnYp1Lb85UDAtgZGDJR5ORp/EcvJhrEfVd9aBRU+4Q9Cxe
ws7Z8x9qlel/wIN0OuRGaf4v6FdODo3ikARPkUJ0kZj4ZuqqRY3m3qpadILm1nRuA9CRkMxxuToi
sMLw5tIS/1K2k4kZlCr+0fIWW7kTm7U6KYxoNslSZhH1H1hi6uC0m2OmevCQGK8bOkumYOHp8WIp
cHQdkkCu1dwCPEAIGC51oS97JvCr5OPzrXeDe781aGWWbpdwBq2J6EDLXx0kF2gAgMWa6Gg23maL
cx6TgmsIAhCarTNaGyDGyh29Z369Dce7YvUL9nnTtkyjXkKL2Ygvh2KB97H93ANCEv2rovBnWwDY
rgqJ6r09XS0itXGNUGI/jnjEjlJjJRqu3bmdPrhmGQsbvWWjRJrTIzWCwXg1CaW27ooamRCw7CQl
Uj1SvVIQEK1sVsxPgyqSgCCIQyi0vYc4bVo3xH4b3wmTZCp6dGR0kWsnJ304o5VWv35WdIDQSxRq
80nXseiOryF+mAyciq3LpUhY+RaAf//e2/CeKUecUGSBTzhtHVRkedR5/jJqDuxG9uAyn6j1dxA6
oGLJYvqcqH0xdyKXKd6AOggjkzm1y8uT33VRByX9rG1uSCt6pknt6rvvyNTjsuYtkyH1mO7NJBxr
n15NgoadhV3StHw9eDpk5pp2S+z5q7e4mySTzygp+ZzJl4RwEjwfs1OqLWozPehJIRz26FQTXuJG
JpHPyWI0XExITKsgDzgLC0TGtCFuErp8+nTn7ZwNFOnfxGrsGNoxULjCVRCQbZf0JqDP+IM3QKhT
LyPsF2faNRv9b5b7PRzK0zZrmnIIvUUoLddiNFhxi/yb8VPlVNvTxdE6XAac9oq3YSRorj0b+Oo+
rmpxwm0nVzrkj+M/VQjigdtkf9amnqRI5kP2czuLgnCDxtQDbq73GVPHiz4ZA0d6QVt3MkWtOLVj
Iwiu+swy6g2ttf2h7UbG0yjH3bhJTbum/lGbjtBRy3J5ivfP8jFzs0XM71KFpx7k4OWKx2WEc4RJ
eJ2DdcwQWc8z1+JkAktQgxMWCk9OkPdqbN/FY/Ktt28jQpNIQXXBkP+OebVP/r4War6lzLtm9a9B
iila8o07ZoyQDrmlFp27JbL+nYqbSe1172qdbgCOXkZFdAWjsCWlK0yUrPWJDAFz0ajhZfi9lpYB
E3DgWmNp+HSwLKV82LHKS4Fu+V9rYTTuNT72AcoXHdXdsBd4cjmgrxMOVXAPkljXBd3dgijoZ9DZ
wPFusH7LCn8yAlweoRx5SLrk2TkdL21Vrou7IfJtP8NguO5e1lrZslJPOGvIp+j9XrysaHvJe0vs
zJubA1y1AEzSvs69TDhwcRicKWOIXPpCG+jiQQCRndZ95HoiGhqMIDFrz11uuv5tThDr1QLT5+gE
bMd36Yjg541+bCCnhnogf+/6YrACKAPm9ExQfHpLH9ia0V35GkYkHTUcIVVxme+VyXqsvw5mAhmE
0G5RTjC8RLplWrpW9RVIujXWTQXk8YAKm1OPxMPm/LHEYoySXYMLl413jNMf01ixDVL55O0/IKwN
iOnCk+pGZiCGFSVOlI+LiKDdZe8qtZfQAkMCIR/5CNQtuu9mxLQlLtzXBgP9IUCTd1yVSW6WRYFY
lUN8tz+bnUAz82VOyLu5J1yoDC/Qs0H+5G95UORuqAntZ7YGB5XFFvRu4sjIeabzEHTi/og1x29h
UTYPdbgczacNFVYmV3S3yZJKQjKe4xV8Sfs/N4MhVypq+xBSKCc6x+OToAuBD0/DgRMb7vziFRZQ
CG/Vpnoym08uWqHPbhM21VJbS26ei1A698Tl34se9JbB7DGsKAGGzIG+jHh75tG+XFwIleTzI6iA
2uuWLzpy3bitmUKTNmGvBH1yF0YIivKgqQiwvNP3fj5Gd1O9MinLw0OIp8WqygaNE8Jbr2HjQrZD
JjDwpBBzlGDmvLbZGH8564NJPO8yeUh0lCdQ/3izEH5PJmsVdO3yelhzu7eiarOWMbVIbyJbxzL/
bVJZeNBvhV7FE7TGc9D+GcIdUq/p/Gxx/3izyiupXiT+HlUVFspeU04KkrPdg0ui4HEAIlFJo/NY
WRYzMVr3WXHPhTm6krNR5PygVgoySRqzHRwITsjF+9cX6tP1fZdSQO01kuVIO8Kih0Pnf7Yc7ohP
ek74K2L0aTT/OTI5x0vyMCuc5NXejFsICmbmnlsjMM2YGVPxuyTbnTah1cr4u4KVRNVDLmthm5gE
OG7XQG7y6SMQhJz4DlYcDBvl1TRdNta+4e5CvRtQvy4igXkxt/ruFnUp5M6G4+sCO4gzIXVxTcDG
mB159drXN+Ig+c5FAUGBmQcEkzXdVVrEBhhCeAXisJiLAkS34wVAUVZQP681lZ9qU2y9OhqQSbU6
ZvGby593CZl+dMgE0hd3Io6g7dHeJS+IXNzVO8x3xzv1acQwlNJAN8J7dSwURL2NjgZeTsWgsVtB
O6ttzmF8iuRk8d2tV/x5zpg6vaBiW9YgjQawDeuTDdtbAtrFrveEWvhbL6P4zO2ZmL1blxcbAkYO
xArXFRYX2XKLKE3OFnuqwCDEj+xDoTadXEhy2j1oh0gV1evrUQtJ8UVmGrafhYLARi3ZQl12n4Wq
JLyJA+nECByCC2kscHyHLMHdI6552K/v+iRgc2ue3pUewHSB2L6erD34PbQmo0l7tBDRWQprwFKS
DlE4qJWBOtQU5XkFuR6ArYIRxkvrxtAuio7dliDnrsfgAyCB7vrwjWQ8AobZcjPQbJXdDikDBrPK
6kfMalc5laCe4s1HMz5MBlxVndw2uGtAB4y8eB2AQ19Vu4p3PS7XFaKaXh51wQxQi7284lTnWmKz
VJ+c6mdVWM/JZozIXXpYVoSP47JF1TstcbzrLe3IvKOIGc1V8IMWMR3mff60EzDLNDosqHQ8ukbB
n60NSQaficTfgNXCovpCXOFwx26EuxCSRm1WVdCbTeb0DcqpBu6Sf+vd0ZVFphG2Nswt3ZkBXeeQ
taJ4sxOZ7HA495650NlJfRB81aq9CE4AUs8dCo29UxCyGBWLS2Ebf1g6cZqCPQTvYnIlaQs9q8FK
E8//I5CTqSbRQpWa1cF3+sN+HuLCaL9alxCGQtq9FJb36UKRQYd0OVab8onYTI2KWIxTRHhQhkHr
pq7izi4Lpyc0f7iLhFuTj4GBcE9nYDKqH0+xGChEp7J3wa68AEcishbPkWMBE+7GhGyeBF564cUt
gz06eWwxJB+3e+fhab+1zjwOC10Ymobhcb9T+ztTUklYKkYHrjTjGMS2fP5NJoDbVPpRknEy/hnp
lwCcOesRB5pqZezJ1+fCZq25w+vRKj8VVT7zeCRrfgfQIl1f4bzl539T2pnBxn+nD11A2aqeQJ3x
qPjAI/5eZFBe3Bgejj/eJxAZnhVeNsnv2ualwc6ivUShSb0QHX7+DVEljALhnmKxx2uQFDO3UmLQ
hxsSA5CmE8DBNJQ8s9Ps3xJ6jbQnoTcpLz0r3LcyQrH7mfMLacK5nLa+6i9kxV5guuVNsbbh7F9Q
JktjnjPU9Wu3LJCcoJ+aLqGEqhKYivNnVEHTjkez9i6RrH7RdTbGEYiZRhCwt9NLVpPHN3YgVj81
ppj7wSpfms/EC76DpYIvUyWC20koEUjJg+oHFIVKtkcdHN3yLIZ051lrPO0Nxg4PRTaAZeYIrFrf
aEQq1OH/G5A1Me7gcWfxEYwCaIx8FdJjU8s/Lub0dniaszSO8G+hxC7Cd1XNdohGyw9GlTH/83Gq
vkZLocau2H7uNbBA194Zihlkmv+lxLwDRSx1MeOcchyT0Djt4H52pRaS8XaQrdEGMCA/kBvw1AIx
X5+y09nMve4Tl11pYyVOTDzIjWA2vjHZPcpb19FbYpJ4qQCr+1sZDE+QPoSslWGB1bD2CXbV5xdd
zwx1WyynadFNih5lgNHy1jCjrxwT8TjcHKbIITd1D8qXZxdjKcRMleL9uJPIGrKKZBOkpd0WcrJE
Z/5RZ1siTjGf74xIXrLYtx8wA2oJW1BIp4QIfW75IOD7R/osIJc/l0pYk3zYbbkk9xhQlhGe4UcA
KCfSnvjHXNgjI4h90QMbkvzywaNn2YLYw+GFHuwaC2/wywMgjfPXKnKkeAi0yDD/ZOY+q0qPdHxv
SYBCSlZwy2ARVTHVhgvt3kVwm+FUM30UShmYDSeo9BAKcdFVb7pv78BMYLURFacfWYh9pKnyX7lj
h+K1H57SwbFnRCTQWLlmO4OoIHR+wuAT9DlQ95HX5/Ldkk7j5wjrbDLI00D4fyGoPR8qC2jbpW/W
VoEGM873I9ScZUwV5T6AfzQSQcI+8lP+gZ7ywwlUe35PWVQLCTkrszyR5cAcDI6mzRp94mjfak2L
wn+c669rWO+21jHw8Z60buC6V9+hsy9xZyQSul2GxCpxR4Gu/4d0CA+czJ7tmScUDHNjLNIZLlfG
KZow1l69lzzzbT+0+Ntj0YfmKZpurzjckB9TleHt1t2UzskrhhDb1+eMQHsa1/RontzHq36B4VNJ
QPxCwBFczJLDnF4LQQ7l2W4BfQsK5Sb4IySoTOgzolZAbekm4onEcXz9MYN/TOvohkytd1dnu/4m
ElcWQLyKAYJ6Gg+DGqSTNH4bifTi6/c+YAe9merJZmT5YPtbhQsEia4ScfEfqoaGu3XYPILNlspR
+D00kmbslbhNQh9PP1NDXF5vNDwZ3uKS8dTSLGz19sUzw6JgY13VjEDzm5/YGnUyWL5yid8NKZSM
oK3WQba5m9y0NsNEa4rCWnOvOkmS4vEMFUhoBBn2Fu6WctphuUwhh9LaLInMrBrNi/tOa0iaW6Qq
BRfF9IOLBLk/Zy3fd55/YjJIkIWo4VWevIqts7kjH1ycCcFAnJl4oMLxTPJFrbeQjOZOZquE4Piz
kKLkYDUoFy1dQ9ByfaPfhLks78Aja+upJZ/AeqlkkfOhM/QtZccXxS8oEp0WFG1EJsn3m+o7VXVT
/7c36eGHywopf48Ab7MuX6g+Ob0joZQGXhkyhUzUTVBB+/UzYtz5n8bO7ylQE28Llg9z7PhR7sf/
1zY7ApscTqRmjiUPmX48V+E44E6lE0PbpYOIyuv4k2EBCm/lS2sH65+xIVwG2q4DrGr5gFA+nPMU
VTAJurK8JtY48Wrdff+5ica46a0/eAA3B9N4vHhGwgfSz578R4HT/hcUFqNmTWwfSO5Mefb9ciwl
m8rXhG2bXGlwtJkxxo22fMtn24Snu9zG86lC0nAGt5qquvfgkT4IxYwD07LHUdxmdcEps/UiIZZv
uj99x9W8TUgXYs6//VwDyKzqrKSqdISkXiSOqaPlcpHbODMc1jY96cfNrc6dpYceUfKiOC1cTU1P
HR0AeB6Yox4JA1I4ORTKQ9SQWebAZbhkYaTyV4WIRvPHI2rULO4upHeiGklC/UdOvNUWn+vdfleL
zpYpWoynVOqSerHAgQeifgOCnkZd8CYQNL8V6qG5LtXALwpS/ikGTpCuPV0KuIoWv/xnapP2IuOn
ZEz8X+Ng0hlXKyWrUROoXBTSy0urEj7bQe2HJnJAzi64wOCx7bYwoS9nA/POlH9SKt0pzw/d0bEU
H+VQQOer+FR39yf7V6kiXhHL+rv/WtH2BkzpKciQSajC391WUZKYdmufGgyNszLg+CTnMjjrJ8hM
LBo8QgdpjQML+t67gMyEqv+oZvoqZbIb1Twiy+M0M/ia7gIHG3T/x/xTGXE4QKMZWZmesHZnRtH8
miVw3iHgf1B3KJLFdl73qf2t6oUYZzLlAu4kjYDI+hKFW8ZwNIAoSMoZG22CCUSi9zMpp2QJrw4H
YFv2jDqxmRH38ydLE8ySYp/hjlIkwpIMLkBDRYw2HxjAvYIqzmqwC3hzdpCKSlX6wEDLNb58Gk81
eICihD9oiya6ACTgSngcL/5X4N0Y2IOsxROCARhUsx+s0HmolD1kD01Auyej76x47C/3XfKC47Kf
aAHJ2qKFnCdxgzIs9TEEX3v7pH1LulL+pTFfIIUPczMxLVCd4vdQ1oglr5HDU7kAOpzaovP/Plav
dCdEuhEW/DE8lec5YqkG1n1KGgOe7nVtH84LsV/+gMjP/O5EozzTRxoPwvbFWdTUcKV3bKvciFVd
gVQQC3dX5JGw6u3DFpjoWSb1yoPYNO3VHtVHgfz+k1gTlHR248Gcyv26yve0dG5nqn6itXq6JW9t
mkWxiB9pgyIrVemuVWiEvgZJO8pbzaNxDMg4uES3oMmqgxZa8MB59zkIl8M4l53lXx6+R0B17OU6
dT1vhbXuk9wM7rCF9/tOWBaeEUwJkmvlZtS3T8K9XvItTdDwuVDuf4i0EPxKv5sH9KoNTcMCifvc
2H+MryzqeA5LNPQQEUdMzgJWUKIFMJBFFsrrPwNmHsEfhRDObKwkv9XHWYR2oxCo+gAPw4dNxvs/
TwLN+6hfjGMn/GAsCP7CcdJktIv1Nx+P3TBFFBDokeqI6KbPy8wM/kWFuh3WUZjOfxvbRfuwwvvi
ubi35Q+FKqkMWtCi9gwKwpw2ppaUJp2zZXIbXXKF1oyd0DF5IsJ77Mma0a2EUxaDBQUp6mDuLJnw
VDTB+5uqJBpgHc1G0v2PcWH/mnLKW2b0nkuGCMeJ60wKpR5yYmfxkUZbsNrTjEOI56IMpbgKV+x+
DTBif4hbcLqWepttuBK/hszY1IZWb7s3J5G086b9CZ5Wcb6X5XormlCPYeZHkCIDBEttvJUSjTqz
W18iU91c1YXXJzAr4LxMwWqgf8j9zTZecSV7tNoPAg13116u7m6mKfQCWMaJGgKwdTXcwKlJn/oc
vAbcK8+euqRPikN2kUnP1dNrpBkeR6iCufH3rsBK/rF/Tm4qjw3vmABv0kEun9s1d7pXExkuor1h
R3FWcBx/Q8zZv5KxIWZm0kMUrGgHf+Zd/1J85zivZ+a6ljvLLYv8mvFhLE1dT0rxL662k2shwo0k
B3cJQzMgNdao24oKD3MX54LZNxfxzo76h5+yuBC57D3yxcQXeJuX+FrpY64yxuxNCjz9MmZMaz28
zB8Dq5mvtTLO8aVUeeAwr4GP/0ysKZsafyJDkpa3/YKbsr6FmxrGHih46Fvpzf3FyhABKGznYfeB
8NxTBCOJ/hMaaycLlO/XkGY86KZfeBqlwv/a2v8K8pU53Lgph6uvouNT0637uAkjJA+TuDJHv48c
nhuAD6+sVc2spK0PLEhIHS2iTezG9bLL0KISF71/5DFWhWLf47srQK6m642inMlSvGywvbnQhqMv
JjkozQhi9Yud0MGq1RUcIdKMEyVuxtAhKKyzInb+gQddTJZz4AZw9TsGsAPEoNpE/TMVBPQu0hYw
ow9DdEK/TLdwWq+1282oVVHKsiT2t1y3T2t7Nlb4jJJuOdSKS6OJREA8FqNASuUH/HBXjpSL7ntW
cAn42ivLzNZ15vShQi7vFVmQQ+/X2q7XkxDEqM7U5/uqQXqAoL1587gIPOLMXEaOnxDKsC/HZLXn
pciyd0L7vMnR4mG4gS+1wKnm8um5oKOQKgqCavN4KZuE1Hc7phYyCt0WQdg6aKd8DD8Ic1MT07ti
5jhwlVVWar7Kbrm9aObUADlUzJGmQbE+UadGxbJM0QWS+qRbi6wthoEeKQPZsvDiPCOX3EmVjjsl
hnv3PUGLWfuPLNUlROArx5waRxXDDncV9u1DMlNIk9BJXUIfmvBcDHpYrbyS57Hsxf1UlFQ7fx23
gaKao8XvTx1/LbOuR0cK4N/dGfD10/2D4UWjqqqlY898mEN6aQUQ49DcWh1kZ6NAU/vWwWvXrpNg
bTetFzcqQKqFvSv2b7noDoQJm0KO0m3lsAP3byuqQoutJhaGMtRITOOwz6WsuzkLzRPqb9aDqvHs
9VLdR1gpnc9uqsLr5Je/6171uNSy1+eCWwJsjaRoi3oeRoDz9OMPu2ghkrdzCqt3cEbe8RYDb9in
fpjwMqAychxBClYJCzKYlS8XS0mOVQs6Ffw8XEt/uqorElSc2qDmmKwxs6q7mcVEKTkuKEEEqsYh
w1BqS822ZspxviEHrbJ1rhSOGO69PsRh088vvom4kudsD3ll8rt5ocN6wGuBtKf/Rl3AhShkq1n5
QXGSfzFkLZG8rnTgIih6iK+IE8NpXXcBi7SOA/Q8gWRtwjR/E/4XnlBu7jc6zs/doXJVowwSiDv4
InYrOtvC7cnVb00ptyJOxKWXw8brQX+G5qCmdccWaZpsG/knC6pnSIWowMTNij8Vu5EVsCzyhA6h
bcVMplgtFt5gkWftbJ2Qhug8BH0N0Qa3eRGhGOs4Z4Lld4qEjiNttsfqxRDOrr1gWNl0K/B84CX0
ugNeOfWf+IhBGXvxZ0aodczJmguyJnHDvVj+b0N4r6/JGmbKr5iscjEJkgi4b/vCPwi5LK4sCj7v
fcFU+V65KctmvIuya5tUX19QZEomHwp3panpIzPQDxoQo8Tj5eatSa7CfssDsNJensWiduEBFJZJ
gAvfp70IOhZJiLM5V0EmMcp+LJxccIQarIXWd1j9wEDwW6zN6gDFPeDrpAigCEGIm9ShRmQhVaH2
7gKBChokLIwuDHvH83jIgZkf0TZA/RG3dLmZ8cZnjAFn2DRF3Fu5yHBOR0jZ6tZx6iOwb+a9Hyry
LsaBZRIINLyqIVbWqvCZd4GOBCbqF0kznw7VyvaUqbj6yR60LFcrcLEv7k0g95L670j2GAAdjMht
ZQaJ6FO/G+CGK2kXOmwAyzQxSk9XWYaZZDDHJaeYJKGfdMKaTZ06EylXxeQeM+bD/1Llnp1d+l7R
VdymWOwsZfz2BlwUgYuLoRziBP0EIOZHrbBCP033vGjEAG8kEUSnyxqZH3i8WFW1coBH1uB1hIqc
5SvaXNbef8JN6WBtaXoI06+SGXYMMU5rx/EqF5FGytl1C45dPLxf3fdMaT7tB5oCJXgVWayI7EYl
zKalxlcH1D9ZopHPzHbrC+wF84dZunMEuUyWq19R+v6GnmPS0Wyjay1BBuuDZyn5g7oA5qE6dBRy
Ksm8pcWTqBIG1flCtHRGHUocYvlcG5AU9ogPF+w1liqvmO8JgPohuNjqKwskUy14GiFkmuhHcZj1
ixsZHGe8Ob2zdd/ASgeIWFbGhiHJxY50YCgWdU72bGilwgVcTPsLgL2GK8YxG6xLKv99mw84qASf
eoFCIkWQRVhdG6w91458h6kkAFvSVh0VYsHJT79f0pBU+U+uU/wsSTjaq24F1lBR3Dz8KpeOzeBH
qFLileN7QxR9lDFU/I5BpRy+Y25cjRaCsLXCcv7rZZRefHzPwDYH7dh3XamEy+FfJyK/WS7Hbagt
wcfkTJZRcz8X1uEL3pcoSzlQxFGH+PI17iLQ9f0A6RDue5rPr4jfUcXLQZqc0N79xCIQhUPM7Cwj
KBiO5tvvLW59AAoqJo6zxtdK3tm37LZfm/xM7e2mVZGmHukPuqh4o2lVnqf+POPFoDD+/Q8V6vPg
wZ/B1JNB+uoZMrmZdK79/MYqbsR+f1V3oS45OcSaAp7T3vDH4V5tZP+CLQSu5lW+/dW2Wy90cWoX
V1rNgUD6+fCAnEXOIeWvhwqr7sb9QHGUsbUQE6MaDsQ9uOGjN7aisQg8Y+lj5RCZqASbaYHLgnHJ
MwjIk4LR+QJXTPKi3wxDpfFSUL3KWavi04VFaXRHvBPr4hINUbP9QVQjxnxZA83j6Gk+6uBEU86V
mpZ9Ed2h2B4Th9RECmfYFMqcajLHi1zje3pPEeLaJCKNNH42+K07bYhv91K/FkeeJ27IIkGGwtRp
o/8M/MEZ/rOux0GhmHzACqvRScTddJ02gIekvarEhdsenamSAfIOzAIfVD7vMuTvYrz4usYlVMl3
XnOgX5z4hpqnLF7+hyeeEyX6ht/EyhQkbFsQqB85mjZMJPoFFQYNY5Gv2qXMqUaniPvpPELx3rHv
v3cF6oYv2UvXw1Vu+neOfkj+i6SgYuxVUDb0HEfxz69E1f/gBI0qX+QPj0AyWcwExe5xGW1piinz
Qz474V0zEDANS3MYrHgo59lRIA8M3NvMRRX5dy9FcT42gX/Jsxaz+92kfqXPSAvuw/EWcrH4qhPd
YQaoAz1myWBUNkljeG3Byq4Vr2errqmtCfNVirvotnMQNxsBeiXWQP1ILZf1iFDjRv9WtLv6y5ZZ
6tAQBvw19AP9NgzA2MXe375/jZx7YAEjBg9HGrPKr+dJPdZImdiGER9YREsltZ1/THQjdfLqsQ4T
WixP57D9jT4kKp1zQJyHsvdma63moCOvnt0BP/8HIyqWStAySEV+a2FdwCARHBWEt9+Vt4kTJATn
f1p7qiKdSnjrcZSEZOEoVPaSNSUhwI6iBAjWAXxeiC5m4Oi+zfgAcTA1V5Ka7ddm//EHZvkH9LnM
LDxszED3+6hPsVCLoXgPBUxLhVDCD+QNU/47Rv5pwGQFonTfjfOxf4njjWP+8i8gFw3kdplfxgtR
BU3HqWvAUGJnXw00MpyV3DgMho6w10Yk5Y5VZPC8Q6FZhS+90ic3tSx7yQjkUvrFR0cPP9aBlJ9x
OC/n1fdwpn/OvfAfpideVydlME8YOHCImBlj15SeskjBreqnEhaS2xw8pTatA7CL99KZDfIIuzkH
ykBI0SUTtMCan5oYbTUogvM2W9vC6r8s+ssAyI34LE8TH8HyEgjTx5GYcyXovvp5IKiKiuPn+nP2
pf2XBal1e+DniNfP89k6x5pwUbKeZVHdhcPlNbL6unkCW/zvzI8YyjtQW94tqerA/NagLJK4UtZi
E027sLz4cFnSvBlUVMmEVXeIjHRaBsDAakTSUz7xjCCyTtJeFOtqRa9wiDFnKXTMD597/uIipSw4
J/mMA/YXjTBUcPV3Q5ctxxAZUyng9r/PgB4nWKcQyYMB/W8veuozDkj+rAssf1FxpQCQES7q0LZ5
7i/0SpJnCpnQB2ssQNXaz1p85Yj8926IrRD3lTgSZgQ+XKwq8addjaK5rIwrAALPH7AdD66SFAvS
SiQvqwBDFywhcTz83LQlD03PbVdFWLrj76mFhIbqt2eTwIoPs9UNld/+NrQN1anL3xnvkUFEr0nE
qifiy/REqQ1cug/FQx0nhl0ODIC8T/8Wh8UWaXVS87E21MugtzzimZy6z4BV4SH9AjtMRjMjtUDs
RjKms1w68dByRD/Wa+BE996M8rcNFPQMz0uvjkKCduvW/h7dsApEPyQMaW6r8isGmyZ0U3lx139h
HRrl/x9gBmmZY/9qmpxEYg62HqLTN4ZXK1V8y2uaz8+Yw0ukkfm+u9YL1c6ILLMaFyyQuddAZG8B
lIgHNUMAO0cU/Mgy1/hGfi9bo0IWGB3hY80K1T1XTa09qL1CY2yaD5iul78jDUxlf0gukHY5r7go
Dpxo96ahJtjostcLhhUrbtJYh7DkayDxUOCuIx3vNGIid/5z9ePY1qTJqMMeRtgDs19HHMG44BVy
pBZ3YV4LyOOp2VMU691uNhDmepUrFsL/1XVeFdEvX1o5QgTeKMj6Ei0/j/wM/DObkTcSFLvx2bnC
3uRCkPrMWVfJKYJerZ7lu/GOlu2x1BOPEhrosTJtn7zaapEXP+7ZcmB1jjjzNcmcDtJ5rKhU2aCU
kFakbFA39s6XDKIh+la6EzQort216o9nA4hWRN1X45FZ2t9iU6jTSbq52btAZaJNTLbZA5r9/vqe
TfwGKex4gjJsnBNtwErxM8238+lRR8zGlSBNCN59+i88yWYmgHdI494/IKYeqqoIKTIa3xkszPzQ
rH3dZIgb6r0XRpFpRrHs8hfgWkye8MkCPxkqR43sRpaHMnLz+OPbAY/gBdM4wwIbH8osHDbH2HrY
MXO71V5ybIylE7RH6wcTMp+u9dhPJ+F3xBlppPW3eCf3R/EykcsMu2fwgZVVw0cvereb1H82yHuQ
tW5XXfsf7C+i9bZX4gvB+kEwHMS7IojuzzzjiaoaBNRQMxcaAalJ7K0FTl95fGqnUI+ok30hgZW1
nwPNHDywFp0HEbhqojp8cIayQXS5gQcyLKhzisuPKgGE9gfsr3dwcb7VkdEnIn9Yg262wnU/JhQ1
oVkPiyqxZq3EtRlVAbbF27ZLdLyqgVBTf+5aBR5nPwQzMr5/5cZsbClSTLPkePq0buJee7zM6+do
uJVhc+WFCvaF703C1UjITc/kG3L1YB5v2mT7NzUBheHcGY8ZvNhNGszWMgreB8WKsgzAPRi8dDox
vkLv7x9J/ua/bjJ/4LEruQlFuaoBQblRl+jSImegRfRBicV9wTPRxGxiBBF+E1lDmTdDnQrkb2eM
WMxPBNnm9PVthsLvhXtFb1GmWyMO8Mlm0ifOfnh64NOfqotqEdlIwR2KIhW4B0vdFLwHXesD0PwP
m85WljWc5qmTlTYYgOsTO6t41ID4+GeDjthC598IhWDZkzwytdPJztMJQA5VrLLns2JCtH/mBIcf
hYKwoiQC6gizGForZIBH8WOIg2JPo/YSyEit1Qbi4cZRD3PhAnGH0Xib90AWPYjo0ELSwRwwAIuS
SGHbq3Rjabd7bfKBnh/1h2GIhIAbUbXtEe/CX1aTYbAyR13Bf4xewNV9Zxpd7Y+etNV7n5g+5eVu
bMuUTaIJXYUqTkNvwkurK1nCWvE5HH8M3F0ntj9xAaOkdPiZvIy/BGhT83kgzNHELifAkoNpCTEp
2aTZvJIBIsr9JgkJfDCfAK31jXGPoiphW0OA/vWQmwilm1zDZaRkPocBFTRH98lGMgrhaFtNpJHn
Cs0ShpxIthAQvcLSDY9oTXvFcFEqH0S7LfkXDUq+zs4mZElLY7t2x7ppPYpIuLrzCWp4fP1hIeoW
AL5vHBbyszWEx61zUCTgMAwcj5XwL5dzdKTpa1jv92Ie0RpMohtL1BGesTuVGemmdrOLRarSCzO7
QXOCjf8M3veMJCGPkL6MPOuQnYElwBr6abcrXmTn5lhBifDdvn+FAS0HvZJIqgtphB+Aq/DdBbPn
LUQMp6L00QuSAMZpwlI/eSKjgxGkn3i0wQG1YBIPbYPv7ADjagrb1GFGy+0ASiDnxY2t2nkA7YDn
Cn/Eb2ovVb1MREeucqL2Dt43RJidgq2vj55BTYWKh0q/vIRNSThFvxY+yAPPWTQuj8FSFhZalxjX
hO/nsloB3svxg2upooKONcnMsCjQH4g9Ru8Za9Cz87cE28Xq1pfZJj5hinE9LZ+pcuZxUC6ZFG5H
zc8Qa+Wp2OmhsPLMbCq3twsGqhZpxVCNct68wslGfh901rkia+3AFiYJavkawI7p9WAq+BWuu02p
py4cZkOnmcF/f0a8bgTICtHuea+j4ln/tQqFhVgPAbVr/ATZ/x9xG9CeY5EqS1Itxy/EMfwf6Sua
5FEtmVBi09chL5zRGWTveFrfm8rgAgsmnrZabyXvFmhGZO5T3Ur43Zz4SsAhQed4JUSAQNK+rGaq
U0oXQhMj/+J4b2lvtULvC/8OdjLZwkZuXdjWa16x65qCbJ+y6DW9URH99EOUweziKcdoURqPWNqe
hDwVvHmkMciVC2k2JL3VFndgHL8Lhwa2dCq7yPbwiR+y3zoIcKttZIsgnfPlaZL8UAKyQD7BV954
i++1xgdacGBtehW6U8PvM3H/Hw8b1AQTqJzc8WdCYZBE5JqCrHBX7YRzghfiCPmh7T5LD543Ej8U
9a766LcYHgwI/VukK4i7McEDlNFeYsXZuq6MUHoHEN494mRGpzuwmJsCNTWxEge8Wh5KmCogw+eS
7equqfqStw1PCyKcY0Z/Y3JzMDgm1aJoVHsjhujvUW76I/Ips8xz7je17jBZHND6AvJEvGkHIWP8
G7OQI6wtHY47IjF5NPn8RdKQgzKq+xiym4JTJ4gvXhLeRyW/LvmQiduomyD91WXxCRXl7yli3Dqk
XKQg8WL5x3Hf9gFVUIsAlBIrqFb2a5Z5cWPduOrgIaljuHNFF7MwLUnT3GBs0rwA10YEeOw7wQyi
UryoLjXamH41uxozg16/oOjru5Ub3CKMsEqp0lgoTdaeNxUef6awG+CoCkykCJ1YNwU8Ygy/PKlM
SJHntxMOByOG9OqjM8dxgcSsYB+1ey14objE2vECV0RR4sk0TlL3DHatHVWlx+Zr4AvfLZ2qDqSW
YfJ/lami+DCx4uRzX1mZeQELUKNQhRJQs3nSsvDlbv5W5dmgWkwQeVSoPA4qJrXP9BazHpP+C8I5
03IEDsNSPUzsNtCDw1C61DrUILqXzWAeN3csFls9ebhvE883X352JDS/vV3ZG7aNwcl+vq4r8I8G
1eWd1hzy+gjnlZnVrozfmaNrJoNsx8vFI3356fsQ90gE/wr8Ip8mJ5xHk2gN1xJFbK/vsLvOJkn8
eGXin7+2R8HhMsUoopUKu/S741Y36vfs0yoERpDTfRRXzz3Z5zHWUa1w0adUgn9/6WtYJVrtg/M8
tD61QF9S/jZyX1H7EYFPMcPxBugx7XrzEELFCwuhmU3zYyji2Cim9RIQGdmjc/ovqcFD5uWM8c+G
gAhY06zhlC7reWWvg1fT1JkDIcBQc2sjEpWCc3BcGt83Jb/FAe6kMnlNL2w/QcntLBq2oMiuf8Y3
aRDuRIrHkp5a5jnZIrnXx6ebtbsJ1fMp14W9G0Ge7bc1osi+THGG8dko28ytzrn5MARUtPap+Ny4
lcH76XFgRDJYJjVmxHYCVjTi1hnWE+6Z4dfa7x8i/uwHXRk6emQpwDW6LSMOvCdUTZqvl4GC2qms
FrG+aR++gjv1bDX7qnH+WT8eqqRKPpEAPFZuOwPzlvxoB5kipLcfxDzsLYMvNYPB0u7gEGLpndCL
JBrmyUOplBE8bXZg0VAqPSvmlzPgbwQ1dzpGH27/v28j6Z1pA6hK6wxOUauixA8wH0aSsfaBJYH2
+P9oWujcxvb5xH/U2jISsjgyiwuuSn+W5WAGbXl0oO8Ba0frcucVNJQtioi5ATMidIUni9lPdyfQ
uoxVbR2MheBevuo652VYE1DvS+FotHVpf71pHmeJrLWsY4A1H2zVYNjjkyMDISKK88f0IjJORYwL
2BSmkXjv1cUVpqgfO319cXwu8UuvVpzD6mit5he9wOBftPPcAuL6nt6wLGRQ7cbAf67uGRxVTMNw
Ifv9HN9wcwqpPgNJ15wNIVk+Km1F9BZiWblq5gxml4U607ri+CjMDIp1ank2EJQwzYfITJ8NrT5H
Q2hJCDgC7Ty1x9BH/5HyA53IXPw1D694zQTbPdlLB0o0+J4o5RTQC/44WJEXC6ZooWZnHgA4rB4q
rTm6dG58OZkPSNeFuIMDBlBlTAbAXNSCSkp4XBmEq2zw6EhhIn4u1qVHGUG6bK9Ru/onnfjdt4D6
Dd7f2CFuE5B5qzsF3b44+eXKMbAIJl/QKI+Xpet3DUQUmP2nTBhULznQro2suR2XFSxVh3QTxbjk
sKPVpHFfUDKbP0c/brA7ATRv5C/47KYdlIgbESmtQIsO0RrCrW6AoOC2PaEF2/7eBuL2P065ypHl
NmP9/OVIDDn6rGVDYXFWKfeiDam6dTgrtLTeyaBqRgoX//GV31QiV97kwxOsWYRC2MXqQ9ifrRnY
nXjceUO7XDr55vVCiX8dR9isZ/jMEVI7VarZuEo21TX97vUiPeAuGC7EcMBWsSbsQbOkwZjuWLEx
ep6V5uBvK5gjb0fYnmS27zufgW5RRT7MMZ+l3TwGpispkrrZC08+aLXpP7nyy6exL4jpeqxpZ4Cw
sZ564YtQXK3wSBeeCqHXYHA2Oyk/u+whU0Q6wVZblKIQmApo6fa2vr55di9nRPH2txrfFcb5H6G9
OP5nd5FY15+PnXoVKcFq4aZSYxM46Y64O1Eev45cY39KhaepLbFWQsdTKlIGp3F5y1LQmvsHusmq
GtUarxs8Axb/2Ms3Q+C4R3mqoBiHHGxZIcuc1B1G28tas4WINSJ5q751gP3vg4P5X2sWkqYCGOR5
0ZZ584vPkrhdU+c3GThxsQRivdEhaWa9QXheLn6nWvtIiwvzol0RHFjedsP9lAQlm1A6OjkWjrmO
PkLCZFBkdzCVnhsgxyonNaoyFMw9e3pxxPAK9k3K9kPuQyEThVSgXRswxWINweU8Zs6hc3OpCKtC
/03Tp8I6/YBLuphYq3bpngQeFBmZYxoTPrSW8oT4cm8j60hMMHnJlnlu9PPzslt5oRfO+Pt1B40g
T+N/GzO+nsMdbnqMMoXf7IOhuld9ztxGghmeJ4HSWeMCQfVRTI63EVqk59ErToqHs3Ym+hsBIPR9
NC8TC5dPEzPy8OOlFS7flSg/jxWOB/+OtbpnOE91JPNgPiBI3A+NXr4vYBg5LGnXAXQVGD8HhJ6V
rRGStb+XF8M7bPH92wd8hw1/O2h4gQzwQkdpn7Cz7jN45cFD687YObsRdJtIernMSps6frRX2ZHN
CyBRkV4zkZDETn7kCPiMnEa1hIzxBfV2nWfwnKKbT6ziW3fsvZwY6XPBEerFnTnZr35RdoIJ/XNz
9F9LEWb2TJDAxRKIvhy8G5Zi1oY9CpSkRBtR22YIrc2rSMn+cNeRUCBHjD7qRA9bkQXlKJBm4S9Z
RU7DV6wb27SknrQdxoH41JEleRyT5sh7/ssw7DSc+74FZQYCGk8jJqxtUOwisb+27Ew+OUN588pf
/2SVYlpv6N/gGRuZFM0WXbub4Lx6cmHcDlBeHWhvEDsPpc/NFVLncoVbQFWM3c5LGa7O/j10l36/
2OnhhRxPog53F+DPJouD4ppQx6TSZ4nrlbLLzgGaussYkWLJq8/sSjrB/1Tx89W6dFjBTQstJTj/
F0ImAoMFyhutzbyqfE443e0N/+2p2Pym3O2fhsGcblWk5ckKlX4QZ1UnUaBj4uZFrudnT2uewvqS
ZjTyQnovlz5Sq9eirUCf0dUgMAoEALrGXFL71E52d+2TXhMIhkUx/znZU5nQgjMshDXxvbVYCpLA
ss8nhI87VJUVrVNQJu1ffQIlfEHKqQxabRiuCtkq9nnKP6QSEzzKcmcGOIyLufb4u4f4srzaPZL9
iVGFLEs3lz2S02LXOVLlnHEKa+E01hrNKuU/pxy/D11e8MD7PFzS21+PMI7QvTgxAvR6IEK5r9Q/
Euv9rcRLf/yHXWzTJP8ccheR4nFNeQY5yUZc9pvE+KnNyRhauL58VysQY5FWlzO0gPTl87tnqcDo
fZB7xuQvZXsDLKrBDcxLuzIVQDz3nJI8W3o/jYJyMmWfrj1gk1NdJavPwzQmSPezaSQh0VqT6uxS
5bhAZHRIDEgIsrdLEyZk3GgiZS8UOTt+mArngW5ydHATzDOCPeJgh1QU/lbb1YW+M1NDvUJVUB2k
4Z/XTsG8V+5RvE5Yy/8vVt0JwOcTkMAEHXcDLJozeXAh686Cd/4Gzkz3MKnetEezrETTmLJL9Wxg
SWdpp0wsPdWOvPwQWizWNZOn81UgtlI3nkpMZzc+3N8coKGUvYvpYD1ThCd+rw11qx6gkNtC0YBY
C295o2+VDYC2Prn1pV5QQDV0mntuPEniPpCnWR6q9gnfh/RYpP1tk8w2RhaWkeOpflrf1Yo6/FCa
KA/cISRxFzrfZYx5l+1W3QdyWUFUrL1QPJnGr5BY/YuS8Lh8lmYvGPZ/7ev+d49/GnX3UgHr3BOW
e09WJ0f4U7u1govxbrbzTo4JKInDtyG3bGnQ6A/vdzL7rrIQbNYofkd0fJmZevbRgZc/WaJc9tSJ
O9F3uS5IyOys7rT1EYMBAsG8M2VOTyaQLiWdBgVcBNXt6ca6Xo/0N1ovG0OflBn2iiTmZcvNykyF
TiFZIcux+GlupcAaRQziW3lCWjOgpuRYzAoM8u1phouNFbZz/kJmilc0JQkwB5CBA7GHeWpTicrQ
UgXp1gwlJ0opyTnP8xxZm7uztlgdj98WCAjrk/+5NoKab0H2YRBhbHSC4cr215p2gwwMKhoykYwl
xewxaKG8LCVpwLoJq5XWmBKxYyAbRPzZhVkQu6AJth/hMaaq9s56UQLAmoHJyrjbFk5SySjSNeSF
K829Py3WpHaRT0k9KwqsmArfZ9qrVHLauDw8my7VLOCA8HPXYOzxFnLGSOCkFs0GbON+rnygr3gA
AozW65Sn3c68D9pUBdBJssCLz3PxJIqmNT8AJlrsY83Sab36d6Kw4+WUGZs0BTLSkda3BxzLckOt
TDN/eQukOqkRWGhd1I/Fj8Ruidg8Ua5/U4EEwBNEs0kLknmV45H/Vyw5FNz7kIGUzC5XyGDWRMml
AQsN7ZQBZ38zslOQFoB98yTUX6SBXSxVfvmFBhr/3ChYBwYEOoV5idhABacg2OviYJoMkGYG7P5P
qMUm2LH7q55bInut27D+eVNFUYy2th1bEdguj78YKbKDIxdC47lBBwP/UIXVr9C6gxUoZK3UD6n+
5MH+nDy2BkeaKv4c38MXA6imty9G9R5u6qkharNsY60wB607C3eoXJ/W94jivhrUtBPVHck0AQHN
gG61WxQ6R5H8vHlAVW9flCx1hTMt9gZ85n9dbxiEkOqWP16yems9Jsl64vAXT4FjDpEcGfzAqgRL
X5ig9m4aT61f3vUPSrzn9OoucU0KOxQvOIS/2sEwCXf74CitqrZxYwzfT3Ipdj2Zr5HUHYgPVKGk
x/hWLtpRmH82Y5RAobwtVpRVdsutD609GWreKA8eA3x4SatgRaBhqqFi5eJusHcaCsJrssCwZsiS
mr04QdAeSrxBnGv4dH4H8gKH/pFFkrxXS3fZeQU3+xlbFpN3TaHsJ93fLUeGgrIa2wcXMiOiLGus
eW15mo99ZVnSoDl+BRKpnaFLGxxYYb9sai5gDK0i5JD83aWmdwV7rb4GK3XvwkbqFl6zg4TDy+3l
Wq+raTyxlQ4lms6Ksdyvw2m3crLZCWeChtRPtE2Ttzly2lvGQFsCZAUZNKGlXZ6obyyqyMplpy43
7aaP2zSltzZQvUT6NHmz9btnCNC0F2+7EAv4zZUkXmV2XPirOMMHHlx5D5hF45WNkmaZAnauDXUY
7raozxemheG/V1RG1Fl2ioQfYFxlED2/RXjRmrS8fLCfHhgRQq9PIWa/IQFJ2DMWQCHwP7nJAVla
xJxK4+tw/VRO5HRtTHrltO30v9DgM3UdTZFP6yJyIKEksUzBNGRL7uq09EeuIvOsCXg+KzYkKD3U
dP8RqY9emeUpP8YAwgvFx3z2oSblEZ/i/7ReMMlEOBSQ2fKT1stok5PjeID1WlpNqiuOSWhnpV8w
niAbPmXJGrx6R22jmpiVbVEIDhGOlOLpY/t48aZWsT4jMToFRDQ6HKGHedI94qwkvmiPz4g2l5fG
Y17A8sVXhVpwca4ioHfP1CzyJa6Rl+Njs3D3hDP+byM0Dh6wp+Hx3I0InVMa3WdFCa4DShVX5KH6
qzPS8gyaPwzqJtFN9iXynaYpiUWe8JLoCmRFvmkHg2jB4fIzouA3yDwmt1jG1HLf8B206xX0dvxP
iFmaMZCXlJo8cVEv4u1at41+Ndu2dDfaTX3WAe8RqIo5AaKxOacEvWUuM7yidxUTd8zatXqmpaDJ
yeuifwDkln26lDaclQ+SXiQOHrzBDeS7RkWxk38pWCdVmAu35WGiWYhF+669LMYIM0y7nNz8BSQ6
S3b3eJls3/bY4PQnBEvRJ8l9+XhPq9qqUvHZDoLZt3u72IOc39DH5NCp5bswV9BoqvLLX6deDI6r
d9LtnCn3kozxsmgw1r2WFySZ1Dh3WOWpxgxFh948SiD6LfMQgWXEk6rNrz/3YBwZwMU+E9DWKxM5
Glr45AONZvUrELjPmgAahTx9qtgDZiVcDT5TqxMgCJl+A7syDhSKQP2DqhCH9VT4T/IqNxnN2sUl
3opaI+ct59VH2r5L3Qbwhrw4FxZFHDEC3s2qtBx+4ezhp4pSMJfrDhyA2uE7t/mUf39ca1DOF98n
0A3d38nt8gDn4IiBoxYrgCSTM173bcEsHrzhs4wshpas8FU4DKaWjikoDJOmmauqpzWzohZf1bzJ
8U/Ykt1HFlTISoeZS6eMgDffHNz4JX+3cSoOw1BAvSbec7swrK12+YOzRHZFmULwgf4b3FEmitsF
nT+Wx6JZUI4GB+plEPK9WFHfkF6So97jpqPlQXVrP5yOFksPErVK2H4je0QlMAWNAcOlACjT7ZRc
P93XkmLzfYELbIB1N6E6nJwYD7uNvi5F5O+8pNacLlHHkzWcfTLWbinL8WYK0a3dwGSOygPamTYC
Cl8XrIqTWhzvODHe4ez3ruclrt68A4x1/bgIshQd+tCfzK/syLNFOhgOYO0s7CVK7Mj4VIUEgs8L
aTH+gVHJdHzlzfJsEkdi5iTv/bM49/pyfs3H0y3QYW1lT99NDE6aGHcR/ZqJgZE0IBczn3rYxMMU
YV/FKQ2skqJ/GKHKhvzzPIChNqvjVFWZ3Xgowy4JdD/VogerTw3xjrKtkOVpkbnQZCLmsdQ92+nS
dFDY5fTquTeTlGG/3vjog7II6PObH81KJChrWSyyb4KFvMoKWZBcPW+nUwp0dp/i/sfsL0HVw2QF
VV6dR1rUi7mvsRw6be0599mCwBH6HlVegAJNx3LhLQq1+tW6mPT7NCc1ALh5z3lYiPWSCVCwHm/G
pzM57bH3MxQZJMeDFIfblBKiU9J/QSzPtLsv2oxSKHf+HApY4TYUY/9LOd/FtW5IqvQekDENVh8J
SiwUhhLNe297VzwSpVC4OJTMaHM4mdByLbOCxluL2YzTF57JXDy65ONkXRmGRey6DmCS1ScghnDl
UisWRmGM1pH6KGe9iO37lFst4Q+/wtPLyRoZXfcgjbLpSYpQp21NIvuuidquD3smoJBBU1JgOBts
mbaurcN3bMKSQkZrPepyZU63BgRDWKdCR2GtuWOrtboJdwlLqxjQG+c+mDihb2jiibHL/MfCycri
2JtgVelAx2qH4VtTFEw0fJXVUQC9kQggLxWtL6VlX/gKYHd7Ba7J8aw2gxBn0eyUBmaCieHoUFo0
GWRjTevkkOCwYfUaIxVCgn9TTCSztCg3XkPlVs/6YrN7XLvVHB1nbuub8HeLtj3qlxnpmDi0/DFj
sAWe/GLNDyQHCTGZFFx1nMHskKhHww7ZQhLefWjwddKxjKgeWHaYUCmpOXjmoNzyxIHOrXAMXiBr
jJhCWH0YVcYsgvhkaKyE2fnrTWr2vIm68vUP4sZQpJoX4rZo6JJcVnoQ3BonETDLMV0RPbiDoccp
VPV4lvsqVRyugXGnKngJWqodEZqt3SCcapg7G40UX2ZvpMVJm6xfBW0OcfNlurJuRRtVGmCQJdey
5xPZRspXaL57UpfIZfGD3pCinloSyduwOiOeo1J5+vwBeH+xKhyJdSiqn856ulMjRxD3W6uxFJr/
k2DnjF83zU+Jlafu28Oril9oGZkqhq4UIHKseisLFSyHrKW2E1iwnWPPl++XXn+U/2dSfhyCvT/4
4DtTVOWRlRcU8+z71/fMKvV78+l9ml/3r83DP272cFOZjZ5w0FlOEfS6mUFEwAGmfVIeaH0Y8KSY
e1FLyXMHY/nscNI8vCdyOtger4S5xsjoxQs8TWgX4J51iNZUhbBvNUyqlQiY7tRvh+Ue8UoehUeD
3tSwgqB+A+JEPvoWUPRTFDyHSLZIvBMt9DRQcnhZpW+6Seoj5aEE12L6T8vGlqUA7zwlQGrQI6Py
JyrJNF73OuveICZjZdCF409Rp2NtaOpcKpTxh4QRw8ducp3QGjT4kmnd4DZGiOgTqypOCSU0Mfbt
mFoCKdVJB/wn994oZT2TLvyyMYY5ug4KqItFFjGzjfr+/s70Mc8vvgH0XV/EHp+pxwGR0/dfLpoe
yW3wxoafKJvQRhsWXfTTzebl4PV6YBRvLGXuJrwVc6v8abAwliNb0Cg6P3oT8bbok+ArxXpykzvw
bbtH5fAFdO1e5o4aAbCspd25GkVusEP+4su5BoDFWon/z4+JQr+kLOWrYAHBK0Ef3mpr9QK/NScx
D1H33XD3LMPCSeDDw5GYWcs4fdU+d4lJfNZM8B30Pnsy+5k40z1K82FyFRTPH/pm12rQDCdpAzQB
dZK7mR1HWF9XS5tsEF7ggqW19lSEwl6NwKsYdvHabK0FEWtuEBU5HDm6Gz5fTrhn1FWyu4DwqTFP
LBtEJZWvkE7+eLBHmbK15GNvC7SOY+nTLF0R6y/e3R0kg/0XQR8zbEuzUtnrVdaz7nMnZcTdqV4F
mBEP9NscUjDGkVjSBEfKBaqIo9TiqVLWYpFZWH2jgE4Q9aQQpZGUYs9fnPgj6kedZNfcy2ZX5E0i
BGMBBS3KiapMpc7s9/zUj/Ei6LTB6Mmwg8xpLPdHPLUdrsVlQuDXCBhLfaeBplCn6mZWfT2ogzpq
Vb0GAj9QrXIcA0eKjrHukenC0k1q0TUl1y11DLWov1RrmVa91t/45hXjNI33543CxeyLWzyrZqBY
1rs46HgYMHd1Yjsa5SnDBWUr5CFU2sUySOgr4luwKnVSlfjjyjtf/2x1MziWnNs0a7m2abLP1GI3
twgbdrNyl1SNPBjawTKmY2kQ3pZxekfOGXZztUvT610kt7OKSP+Y107Bb8nfw5x/vysMKCzPJY88
s1e8EHck+M5sjdSQj6ZSyLJSZOncDKAOilclqDFQPKhYLkBl9vCXEJQi9Kfs6eksOazR1ctKWXTZ
pi8ANaEvb3JZyjzJeOIGvpuAfG8NQ9NmAJ4oO50wA5C6A5NnFQ2cJWWhHXl8gDa/fUoD1/Ea1h54
WN697pGePoCoA1HGhmC6sYVglXfYLl8nt3YoJCiuU6rQEIdklA3XsdURvh4xhf6+p6scnTGuddKU
7z9q4hXGowIqqH8QX9MASgSIwx5T/NyBPnVY69czIqM8JgPe7A16yVPXhdQ8cx6ouKDYOIslV/TB
xQXab2myRN1PYGWZQCU1ZOwYSU7/XeaLRxlKheTRG9yHL97CDRuHHNkNYbB6kine/d3Nt/3xbDUI
36vYJDQpuDOyZ5ND7Fhk4q6qS0twCRI6mIzn8fUM+xq9G2t57W7rAIkh4sYg6teUKgfPXPDSM9OI
Chf6Ivg1zr6SvwqnindFuVe51kQO5Fv2t5Mz5CilsmGD/pnjfn0xxT8HrcKgehj1nA5bBgKKYizW
QFZ2uUglAT2jrY9Uncn0DNqD9/pqrnL3uhLwutKMUX1hEWi0G7y5VP4660twFxjQ1JAT/4an5vWH
HEaNk5lj3ZZN0qK1pi+07N+QQwkYHujhAcR1QmcIlMVMYyxBDeDk2pgBdKKx9BJeRbcdCYtFvNbk
HV7cayckS0fN94pWjBtUwlRGKo6XVyhk9f0epLDccTdfFt2rCNnBiP+wOB39NwE5y+Xnqf72SaXp
iQoKYIW2szymu8L86XTXee3QLpv/rVAkN3zcmVyc31C2xSWnrIO8qG5R9GZYBKJkxWuRDGUY2y0O
S1FrRMMraPlXq0PzBcRPYwR36bqm779aiUw1OJBBKD2pIw2Dir9SgDYDvyu1PB/jXYiSLbttzmWx
wzwZq6i7xjO1KXPvjG5jABxIBnvNO5cIuG8VD+DTKt1QzLPqmoyCnuG/7N0Z21P1Eu+h+Owa0lCB
GzIwdI63iCzl0a6cAJzlqdUGsdaO8y1AZnhAT1Mq777mm8DN275V59nD1e+yrZBi/Om8/FKJpXTO
2Q/8zk8H4f6LWLCpIcqfZMarp099WRr04r+UEORvcICYE2NuLr9EVilXjNJ4vnAQeA6ejvAFKlfs
s0wla91jgyvEkRxhwXJS1A1Qz5zJ3reintupGvII7jPMMbGMwjwhFgtc99ugOBRSysA1DdG78HDK
8OCYsJSy7eljUt8uNig+xTbWgHusKdtFXcrN1bqu29CWER3W00351fHIR/Zc1uOI2K/aXmAZsCwt
X71+YhpOsqFN7QZHjpzlwtJ/Jb0W2pk6a6xGavAVVsP+vrBbul0mGLzVc6/2jJY4Qt3VfSOrR71P
BxBfOvUuiaGO92AhzPv3ybQSy52pLPrKQx4gpUF0szfOnHiMj0JkH5LAJq0azglox+9VDOh/u/6G
Hj91eRKn/dgcqoinJdvt1ZrcYQpY+3p0p11zlVVzO+kC8UZgWFp/Mrbnx8AM8ZGM36NHWOdHxDR6
wW/vECSY0PVdbGDh4N6C6zYSbreBKUk2TuVG1Q6CuPRgziHPfdsmeQ8oMkkFHAK6UXPwn5w2F6ml
EtsS7rEGQiZmdRBLgL6zSiimkvTSFK7PQrtgXExvyfm9wRZP28CGcD45y92bUVPDwhB1g7PNeVEK
FnAOG9jm2KYPjX/QVOfserOg9dYSk/DCRFeahpS0tlTj2DnkLBx1rchRvoASAx8w6zt6s9LWPfdN
0h9dUWG+a1qwM3FmxY38Xv8kFhY9kaxpwKQWvmIl1vtSqcUfZ861isGkbliG5MTs4tBDHps0w/kj
zlyHnmsQuIufQyCv0Z195d8imjLAPJb5nVrPSZUysabhli9jaNXS6I/JVS6/eL4q9Chojokue0VM
/t72APeEWtpGjNo1lv+vuUtJ10NmDxxb6UYwWZylqBkQyXW78gnfPK72xiF875GOQoEBZroC/g/I
BFYxmafEcGwLmWT5pBEfPAtTYX99CkUwnZnzfZVKQEWW3aglcLm3e7Q7YMMNOYMORp4G7UvccGoh
YmOGR5fRpLhRM5C/Ko9nc3GOjnSZGd1UCxq/geJ3qJAnGtOZoiOqb0/bSfzQ1DkxNgtG5+3hOvJu
fOsB5vc7nzpL1zlOznmt7/p+XoMIAcu2gDd69w18pN6oGZaIdf0Y8iCAxTU+xqfPAWFH9VSI895h
E8G6PzD/OGDRcuaFN7Jm8kBOHUl6JElhTd5bRtLDBEViSTU1Mk1sQu8cVbnw6LdEdHuRX6Q+QP2N
zV5CwB7HQU8re6aDI5Kv8zLy+Q1NK7Rp8MjeCOfl/QjOK4Oj5hyrm0411qe9rWZXhCdTdN+pGK1y
rzaNXdBsPuk3ikl6uSfmS8+BGSASenCym20MtHpBydggFS6HcWQdOtHSz5qbfJdG88mL3SWrCA2h
fvlJ0su9YvGG/wjk3aOc+4RfQEKCZ8mpPMXrMC8wHw/tDYry+uSaU/E8VCPyntmWnKdLa48JstW1
ZLjQdG/tUQu821Y0ZR9gEfjgIf9pM0tGbdc7wef1BtwWNjK8VPc4AnD8FvnCIKdh50eEriTNMzlm
e35MCojcUNYgfHwYmG7UV43YycZernUnCIA6uws6yXadTka0KBul2QXxIHZYnYjGtRbfVDkXwJz/
WcyQY5H0Hn/Id0IfELGLKltPpAf6wEASLNgZdl5JFPEdaKCbqA3Wc7EFW/1v5BlvseKESf+Wxezu
d5lhA2THnUEHTmv1cTAnnJDXyBtGDsx4k/BrR6st74dXiwHgtmjJoT/6+bSeupuEGMDjEwqGACgo
uoE3+MS2TyjUkxgQQiSDPYFNQM+Y5+mpR9O6hU8bALR9AeOssFr6Qfrmj27/sHh/p85AUttJ51yK
9OP639uM7dy+7BkDTLQkZkjtjyKEVyKvx6iTmMJTOsBciAZ0RaGPGibIXc78HjpSuOPGc+dL4E8I
whXAbScd7TlCNVlpUFtdwpEsjUtrNdEIP/sVSi1IBFugzcnvWr9Qm9SNX7/hOdAmGqKiOqDrDUdy
epaNcpKYKC6bihYb6x2Ft+BQ9BMi70S4m3jCcSPqQMbF2hnogpgB1gwvODxNn++iFa9SdT3IPD72
eLuPvzlPPcCs6vt/AA+Ci6DODXoebmW/mU7u3w5fgJ4pKyq8KKh26A4fs4O8Z3YgtIEmJnmcPwgN
dUIz4CA47UVfSjqy3k3Fe+DCXcWDu18WIz1YW4vxjBMe89gFCj+82Ep4TgqwxioPEdOZ14qmS62w
W+tq2abkoX8KdQ3Rmx6VcAc/S3A6f8piiObNxoS6Iyn8sAPOWAPIR88sY5/70e534AF1GtwhH1KO
p8Soa/OSmOvEg48PIXazaL6neLj7T2fFn8Pe2EQSDfLkd/g0in4KrfBSa5cKF+l5N5FwEPTgAwxv
bUJE8YSt73UA66YfaZrccboluU8juR3dOf6C5VqtvBJbq02IlpgJqLEG1OgeuzlrFowc2oEpN73O
kb4mKUQLDxnABB6cZnfuRrJ4pb+Qie8yEQPJ2vhs5Q7Uvrqd8GAepocwkjyBVpHlw+Ubfyx8juGT
aJ9jiRgij4Orl7FiKl+BR2Z19yNlNvit6SLby2/UGu9NII0Tu39LxWzE/CcbVpBNTR8kvSYz5wfu
yYpAIHuO6mpD0LjJt7TePEQfoQ31ksbFuasUy6Z8TFuAAOLpU04pSkZleVST4Y8hZZJ5AAKWsNqZ
giDvzQJCh3CVIEzrjbCazujerd53DUR+x2WViltd8DQ8xn64mf5ygG6wCy896tP8zUOYuubsKYnX
Y6iWlhbjstyYXubqJxGAmTNsSJynvLw6UaxPWwSHW4xXkgVGK5X4ymXajsQrbtaqkdcPTeVhU6QM
C0fW9bkS1B/a6e5UlGT1/SNUOdSfIdD8DeNzwLNiIScfD6TG8jRSLcd5FjgvSibMQUmMEjF/rQyH
zgMj6D9w2wugcFvB1nhQ5DGBLP9Aeq5wG6PRgQzFpH2G3pcmH9t1kxJ36dekpCsrLSJ9n3u52OPh
JGBrz7tHeIh3bn+gAZHTe1sQI462VVQrk+RODD/EZSXzx8P0z39rdYiW7RL4YUf4fOYprQtVPctj
axk6ViPMndXfron3HzBhbTv9QQWzP75tBSeUhUNUl3V5+dQOilcHqvLyOtmvbbRic5usP8/EYmgL
HAXv7b86SMhhpykODiACGyhVM12re1cF4eXsOMt1rPikiccflNOuVtvhfr52q96KVzToBJPzZBFS
d5IGw0+/Sj536Fs5XnXq/ATlAY2F2TVRDzZq8wdWkq/cIeRLIPgGExvQCZjkERMoOqgzxt3hDBVZ
yNmtkWvaBpmG7SWWQKIUdEvPANj7UviMsvbtF2bXNvNkjUQhy1i0jTywB5NgolxfaXjlkU6bTy9M
a6AtWyz+PMn2xn15L124EzW9ZOKG0M+k0NAWWRW6WF3cjYOisN6OTsgkdx1Tn0d0Qa/l0Dkqlbbs
aYhIdpgp9P+7w6BUmfD231F83hdFmg1qHHtJlqrEvALk8msew7sHBxAjpr3RTFhVo27ygYygL+iD
r4cK56N+uk/q02mmlnPnK/x4jv1B/wSTkheU3plPrdpGNIQ3dZNrsiIC4R2H24+UoTo3X3zA56p/
6agPGPMh8IIHx3a68Bz3WLffFQXIBWe+AyFMrknw4/ByUN/TZJ+XSy01xsK8GcMUu6KoH4aXerqf
yTIguCbpt8K98ZUB4DD2tHmHnm0EsZ4t4Q5LPicWWL4Y7aAhyLleTACAg88Z5E/kKf4uXqvukWBp
Dz8htPo/zHQm6xzPmt1gKqw+JqH2DYegiBH9ibqZBsctmbZt0V6LFCyXNgRMgvNI26hfM6Hr4zUP
VvwUxHUsDdM718h83qwVKdgkhiT7v73VXeaNiFVnTBKRetpuZAis9a2TsD9OLDcfyJ5JF5+DqDBa
5t8mndCVK9iRzmAFJwijbDLXX6rJiJSZKYQU2benj23vyOdWwKFYgHS9J/9t2CkD0vgEpuV8eMRB
hLI3FI+R9qgKXs6VTX6vj6t++QFVTePWy2lSYbGkgvR7TL8hQHhajaD+w6FICnAqDp4dKoPDokUz
jQ+G4jEVRUrBs0UIBn9+ysbrSKH1K2vcQvQTApAfZmLP7oxxahsmDkajbA6YDNBktZE6m21202iK
9JBir3GVyBtZx4K4zodavOFnDFzQycD7dlSc3Slf+z4o/ota2/fGDYzQoPaIznS2rhMI3efUb3z0
kI9zfFfrw5Qw+LGSgfa+aY0g69PKdCfxwop1Isj8YgykU+UW+sQ5UTwGXIo1rm6NWstvFYO/XPg0
qnNI2rfTCOyMwtoY4uxab7D3rLOQPlQdBsFrYPXU6lUFVFAK4NLfIziM3tn4Z4e/+9W8z3VPYKrf
rFcmjogHG4w4ir7Kq7xOJ0QSdytpHExCq0pzDpPiqXA335u4yT6+rpwmgxSvlHTGYDD2XNYmvChg
UBEs2od2IkJ8D8hhXZ6l32t0AHQiGBPmhp+MN5caKdk07agf/hPCwqlx2p6QBKljFwPdYrtalwoa
Qm8n4NmH9MTbDNJhYyys9iW2mDxbVCnYyT2902vNvQY6EzF4umDWEVXadKesgN9kRO03Hq2cDp+0
vRBiDVjuYhEMFFule/IZELNnEVVkJz/HZCHR8xcMsYrcNXN/AQEV4ID/zV3u2YGKQlwKabVcG4sf
5huvbWfFKp0iYsQUvKD3G238qwLz32rkzJg8etwQOkr9WCffWph9dM42JaPRwyd3VhYpONirC9PF
P1vm6ySX9ODdbuZJJIGcyB4XUPT0lIRbW4tU+1CPHMuXPrKhgUm3uo67LLXEPEeZbWbEBqveuGwg
z7EDmVMssbunzsq3aCkrkXjQA7SO/jyCwge+3fOCWVuGzvQ5dcPq9FAMgtcbK52BVpe0+Khsg/3L
154Hr3qFAPdPPsEVaOkPgAwwslhSe68kel/F9WMFPdLgmn/waP4prVl2rGyJn+PbI1zt3Kh0HLO6
7yVTcyWH72L+JE6/4IuI5MmQk9ldEhpGu3OTANq+V0NHl4VXxxuJJdtNUtnKteStANjh2HL29u5L
z6KOa6nlzb/qXCQ0uGrthiHN7Qner4z/QbOsJ5ljs4Nr9dyvpW84amBjCWm0EB+cB7Mmk/eFZ9Y4
VoN1vvI37ZWodA7Irig4qCOr177Igfc8B899SzSNNefS+2TKvEAxQtl1xxMLt/iTNv3VuolXt/LF
0UtA3iM7VRrWG9Ki/Me1O9KKRnCNM+bWadZCa49hG85H13X7xBTSbLgMxLiIfbHy0AfZA+y7OWdI
yQavdn6hYbsxWw3gaKenYI5HtcBc/OH+9PjBE+tYyYyP3XB8Vvl0FeGjni+V2CWqiq/fL+oAR7Uo
3IkB4D0JDXbxdmJQGxqnbzuLBrlkX1MAJqRSdNX/JVR8J00kZCpSXcB+nSaUCEGl1vBjN/n9Z1Tr
2E80EYtGJpwWKoXfNtcp8CshrJOVkj366ykeDn/+bgsN1/XRf1A0CwxNkn7kZB6NGWJf3cEEZkE+
/iFuugNmVUAdMUIFkucb1L35au/up6AbvgOvRajrdKXRm/xVhxTFtCOtpV8lxAp1d9VrjbaIlteN
3ItyVLKP+BGaH/1yNsfiKgNFccRUr4x65xn8pwFNtzdTFPkv1nmuPVhP8mxCUu0/46bJNDUNfx0H
vvrG0IqPxfq7Pok/WE/tSQ5PdaERvL56Q8NNtqmWqLH+HSl/duXnZY31PCHstlNaR5ccfNOPgQLa
C7kAFOPm8H2IJ5a1zBtNm/Cb+meHS8Kg10nV36hPHYriTpsBN0a4+QimjQWHXCA8iasrwY1TCFeZ
fBws4NyiOxWw2mai95dWEZC7AvRfMB5IsFY3zlO5qd6jfXttNjnIeTBlksAyfJxomBvj4m88nc5c
RxhxET3ghXndKRM+D0ehqRE93KGUKZZRywYjMy5QR94hNrlXSbZEqSoqDsa8N41Hudxqoh+F115U
QmKgkkr9ulMA5tiapUKMe1akRJeOsvF6eEs9MTPtyXsOvwXIUQH/nAj6oPIPpmyrUyC9FYO5U9OS
9vH580fLN6LiEN9IWvlIBTvRqVLEg28IPC+nT4slBkRSx2XBGdlqnI2z2I4O9CtJC9pTcUqRYOLs
njjxtxVny7yfSpAjakAd7FcMFGwflQ0DHKFfYGoN+hSWmH1JvWy3P2MuHsACBUZ88ZSMQo9M3zob
H3MgsjZWmmJd6gDb7GE20vt8spUCm/LpZ89ScRChE5f3zhV1zV5LCSyCUm8A66Nj0sGOGao6m54H
/z/6htkkoZhergJj1vEDop99DY5rJARX/HgY7iGU97SZtTlPQNZK8zfBrqpKvy2uTCyubjxq/rKL
T5x7TMBRaL0Sf2jXYWpQbt/3WIrpSHCy9N63SHUqEeBCXNWmaTc0sGamlbMW9HgfF2oI7lHqwtBM
ML7lgCFuH40ktp3KzCa4Td25SxWzeeJmvgbVuwCY5hmO1O/pg30fkldQDWVTc2eXA6nlvA2wVbVK
Mgd5guqtoAUmNrD+jBcMfcmr5w2HTbii47HK/WJb9lx4KQFytB1AxEdRxuRcOEJLLMlbqPtFxyQw
N2dbi6agfB0MHZgORcUSHO8aoVh3YlxEMvqWU66WE/IrVjuj6wvoB2YaK480MPJYywnH6GVBhcN9
3wBvC1zrct380rGqR6iQYbF+8z3PrjRKvug4ea5U/AfmLrrcZ1C9Z4kH/1S95Na/QHQGD1gQivS3
/TLHCclJFaGxfv9tndHjypzR/36LUDb1UXlw/2eAzLMnV4pXfgNmwHQMV+L8bcZDodXAhA1jREuQ
hWoGI409JMlz42+vluVAXbXG1C3qT8ih8CW7fjWakI31cB8g8kdSfIYD1J5VkWbTnPftBXabWHKp
W8zeyC0C+dFhdSDuqKT8DrrdgyFBtSea1EORBB88Q+vIuy0fWlhvmZpdd2oCBfycOvfnJulrMKJs
CUmeG6a61YpNeCNfUYR7K4E4zK19iW5y2YBaJshTgWOGyRblSJJ9LyT5u2/0iFncNxQ9p7p/BhgH
WOjZOcSZ3aCOdqwxQYzBoTStU96mHRkofJ3HFC9Er4cTdIQg4aB3kgySOJgIfjKcXFVQw/4yKwyZ
MKd4g8A9r4d++Mo2TZm/W+HUSSHsyasqtl5jJ2r1+bpzx/6CWazmk3vltM9mYIf6MY30fKi94BMS
S6gV4dT3yey1nqrGpR7lp0td7I6X1ApeNefwQEP9qKk+6A1F3amv3wrS07ZZYLy5e0RneOXi3RWj
MXmBDNnvVne4Hg1QGRV3IoEU3ALg9a6qparsOoV4Q04s3A/l3g23/Zbr0hAv2Z2s6ZK+aLs8Tb2E
zDEgAdJhvyOBiCSsysGPbn6S5t7XNQXThG5tUrHlKvDEdXtIuQVTbQ927SBHBDX0oA7kR4GXRgoR
XI19KZp6MwJQL+ZyosF2Ro4PzqWO6wWqOB3NCDVqwfTuWaG3I1sIDbYmjYOQhuAhj/OJ/Txs55q5
IuB77DjJeDBFjQ6TwhRtPfCCh5Uh+aqGQtEKpVk7EJt0i+ZByNiJX58/Hdv+1PfDlBbqvoz5GAa1
Poy2WkqhW+4CoSAvOVwC7dh90wDCp9zlpMcW+e0VaNxsy+qyJnKG0TmHqUdyjCGOMvbwFTQkpfMM
+9SFS2kWd02dtYSENATf+PR9Z1lb9yat6KoxSc9z1ddp4+Tw5KjlvmeCswR0OJVyTdeUFQouHGmo
1zQlnoU1KzQGogPpwTqgOpix0YPy7VWN2h1/UdwF7M3OYoSblMtNx7Jrupko1rgh9w9/zrT1zEjO
ya3pdvxG/MOpaxXiY9TtdSBJ7b2LlpE2ACIyAbbuSamtqjs2JVtWClVLTGTtLIRaqHZeB0BdFKGk
r8NhFhHmKo4+ALdQ/uQAO16xuWVbNe5xqn/ru0gL8JwGpmsvAW7K51mhgZluuhKJBgKdgYHvvay3
36yT0Ynetq7e0qmDrny6jCOXfYOlWouVAW/Bm4id8n30vere1GQvavtE7oPVxrLQRIk4wO8MkWgP
WcynmULB7iPCmshbcKMCgLwM6xujVO20ogzy3xn4GuRMbD+pgMbxe4nCTGeBzMArfPVzw2FfUF1k
oHwa0Ow5mS+x9iZRPUESgCX0JuUtHZjm7B2WcsCWgcLnmFHrQPhEEjy9eI9itUyS8vcN9S8Alxrp
+Jwe8WMfUla04bd/R+VlBj8L95mKn8BMGXrdetFqmC0OivNLJtUJi824u/kCSpo8IvcV6zSE7z5f
6gLU1y2OSIfOm7TWnzybrrDwN9M4qZQF+CImWFywwgsv2hDGvFcii8N5Ck+G0G385rnYTYGzvUjm
AaqwXz1ubN0toG3reqkA5opmg7FeV0OBGKU5zfl+Ef8r5WlBw1BKcQNLBCVZz5SU4BzqobDBSgYe
Zf488xA9M/Xxn6F4TQ4hG4wmbgYeVQ50RgEcjTbMDKSxbiz+o4Dx8Lm+jewr9OQsDTWyc3jDu8SU
YAKiYOCulxq6UgHOOmXP/1UtrUv6IeEzf38wpssHIQaAps2bGUMMAv4u2wbd5SLf9nNMWup1I3rd
1R5t4HbfHTeHaRGPgNCcfher7TgsVL+sPg7lc2Rz7RwcwjwPTREEXXv9c9BRTIPvexyzPGmJbKmQ
7NvDN3jlKUIFxYUh6HbsGRYj9ujyW9W4iTTMvan6Ui/HONsfWdqKW1rkhEY2ggzik5rU+BDYFQyl
QATialakjwB8ZGGAloJeFVM0Ix8Y6rKQwd+nb9TabW5bdu5vVzLBMLUqJKocpr9Pext1HiuFJ7LW
txA4C6lgTS5HgtvuXddr11guH2TMD2foZKcsE9dNbEaMHGHrVpgTpdNBDqDx9zI5G/yBbWexQSeJ
/pVfwWrsTXhQz9OjjiaUi8uOO4RarXwkicdxTE8ayY/xswNso3nbn6eWOYMpFUxntuUkNTTC2/0d
iZ2VRewAECMcoGDiFFSr0X5qoxcckPIUqhGQf6MOKEkHYbL8jIyH9rhD9PUDxlblEY6K0VVW1Vbq
wJdf0NzQFa9UTLvQkTkY8IivFqTzt14cp+SIJofN4i7wOzaLJ/liwwdLuu2nKrGdjwaOyUSsrZea
+vkffASuMmicIL86955taVjoeHHH678V10unqYnxnS7d1VzLE0t0/EApca4fKsE6zoW08mi1IraS
Tnoj/R70RLuhFo69fjfzulNegZcITpJCkx8OPMM7SL+QXYl6g4UJucEcyOiNeyYbsVOhzGLNyPyz
2u7JW92CS+iM7ZaPRuueGYIk9lpsoWjdOPHCHyNe9P8AOVhg7OlFQitO1/6e1Ry12LwIKQP0rwR4
S1HydydJZjnVmU0Qsy+CPuJRIsaRcm2EZRCg6tu+umQjcguTHvjKrV0gCA5q9M8y8y4oVQHKMlto
EaETyTsjWp4+h/LL5GHKlosi2ygV+6nKWNU6pSOP/dT22B3BQqgrOGU1hbXoz6KMVEcqZTO8wlVj
BjmvmkZdw7xhjFdlBCVEhYPj4wrc5o/1bbHkFW6E1HwjlQ9GXbqwo/QbL1G+wUlgWWF4UAZUO1eo
K4jVjRJ7rXZZBa+VKcVfFBt/hXpky+7JLZPREoeQmqqarhJ0YH8zAy7Fy5tyBu0IUx87LdaB8tfg
JYD455oItaLd3By9fJxu7OsZmBtgPdVDNcFYF6k6iaO1TA21FCMiaXI3BOfibu7pGT6bCF6CJTve
snoHVnTcG14DBhJjh8eF3ZKjZtjSKd74AiByrueZuyFGEkwySF0b3A2fJws/JqL5xzjxEK8wkcQR
+AHoFvj1G43iQ5Pqv6v6rsC0iM001AMiG0HLD/s2nWzzZZyNL13qjJDhjRiW7FdVlmPmIJXjChPu
gQ7XBFVCyEO63aWLFS0MRx3+5LScjKXHeDO9vIgvh96HJCn+tlfpp2F1gdxnbUD166UkJdW2UtvW
PTosmX1giY3FPsFBEm/Bz4mDdeefCb5olZI+1snBAHmDKa0FL4pQaLJS1wH5Zd7ZiYt0FnPojc58
Z7wPFYJdHyWCuBhktzhyUh3fkOz36Wo/DEyiOYl+g1aGs76cfwqZhJdSujI5SyoV7O541q87npc4
8rLFWjus4+iOd872s56lmOriXdNBLsN06YwCKTPspQXVxYEVyfTmVGzUt61v+nAHujfsQC2ULoFs
YiIcCUi4MlGrVrG9VB6IuqCVojbAPldNKMKH3filjiqxTGTZ8+I/uX4QMG09ro6QxB5f4CrbclQ4
d8dY/jahQvDCe2mf2cSAOp6w+otW8f6iWkmPzEbxguIR67Y7/5bZdNMBoZFoThE3iDWcGOnUVuT3
0OosNJHJlmCtXeJ8SP/HVytgn1zKM42XRRkvsQ22ea4bJwe9NxqzkhEtuyfe4hzkvAMSP49nBtzw
wP824eO6zp4pMQBkW+xORyqhl8KlBxQWhyvKEEVM0jB/ogDo6LogFKlE1lOR0spVhv/JvRbkY7Cf
aZJ7xagDKuhbrhhYK6miSixBGsHTyuSZ3SLFYa+Be0WbLS5hSWsjv9L5ClnFYg4/x7nyXGWoJjUx
xYK6HQj/UHfccdeMf2C8+rrLxk+kXZ/2VlJC7JlE6tbhhFPGumdPMDqNp+iSrKN0S/Gq1gmql/jc
jallKgupm168p+WC1nx6+2M8heRdobo8qMwg+BcJ6AMq+mIt78ccwFAhX7Fv2ypktumFS2UACrCv
dIxsDU5L26inB4NhnoZ1fADhFSwz/exj/WYqqqSg31+4urPyMJz9crGEdvY0HMGYaWINeun84WnD
gIPVWKoqFdiK7XNi/i0t/nMysCIklLHvTvaDp2XoLDt6fwyNb7CHgHCkQqy/9zrMJZOb7AAwcvxo
JZuH1CwQ9hKheDCidz4zg/luLpCY+LvfTc0X+qTT2WNXUTDSsLWBR7kvWD1jzfsFbFFo6/iR4ZGX
rQ9lRbyiAegEs7cuuNrxi6AUJ8ZwkiAV/T1lZ2WJiKFGyljKJxBRDR6HXwIKMohrV16D/YoOldKx
d08wTOQowmNgEb4Plwp+D1EJmMRXm5Tnzf5MpgnGKU1WO7HfwPo3VCHXVHi1ruHPzL1aZPyECNZP
EY63lfdusd/YQp7wqU6LlPp5AkX2n9TjuNcL+KRcOHlxRqgwm5fBrLh6hs0maiq/7H6pf2pAn8Y0
xPaNLDR9uAw+/sLj+Tl3nnFNVF73ssYytBWNpeZKyuHJn9FP4kYdBE56oPsQUAkVL2ZaySjWlAH0
MWpeqVXTBWK1E4t+xtJI1LD6Y4q6MuklwxobhmavC/5NK/Yri9rPne9SP8wyeSgedJcoPfkegyoO
aaVk7d+kS39/FfB5leuph2BYAnadopJTLslT+v2uAT7AzC+nPcloqOWz5+JXXFhgyieS2SktcUl4
fTKUczOTazF7Ndg+Qph3T1X2BWwqScip/IC9xR1MUz7b2/D6OWdBiWu+4zMTS2cYkbCW/YvEQdjC
3gZ0LeJZTDcVpZhb+pdnNVL5VgWtiptuca4SDq1HHj/4+aaSF9w1XiqyHktn8ApRKQLczQ9pqW+i
Lbyip2vjl9mWOOwsF4jaLfkM0B41giw5hWFCbPXTaIz7vDON9UV3IWmzZlrr0G5GZ2S30LjRm8sH
JFmG/5dwxZvfy4+05gr0sYqAN+90FkXIiWbS4ChmqMkYhry0/UqfA8mg4Ufn3zrNqzRU9rp5i14Z
CSSFFvyYR76EdMJxQTtJg9lB159EhN1JFJPwIJz2bv7h0W/4c8CP7EwLY3O2kIx/ItRE5aX2d+Gi
FgOMJLUF2+vQFknXY3r39f3/0QRZUo1PFjuqmGJ5NOHeL018tLiWwGIVv4Oo8QeVRQhaqeMLU2Yp
7pPhfbv9MXFma857YGVzLIFddYIMA2vLxSs3YsSXRwe1EreArN08FdTWKZNBlznkx11x6bMe96lT
+jOCZ63XvS1f1fnaYAvpTs5utiMsgyUBZu46F4Fw+MjqtdGjFg0xvbjW9aGzo+7Zae2xJlHGgiHz
nBJpr9hQ9CEdb+AHKATxdlk5mUt8sbTnnOWms7fIgYV2Em+syhqsRgzDW9xqivq6YS6qvP+cWKO2
KQxg8QOUkt0AwdmY5ADCj31V5GXdmMTfu1o0yU9ORmtr3Ii6OWLiyVklx+ux1qEmXm3OpoftyrY9
Dukwpv8+pFYn05Q1FODQRiQ9RG9Y/fccSqwJRmKJ25RUrKl4ciNmcU5O4xgLouHXueslPrpqxLps
1751gXYRYRkMlmcfpRF6nsd+SXymMT+iU2w60pfAI5lGGnoF6Jzdiz6JA6YkMOSmHOc7m6CER8Ct
TOte7uUMfT/jlMwa+y0DZbvzRpEY2h1x/FEd40N+Z+pCx73bc4TDG3h1hjQf7k3bwF8wD7QRCF+r
170eGiQIYADzzyuGW0frmmof6ZSwIOJeGArEBSthfvzhSCH+4aXEDEMTt9eoNoELG/5q6/hfI7Tu
kDWRVCof4ebKV++JjWfekwv9pl1iI6AUzt0H8icmu5JLoBmNApKMbmCZhe41VcSpafnPQboDsMgo
VAMcHH07Cni+DtUVdogG0ya1arjVa5PdpzmtkP2KbZ6B3/li6rCvs5/bUtj8wEAmFdvJZYYVvCfg
or/9NNPFSalKNFY9ExdfEbieJojVrOt6uXgfCYq3VizxdmMexDM88IINl/EpUJ7KXDJFuesFpbML
bWGJuzYdqs2xFM+qa539DQx3KPbiE3a9gUGhLVBzI5ROGDkgWU0ZBilJE06JEHlNtm96fchFf1nF
QbKzHWmOo1ZoM8Vyt7iz/xQbQLxCD/3kRJx3okGOb/StS8a/N/11VRtt/b4Ru1eG28FI2rAsy/ZT
ywdFG+t2SRbsXQl0nX6MFtxzr7+j9ZR+rB/5YTLyun0qhvEy309W949VI1EYT+Z8vfducLi9EaEV
KjGxJIcPCkuf/jS/MAOTyK0PCdH9ejixcQyuLj9xcacwjHq0dsige25HigUO7hks01xrzk8xTk1o
JDSjCe2engQacOZ73c1og4r5mrYsysoGKl3p0peSJABUkop7vo1ejfyZyKoxB7pNl7MkTVjNGil6
maBmA/9eJDTQ5L7QScWqGkbc9RtJn3kyZmddEj4JlStDzz5M8UNJ8r3G5s6c1Jror7hLYQPuJl0n
nIrAJKfKQan4prY9UPDcus9HhkuqsxW/PCVNd3lzMHb0OYnkw1tSZ20BisX/8vj0NjJgPlvII+rz
kDjVUC8+oDgk2IYtr+zUT2brd8SCBZnqofwJ2mbJMI4P1SUHPY1Z9fWyELOIWGvwnN4pwjY4HEGn
3Unr34qKjnbFgl31/6sxeWGtwnjoT17WY8XnUU5zoG/7iOAlOFUfrJsIULrVn+qOQ645aMzLdVFV
KNlEM2J2FoIwBo8gT46G8kl/rMjhQtExNzbRZoEkxHcXw9zaZ5u8JX5fLxRDB3QuNZW0XQ2SR8K8
VM4upR/xDfEmx8nWIA0vY4Lz0gXKgUqxVlkd/uKa2mNzehbDY+JbV0++udSN8Ezx3mmgdZC008Wr
lF1mJ9sORSjXn2y6k7/fA6Yf/0KxQZ/0IDzYuIGnIj5BenPKa3gLe2QzTZ8QjSVssITOHacGUkDP
JrfAiJgIsF5Mty3K9sghWhkKKRuIbE0UbxMf4UNpWZn09LmdqVvmOatwP+4BDvGoa1W2/MJ4Tzzq
2p78dzuveYaV6cJ6KRvnAD/g917qT2G02U6u05QdFq+WgCTSMhhwLS6zZ7zo7bBpj+avJUwqOyHd
Gm+Ei+pkcIq/i/Qay8zJHQHCNo3mvla4iEYj4RojNhPnIg0N1/bb1vYYU6W7wdjUqP3b9IrDsYDV
OchM+DgoM/UKL/5CagCUD2UitHKVT5FQqzjdGkLFiZXHn4V+DbeIsuzxOXp1CRRaxpJQa4O85ZPm
F3xmAvuojhPQwWjAGINP2CEQh5Z5UFyLkw10eHdlLxiJT3lZz7X5hi/dzD8sGYvMXW9pCVDdANf2
qC/JYxv8YDDdMGtItLrvMnRmwGPOXfNEgavRTYagjapFyKLEzfP/b+lzjxlPnE99nu1Nr+IkSZSi
AdXfu6GmLmgWe5c44+T6uZP9pX7LaukMt5Pq7ozVwZ5DrK+OxBY0hebj+zCuqW2lpevxeGkfs3zq
dKsncuxQIfFFc9XHeJNcv/s6nK+mL7UXUjjP56ja3XsSM4Kqht30srvW+VFG9Tvxax3lMiBPnyev
jaqzlOgjPu7AVKYqn+T7Dsuhe0ij8nXppY3SgZZ+s9qRX6aqXG3YeKgbM0EbOZ64/8fsSbYdaEAA
xsnXlg/6nmWOqZxMkwaO9iaTxIQBTEOiEUDt/q74rg+A1z8sc8dj+yZYPfTPjh5gBcZJfdiF0+D8
ca+Fieja7OvjqeB8cdtMCNr/TaUZWhaazAgVMciqwck1NE0/yubL7+z7vPEeimpzcbHuC/5tY4we
4L/vwTWGU5kTXFJ4cPVZYJQAV1/PimwQaq+z76YLMR65nrWqMBlt0swKrK7IbzTs+k4h/B3Kn4Gn
5DuiO5dUp7Q9H9k9eao0xNvA19C8azDHXAmybXHnopUydZr7xpSO+j2CquFXgZAlMR1zk+YH+R18
hWj6ysGx4yplMOHlCkg1sVkwoudkIW3VLd5ZcPAvMnjpTQ2X2GLJ1RWP6Vb+S6eXbwSNUXQkAzDf
JMnWgnZXxrC5xdB0rPGfuIVbbsVhA94ldjK7qXj8oeOKirNVKh0EC7/Gp4KILwEj/65VDljSsEho
PziJMlR3rpcHgarCkYLMtsd1i3XmR76Vr4YyC0VGMqmORENx7XELvBCLhM7QErB0X0jPY/39EIC8
BEBEejsWTI1AOeuz63VRbfns/AzOxAPawR68HEcOSd2a/Xr52MyN9ASg48JLFs3am5zpWgLa+2UZ
tRq0fYLBBEEzKnbK9XieFGB/PoVPYodWRBLPNj6tFvA8XyQ8W/bgkfqYDVFuPeRMv3cME5zUljJV
sXY/CuLEtDKnbo9AL6XNg6INQrS+gkIMdATyPC8qIVz49+B26/E3gyPRlDZhc1fA3PJa9Z6uTm1O
S9EzKTx23MTOetiLHM2kHmJRxIycYXZ9j+KbC5bKWzr9zbxZilej3coJdtV5+1ChN5wBN4lrLFcg
Zj7bQIT4LPjkJDQ7455bSYQbiXs7e9wCjNjwpeinkJZeb09L7qYQLcITxVxrvh3SsrIIj626dBd0
jaTDTg+gONJ7BOoaL8cPrc9orGL6P7bYORs4xQz1BKhypYt80K/+phqbm0vTvqixf0PwbmWYs3VW
t9c99y5ScCMAEzWb5xtbtsB4bHpqDynbCIMfMmojmIzP4OUgts4oKTrMD+NUVn+94g9F9tb6c+OR
CDIEikbNptupXHkgjxJiiUmcyAzPjer5eyO5cpT0uUMbvfL0uQMR3gCaBPigVwOvZoCvRoEXRFX3
GIP+rmXhJJYQKqvRkLI9Gjo+JUP4t6pc52TZR2NBdScm5o62mh9YEvE/FS9wc1SV4ivG4FR6s1L3
+KOWMC4p5wtLwWjPyIjQSkaNXggfOOLWoB+5c7KsuhMmz0zMa6HT7iM3egYAlAQwXCK0ASyplbfs
WeUVurhbYRF2rONJj7rHJdW9hPDeT+4WbbAAQ0cLhd+cLGYgRZ7Eol92gKMCdaOd2+81jLchkL+w
9gKrN9Y+/tQRBbuS+foICHPKZm8tHSX2c3om+qkpc4Y5KHLAjYx3/gI4rfKbS9JACk75fVhUJUN4
6f8kD6F9zjfc6ZfNx5o2/hNXbG+TjykdtH+puZwWvmcAw/2MNkLNdrjJeAMKivnElmefiwOz4OFp
95g6AGoAdRsw3UsctAW0cDGpoEWRMME9+A8MSHAOOIWEB7vVV4LEe+Iopph8CAd/dhwzxFDBlw7+
tiPH2Az8Xwm3RMuAoGXpty06cxKOcfrq1CtiSbQTyX16E2GRgW/HCUtAsIu/DuUH4SJydi3JRH6M
IWDHQ6kFMvAh4uC7jomJasrt1PsYJdJg30GCY+gJ9UOSouv53/STF0BYpZtQZ2BQg8KUwQ6N7PDF
HMMZobCbepaMBBTkWnkrUpfhPPoBW2AyVsIBN0dfPksjwFxDEdmoGTSHPLV1CospZaTCxuIPvZ+O
iK5TF08A3IbTmjNFxLP1jp1297Q/LPqIOsO7e4ddFFNRzyEFO8q7VJxpoGHxhu0mNt/dIN/n3E26
z1HJLEH9H6W4r5nikm9BvYYvXBkdwNUcJjD8niWLzWzKQZAzyaP9YDfPAjpxF5QUrhStuxmNkblY
fY8M5Ao3HNFyDTdRyyQ3JW4U4YAAhcXrxojlc87R4x7bbItSNewVJJQaJXnaS53JJllLddFC5Vpq
emTCmsuVIda/UaRiAkO0/NKucIqe/lOIxtBjApp2MFuj1HSDFbuoNH8TX2SZX0FgErExoTyc9Kl9
RP5govCSthLqVyKyQ3ZGpeq0XfgXetnLB7Abe+GngoFOobQEqHm2tEsE5lOgCfRN7RL8Nz4mdUG+
Zze4B2E9bJjN6NJA5/CcPsgeu9bMJiJ15/S2rQhRvBFbJMq4tPMBfreB3phJRXxEvbhRMU2hT+y3
VbEOqQd3H2Zuvvrg+vu9sTHCQJ05SPpQ9vUyDe7S8/60/2z1WjI/Ir3hqw8ziSGLuM9gAW6rNRzA
Vatl4gOTMYS7EZww/0iOd3dgE5bnJw0hnOqMT8wOUML0E4VcHRiAj8rDXzSgBzsOVpA9I7M1SS1H
5PSoCjBgGkuv7BjF7zhFHhnH3tc1Vt1gXPQgHlhnKP8q9brQAIo98q96uORzkxp53sjj2xScZyKD
7eSQkTlb8ZcF1rGRZlg3iofNj4uQsLkC9MxrKAL8xHaWCIfahPo04o1XaZd2/iJE750oRzA4xP6Z
22ju8Jq2oHgbGsyjMzjVBTTnoo+B4X27bfV3rvA+AN9WIy1b6aR7G8713F+4fthm3mb9ncBvgPqL
cjaSOrksS5JkmdTqMbnOy8oPg2EW8tZDEQgWxhZ61OiNC2rVYm94zdXISPR/gqxs7YUr8LX4wDgO
CggOW3zlIxBsNxpcsudz01rISXLzdD3P5U2JmUOQlmk6jCKfhITDbgFxr5Tx8qRUtkZBSUMlLyZ6
EIwqfpVfxK8vv/GbWH1kwN/j0MyCdUTGW64rwn7e7xV2hbgeBlf/4aDgCB6ZF8lezhcRQVjSLegg
q4GUgwTS9Oy2Y+t3KimQRmS4UMt3mY1FdWl6J/BHiMFdo1yJHSUA0wWKdbA40ro2gryUKxFA+Y3a
N+eATDLLDBtbPInpDSa6XcDA/AV0c+TOlVK0fmbn/nD70pHgxf3AcPuhrUHKYtQYCxPIsSNZsjxi
XWJXtvMqh5YttuxZBcNojPBFxnxp/ZQjeuhHD87FeJP8H1hXKjRL/scQF2wP5iyzFDeBlrZGlOfb
9+WpK2eYT3Apmlpwp/coSYLy1pcsYYEzg3VTpv8VdcGYX7z92KEHsyowOiRghsxK3ny727C3HME2
VxOLRIEQ79DBTNZwH7uBSUjcgfFXTQFamHZsQeLgoHi37/bwEFCXQhRLN6wYLZ9DWAhzrD+hB264
1g+p6374B/QsYM0pgva6T73pIVce9x2u/t7tzm+TQUJY6Zc5zFfh5rJk4QlM2tbSm7e52Q1iFVer
5kbfyEIrxMmwuTnLCcW2ehw5zD9f8wbocXBzdoyh8bGqXkgBKtkId5LNElfmmkn/s6QLhdV4f4z2
2n8jme5NQH8J3973rM/tB+r6ob5aJQckwmHGPIqqsIc2N848+SEjS5D4hiLq6JuceuDtigeVo5LO
74FWUJGzJUNhWa0gu0kk/mKpNI7ATG/3A+loT3O0fmAt5AU5D5FmkeCUkqHODaJqLi+iTpDekBxt
pus2gEcv7rg5vded1NdUVeNo1/MCd1mc2fpVMYUW/PJjqzof6E9dTVgC8rjWGTuU6O/9P13j+BeE
ryxIhh8liKDiXTHP1RtFM51Vo0mPcTAAOAQSkUcmNhQ6w/+UMAuB7MqzslofKVdRfwNgZoqJZvMi
IFUxPICgSBOu/FolyDRHqt2Ju4xtC2hdw30PoNJ8Ea+IIN/H+ux1+anKu/wt9uhdNkP3A7OKgJ6Z
xne/dDosMKrUT43lKWbkf8deAkJ41+9K2xS9dKU8DWgH2cz+GJcA/K1SB/qRRRIkq+EXtOtzfWhT
pul2bPA+jIdfiLoOgYLmbDKTG1QYnZmRGST6yuKZBQXotY7IyyzOWNuk9Y4lF0q3e9jVvdqjrNj6
pVyaT+Yh6oXNHX//qwcG/8JAKk3kXNSE9VQ/QcS62U9THaeyv+DXM7P743y3tiOEBJbvX2SQyZ+m
SJoMx+M28U2H+UIv0hN/cPck4f/bkzizSYFrnigV1Ud2h7tGZ1h4ud2Yq0/6YNv3iMr+tBZZ+qSo
TM8OtM7GnMlaLb+TrBoFzR1Bakmq6z6WcSeBPf3OFPMz6T0WslRVizwItGGrAUuL/exsfLAGU/U0
oTxXUZeSBC8T/oif/5pYj1EwPKhQiIX78h6dbNW1ZLbNGlY0dMdjDbMniqRltnhbfZjHHF9wfalg
TOHME/MinFGlWqLQ0SQYFKtgeRYllj33jYm9fmB1WRV1vvog8c/a5JamqR9brLd/y4SwYLj7wnFa
8MYfKKmzjTG4MY6XloJfsDbWfQmZch3PZx0bvWm9ve6QPMQ+4TxRl9+WrhH+SbKNUUkf7itXfkT7
LiRF+0NLoeHO3IxIx80GyS7jCo0sWiZrkxAJsehbKgHuLErHTv88CsBvYgmgqdaQRS9ukrKpNQjo
MpZcA9D+4JDHVv2MF29KR/o/CzlcILj+80d6aVrVVg4ynv+Idok/rvaq6mZ7wRcveELtTNECrKoY
okBC3kBMTOYJLruXyOq2wQGfiyjQh8WNmBvmZN69ZfLjxRVREDA0d4lGXkPbUE7npo/bmPKXaxVH
BHeHfWpaw7MSUfJl/m8PYbfZ+lm9z6wjOdKWlY16DyetxkpUpSpbvDXrQqhqoXxs87ZcDAlElVKk
wpMpVT4Fng0KGdLNNYgN9U5fykM5gMq8kJtqzAkRCCMstJDmu1SCvaX2F0ZZuj97dXvrvLoFhQpQ
YKtDjsuU8a/I0j4zWVV5si3z2MTPV8LuvUoFMgPdtpo9/CBQpODwxrNbqiKX7KPuz91rnv0wpdMy
15VtQRQ3G92DtyuaxVueyz+6LhPuIgPkNoHvrk51H5mVXmusMRhlpPJjOzmnGgnyN+b8THlQCYWF
uyGXSRECR1MxDLSzIs3rGGbwveebihFV1HaYyY1TwljKh4b0wrdXzzYnTDCaV+5QcDtrcozbDGUH
lcr1ho8e0b+z8eUqdTZA28YbY3X3bbLUnhLphcgsN5vhZ2aiQCCR9YJJmWctmtFdUWbVDrS01WKP
nHLyvjyyBZKnBO6AC4a9QsK/Wdu48Qww5SM1us4JVsW3LaRSnRkAwDxajt9w461yx5ZVbIQ3C5nX
yNwpKV5sVrTJFy+WgQC6+NFo4H564WM0Fd0JK0mbr0TddL19g1vhFy9ZIm42m439MBYChrTVP+Nr
sy5Dii5nKXJzF8VxUODLYej6wV4IOLa3Ju48VCwb16KNYiR4J4Oju8AA/turaPPZK2fMC22evhFE
PZTn2hBYSJ6s1X9irZcBOn0Ws16nsNkNhPIcMt2vkqe/nycSsvrq0KmgAFiByJy5aWZplglavOSI
ZmokQ7/K0VUAHEgyQD/wgvDGPIiDM3Bhp25J9DrJy1T6I3LJJ48pC9kBJHaYby9V++S3NssodQ+9
Sst/p6L1N4+Os0zH0FWoU8OOxsNRaeJT+EXa/JkCVm/1mrbXh66uRJJYPuVCLgdE9El+5lhNcGlh
7JZm+UfnvHz0s4HZr0VAq3A4yWRm0ymXGyyWxAe33oWuqzow4O0S07nuYgsUCf5v5w94veXboWQ0
b/cLdwz3N2G26Hzu2z+ALg7QG77m8OXgzDqUkdeNfMTmNkLGm81wPkeE23WwuE5yaAiYVqz6dXPi
Q911Y6/hOszS6eveR6v/kp5AoOgdvUY2HHER+KoBkc8wsLylWIy9YBQ9PhoxjrQ3MRie2yuLLSDG
TY3/2ws1g4DSKan1VrJJy03jaLwR59COCPT507164L9wQ/W2Iar4HgQZEwqR90OxBGnRVCv2Vp8Y
wiZ3o5ItmRQsDSu87QLTb1JKQRVvOHow2VTNZVyONWmkjrRqzjdlaumGpiPg4r/enhV8blnOVAuV
nHJ0RzlCwi7t2iRb6UX0rXZfaQ0oqPmxt0JhhpuqDOJLGSZwSLYZKxQjfH2N9DnbhLOyG40qCuHJ
Vi5dX7g5rZKjyNCDn0jzbuDCTX3wbXWk4kg0e7ocor9RtlhT2JJzWp1C7Uir9A58cd+7E74jvld4
6TS/MkPdZyR/X0VwajVUAG2kRi183rYlI7n4BAQt3x/HWbr0Xut8jw0ZI7shteH8l+vUc4uJ3RaT
VtuSBP/9Y7nLfiM2S7RuN1Eo4U3TR1OojZHSwLsbvpS8Ba5cYy28YibOq0+c2YYg7xzhH15rrRG1
s0ymcbH5WVipJmdivuDIANDgad1dQkegQp6EoLFdJa65oXi1XB31/DCZuFwhbAQnwjYIgjEI7oIJ
CHFaAl2u+gYy0npTkVCMgqIIDXtmIQjD5EtX/jg78rVE3YZiMU1k0BO0ho7L1Cguhktxrc8D8As5
pHP+SOonmWqVq0wKaD20cn4KgsuBCK0dR4Ev1az8Tvj+8amFHfse40Ei/TFm3qxEI0RCbpLA7B0p
WwnsABQjD6AnJ6Ihc1QBK2TUnDPM1evndwDpRiET8Fu0GCNya0SsqepgFGTwTVtcgDXXTDkdZ6th
B+hq4B9jqvmvHnHvsix+m+NUWCuR+fRfNgsjccsKF8evC6NX0Qalqq1oFvv5F/+yo3PUdGVTypw9
3THnA8M5NykjYV2kGnfXGHk0BDZc5RWL6coZVOXnL0+YaFWE6dNXlMZ8J9uuJ9Ly1lsXVhvQ9p8t
bhjVmcHCegZRq31NF/OtFh3zO3PWiML3ay539KN85kumG8Dgbi9cZn0s+a5yVgnY96mn8DhqXDbO
TNXqVMxKCjg4zur3vCMgD155imNViq9iEX1trw5K9My1qZERnMJTyfUhtaGPiyvRhvkCzLkcHQps
nzYGvsbaYztm289w3kY3zM0cooVl4LIz/iUi+ZZnM4rIn8p94hOL/V3KXB79FIZuxanZRLUJhHwp
vfjwLjJQiauWZMkQ5BJpKmB/q2U4U+VJJNPSvyQgs9DCde54vwpUXjMLFiMwiYNNoztjhEAtIJSU
chtAU4za8AXiCDmIqv1g++iEOUcNiNCtV7YRLkleETwbJVuCEGrE0tBa0Upk/VeJr5WWjPbCp9Rk
VsVWIVDeLVGyn07mXaeiYITqCsLpYcvTYC5dO/jzIlD/n3chBBUz6y047PjqPRZ63DgZz8qe1wC7
7hWG2KwTZvpoN/+/it8apCLjwerT/3U+BL9AUdlSan75S7Lfhc6k/ylTOKK6W6KQ5pcwIAmdb7jC
Fq0BjhzXY9gstCgwH7HhcJD1ZqgSVOAjMNNFMos2OYrsPvz3Egb1vEjVlC447Wn7Eu1PTR0jvP7p
tRrnzT1ne2koXlrMfS2DlhECe66LnEpNuWq+bV9m9/iRnjmMg1nvE/55SRuAPOKd5GAp/cex3i/A
Lm/Y1+vHyoToSHZN3nCf1fLS81OfKCNSk/+8Y4turP/rU7q0ZSklq8ISCkQoK7zhh77b0PAQJ//D
LHEwWOYaCfskhSSc7bVoxbsvWZ+Oxpuh0LEduymi4k7NEDiegRsZHbIwX27uS/M6a+38r9AHc60w
e+3AmXC5NP4aDSmrOIYSB0syA/cYDzflptOv3pRifrgyEbbQSRSoyvdIlfQQMvhKk5ifS3w79j63
Cc0ZlYdo5B9i6j6FYecL2HX4lUDW1YYWNFYeN74GxmzVzDAHrYIeu6x/HcaVql7781Juw4Ygej+N
nD7ONiUZPFM6Z9QDcpArbkRWVcO9hAw7ESYTNPCAhJqw4YVPtj8JotBENKgA1bdjxmAKGjSNTrJY
4/3q40wcvMhr6Xi5vnz02vx/WrInV9/dsVPJlC0nc6JwVST6QUIeF2HoER/2zSofL22apaxoe2FQ
674PIn6Ktw6oGXXnJRnSDprRwa66eHpjCgj2fzy95MwdYe+Wskun5DW4cltNzdBhYLBUTNdkREMK
aTVIcg5pPdIEPaF0KHDU3Z8O+/LAj6AKgL25i1XoIBkEvX4r9Op0vwCVJ1cww7ECbFM0dUiGHZZP
5n7rlKcErHr2FuyFa4VIUqJdtH4nUsUbusaMBKl2R26VnOrYFEoZ85VoRhXrWX/2IWiWcDkoalF7
O7l1wBn+GyDKRPgEWx971h3Twesxc+KLZCmen0G/Ydnm6B8XzKbJ4jtGePsBSbxsKxisO+ArFQJT
stKKvKhloI2Lamij1H8dxK0hMvRImtmREzeD5QJXkJ2TBiOZx54UP3algBI0ceA/wkT4ExwovXVT
H57uq8/PKBwgp8R/JitxqAG/zX3rBAmgoAsAWxKdOt9I0DKyT8sj1e+QyZGasqIi3F2nfeBZ1zxD
HhxDPEicKWR2Q02c99OyH89GD44Sh17gUsvfJUrjiWErk/KUmT/ec/jK1VDMVn5jiw0huCYABPW4
RxSFqa5m31dAK7zpKfDWBlqVVL49nmWgK7nJRd51fsc50nX2iL8SMC4crJLVB5bmmV1S8i9pQh+Y
5mW1giXjZbqNW6zYQFPZO17C6mIbS/zAb49qT+oMd8PV7KLSMKEX70kdM2HmLXujEQLZKleajN6B
2aVes5fUHxlF++rsvHpcqVDoxx7W50kgp1Rop6zoMXS0BDD4I3UvMSyOUHLRX9OFCadQe4SnmK9Y
Te3dOdfdHSvcS50K9Hq8lkh47XsFGKWexBZ7rahDaBO7HWUfcbSApU5fJ48hhthcmy495g2kh+5J
7AIQG9CEpfIiXLPZXy/ciTMZVr8/eOSKvI6d96q6Ggfj2jHsEO/E0nE4E2DauR9DtKNyE5Krup6H
PxW47m7BB3gSgqyWtdiVuJ5r2Zj1kQXete6nGZuj5jid9D2hhYBOmBzZTAo/DpEuChAaRvAgP5PB
GPYBBxTUdmX2uKfSGPwMhDp+s4snvStxgxpm7Dnn39Jx8okbNyBn54EbaWC5i1Vqx3FzsbQRMqIb
yJUwqz3IWPHG4WxPYFIoHZUqUVdq1tNjRdIdM8tNP3rUZtOFn6HO1/HTh4tKLj9tnT0/O/VTfOln
txtrwjfQUswDzyqRH8pbHdLdWFzYqol4o7h9B1ddx4cwvaZVVxSGMYDollmV14kunopZ6G1cqbZz
BpjRoJoJiZOLVJ94mVTmMU54jPUATJVfisyeHwI5FxWud75W1DtQDLWJ/OD9e9PL7BGB4twaddZq
53gDyPNUgRT9lXUbuk2xQPedbbZ5tEDZal3K12nkfsqlKm59ZqACApIq2B8Ia+B/395k4JrxPjfZ
6iX9kgi7pOweV84+YcgRll8AmbY4GBZd5++cgALxAGlPIEqYZO6wHSv76Bxm/PGbleO5M4QTiqoz
KPN7uLU22cHg6g0UhotZGoPA9UwpLuDf+dmZoEv7GLVTravhTXg/a20dIg4Kpvtar0CzG6wwl6UB
aRSjQaf/6rIz8Yr2uoC0jlIEi7A2CFelKZX+EEavSrGPR4Pxh5pVvKEbBygXB5N+nQOIRZW0McOm
xk+Kmt+4vyHjgS27PPxpMC90QIueaE1hZ20OhbBaU6CtoiunEGbQN24q0LbYSC9nprFlpm+1kY1+
pfiqy8LV5mmhO8+9sT6BsRTM+1zy3kxNNKJ7RJn9xA3nKpZ84A1vOKXpgdIwIXZhWD3RHhBp1etI
uiftryUoYLdwW026NMb59d6tvjMqdxEWVssFpmeiTNcrV5vQpjEt8cVbyWOMabNDMiLhq0wHeEmp
21RHmtuO/Rmuhb7HHLbWh9grVx2+MRVbp0hAHRS6CJQvp6Nc7UeJ4BUNsiw1KcnqDrYEhndmRMSk
jt2OMRrh7Tven2ETMARQ9tuwNh2F7GepiAboKPlfk9H6Oc7qSfALuGWjw+CVnLbsoQqC5ACmSPmV
hrypHDneZah0bWwKNagBTBO6jYey/UymJlbz7Rwn1IPXGyr9XN3POaIjZKM7VvyIV4DinCA4JyE2
U8yGOoYyG2PQJw9LYvMNKwdYkxqa6h5sJTEjTnfwZyiM5m/7spK1/e9md93sFx1yuLEyNprYV77b
3lOlvw81+LiAO6AkTHaau8ebG9hUkZv2Qlcu1g+dsnfIGjEujbvendRc5XaksEqc/xdXpDRCq2fx
Gebzeon0ScC3Lmc3k37vNB847I/fJXCSADCa8uKp6V0Fkrn5rP3yJU6c92aw3w9H8jawrv+vsKz4
C1grDMZZlY3u3/0nHnY1a7L1zBoelapVAZYpCTv4pA3Ju1LsTvD8aAHyfw5EJe6hNO3Sg/K96sM5
INk3AZGrLWnWT47h90wyMeypTw3PzzbZ0MEyQ+nAQpcrE/aElpjwOGMXFysHzteqeNAl2FpIDvXN
b7yCaMJ7lrB/4+2V/HrWf6uSIU7gyPzeBUJIyAIOR521U38gpSzRS7Cv+Dq+BgOCGCTK8KUrbHcd
3mHwL3eB/St8dkoSxcTvs+XIUOozEa7L5CxQLPRg1bAzVBOWd2PDMnDM8R7g7rZgB43zWFTwEGri
pV4tkSgKPA6umNmqzoJq/U0Sa8EzlLtcF2Nsq+xXUcVTy6PnEtLxWDZp+dEBO0pot42jBOxQoOiE
SLgKuM6AXX7twrMQUlbhpWeI79yKuScjBev/2XU+sEcRzn2bi+AO1GqocfBDZNILOHYZxpFN2Ui+
kFDGhx+vTJ/CwihPEosil5JjtrbH0WTFAfa8QeXT9o9wQqmvak8kZu/QHZKL/mAGrJptFs9v9abU
O5fIHnjYKQeg3G8VgurYETWjZFG3n2MbQhY20zvaigEwrGTteHqkvURb9LTSU+qav7ouB+ucRTBG
XXQ/8K0FFSTitOxqpuGHgqdvPD9gMzGlwo4FShZZ+dwE7hl+Db8udeQ20EGbxG0aXbn+JKRqMr4b
Triv4rdMfxM3xcfEVQf8CZj9b1ssYY3v+vTF0s0WkHMop+16iAqsdU77u+jsKX0ZciHZbkCT8W4R
qewld8m+7MMgUzbwCTLLN+/jl8RZw2GidIPGhqUHCjtqApxBXYB4sAtFB4kqtH/s+MLRN4Uhbblc
TzMwaNC5UcrprR3vArNda/sW6Exmc2u2qLQUFjHgmmp6wEw5AyJ3c3viO2KMcO+97SrcF7WfCQRS
0Xcgup2jzEd0JlWzF5nq8MISoXwDJK1+vtvLjpaEePV15vrzE+WltsneRr2Yzb4DDhvnclqfHCMM
Pb+A/o9Y8BjHhbQ0+0C5zkDEo7mMIv7dphfy9o78YDRZyaT2Rl8D30GSGGUui4mOCmmwXOmehEqi
EHQIVA5RwgBSTQN+HnseP4FUtHwBYE+6K/GbnDQS2I+I8TSKVU5m1zRdQT41nJbN4wdE6CvMZWcS
eyVv0Od+S3PEq5Pdc6q9t25v8rvzJZpeNBn2kb1f2EIb5zS0iNaAqktTUMGq9g5F8Ld6SwO8Z6a0
J7gCX+8HY/2LhsA+1UErnWVXB4cJNFbK1qmt/70WeyK1Vq9n6MFWqUodG2IISr8C3+OQO/bW0sY7
aX8+2BxK+4zumrJKagVSBNdTZHQDP/DFMZ1MrePCLT6eBVWhBdsIqCKPXe/OQrdF7caJmsith3Rb
M8zP3QjFCmPyKsm5TjKF5xBemVz4G7SfyAjtpGqLuY8mEOoW+XkqiCvh3l9ZBllChxNST/lH57DF
YtEIB9P8aodFBOIicgLGkxAGYEbXXHyB9wd97AIvm2LxoLQq96fk3YDU7xupNstrDVYsifE8FDmg
ZiIJh25HMrNp/3iKqUqSMPYsDctMue7WsWYfXH2L6zumU3YEaYXjVto+Q+lNYerwG/fcIk9vH571
pDa6I47khXNLoBP4rD7QbBB+vIui3VyKmAtHyKvBHPpKeiKsWq48A++7LodWVeyppfISG6mdoTyK
bbdS5y0ITsycN2aneLC6GPTPlM6CgS+3ZSD7J3zA3EJPj7sVzoHJB4cMo3Qj8110azXTnWvHIQNJ
2odjgo38HOPdbS4n5xEJulcVyQALiJ+3V1gawYPQC9gCFfDxB8OvnTiy96U06L9LBCW/civ/31x8
Q1EDooBLrlnj3SOrMhviXuFkFKq5l2lmCsSZI7gC27TIeZFMM6JIwwNsS5cJX/CcYadhXJxwQMts
d2sJ+GKTPCMN4s+7Ijfv0chSb5QwkukEQ1W5I0gN3dH3NSxGKQ/JKqnR63Yrg0M3EkUeGtI3K+jA
GHfFxQei1f1uYAGRLB5H2XZJKr8mQ1ALb7wiMeKpIMmZ1eIyrcDe2/PJVBcx2MF80r4wj2WhmzHf
skiMqE8YMXOHu4rA1VKTAIstZzQo/VB2+Q4JGFQ9v41JuMPsxBjMxr5nHeE8h9qsEDyntJ/u3bPL
280V1JumKRs8li8gsfgWxNYY9NZ+HisUjfFlu2VSwA8pUjLu57fqG/EhX7C01+guFjhbA4Luh5NZ
+FC+c0NTTlPE4nsnooaVoYxIAoWFexFS4rPaZUv3mzklXG+E3KZP2d9N4VJHr/s9GQUjSCHVpPgq
LACvOQlGgYiArz3+8gdH0RL+7HWrQ3cx13Nd9ZG/y+GG3lxv4ogpzUrQ2g7VgEwa/Ym+6PTCYfeq
fFu0wIju+jA/fZNEDeoeQqI5xaCOdENMHijs0VZlL6G2khz4FFib+f1TbluA1nrqgLPbKCVF0zXY
W+Vla3zDCTU5A0rQdEcEdsEr4EwR9a+gZfWjvjhknV41p1lJ4VLf5aP5Oio6VImsuk20Rp/YJT59
jO0NZvfAnQk1Wmb4HsMIw6b9UuFCHnXTBogo0Bat9/DQAHPNmH/oKYtzpqA0R4W2A6Z/nZuUPk4k
kzP89p2gA79RKF8dQKC/um5WXX+iXtJ6GAAKJ82FYzy9zKzwbjdA74X4d3xUZGPqcnrdQuamMrQ3
spsewN6KkmT1YLcokK1am8soDyFZDwJdYf/KHaUmOBIofLnOaTPiTiSlDyDsw45Xq24sL6cNygWs
mR6pPQhkXZWEG8ZJJKLCseIp588ZiT0XJrsVu8ujNPr8xaAnrqOWqK2Gei+W8Da/+txWFlvHCXe1
VCGQVULyKxi77oUq7iu6XDijBfnPhC0EALHuVHkWnzbEkE5K7xINvmkA5qn24ejDFLkwE6NfWscm
BxHSzEAwqwPozEXQgZrJ/9M2mDI+ACuzigUl8GcqLvEcBIYlAEiAs1WZJiATL4sQ8rQzFjoPMOy6
XuzffEtHG5Eo5V1i9AHDeXo2jR1WxpJOR5bCF9quZ+Pda4+XGTIXKLHGf9tUXyUsuqFvAQY2UkFw
+ZfUH87enPwOKa9pEIx5tX4lavXVaq1L0oJcGdJ178Qa52D4D8bd0NhWwpGLOlJwUpc4PYtEHXSJ
Th9esoK8lEn0/tiR0J6tVeNmJzQWq+Nb5NKLXtpwuMd+2rR4HAT6jvm2IBul7QXm5hxl9FuGkqRG
cPFkxFjB5zc6LZCdTxaCz4Fvrwvr/O8k2S5jbPJUl8kwxHTHu9BkHF2jIVYvuVpNAlwkw7gru2k2
/Ose2F3pP97Q0N9XLoTWAliSzJCGOioxI7oBBp3XviEIGHlP8TDw7Uuk29Wrv/E0/zHluvCZMtxB
8g8kbxS4xjaHns2PPkRYYXSikYJDXC+iq5N89cqwPHeii4hkvsvli8tPXwSW1i7V41BIJOh2MJNx
1LqXoeerEQVytkZZo9JGNjxJcgWTMMdpiCxoUKeKpIqvC/7PGryCLDxvxgFpn1hxQmNsFbdw7abA
V2CUeYluHII5RjLKnEbMJG3KWQJf8tODLLs3Y+g6NfivpB2XM2sns8+2MZRXS8P7QpL4Z98JYS3u
cKhkLMMCXYTRwOaEaRBUgHoLNYR8ZkXZzsCMwmSW0v9fXQIImL/+Nc5F+JvOm3CDJTATZE7XOoS6
OcVXrrkbrbFRJA2aUTVKw7fDq2hDlHjsqpzW+pdA8qYqVsbmzlOx761E//wU28aAC2GKzJ8dglVs
q7goSjMoFkUPm/ujQGngeLmpGXHTA46lmW6IJw1Gwrpgpucr6HFOdsfXkcZYnDpsYlXGhZJVX2jF
mNwbS6WF19MFnNU0UtyRa+EycLNLIBWYdtC5wflST10vfthpiKSuAwcGlHbSZvEOh8cTTpv6aii9
QvpmtL1UQWSfPO0Sw/WDsIaXXEe3WCT0yiLGts4NXBOD0Q0WTvxymJlkNRMU+jOK/kUs1QPVeW3+
RSpmb1caFFSnonEuHU3B5ALzJpL/HT3digjwHHgg3Yeg6UVXikLdVOrp8AP8ZRWP30zBiVvd1KT3
23SdsU4CS9HzbwPYj9DOsYaBixJroPmDuEz72qvIl58EtCsSY6MDLrXqNsYm0ELwNi26l/a2C74r
xX8I6FJB3Ve+Hg5Q+37AHBJAGocqEH16M04sXsFh79xYAb8tlHZ8pBf7Ru4GHokmTHTnpKT8Pe9T
dV1KIV5c04ThE+JP7b8IChgCxyz145FmqLLhMBcE8cRa5RBhuEJdWAaLS7JeOlW8OAmqZgiZTCaq
Ptc/sYqsqaOPiHDpspB3/81ia3RvX7hhHJSyZZ/FkxKShKxznmxSIQcr/EoMhpY/KGmJ+QF37qmX
SR9de3x6mYw8WYFpIFa8JMjtGk492M9BlG6uEYIHEB7wMdyGK30C94sJyBF6lcViSIPZlLi13HH0
RkNtBBjlhFetnpVhT47BNCfedAgs8HNk+vvAYpKtzBNjv3o4XKpdx8Awp0zzUfYXmMdJpNX1MEcn
9TSjjpJpMDXjQEDazuzgzmLdvIouJ9GIDT4lhS4tGnExFFVvzIlyiKO8QV3OteqoAdPA2xOl7ZMN
3j7I4v37xNdDXIb5nU56CBCsBggmCQws2QEiQKCzOlxZQkKAQov3vFUwFegxiCk52TItuBj4PX0G
T6xuRm5EYbCAC1euu2pSVMob4BH7y+kmZqkqh4uigfLM1jFuHHWSrsQoNSAWufc3DEdySaXDmo9T
QJk7kvDrDZzgnc872g+Z+w4FGNfjp1p6XSHAELLy2SI/iXzsSaBPRMJPobOeJp1QoAifbvjtB4xo
YN/Pbn7IQNnA7ht7BRgv0dJ466D+InHY759jwKBUciwFs2r1LFDTedxmDGMHVuhl8boFOBI9a6oG
sfiFTbyrc9fI5IhNwwxfqZ7Zjzy0zgUOFGX7Y7T4s87rXJ+jTCO8ZZ8GIMFWQo+95tmjgkCOqpVJ
iM8kicmteLNnZDxT0fMxtcEwNOXU5Z2co63L9n7gn3hsK0624q3poyz7w4WmGVmFue5CVE2YZJC0
X/HwzarwTfFaAXUOhsZAaPEAWURceQyFaVy2HAtG3Me0yWae7JRLkFxL0y/3z0ylMGFUjbysm18B
Kiy9qooSlHGqh3zWyEb6x5TRSDJLjp2gB6zUEv8QlA5ArtYYjU7U/88S970qdk7NtyukhtE/DBQq
IjiAvhQTvj/AxGL/kyrDINE2rxZYDewEqCbp6xYYiPjBZAQk8sMddC46wGAiMOdPonD1VO405sEa
RToXYVEADTkM/HRVdRSmFosCJrb0HP0SKQ75IjOiG4MKJCgt7jIyuurZm1zYk71SX4lbDNXD+ROa
vI8qLj/b2rlBU5hn13GBHP7rg3jyPMSuy4JbxEFaFSEC2gj+ya7V9QR77V2H8pmQDDWuf4ZE5M/G
vMN7o/eozrEh3fg+kOVzyR8aIEvASfs8y+EAMxcwXvzPxWmzp5mAyGa25evwtAq+iZaRVpRyfbU1
/6ZpAo6K0HOUt9zgUk/bVMg+KRE1TTPYz9UmqK+n64vZcfz6ZYbHk1eet9w8tiQ4+ddBVMM5a9gn
Lxw+mdVXCpjjBvN+upqqBBpSowg2g3BCfhjOAtLre01twvLEdskPNqZ8Wxi9B7oO/KU2fzIBwc0S
uCiu+LKbDI0STYZOpJTnFoZlPdV8w+37SEhRwkE9sgZ031qHvqxPYeuW5jSV/FM2nbWAB7pyL6Yw
Q9IL/d0EWt+RPZlGfP237xRLsKGrty9N9NHJ3UiKthdyo5q/vcbO8vAUkodDwq233QebN+6yqS0J
1YsexBW6ysLqX2hHpLjsInHPStW4j0r3/TzzcEw4S8yuuAfAEtt+ep8r3PvJcp9th5jQX7YTAcZ4
LrxEA+iKEHeCt9cyMUWMToy1nxNwyuaFmeQQxffMR3/dg5IVl8p3x+fhh6/RriVaxVoKIdB7uciY
m4sCB6fTx+RqR4yIATVIjyUigdviIvN0kCU+qGhWrxfPIl5QZc1OZUmMfJxnIirwhOHcDw9A0Ywl
HworROjFrgRNvHFst3Zf+tNAHzwHBOXa8qZJnxNOt+OrlNMq1xG9/nQkgKfkBgRILGZllKXkEHo3
UxvbMpNP9HLZwixTBK/gImoEjvF3dMwfF+pQDxhq0Jm5qZuFjvHMQaf3saEcFOT9bUfpIluEH+OM
iFHqDTvYXLQ25cgb5YXQwEdWC7IAfPWdHN2y5jDAJsDuuUb8KwT2JvvhVxX0tBSM6lcNbP9GkWuO
kI+2hvB6KUG2dtELgNiCEJjSq4MdEqLrZ6HhYAYknVQqro6nCSzT2uHzZRAQ0ceCXFMsnBpbxZmd
4SIemFcNEy1bW8gINk25qDQpqlkAkbF/mUjHOVfxG6A9leKb3qhohhZJeXkyWH2GIhP6LE1XrbbJ
1GotbyzDp9KTbCnIgef3CkNUPaTZx2D2Le3julNlkLihOrA6SfZlT1RsWjzqyWx7sU32srkUB4HZ
cB4rl3p4C2BUTQYhkzgBvFS2g5dp1iKPrB5nYStxB7e2njQVSjbqPQ6g9eDTD0gUr3J5nZeEW1vX
/gWbVzQxhq781YD9jZtlMU5yK1vLOlmEyksQoB4bsoGl8rOnJBXS9Jmti3TGuo+ChSeUid+Tokgz
2q6BbZCgfid75ZJw0OFcZBhOPXQIoc8gXb9l3b4OSgpDbeYQIOpC6yy+A2zkXXeL1Dpav71gDr9Y
Z52N3qGByt4mVhC7ZZ17WVxHEbKoMuRCJ24geV45Flm+QMuY+PlA3dQPUa28e7EGL5EX3AGBusNW
6RWMp+w1iPY7KpLPkacos+i1yzj+U1saqK9EA66OkzwA6oLAdVkFWlrulpK6X8+ItP9KX5cT6wYI
JFLgZuS4oxznZsu/CvDII1sLlEREbWUB1XBvuw3GqXsZEmc28i0C/6CbI6bmUywGU5EJ1VH4+9GC
o+om6tWG3xCQRRqFZEQa11zqYyvRvtXzRbGuq7ANgIqC+mX7O9sVTVKlju/OQm9XLUYs3nfbyzvt
MnoAZuAOta0qv1YpYQVAlewyadkia9k86B2h3mjhYkMRUFiuAik5koSla1Mn0wpspUuEu+y6UZGE
ZT6SYDDp8DD5ZJpLD89/T8O3xW0CGmbgiDLRsCUqpKU/nr6QXkW9tjGNtNXEPHSJmTd2IbWBZPod
+pmoxbfKoBSkEOOlhuzIqIeW9QjGj6O/XeYEg9q8yBPt6LYlbAPWA86dSqFR0MT3F05xwWgsbO4S
hmwSv5iLOG2r1tqF5FwNOmtqC7Qgr9lopu6UbXsAWULwUKfF2yt5CpVMOGFTA/W4ScF/9GMGsGgl
L6ZVoipRxV5/bDg3BLMv3qw3Ct2XXPsGD7qwhUEM6Bd/BYN2V/VdQ3pcTA1QN2r2WnWd0sWz2p9D
TkS3z5Ts/CKavu5Jc/wgaocVmXocSTSKgCyOGiWbx0LmMDlJW+1HAKMhO8prYG93K2Omv2vSBjU9
aID1KNqf5bBUvFDT8Mw3CDGmJOM/54qRvaq/lGz3RfddShFFVA1XVRRIOc4dWVF0Z0JOC2oF35as
jIQ555wiFn+ZDJYUU0adg3HbhTXT+TGIWqSGIBl1vmqIlMZ6ocrnlIjaUG+W1lEUSCwg4k2Sv9IC
XrcONZI8rMr3v5x19XCbXQRMRtPf3zNTRQYjbrtdkOwhEkXwMZJMomuu2/bERspDCBci82fqKZhb
dnz8xKwpail0y5j415LMAEb5AlIWjQlOgolOnnCDjLKYMgabNQ5yzOFboeozdHgHHMMuRwW3hSNU
30jnP8xikekq8Ir56s4Y8YOoawuVR+cLX7hOLCU/NQpBhnFZ5/8whNTJGMriCSqxLWITjJwtv/D4
n5JvCoyfdzLDxmBX6mvzIjFeR+N5umryL3o3eTYx3TQkC/yqUjD6OKJCQG1/Nm/cu05MUhu1ug9E
UKP/jJYeP3Rp4qwLDiWM1surMh8WY6pkkOMDgJqQgOj0juMU2BD4Cw1Tc7APcjNfXMFr1UOfEDWZ
L0QWik5trk8EXnPxLYmgW62iblKyNosd1krzUfKqFJKezhlk/bo+Bf1LWngVCsvAHf9dh/eEapbX
EZQtoXoDmgBJOLQRYUzP7SliybaZ95q7OnBFNgBlk8OYn4Lyl+eVk1cpx2Di0y1qWZGjBIPyZFgD
GaZISmRKmwvTONAYAfigGGJXbOY7BF09R1RJ/US3OKG7sam9VOCUD8ykAAZxaZvHXaC/w3BFVkIn
0a6UGYg7voj5DHAfAvgRTMucMIXtjozaNcWUfXt4y9PBCUds1Wp1QNxO1JtReFj5UuK5LMaJgXJ7
VB07pbe35pMflMlQq0plcIMguvPD0oiEx7NikUQIgUZwoaDkaeLfeNscZRj2mRM9JWESMfdfocpS
wRM5uYbbuMUh1YgCRGQJj3xZWKe13PGslvYLwRX7TTKshXtd9F9hs4RKmBPLnTQlxDorL9gacr7j
jq2UdwTKX+qaOgOdAkK/DaAnym0t60Yt+jqUruy3z95G4oQZJHZrDaJcJAxwN7uBIDxBoPkYPJUI
eZMfUPNHZEun+ddTiXGxTMRkNoRGt3a3Tq5qRHL7dHj6YaEuHIOc1rNS6fcLWTZj60IfIFcDD2bj
jr1vuVrQXkFU5SygLAgWnq1GPqPBPnVXylCz7bjpFE9S2J0OpzJ6gIoMAUQ+b+h+YeWFr8QErdxi
dljucWsPzGPp8JADeky3pSNwAPY41cNcj7SjUc6GtYgOa1AlIL6772bXMUvLPhmrfV3xKH9mMY1Q
8j6GZdsdQoczoiSZdKAakM/km5MWH6rqERvvdugJ0rMNhhzDLFGi3kdsy5LrdkcqEX+3aFDdEUfc
juNr+yGSFJo/QlrxPEyY/RObBaUM01TEaeFL1kvarUW5QLu7K5oyNv7XyoMRMtToVUEka2s20K10
+IKipgSBJnVBojXrwwM53dt8tsnHo5osHhvofkM9xMbg0kNnDexlTaIZq+9XNYLhcXetxPfAehHC
EU2vVZKFoIIHxddQr9LYzkLT3OsFf6eaVQp+rbENXeFn0pfkNRXF7CtQt5EKUnbdJu8SN1/0lRvG
CL4wZ4fmdFRNsRcm4QdNNZfPayBeNiRQj3iPAGz/q6/ykUkI5dJbOK/yqvYletcc03VoDhmoEIyH
+yFLrPyUaVxbpjYTkOkGekRlTu8qnLmYrszYyeKlCfarvTEYFGGWBcqx0Eq7NUq0rGFr0bmtnT1B
lSsndQgVuEctB6CRtn+0a2hzOSM0TdfQ1nlGevAYbrT2g4swy15n3OgKFMpTj4Tt3aflVg2EMGWO
zAovK7+ihmGhdQ5R/tHYFAG5pbYwIumDV0cCovDfXxfLQ1UEksLPlmh+y9jUmG4raRnoYdAdEJjQ
M46VFpQDzU0nUl28ab3zEgqDYsx5DJ25hH6bI+Gq1Bl5jSAmE/SKnrJqko79mVaKC45zlJn3vOOc
klL2xjow9jo4izrX0dEvH9DjsVQjHdnR0tzjQJ9HpuZqJNWjQRz7QGByhoX681tLrpa54dp/Vf1O
Bd132pBpPbzfHl+Y3w4dkqzHg60gIiZ0Am7HbIGwsEv7LGF81quWO6isgYFxydd1FLiiFKwxYhDO
QBC55UsbQgnq60kXctGclN0XaxMGE4Edb+n31ANkFbhJ00PiBC/HHAK+W83bgv4I75loQOwEEtc6
UPqP4PSj84TuyeA7ZD4cQVDkklQYFDXA6ykjn9Zo4R6SSjdLJC5ljVuG8XvmgTPmrCzFcTXCUOcq
jmePRErQjGyqr+y5N22H5h5tJjfRXmQMCQpNWJYe8hB1zfHcZBoFhrLzgCqGw0PK/sjiMxk8nFY6
zQvA3rWrEP5tU48x/OVH6C7nI0evj38AB5ItbU6CXLpE2otDfqK3/aM3FI41fK3YjAhkyBSdbwsD
0x5NQqqfscTSsiGxfTaZuukNerk4qcE1NmBDBiChShqL44GstLQap28NX3FtZh4PYhHldMOa+efq
MsOXcwup/LOUaMSiQS5jHlc1NcynCM/MWfeY8IcBl1SlsjbbjFWk96AeP7lT9/vICP635wvxGVGC
kyJSefKYZCSLMKFXCdkebcIDbzIa1eDI+p8x9+uojJvBL50/EDzqUEALPUK3Sd9fTCJMPtnNMRCT
GUIIxOunyGak+HmlOiEMAaR1VGTbOKsvUDbKPQdgNayB4oAFdYjPF5tPsMkmOJqA+2x5jMNhxlc7
6XeRC04PhS3HhhH0pByeiaDBCmSVwuFiAafh42LmQgXW9sY9CtBx8/He/X9DYZt1nHl98fojjSTQ
wWs2gIujrMbOZbWFNTZTNx1Y/4puTnGzPt4fIcgW9+Vp1MDY4AGgjuPrtUhkVM7uNa4groH5Tgz6
FbJ5kCEa4rE8Mg7nWkSSompmNJDK5ezrgqii9FunFt5/iUjZlnyEv506MNcSyhHsMbd89vcQRRVW
WAF6Tx1YFsUGRn3Ngb9SBfq6Q+X63wjpNwz1OGcRnI05FCI0v6eHmwADT+dBX0lxzMiUSrCH7cKY
uyU8WpLHfhyyxWD1rtwK1jvIcCSXmUO/nBftbIDYVgTwBIidKlc5bMV3Qd/YPZYivGYdz8rm69yL
kfckflqRW1e8PzZwysffPlZzH2eGlhnANKdLdaWLvTZ1yQFgdoO5PQ5oqq7Gt62ohZwZexsch0vr
Yoz7lg4HUdGo39nyTwhTnFXVthM4D8RJqJmilnxKHOhVLF0ExPTAk341euOhraTxO3S8Z6yPvCWU
gIWIz1Lk6gZ+0/YdENgeT5L9inP1odlpOQzoT7eM/a04z89pumFS5lJSYsLI1N1ZjVUJ6ot60BXo
vWiS7g8sRUpNX/J6V4sdpnr3K0yA9JCHruH6sURi1N7AXZV0tMGSPhYtNNg/EZThlZENkYFSh8dY
qNesXAVNDfrTc3+b2IfYOK7RLPzbKb3KQhRTJLUjpDb1w9D4BGVRhoivjMYy+TCoWqEmLQQ72pK3
o6+t2HU6gw8KnCF59jdhwQnFqxR8RJaMs2MVWjcV5Ao6r81uG4q7CvM61hJEAd7uH9t3I27Np/TB
RXOhQ3MFyopqOHN0EgTXr/zl2KnJWPxMTVZnqsX0ZimZfOB+np2HvVzo+dAgcIl+mMVmB4wUtt4f
AfUtywWiIjrpMtBXdH5wimyExlFWkY0oB+J4Fjm28R+uR4Z2qp7Dg4AD3TDKFyEaaVayjcrVpuAK
apbTWD/qnWu1op/6DUthDsZGQYh4cENROz1ynXixhGlpUZXu8UD5OhDtCZAuWKkI4UdhDJEPABUa
8K6Dtqg8OY3ML7n6s2zQypBZhv2yyIw2eacgCfv1haE2DHK/xA4OW0kBqlV/4Na8+iQdh/50WcMs
xz/2u86g+iGNaJZeLsNFfsBNcXaIdtZd0AhrvfqaFxoVjoTAjb5vgj/49oVKe2lvOUxFO+Q2+NUh
Q+dtQMqMLH7K4z8OjQVgWm2n+dj4Pioot+c4rSi18ymJQjLbG8tl/qY79oMxtjAtN8x9ipXP8Xes
ELCLyvM1JxRuK8K8veug9hAY8fusdIRMRZts4jPV6elelhr4K42A/1hmWJiZin4y7jKd/UaSivYQ
CEkpaKYDkrkqnFDvoTp9TD22VQOmy1clMgH3fkzk3H+Mzadf1uIZTV1EXfK581kH+gLplHSArxqS
eL+nVUdveMX4lf0zk4q2ZbcFfiETLJzkAtnDk9DQoAi7o++MDqlAOCNDrfWY4CU+9Z+ReyYWsqhq
ceB4/sCc83/LHJkd0t9ZPk5y0I3MGQhE2BRfsH8R4yx71D2DvgufdCK9o+f3mawR2TFtp/OM3KUK
q7bBuYomwPOB4QY/pnqm91i+rpqPwkyjTjbP2Mw9TStGS1oQjX+HQMMWc9Ooldk66W/mZkJvbOUO
/ewCy9Ng6geUcfaNv5HAxccYAGZcV2X9YbPKwL/ZN1xnb/mCtQmaZz88Il8ua5ET0qBI1eNYDQtx
oeLUHPaeon1mkfTtItCpVOWKHlqfUPb38LFjqaWRhcSkoRrd3kVH7fSpiNWL0oxpI8d2Wmgcfw3a
aZbDt1GKdA4ahjdOVX2sjQcsQvavJBp4xN4sSZlT8nNjgHDqqYGXBHL5/XOtMxQhHz6NcIvA1u1A
kj9BW7dlfuW94VOY/nLXvlbphx8CHSOcKx/5Qx/8cY3I0LB6LiTCVCP/rGLyvQwroieFqQ7wKWuO
7TaDxs/kFhb5I9fmCxSlj0F139+/CQOUrjls70U88BaHdpKf4UhuHRGWRrVnJzFUGLT1QO6OjwNJ
d+8zWh/+om/l3CHXNGuVoh/4cbHHL+I+Vjbd62c8eUQzvkmsPQw2bk6n3FjvHsyqYiULekhITQpI
C54oYKTYM5HZqeHYHHJABgOXWGzw/mtbBx+EWSigeWxC6xFgMfrdh8Zl/mRTQBUrl41oXMpZUPmD
VGp9VxuSlIbbiGrXo5IJpBubNMT75MVIyK9Q6YenfoWnw4wLsFFy3mxVJMagQ4Pwl8QzmB8xQ0q6
D6awuB/Ifg37o/GBoxfdE7pgg+jvz4kZj+WeFOPQHkB2RuAUbZ0QPWoxHIq9F/7Z+CcSMSYnLi9T
wekDf/jWP8FN6+I7tCKlJTbXVWTR6hpTRPCZPZnWJkujM0IKcSrT/VV+QS0xl+TicG27O5qPMIPG
xp2U8ZuObqVckbZ59OGn1VB7knQwnx2MOC0NjPGcww16FpziJYvhqR4Rv8Lal9JKQukoGAtjEZ7Y
SOHXQxHELhyBIxayqkwQ0ykXJd8IAPvetBzSXfig/Ca9nt1utdxiuLhy911S1oEyPbxXOmYB9BuJ
LTivSsynAU50s6RhgezsjsqBC4ksBWWofwMIThLgMY0VV+72fV3BbFT1IKnkxkfh8+QIH3GcmpdL
6+16aeWcJ+BmYZ3xNe+6yunRQqQ0IMoDit6GtPZeAfmbG2MiL4MnRFly2/VmAzzeu5C0o1sSJe9A
CjF6a7qNbPBIEbuCGnovKoyh58e4uVMI2N2F6cxR6EDkuoHinKJ2zkgxtgJ/eLKz0HNCptxrhBKj
k+F+laNaue46VZ8TTS2OXP3OSOOshKjFnbYjhTxSkKf20ZCl1+IKTxT25hhqXXZMDDSVYooCtWwl
Q3loqzi53gHomxmAled5G4x2v0ZKIYftao4oa4syrP2EF6BNCR9gvtPDXsG3CfHnf1117ycrAdJY
yrYsV2Gzs/CynPT+IlDzlzK7zqQ8JqqzJPQ0mlOmzhOs4SOMKRHP7M1lOLwNhJcCOKLbsqXIT65R
O4k1CLj6hdgBhgRJkHaXDt5e3txWhYFKAwXCOQktOcAVOXHd6c7ugQWNEPxtLtEjvWaJCGqVwfoa
FfixaHRopZD7hGBjmwZ/ulQjWJBePRWRPMLlm8rSeVtW5ImJQgcWjCsyE31Uog6j7SaBonjzt3+K
/p+9E+HYfnYjVZ6O11O+m5q8Oe/DNyi6OKtoEonl+W7bj2JyVtEHc6u2KT0y86a/cxWuIXm/qSFs
s8gWDWTgUVLbOnXjzqcOP+2knY0stv5c+IPzYka1ZwNvYKJ11+7OPqlt3Qt9KDtRqwwsbWu/tkO6
b++T6uSJddgdt1g5BcDSKxiM3GXU7xiV/Eqg9+6DLCzhVjMOMvHMzoTN5ms9TiGXyX6QaPCIxxc0
zjchBMM9L7eB5fnFPAi07gqOKVVYqDPaAcEXnzTTYRREKzszDRlHN692phJSSkRZvJaIXxgvYX7b
282M5WoM1QgOuliAoDWjXHOlnLcm48q5E8jMMsAkxGF5SraJy7O2KixFDBIzF3aSZFTsPZBwZZvp
zGzik/NVobWHS6Ykfk+aa88CeToZa5/sqYNEOhgl5BwPsAQB7atyKbZhmSy8UW73KgxYseunx7kY
90XxCCd99elVUN8zBLok6Ib1tqnD5ybLX+IYx062Pw/8tIn7KrjMocibikaCDpX1T8+IhuErctl4
rKD1LVQedt5bvKEy+D1YvCBxLuGJYt/g/9327nYOrY9xy6KZ0LZuthJjMieZUqoX5701HkGYZZu/
HdlDhPZUwbRo6PesqYGB/aSYI3UfUz4o1xflI3SMJYR4QMXW929HzWIHTfaruPBrONi9zNVfzaCE
89V4gcaq8sRWHyhGa45/u0oz3uS/8eMizq6EX09zvCNStGSseNPGW6qVRyyx6cegARjTBEPMb4U4
WeqmFhIPL+o5O4UMPhAEtH4LvNwrMpdWG9bwwxpkLplajGdTxp3GsG+P43ZclsvQhKxKB4aBKf5L
9JssUxI5SXCW5YbOBSFq+uwQ/TNhXurGbsLI/O4+x41WAHPwJaCTfI2kYOiQ3nNToQlh3ecH7ZQD
Y9bTm/zLbDIq90gMRFwNdYkURLTKdRcjivQBMHzORR7iTBb8yX/5UsVH3162gHlxxzfhxm4KGj/9
3/aQLjvZKUWo/G78Ln6Hs/KJkIM4OUUzBBT08LwwiNowxxF3HZ/V1F87e3kPr4PeMZz/FOEZFWSz
oMaT4ErHdNTCglZqWFdJNF5Rtakxfa/ZWpGljX23gMWbD7kOEWr6Q9Sp7zvzz+A8aAEgOi6bjQmt
rXiqPtgC8GGwFEWLZscPYSSKTj+il685N6O4qA/+w4t3qIKX/dUgHgd5RftXlCfm8E7VFGEhLRYs
ylZ+qS1fZAhansKyrsbnWFMIKDYA3Ltbzh65rzoEao0PcQhHDBKf5l8igNXfWozPIy057iaThL5f
y6659QRDSHzdIqWcEDgNA+ExhOEyar57S7Ye5l2ZvOkaoswyr3VrDBtIO53uvw3MfOZccGFzxSs5
6lKM2DQw3OdLaqAConsIS1uhfWyCfKnc8vBhk2meF72x60vbGt//jPl5pmtqkzl6pUtAAiWKHXRY
iSxLcZwxC2d5TDJqgdVgKOxaHrDIlT6tpXaKzn0hO73vuqtEhM/Y0eL4nBhyugJVvOMmb7gYMHg4
WyOD1Z2Gkz6DY3ufZPxPDRPp/8Htux88X8tjgqGzkW9kjxba5mflnG/gMyZ0EfICRErQUHuvssiC
+Cz5H07mzxSSliu/2zW9U37qctHtZ757ntkM1S24pOeaBDZJhyq5Mryd30IVMGTOyci2e0kpKeEs
PCH0KNBwV1zgz0NUY+UggPr1ONkLl/FTzykxHsr8kKu1I9a2LLMW6CAfzlJTYrLuPxNeNaVJ6EBI
DaR9iFFZdgrd7S6lDpmjThuYZvZJ94vdLRaKbb5x3hlgDAOcQUEfni1lvFsjuI9pG/7qXI4w1QZN
BKxpuiYnAXtJItRapX5vcwPW4Fm1yVbhcKEIt2oN3XUJUkuotCkJhzm1pk1oP8ntPTstGFmmsTuP
oUsnPadtgEuNIiWdWy0aMb9TTCGsksjA2Ofkp88pSJypFRtdJVowfkJQZqkcF7XuKgqfG2eu80Kx
erqAPYvDPi8Iqmfk73l7PSQl6KktbGyGym5YWdYS5mNGRmcCt6eazfoDhaN2ZDW57Fh5ROlUNMKU
TlcvHdZ6lhcp0b3lWZOL+sZ0DUC7RjG3SreoewHSEmRyS/fJqSTHeegBUUdXDWU/id/W/7xmwGAQ
7Tys80jVygIoriSyzQWW50eadf2Wh9DhyZy7c1gnLDZjyM4W2iMyRsAfQoOQmhvPMHJF/NZfZfLa
r13mHLQSNrlcO6YLWLPJxsPn9QhEUjmuDnP73OG8CMFSaxQAaguGv7tp65trHlinwjj3CC5F4m0b
1ovdjMc61XvlhZZ0OSPetQTsdIVKkRiMzfqEcAZb0+TZjDWEDKyf9zuHx1ykFBpj6XVChssCDZ/l
aR5r/EwxY4kmsLVHtB7HC1DHUylBV3oanJh3g9kBDHH5At8DAYdLOxR4GcR9S9F4Pi1yTB806M5x
XSxnlIoAwsRnMG4vxi4+mhfS2cWOEfDuIGbDEMoPTKMnzs2KT68vmELijZCKCyXImFvh8thHTHK1
pPFUp2mOpE5o/HInpAE8zKsAc4Q2csLmaq9xJV+L22ht2Zx2px2w9tJMKSG0gB0hVaTY1hN61aMs
JUwPSiP7a5Ej2fX/4toS41SA8cKo3wlS8yCdT8EXULtxG1UPHyWTjdtZ4Ht0cDBJmsvUb2kq4vdX
NE+ZOWw7vVOcnSzuesLrY/QLxA39B6Bke3Ns76m0pvnCe3mpWHbiVnFTKSFsTqWygbUQH8CGaS6r
hpeTgaXyIBx0u9Pk3Byb4pBbamoxLMLidgFo8hlB+6R5jZAt9oMBSbmT66umkABpqknTpaOBvsoc
iMVxOcIAS97Bw/EDrTiJwBWwx0Fn8d7zyhjq/p7sTpLFOrINkfkNmSGAIeTWUjV0LpSFx60nJfhf
18uXpQtWdtw6UGhiKnjgstl4pDTfolV3eZ9uVyPL4B4bNgtRnjs1UV11gP6a2BNCbe8NHCn7M78y
ZBT9eZvkBDX1TZHWhff0xzzHZ5rMc9ORXlABfNb49NRvV9tKaVkS27AZVKqVAvLZSzljT9X4JxrG
3GGdP4osHLfVZ+zviMffX971TrDTxbflrX5pqA+vJXpTSYQTP/mzhPJ7wffivOAtvxa0zPo6THZT
Ywb6t9YaNGZhH16wFjdPNoatcHlB+imfp9ZjFazXXoIfVg58VnpHyqMrmJT6ZugZEWoQ7Rngizbr
O+uxA2LPlKAjmlcA5CAbXG3zGVW218d0/X3vzlcXgkrCBX6ghzacfPf/lfUo+/9Q8HXjWtqhs/cx
cyk29ayl8ntk/fnDQtOfLVSEgqt5Pi4U+DgkPz+Nh1KwAeaNadniigNdGxPhcWNwRWOrEHdbL+2O
+S4eCMoLqQusRZ2QfjPhGY5vQN/gHg0VFFA1HV3h3NiMvZQDXkuqO6sjVq7GQ2QYTJhXo7fN2c+r
COfLgzDFBZQFqZD9z5S/T62BLfCdY5f8cyueZmOd9vJpjxYr6kpEJM/wMaRyFCblAOWnCb+oToYi
xRW7V/vNidXUqIdbV2NR0N/HCuf/ElX0+dsOC8cOd2LkPlTAnLZ9SoT8Oqjy9Vo5uGTmqekKFWdL
As+9tnzsUR7REiGG0e7xK19yqW4VbUn3sb6hKpEw9QcwyIg/w1QV1dAJLfsOjti8g8RlojrMoe08
UIB/CxC8QaYHnHnrJ4SeVZIF6fC3ayuBAau3utDS8abGxHRyZDIFaGpnTEuFs8jGqnQlizt+KAGD
cd0eJrPhbPVbndiCcbUJJ1e6o9jfghyWntJBNtAwVUMxep0wTpQnHrXZTDLLVjGzY9hlLzPsSpOx
/wbe0Vlgm2QAsMX+PMhkbVAl4Q/xMn3eztHIBio6SERIbxjqI7JsgurpGfDR9KVLXv3a4awrPMhl
U59uOrlwW3rvOkmFwcE11QjJa1Iqu6fNHnZFYjvMTt4LZVXOlBYEuwA28Enrk7JKRE4lidR0t+g4
o6BOfWn92JaipAXOjcKWaGDeU5qMt7kGbOVookd5qqIsuj6KoZa9ls5fLkJssixIVimv4rOIzdvY
w6coESqwKcSu9j49TNPYgzENffSGbsokO3cqVefWJHC2Ay0DvhSyhWbQ5HqAUidd7MPTsJumEUu6
KgYGZ/2YadJbX6Q1Qcoh4jmL36ei6lq1ThSGfsgT16qiupY+/QS+xXrkKNDTgQsrQ0S+oxpno58r
22Okd/MJuYgQS5V0HO33mPRtZa19OXefcyOPwFU8WV23vUqUzffmLaaN7gvjGL0KpxDXixDJNaqn
cBBNY3E8ifFC7/ViGsChpTqzdwcx7Oarg2+7fHbEhS2m7PxCLsq/8KxK9FgemCeqkC8tf9DEcmd/
QoE/vmwGPQAbtnFoStrVvd8kpJRCKySEGnhiYSqhoydbcIbjKyqvt0jVk+0eT4QHQRAM//b5J2F9
/FYnVzdH/aR0wADqw8LazQhbTXuNw2bROXJcxuq6Zn1EiQTuWk9NJQxtm9kIA12gG/5MHE42kmNN
AhLeFv7FM9XnarEMT5LXw6Lnkq905VLY+mNyyjahPFdU50KL+Qrc/ge6nxH7/dUOCvRzzDT1J2m6
d/ecI5M50KDghk8Oo6WxG5uxixQhCslqie6CKJRkuARQi7Hy0cxbgqSle06sU1E/TsJOAKt244oi
F+5eyzcOq61Pk41OO5IN+BOMc6L4CeMIvnP3NnP+r0MG3likDFVaQ3CKzTpQUoLZ+t9EoyD+kIVb
8Gfdhj2zPUe+WILWDw6iw6c+3H3ENXrA4LvICbFIamJcSdF9wJ7LCCPW8FwaApNe3ZDWCjo2llGS
zuDOFYCtJzafZlUM3As6rHiglT+9NHWFqMvP+7U+jaU/qHscbiuaVztvh7uXmKZBMn5kUCfh99dh
owX5D2kHZsLhXP64lsPY0e/9IP1GMxO3CcwA1iZGsQdeRcDuTAFhlp5tKFuHFmMEL77JatP48J33
J0SVIilUTFXLZ6EkoKbyfVTg042QY1/ojW2eReWvBZpgqc6XarJnPTedXQC3Jd8Kk4Ux76stst9C
+6knTeE854PdyrEIbEyPTOEhXgahn2sSXDJ+rGpHDtkZO305hFXi13QNnQSn+c8EhYOx3SOGl7Mx
0g8qRPb/Zv3AjF+DheLyf8uue+zh6jhL4AMNrBePfaYiHb0QYCKcrLXqMuEPskJxjLX6sM5pKwOs
atIGiEoW0l4+y36p5scQx5EdszWtF/yL1RGqxaqr3scpsOPkw32F0JoXssGMKh7PThJ5VbJvKL4x
MRKIgC/LnCj+ZJfHDZ5PsUjOCpMyNYNzO9Xj/fGLUBD8aI/jcPJJITKIWUeW8SKnY29iAciJ2mMh
udVeM9QKLpvZ9QBzlUI1GEqmSRFJVPrq73QFtYPTZmWQA+eF7QfWFDc3vFbV3zaATX0lnsxQvgT8
zqx/JE5A5TTSBG9igwTi7DKUgMlTQbhBxlZr2eAJvQ1zdrJfnbLgtpFRCV66Q41gVXYT9WQK0M0q
2+7zIhYdBSMQ5S0DG05n3uiczmPpeGIPkeV+O2yo8iu2/lT/kMWGmMWuaWuBuqyJ9oLy71ZZaaL2
4ikIQ2XmsL/9AnKGfR93N06h9ZuEliRyt5HPoy6mzstmHrK6g59BSyrP5YvSzhmAXf+TVAE5ov4s
LmLArJJv4xkcENV9wsVxyHF9CaqMpIeK7wRzzr0adbKrwlwP9HVPrWxgCizJNIESVnLfzUGzfxJ/
4uiCjaWJLb7SNFepNSwpdFRB172BBW1dOccx/pc1+C49d9gzJBWAxokJM/lequ8n3ulK6vO4oXzH
7MuxoYpQuO3FEoZZne7wIsvjT3Jr2t+d/2F8bnPJm9Yih9MGkwK5LTqCO4Fs0L0dWQknu1ObvjsR
A1APGoPU/+ArOvz2bUIUPE9qzBvrnXw9teATaysEjv5d7x4CWuYILvUfTCdO2bAJ2MLcsNmJ6E1j
ADvmLv9xM4lUGtdy0LxR72iz9oD+wv0ILOvPms5bK1ASiUeKuUB9Zj/zSkDBI1g0UVs8t26DKUGU
O6S+AzsrstUKr0AJvw49NfCZAEDwWmX74ArlbaasXu5PysPHZ+1MiTZSqsiSUhhzZ/kffQPaD6DY
xOV7012ZaMqZmfSgKukAv8WsZrtG/VlKW20PCaEK9Ox7UPZ0IFg3uKKHN3IQ64Uk83UcDq9eNPJV
pRJZ9Xb2pUYvZlXU0gsO8EtsNF8D8fgHvBjROojGvORq00vYDra/BTYWzZPHZ3gZOY3PcYmPm/Ju
ji6RdZye5/KDOOrcaosbuG0IOPmrIRi63uFwO2t7fvRIJvmYJ7YyRvQho0748/d26AA+cGL5pKZ6
mkthY9lCaLaxaUnDoZRTV6AQS2IweG0rEPGRGaRRNVCmPqnKJHINo23/tJMbQXsVBzVE0Mp3mRYx
SQKmSDfIbylw+9MkF1cM3BNX3ZFaRsOAg8BfZDIKqj8Lo6lBOf61TSOJf/FrvlaV9zXFjsh9Uj5a
YJJ7xNxDwDWmtKJcqOQNS+c9uoHthB+ZVRt4DlbTELlfcVgEDACXxlm8Lkv3NtVp8vmQ2XEOpKdT
yEXbk40hkxK90eGBJxkvS761vzzoL+qCz2xF1R7lGjP9vaPMG86UoMHxvmzCIXpHgmAR3NPxp64v
XQBOwDEB7ZL/OQ1ybbbPDf+cnxKuWDteHukoPpxVMX2hZ8AZPwT3CImRDtVas6Egbqk+QCvY1fkj
8fPKa+bJOFGD2jVgo8j2SMKEZIvPbuM3MjH4VMNKuyfYVhlCEIUJGZURH15G+TjozzJQf6+zh0H+
UqEPZJBfMjxJBdXmicv1UHSr59Iov/+rWWSzxPUyjXdbraLxTcYsiGMJCkOaaLC3h+ZFW8EUA0Z3
8BB73U9tr9yxDPnKzBJjWMEf+LMYATQqIllKKB/h4TlL80hCNgkCGZEWw1cxsK7XeOak/UUMMTr5
pjrJ+hJWYyX62MI8jf3Ogm2nP88RGHraV3P2BrgrxNI0vUMDeX3Bc75vTayzLsjEjZOpsxSuKubF
9wp+eDoFG2tRax0brRz5y/yVE0m0h5Yp4vyXQ8xYo2M18y8fLQqbGCP5zRXJkMVHNKgtKJvsyxms
iZQbbgqYjJaxEZvXmn8U3Ik3HK4M4uNjigo8Y29NrAqOcvDpS7pXx/+rJYoCnouzQhbvTdBFNcCl
QWPPiPxN85B8dafCEL0nlplJy9dSkEREETWuO8EGZYqufc/zVHNVBDAK0F4pgUse+59wZxWunb6x
PLQRXw1tHOupBPNVxjtErqdHfSpOGnxr8R2YbfPyCRiQ4W2pnJzR+J4ExyikDJxi2eJmVUorj/J7
vHq/Ked44WvNC49JOMRVprxyBcZDkfkPyj1x2/P4O6LjEo3moSDxeLD1+DHGvIfsKspZmRDbJb/k
k4J7L//9S3xePIp1btj1vXfVhJH0/Nr9rrTrsUMRZ0dkc27FbMxCKT+GMCF4Ft6j4PIKNhh58Rwm
mNOviaCUPMINYuYPrzyZc8oApvK63GHkys3QT/wiQzs6hZ79SnG8lDaB6hp5drYWXe1bSblOYVFq
I6aJ9z3E3ju/ay8Q/IPVNvk8zK7tsQgcW5ah1le0qrhbrnxtH81T0uUpfyMCYpkFkgsCtL3fU/lK
brg2R1sL59NPWUxI2aaSnpwj3Ch2QTPbgL4rStSAaFPqwlaCFK/6CU5bBC2qGvbPrUr7YznC2oo8
z/ZynihpRbVIMTmjD79k+IXkoYGcjRF4wXS1NWyZ4s2I2UTVdYLkl5ZEekSVLxrVebGsh4GP8/Ib
pLuTveDNNie5+CS+c5mfpLoUQwy8Cd8bU0UObUPXs6dK5PY3YVFhRzbDS4nJlm4HqDBrjrkfObwW
EqsVb93a9fz5q+/IVr1yJud2MyU1KUQnnDQooo2avpokyfn07NiabsuZ0CdhjuCa22G4BIY1ESP3
MauDR9WdBYCd/mfHx38WkPF/AIb6U2iLGjDE8hIxy0pqMwzVeNmQh5RvT9H8lb1il9erEhv9AJYR
l4Gj5Lhv6Ead0nByyswj4NMg4lq+tb9kbcsoBPOQRclo+LXBQig4uTauqdA9D57HGtC6UjsuiZjk
ryvI4jZBjLmtrC5mwTIlR109jaeotk7GaLo1RpzBiE46zNDNRtN6Mi+2MGRDdbR7E2e0gLEj+8IV
PuRkFS3NrZcKwNQiIKca7wFX7+APuQlXMckV+/DnGqLTzbFULo6voxoY+1zHYY9374Oe1oMCHzSm
wNINPS/Fcw/XTfj3JVh7hGPpl9z84SJXhDfa0SX2Vl6ybh6JeIMfGWhAOqYq5KtsQX6U0yV0X5Xw
bzSF2hqLeLQCOVxGWSzwes7hY1RvPNvu/fmUA5jfhYLapnMoN5a7J8yLqDzCJCpx29Mqm0V09Msq
KH1sqX8wAIFdVIbfq8t5R2c2zCPUMxdbmmh/tIc9pdB79GM7wRQNUnBjCwxumESwHUWp1vBBTGcH
L7BACeRR/tqHVz79+D7DOyIkobPhoZd0toTQIzKmIrBOIdTsp2EW31gIFzhvu6gd1VreYHzYUAwq
Po72PYFaFRrRa3a16CYYb3KDig71pHf+k06cMIYguSWcMhInmfSzWChyVp2AAeocqxO+esZF15uo
owMpLqMmKwM3SLXsGlvBYKPO9xW9TfczXNDRM/FRyBx7y5UCt6mVDktu19WX6r97vziYnf96fw2y
TZY4ChVwjWpyvA4UB2eRk/0fmiBdda4naT/kaejq6YuCTF0FjQUFqF+5M3eRoXQHkEGOnTMURL8O
wmbtrlG8+UJBX5NQ/J/4Dp3ZxGXD/1EJKoUetwRdL9+J1fOk8vc5Ktg+tfEzG0v9z8u76pmYpa9y
33V4F91+nXkRcEMUHZkbdWQH4V/xrhML64b30pp83M5J8425V69sM8Q3ZFrWhtGj8QIaVqjpf7kc
X3HOK9eS4AnyOiXGxDvD3TlfY/txmj9tSYjNkDvdFzudDdIF+sQEi1gDjXBCaRkYWfZpGAc8OKRB
zPK69RKbMJ9V3YXHpF4DQu4v27VUsy1diJ9t3S1AaWBiJeg+odanL9Jj3inzZlBV0GYFdMxj5G4M
lkpDgZ8eKN7xJR821j4z1Mwwys/0kEgHbOUHHKjSmoeaDnj1zSpjiqy3pW6nFCuO2hOlovvBv1Ax
j48mJ5mdV05kooLw22Fsy7Ym4aBlUCw7J0DpoqDUEPsRAPGvfJoFgo2XQtiY0SeZQ00anEzDZtYy
30UT4qan1aDEAF1rWAEdEJLloLDFkLrgdTxQ8hZhyc1JbFeF4OAKlJXrflfhT62qTJmTshSul44d
cYYjz4PpTB/DBc05r0BPvYxcdka30IQphBtLBq3r09wSkIdbnIhD1/OmrmJveI2pF8xD1UqAFjaE
LSN4u8Vk86N5UQzQ9VgXIBHRHYxjE5OtFcYo3Vdn9Zwst4enmwN1JPHey9YYUamCERdLpub97hK8
XDgDlhnsoqtl8LchYDD1uHPzOn2Q83/uQv8voSc4hG7QqHrIACK377BdaNZgWTUSBqyLNAp1AnBK
pHBK6uowGGfwbgoYFeF8rWiFFs22NzKes4ToudITtKOQZ1JJAzl6wmkRB4rjLtl+HcWQ7RmiMAV8
eO/mmIvejNP2aQ2J4097zaLCGEMo9gyIYIR2iM0rMj1ii2kaLcbd/+uC1M7vNFatll6cExIwnywL
+Wqm6qTvuTr9YN81c+JxT2DkjyLzvRkDfzGBPhlR07gdT+16ufTkJ8/nIWADW/AGsvUt1y7AQyRe
gZAMHvDcRMuY53LtDx898HetQ9P9c3ojU+v9p5ypEm/h+9dizsqfgxnZf3nvNxpktarFhIxwwKa2
cAKzJmaa0LX6ZGwku5tSdqQYNmSmOcD8OBIIBFUk/8YyO4PoHJWDRe/hMBcCel1QfW2SUAh4NczW
Kd3juELvMuHMShpHuaFEfWIEzJE75Hdj6egMdTBx1OvHXvOT/Keh/FmakrMatImlXpa4dSVUC/SE
WpGFIy+6ztGJgiZCEU5u/Slr6lpHoVOoJRk0xoVEs4A5fEembf9GwOIS3C4D1yGgUlac/0QeuT3i
5shdZZwLjq5/cFq/TLFX/lqiFIITng5eX2XPwNxrB61aw+jFQamxj+RqDOF+GDalElH/eEOtAwpI
O7iEZYRq3lERdKnjHJJEpzbGyWyFvoHnI8l+/7BnFy3g4KhgzbsPHYBr8ew4LiM6iVFbKVO/0MZ/
N0q3rGEPWaJ1ZGexGdZnSjlVMe0ceC+iCxRxR28FKkHnVnUNT9fC01dy6zeC1W1T50Kxy5zIP7Bh
gLsG3jVHxtEJ5pjfgwUZ8PkMR5uUcNz4h36BxCUwaxVoU7xnNuCNwIEbJDaiaHnLJFW6Ld32DMeD
DfqSj+Fn4OgMNmKo+4U29Y9IR6uR1xa7PegHhaeuH5DNzEoj/I1h8pBgVOxlEeJ6p9oH6ZTBIQJH
NwkSSP6LquXpE2zWDGmgCgpt84ocu7LTuF3tSq1aeLmMB7gS8fqoAMHh+b2AGCJeqQbbpX0JnrsF
rl8OTYasmXNAEwVvGcjD9gpM73pGb7xLC47Qx3U6NM1ygVM+5Tdn60+DkW1jwVDWdfc+YiNQUCQi
2s6MQJDtzE7WE/0cZCtjMKoI8owQxxYxHEUyPwT72lOjFN79wYu5pIj9mUjrkkJBrI8wfGD/cRrK
JZHcoD+ylyF3JThRu0YAi7yGWES3TXousc1Xb45P1xNA1eYae8OqIYntxOSr60yNrj8IjVvBWE0Z
seIYVB/BxCcAGc0cAnF0mFwUzDrPoZgIGftkQoQwXZJtQb3Z4buFSFL6IjCMQ4k90+XeESNYgxp0
9kzF1A93YmI63oohueH8aBvzHEElZsX5lLrvTioygqEYK1aK59QWMPE5ELf11W0gTTGMgR6ldK/3
9vxFXOKqSwAgjHXle4znscTRWmHM4fP4zF7cBUAmwJ+zyUtz9pkIsqO5U7s43R05u3nBOwT6a69d
VEEzS1bBJwEuUmv62LYjB5dGBxVuWeP/EDhqlkrfFUdHt92X68DoaYdd34oZ6mNqZkmeyrqTa+Bj
TH9QQTNVoC19ZKjtLQo8ymkyRuEJfu/0tewJdkUAR+WMJ6z16G+Q5gbSRXoMaQ2IBrj28DUTVyMz
M0lKw93Yi5FVZQDmf1MBE24P5mmK6LylocWC1bEX6iDBIKwRSJz+StpBvXpCZAHVJ+t/pZqz7wf6
QsV9gfHP9gTuAIzO9SgNRSpQL7efBEHWiUh4LMwdrcQUchkdNnsUnG/m1C4IYWGdHmEZpQJTxPQo
cwvv6xOLgQ6rSV0paJB1bmGwy34OlmGaGnBCOjMJV7j6iSd/AbdDQ/SXCahc+lhDuKDdisAhU4rW
ApSBd24HPRo/vI6XmDqdHuy51zUV2xvJEYMGq5VxovSZ4cDOydfQ73eSD46RF0tNAkESJ4Ae7IPk
MFy0ekrs+92wNVp0dkla1QT9vmPz3tr5Ib47bDzBHl+Aax2SZg782C2AoDJprm3gWCmK/QehvzaD
EG/5a/gXa0k7D7Ck/GNjjgoH6oGESxTtQ4gP3wqaH0+iLqDrimKGDR8SSmf9V9b0IS8TgaWtoSLP
5MlvFphyLomChUlk23qLBufjvaDIPtAtZf93psAbXxduf8k3gzI1Zk3dFn5s1GA9epZaVwmAFo6I
OfwwOA/ooFh+o/8SZK7ZJ6dMtKYE1vd5BWvaeV88YtDYeNt1Uzj7dmKl28HiXXZ1le2wtPTxNypU
64B3ceQEtdxYH1Ux7Zfg1C8e0f4LCwfGlkdQPN11NKG8sL0at/Qtn2ioVOj+75ZAUirctmmdiHW5
MT6ByZ1C6xFF//uNAD4MEw41eGXa4dWRubBPYHSXpyOvzieWzxYe81WEk46yOGGlZZkd2VjHMf4B
vkykls/ebuSi7er/bT+xUdLv0Qxce/FjBOfvohNLUnc8I0TXzLF84rf8abS/loDrBgTIvp37mD8g
wyv3iwSBi+hz24jjWd8m6L0i/OaEh2V/UlrKhUJf8tFPY5XPMUM+Zr9HU09ebc2KQYENRW1J9s5W
VmtnqwlgspGnFB0oaFddM76sF0EsTvt7a96d+GEuXctGmh+s7+qjpPFfxFPHym1FCs+ouBpeQqal
oxdAmgS/iv4iuitlWxAPeg29QH0kmzbPKLvhTvoE3s5Eqj7l8j96F3OIixmNxwy2qeDjHsvvs05w
4+H7HsvCcGuNHDLGF5OIz1S3W7haCeCWEHyZNCkB+CIyvQ9nVP6kxqd/FdFSO3tn48lw9zD0id/J
jdKqX0Ey3D2l0rk1JMNRjqaJ6AKEIQAEMDseqihMwqpjygzE+ni1pKIk/Lbr/TK5VmqMRBt/FYQ4
1tazmnieJttyROIEwcbIDry6kTdblONyj8sBQ8TgcGRnZgKALUzcSDfWJiOKGy3oTH5lO8yXPl3y
9ySxzDIG71HJKnCUfVfzWip+YlsGIuk7aDg/HSn/a/y2e2CeVt+pM2E8VLQyJloYWtjb8RjOPLHQ
XApgTsOh152H8GGLi0MkQqG4bHVpjEWLuGAcLJdeFQNpiPW3tOTBeWjVNCFSoMjeTs2YSoG9I4QF
7JF8G32hape3q4pXRDwU2+nDMFiXFGGXfvT6Jtljf40aTWRJr5FE7NNiARZj2/6YTVO7AELnAN2/
4wS1LOzy4ub6WOg7iSIoAIFwT6GiBs7YB80zs+/mvK9qj1kp3PG1TG36e2cEbgDZKgBfUEqHAM+j
i1yvq+GLDUibkXxaH5xH2980rJF/svL05KFqDt108wBBzTZAL8EYl2ZJgUF9YPCG3HHzjd53y35j
2w2XtdHNGds/NUwcdpJ3mzFaXwpp8kNS3dDyPR7PRAjwVHhFaq7yMUllKtjtkYHVZqR2dL7NNjlV
tj6PkVVO/vlwzOAcM8hQbDN2MtUbwwGgazO51egYXBcts9gstYX5rK6G2+JbVxqgKxnClzd2Q2SE
+QhiyLEjEZIFxWoBGe/FYznbcyi5clT6Mlq3bWagEn51L9n37mSxB9ckYjmVBHb1uWDwGNF7i2wl
n3T7Dqiskm/lKQmAMw6K3BczBDe2ChJ/UemqEVR3den6MUEtCkg+sG99hWVp9oYD7v898hVq6bht
vo5F5+ERUCTlTJfk0QprcNDUVkwiWHBiFNsyM68EBZ3XCvae1Pgj0Czl+0ZPCMnCIBrs6cGtvlGO
l41OFgig1csT5pza4gaa2iMf5tn8ZjU5n3MMXRiA9UQDvtrKNZ4OLESnB3bdyLzwQA9ZMboC2HC+
uOPF+3ktUaSA3RY/oz45aYzqBRMMC2moJhkME268k3knD6sj0t2j7rSRs3IM9i/8a2whW/iv4tJB
1Z4epnQDsoLjCaxT+vTJ+pjG0dTFG+WkdRqShoxR7Sz4gAqDNsB3rwf78a7ZgpfwUaPG5l6IM4E3
33OY3rcz6bA5yGhZ25J0mUwBHn8aKcqZU/bh4kt/wxQZpzrPKbLKUU9QCm4mCPX6rXsRMsZt0JOe
iBlXU74/nbEUHfc4446v9m1HiElrUva/rz5WKHNfIcvwdfsd/uukzmkBP+LtJZHo72ivEA1tebb3
N7yQZGISaT8dP4pIGsLnH6y9qv88gUpESdo1nS/br1JkViAbJWjeQ9LKd6AX4TV5YpvV8I81CHlD
slq34rhhoXi2rT8ZH+wiv6eewzBiy6/vkKgnrChtKsXlC/o5AJjTnJ05QaDJres7jQxggx7LFDRZ
Zb71NeAbAP/xnGENS2ea2tGd4+qOIgwTdZOYx2efbI+RfgFfus3on4qCeRV5OJvJsbbaQQfCwE3o
Xttczl5reolxHixtJhuW2jfp8fx63fKvpL0Pfvw9l7NOj8TT2DXau/jzKQKJHcFMDUvxs/LxB5wc
JV0v0MOiQZH9cZJjVmPX1GlJtMa2fJzD+7415cqPKfk3V6zK0P/dyMWvwTFvwgn43rdqnM2WJjXJ
CHbDq72RjrNp9qiUStdZeLjz5/+p2zPNdT0imP4hYLOBIzajrwR8hpSnf8yufa3nvJsQUJ1LvXcI
UdakqztFag61DM4B5kcMVzggmLTrM8IVLQFjxQ4wwOCkSrQWN0jRnAnT03dGupjR705UWFjZp8iv
CKstOV5pG8RwDB6IdYe7kKkOPANTQ8QVyjgGmuQkvVJS75MYBAHrRoZjKAfR5hgXiMF3AWAi6quQ
SI1lRiHWl8a7XBAk/kaTAhCnz/rOVeaeZdCBUKrOMDg9z2eVlKD2nLQqXJeQz5tSoDDtTA3q5HcL
nrCjOdYPoILPP6+LPRTm6Uxp9QHMAJaFBevnI1uByIwMQFga2Vpe+gbOB0qH9Spyfw9vpPYc77Ck
QC0oGs/pFRCGAmwLYN5wvgDcx02JWQfGVS3DmQn/4gwkdN54GdMtcU+JxKb9bIcNzsqncgUhGLLs
2P0b8EZgEL4ocA4dhe2+upMNniBhVwC8FPrFBetqIPWhADQJ0wYkgNcyamKGSTvFq0cnp9lzVDlW
mxPqXrtASeaOorbx/bpxgfILTiHFdFPv6y7uYdgfxq1wzn7qhjVd1AZhC/3SqUbYBv1lmI31B7ke
Xp2Hrtt9KQpbp3BC5sn9aw6xZM8m0hZ/eLIvE0yPv5kyrLI5Y49x+Mp27u/gn3jhXxVBG/Bfo2Z3
xSH/7LvgJgHP81fq62t31Q+6GT8pyaJaUXX1NTppafl9PkDWrX99a5gZLCij5HjN1JSrp8asLNSd
tyakrBYe+stW5qRDDTQzZQvovOtfR0gQIn+hcxfa9sxIPqdvmkyPU/XFFSqxBGP6bCr8QB9ETrtg
LpcY9Ejtx1EZaxSJtAUJsPxEsZZ2bcf03Hzu6twk9XOj9gJWb0kXmKxSN8/F9/KIiF9+6X6Koe/F
uFQPOsGygifh9jtat8rzCtvFshUAGAOXaIF6gLWoYO+3A2BGGti98U3W83YftApsX5z2Zeha0+4f
WbkAKfVpNCptlQrV8nSt5A3RxvvhEspKMGjitVebuQFyGcHqEcsnlysJWLMwlkzbQybrLLioaHiZ
63bxgXxWjT7t3KEWWXbMi0UO+4QuVMMtCZkJRxDjMuMa9XF+ykUKxkf2KqTnZ0vtXW2ZpcLYzKVo
EqjdN1P18T+IKO1MuIb+EPVfjqY8E7n94wD3UL/YbtwxkOrxNASio6l7EJEihxtnkNIMnPn/OZnS
50IdUub3uN/oE6ihODARLSGShg2igNR4QLLOm9tYwMBR7s4cFzJBEGVB1cODclD+OsNjmlhK6rGj
hzoH7gRok1hfEJQfb8qiydhe6fXjG1Wx/krZ5XQB6RoOQ+zAB4FcA7YmT7NZqRWLpqww61qooDRT
Hc5Lu9RpIGkBvx7kdgH9Vc9nBzFk8nEo45wxuLAlmF4YIhjYtbE5/EUO7SD/JDQF6ft8+BVMpX8z
yvTz3PQ9OmsH2vvkvPHbalSj2oomnL4zI4/pgxi5dIi+DWLT/1Th93bFbTAA8JZgdlvBmhK+9mi9
AClHLUY7mtv4mA6q3AG8rWE77eP5OBbK4YD8q2D1XeYBxAuGQ9O4gQLZHIZv8Y9oui4xaHbD84aS
4Mmjxxpfm8VLIRWdIMN8vjjZcMSmnlajolLvd9HkT8aaV7FRPpW1sltb+ADOLP5tLh4Ew3JjddOo
sUq0AEe+uVXNzsaBwlU/pA5F58c84npoL6rdTvy4WhxJh1pM7qhZNefPeYfqyl8vIwMpeYnyaiw4
ylj5VY6J0uWC2ebBt/beAKrm0MZydSgL8sbfOMyUbrAGGtAe18VxMijzMJPBDCR83I3OFTZuhtNN
S4YsVD+UEWOfT20zVyU2oRt5eCL4eAjZH305+y+JssEYYPT4zFwe5nFyDfUpCGV2ITFKreOlMAyq
9MrEDCs6Caq9ivUwg/Oh2OR1PrhRcZFWh9KGld4/efyoLJzInc5eEgIhWTQWAkVYPHJCTuK5rgWO
0LGmsJPUGvrgN/jHBrTFSAObVMZ2CNNKA6b9bo7ax4tM8wRdC9ZoEq4YGoEujThHzP5BmJ4y+eG4
+UXIkRmRoNajo39rz9+L3uoZdGyyi0bUCRSyzFlGHlYM4GlGgDs+Cz8tzrIBRIOVzIJgfDeu2fBk
jVb5voyk70mNT9zfKL+7jOxrU97uv0YaBDjdRcrZHC57QurR1qyI4lZQh2LWKpGFGzz6iOhVHaZF
UbfwovTDLZaW76DhdaBQbyiR4rxJjE8YbbD67YeBCQrjynmd0kP5Qo6iaMaCs7tT5rL7P2mogkCO
OXOiveylHTz+6zHpfxdcP1Z5Apv1QhxoKWm2CIJALrhACKeSgIvgIEUqmiJFQGZv9LLTF8WekpJj
jaHQe6jMvhTQhxDbEnMOCY0EYYBChvKBcOxuuLgsgzXlzYVxOFnHR9j2PQoBNiJP0VJ1eekGg5i9
0C7TQfvyHfdd6WjxdnjLZY52t8cud/YFICA2Gj9Cs6oIh06XGNnOX3OssZQUqYUWCxpCYw+9uzIV
EbKAanjXQbWsrv4qiDxbTFWRnYdsVzSlum0FQDs23ThcshAI6QXg2l+aNWZeTM9chAf5t+vuCDqa
Xrdhmbf5KhsKeSbNu5LDk0abe8vqNa8NImqVHjlQa6DQecgv57Gw7C43kbVf8KnlzYbEwARPf2BN
6RwaXAZUCVj3PzWvlpn7NeriaJ8rTbCaxYUYr96Po8D+fZ71dl96qdAWl6CykcY0WJnCPhklG3Yt
/LrlCSvvbT0BCm5wDzZonrv1mwPyrEIDCqJEG47aOxK7ycgnFvPJWQmfF8yrBdzmzDLQPOwmDfVC
qyq1jj5assyKX9Ab0eylX9X2OyRqLvhR/aeLtydgwLKKOGYe1zXgFj4Be5iDfjcF5kcCNEZXz8+O
2hJximFpv5+whcuI51RWM1TlAvsJKlxT6hYczy5VIjwXpFzIayZNobqk/g8kvlQ3FHfm+Eu0RDeb
1sz+RCt4B1AdJ03vzq2p4ZUJZ5FnabndpWpLcdQb9kGpoFY88tTRIgPpsF1TNU2btJHgd0xO4Ey/
zVqo7ir0P++mgJj7nd/Wn5rQigkUNn7GPlP7aIyuMFtUhNX9xxLxYLAY6nw4luGm9RjWZVOTPzGI
vgq8Uy8HzpN9fwB7G8deea2/QtPbBcvAJM6LS874JJ5tb56WT2uVymcdNuCn6Hu3H+9qGx5hoOPE
EKMGNSgwUgbTXim23Qw9JN9lgjyovf2Jz1Wo/ChwC2k1CyFXvQnTNwteq5xRXTbgR0Ks7AgioKz7
XdE2Yaly+JJ7kzQJpU1zzvTsvoju8pWR58+KIabLDrU6WpIeoiMpJfCrcIM6IfGfVEoVMjE8FNuz
CSnBQgDcCCXhjoEjKobx/GiTNixQdFB0ascXS2TUfn97lOtYli8e9xRBlbl2Yuuab6tYtVsscOsM
sv26vYaJmfigUW4ooHGLsc3IpTnFLtyuXTzsoeDzrV7Q6KG3dmB1I5QR5gIAsH0gZXWZJRkJX4Qu
Hvb3dMBz+qKF603cfI01br8k+AzWyUisUUwschtnDbS3gdIWvQSKqMe9cE0W9Ifei0UuQIr0omVb
X7o7Plk63U/Kt2iiBhhwAB0xYH58NwBnlz+71YuNS64sHZwo9JDq2va7VVAZOAvMTfcz2ZuKxH29
6LD8N7p6WqZtc8ZPyF0P7XgsqRVwlNLkAP6wymrE4Ag1STZstAeFhhYAfGE4oAJ/useOXLN8hIOT
lwStxl0RFO6TIPc38KeFip8R+w4fVj0ii6htqZj2h1ntxQw+nwEfIYK9YWliP5dCT6FE9CrPvL06
nDV/kB0tobcmjer0NOZNhzILX1/Ip39DPLcCtexSPmj5pZs3nvS+d4mUwECQ1kf2DS7c2ENnCOFi
VBPsP/9KESF/F5hkyF0T6oKUQSIyGXbHqLDAjdJuE9Yhm8y2xi2lgOTCKa6+XwCtOkKA7wnrMI/H
QgucqsnoJKrrPWSSvsDb6aYGFcGf1MkePlb97eD7mTaA4hE7Dr2PpOg8ofgO8Xtn5NQy8C/KWCxR
ig87QxKppULUXx/exK8W5kSFideaFSNQs8zup3VF2GAyzaN9PgW+9odN0PkD2dLJ2Tq73SsS/zdc
W1OLQsXq8YgT3HKUQhblR5Iq4o5LVHTbS/Kulygyvi+y35INzxGY0mZNGv75NWgFl3vkQkiPkxb6
j6GmROLPXNzG6i8/njfXkT/lr0rnsnzNoOZVU9GUaSCaEGNbObDDHwGVFMinXRKIAuEdM+1Gu+b8
oa3do1rXKm/gmWYjObZAvgAANTAoxcDiYUaP3pufrP5xoCPbkB/eySomWNuT9Eo8i9PBtr7UtuO7
uDtEWW7vsnCTOwnTzjku+IRS6TwbaedvcRSDP2ZJsmTNwRt8ff+mNWJFnab170FKqB9A5rtLzie0
7xDpMd+OSoE/uaOg7UIf15Q0uNhq9hoDoEe+8wK32K+fstFDPphaDKvEvJKjKjUsxPJtPy6PiHEM
pAKFrLEyCoR2cPNNxXX+6L6Mf6IetylV+iZD7Bw9pniCKnqvPOnglhlmHx3khC1gzWAwEcgx0xWy
NgOpbqMIi9bkt8P2HZE4aHWt1ZORzzEkLNr3RwQ/1JSy8NB7js1HjgBPiY91ecEs9k++jq5eJME0
deQoYZABvNyyDdhmxMx015nOF8fqfIiHTCql8AUdkBH0GNUu0IfTH3pk8JHv1HVPtAyYtPnPqu5u
hPAWxcrt9JWQ8GZcPY3RJ2b7HoEnWS70y8k+ak1SoFHcm0bYr3Pj0/5DnZgbx2I1CKuugdxzBwSZ
InpNwEdBrucNlMSc3PVqXY20zB2lJQKeZCRXpnK16ocvbltHmPXbW8zfw82XO57yLUpmPWjcMlG/
aiWxKh7HQB0P5XTGYImYRwUvUplqAj6n64D26eY/xtDW+b0BRn553PXhiZqAZW1zIsdjlDS+4eBC
6jO8eqcP3Y90ci/GW3ywhulgJFlcMPliN7UyklRGGasW+CNApXGtNZ4/NtBJ/NY5EF8qP89njB7L
/EXOBegKzXIpBCXWvh9wjDNYp6P29cseUeaDUaOz/DLLD7S8S1iENToThpjkCsHl9V/+9+tkyhOE
wJNGxa3GYbm2grx+t5aTZedYxP1iDfNHK5CmcWhvc53dQweH3HV63hLqQE3ZC80XnmMFHYv/Ftrf
7n1s4rsphvKkRyAktIjrAFw117zr+uoGVdRN6VzF5CmpcTtgLuJiZx8Sw5aIxKB38Q6ZDxjjwzb8
8Re1ot9Cc99toV2XuMJA0eKbcbZ7E2WOQR/ersiEnTPUwh6kHmKz0PfWD4Sp1Tvz5IZ+UxaSrtS8
KwTf0YqqgKW/av90lFHPVDZV7rbHRfHoNcDdhfdKGboHCYEGPMN6L/kOVWxvMZtS9hA4tMcCQsAm
7+3CKYTjLu9Vo/mLH3iKuFld6WDoLhEq8gUSVjz1hZKz0jAIqZ9FcfZ4maJ9zVb+uoSF+hA5WbEW
XZBEjBo6esYXAwvUcaDCx7vXaShduAu2yfJc79XC3n55qixO07grJCUi1u5hYrY7OOZtk7/m51G7
G9KpnE7psh3leNJtZgB8P/Op2uyCMSoOQl3srsrFdIfa5cCRCYh9IwD9p6Xo1AUzt2+/mtJ+Bgm9
Q0b0RhGAd5CCS9ZVeOq0Su9MSb9Yf94zCUdL9Ulg5cx79RvWQvyXhLbzBf74/3/wP7xrE0cV/fI1
aDMmxgCTZ/Ovf2LKMZzoo7qvjzLNXO/f4N8QoIvsRnoldTJxieIkvye1Emf9yUhmWb/BRFaz/3hc
oqohUiYzhjdUhKDhDVcHMNzIOcwX/c5C5gvIRsW6B0ffjYxSMBv5XrZSugvIOpmo79QZYYAV/Do3
IS7oTsjmgZtme7uwZ+eBCGS0PUYsVRz05XEY/Ht7D1j1sVjWm7j4aKeIG/ZYR1KXF8F5Sis4ONtN
YpenqPFNztZOiiG5yeA0LmUe6MC0jfCTt/BW+qoNI3esRwj2m4HrIAacU1sSHNdq84D7X9qkhZ5/
duxmDE/pgKqe36sQXRfMyfsdcvWVf1bMX+rVrKoKNHgXvaUttV1jNAFeo8AePO2cFGtyyIIh5CZM
dhR10P+ctMnFhIj0+JFrn1PgNDDYWpphY9acTy+gLno7JF3DI5BYLkJGaW22BemFZmWcX28bfUgM
/WrHZwtJO9hIQlHjfmHZajgTNcd2bMjGoMmngaM50LtDynn8HqFLok5dHpm0TQfxC2Ny9Fua5SXd
d7iF3Skho0PLFm5UVH9GRWmJIWAeNoPPKDvHob7SJm5M1RJhTjM31u4fIOWBp+gW9fRqaPRdKRmf
NWsvBTmua0S6MhcTQhO0R9kX3c81e59tI7gunDPz++alWQVcQKYcxGJ8bKOX/dla1EhTUXQQnnMS
tiQURj98E9SiBa3eIj7xiMp73LJpR5irnhLTzUQtlOBWQ/y2rHX4zo/7/k0gPIaOHALRxuXcoW3B
tx93cuefTUdOhoxULoFQPR15iADf8D08rc0gLcU9P/qhD4iWyjcc7s2b0PkMjCdysnlQLrkx1AGU
bO10isOx8ecrbZJGWzLbMJtr3I+MLgHlQCRbkLcG+XsFuJOnUVghhfLykZ0ZX0T/asUlVBRvVXML
zkec78eZaxJMPqFg7H4zvvYBrIxTHjHbf+wyCoNak//bCTB+BPEjFrBgeFMDU27ueKCBWWRZ8iXB
sV7Bh8Z96QY4+boAy5rm4ryG/JOzuQdoIlfrRX/P/vl9pstRpYxoyMIBGU2x289t+nwOIuhsMI1r
oiDj93umnBT1ComcQwRq80fGdoXMPCkXlqLPYFFHuIy4gf6u1Ncv6vxLtbBHx+1myyeNjF6rESX2
TVM6X5Rkm/ilgy72kZGM0wQzOkViPXAc0Khme8/iTkGIvSJsLM5/YpvDqOP8bH4Y1TkZmcMS98+Y
EfIrhyCkfLxXxbj8qKMF3zk93LknIgI8eDkY1o/PbIjU/zD2IkzoR2N1NY2LtJ5VdSG5HJpBiAJA
b9PyR/6KUWlOn8NzRBwt6/pCMbEwbWSgpGTk9C84wosMyrCM0qrB3mRVcHeo0+U2Z5Dn9V/puWDk
n1hKk+kDO6O6K3ilutsSo5OL452bD9ds1kanke0/2bNwupdokSAcqi33A3NMYcyUyhL6GQZAE/kJ
e+PNsdKuVxLFx+sUmqsLo/0c6NKzbVDRYgd7Nt6ZGgB6QlYEEho2knRO0drcPkSf2rJtXGHlWJIV
qK97fZX4zpemUjhzDaggiUjgP9ORwN4YDZRkO2hrNVtNLqT0lM1cizwvQ879ocBhNUOsbOXESVHF
pqUf9lmgfr+uJk1lvMNUNxICkYl8hPQmI6CFycLgJXvNgS+Yire50uNGvipw8k2q35IG35M98Wcs
Xpy8bHHC+xTicFWNUNiBQ5XNfW8Vl4WWKTNUXWSZq60/tlq93ve9jC7mEdR0uMdEvzjSPjbklAhF
OYfC9NdK+pRhFB2ko6Ut2BEL+tMeqL6mHjGENuZ8BZTue1hiiEWsP1HYBwaplnM4i7udWBeQqobL
Mcrd8GmmKGsQowCLy4cC4EvJWSoO+gH3WMr4WRNY1hZOflijkGgQ6gbfDrl9gIyPM+aHuxOK5R2b
AdUi6Pup0E0ucFGltjqdfkEgahI2uowvAfTCNuOiTcXDfhFVQKcihw8amhl6q4QJPnOMf9664Jcq
2LZnbOZGhL/gGlaF8eclvtQHzAmcovdA7msh0fCH8AxHSSDa27HBpRXlSl6sgVLzZ2Y1L+29FAiA
pC/gQop4CGo/xplJLOq2WO3lYmWOJfsZd+SPF7dGxJusBKqpWbn9l3ZXKjJLpy57porHHn2JQ3jt
m73GS7sSXdAfIlOKrX9lcGt//BCUy04xMh/tn9nS8blCSsqGMxaf+8qD0wSRFjX9FF0H06mvS5Ar
aoiTUNmCrAw4lOOY5sOoXuWWVmsvYoD3KQkB7EV+dKmqqq7OAOpeTJqr3ensV4piDVh3YPdMqoF0
enzcpOv/REB4bNdlAg4oArCOTHc+wDAE872JKIYOwu9tifblVIDrWeuFSbDkKdNSTkRkQ0EWiUNT
a77cXRCHZ/+Da63ytyAFgn8RS2uHFbkkzxAGRpsi/VawK+1BR3BBqhjd81I0l5QnnWp7aVRKthDp
7YD/AcSPrSw6NX9cX3vG6G4IUuguG3HwQtDZU13tiHDiHWdv87Cm2PEfI6TR+9l5G7aW5SapErGF
gAGg7ARC12l+yBF1v/XCxCwEULCYis+N2EA9XiRgRaNSoVct6YwHjT/E5BKaGYSQQ6EzQWeop3bu
FT2F3VJyyDGrIr5OlDH8ZJSIQ5q/8G6V/TmNTOAdWSVrwZkoiIe0jUj+7YF5p2+0nWjhcUMjekQP
/9U6IX5Do2/1RsHBGfnUcVGuoX5YW2mdDlBH38mk7/OdkMMZz6hNhb9QEATLWX7dCDuxal63IekB
KEDMB6tG7leM4h8s5jSsgneS282azcMkuWR42ikC3Si31yXqAqNwRr/isB6XDjAo+GJ4XUQzsjGo
Y+WlKCRCi+lFRCgLjx1cdP/8pDHYgGOT624QZo1DLl+fq/F/Ow/ayqxxgO2fwFjPRVPYGpKesH9U
DjoM3lwxV0fJXo2mi3Z8m2ThlVzZZhtOSrebkohTfvcu/ESVV3GcvExe8HAW+hvAYDkWHeyGrtsi
gH8gktRg7/yDBdpdd1KdBhCLuoGDut2eL2g21SfR2Q1EhI+qK14uWlX7cvEfFOZEcJQqkGYESVlh
X2XwNGW56NZ7rWmBWbKqAlprOwzHyWNT7eV9x6oSPc66NFVHuDf0YNxL/33h5WpPPns5MtnRPQr6
dAN2fPkF1u2O6Uw9DB06BxqK/OXYH9aekr2S+E7yjlS71et9F08DuaIVPPCDx8JJjymyGxrRat/H
3Wx3yP+Gl/MzVSVSE2gPrmVxm5r8vXkcXxh5tTPKQyl0eZgE0mn111x6bdTAw2LhSRF7OIAf2zk5
p2Gi/rTJwWQX8a+5DDFL4hEa1y6KO6Z9nE3Pusdhy8J7YXZdgqP/rT/QSmyT8eNgEvPXDf79Blnb
Mtp7tyolIiJC4H6MHj5W6Trvg/8c4Ct1Hk8T0C8OHyShS64zQHv+KEN4McIJnEGnr9mORkbsNtGI
nD223OM3j5oVWzHYud1NfhQb1tzU4qLXNOPmHb3b+CqOSolsRNaxvXrM7jFfzY5BVFYU2ThHuOtX
Rmoq5FAJqT24msDlEmYSoud6pWgGXVW8aL1DK4uCiWUZvhvUDKKIzvMkxGY+2sP5HUj3eNR5e4c3
EEq+itCPLpvI16LqMiTba61133LdvaW3QDIZe7eYKDwdI9UXXDt9TEdEKShc3I7bCwiU3NPAo3az
nArxY3ueNZ8aOS6q+/WAdiJcuYjELhAK29AVZkrjUpc+fRZKYGQC0stPgvYXIcj4+qVW9UiteAWR
Jf4vgq+L7xP30yvRo7MGq93pZOvKlvg1n+3IeE4i43X96rdU/zDy5HrjiCYBKh4QJIuEhFZ0Gzan
K4D1ndRx4Na4n02plHjKN0U2NoyY9g68Ulq5fKRIQVuLnSxER4ziM+DeysFQkmj+VwX75kQk7Dso
NVzt3DR4uuJiAumj52+14uGapLVgK6UXGAHvlaiQMNXJPZxWgkYvLW5w6uSz64pLT29v25TXsfxj
rhRDlHdLDTiphZ+4BWWAYNQNvwFhCHujYu6xuTkVEUKL2ypQAhn/eYAcTDj7BNFW+IqBkBjRiiO3
5aNlqSiw2gajSA/47cCSexWWRah5CdnyTAvfx58FOV86z3aXaNCMT+oJPG63uwF7TUwAQww8q2qG
7X9Y5xiuKmH6wRUPj7jUqDU+vyODiOZfUdA3gwSwe8hd/KR4BYG/vHsz9CgjeqHqSkNiWF5ncTHk
ZKt9H7GhMDUJlU7YOCMY05n0fWzZViXP20ANs2oeNzQro+lmkZ4ABfQpHCOPQ4Z354g63X/a8TA6
ZjIG2DpvrXozDtx1mJrIO+UgFLdOHLUt46wRjWg8LNjlFi7Mwm7rEH1vnQT1hDg/B8vU/SggzO+7
26DPRjcTlKt+7Eh5Xm4hCqrcpzIXONU/AU4+ELl6YY/iu4A+i/iGBKVWMGZ70zm3BpH2QQan2iXt
lA787BgLs0TrHcN8ZFj2b4QjG3hRKs50G0GIKjR1aQ4vkftfYgo2IJYbUjQ1bPeFOIU5fShksE9F
ZIFBBScJDIufzrYAE2AO63m5vL0ZIdZ7taULiG7ffhRZIhK4DO29bVS0bGDIVMf9bELG2NuNWDpj
TBQHBk1poFQSStOGUR6LmvPjWraNmFBhgrJZQsoD8xLPI1/04SjgGAclnzTkoaq1z3yk9Jm8xG64
XGvhqCi7GehqQEHwMioEJ5MHDk+n1sEVI7+hiAGv7JqJ/Arv1BQJFT/7j75zwIiIohqeTne7NLOg
ueAXhpJ9LYjXaSbDzqS8aJY3uY3UZx6pae+SlYCd4kFqtVfUNJJ74u+F8ZKCVLQ86ORHpR9RMfMH
1U7KHmXH4lrjlJmV1u7LCaZS/OxeAPU71d+LFx/EntDXw46hhKt1JJQkXRaNHNxjDC8aFxCS1okp
KJuFaTR7Ozuve5PGeP9FQhYP2nYMWy49MkTog8Mo1LqiisBO3t6P96TTYJ4eCMya2xYguGBGNE64
JSpyBKuYPT1fGPZ5KsUL+QzihJx1YIAgdNQLoydkxmSso9+x6rjAIYbc+sKuoHvHId35dc+vdmYo
6bTwY9qZCf33Qhbi05F6S3+FsirXXowHYwwhsDiDUody/vZVxcwbiUd4+r+dDFSdL3JVlC4kc0Sk
bvyuNALTKgHY+dsIOneuy/JkqzScDcHALUmK4ycbvV/2YywfHpHzatGT8eXuflut8orhvCoSsO3A
dgoZmf4rvbYcU1LZItCVpxAvLGKF9Yv7j6UQS96OSp6hixq8lbfHOwjf7mH8cXfgdiCZavNxGIjp
1xxMcMYFNIKJBM5FP/yaUKw6SH5sTA8sEB/ZayPrZWWX894aryk7lGsXcZetHZr7vAoZTPzYn4ft
N5vllKGA/vHEZZYSM3BTclgmhlo0hpPA3TWD2C0iTwP8doi8Do4P8jwqrqKqFpQHRTnVX/s0Eroc
iaPQfVlF166O9PNzTjoGWMfYI0KN5V4JfAhAcVXIRRb2ZT9iNAwki/WwYMouuCCDOWSYnKvHyoor
oMGiF6wK8jEsmIs6up7KRuTaBJBOQzPFd+4oiU2CPgFN88KHn24x4eXaZbq6OcMMyDG8WIMSQNf4
UXCJYSi3OfeinZibtwCs0gTUM1lI62HtqA7ZHIQ1AOEI3Gfw46Od07a3rNBO/2o4ah/PxtEvNOZQ
DV0brfr36Pg1pVNNYpdoSTB/FXNkP7FN/K4CF4L1pcT82+1Q+3yyA1na2FtjI32GoQMy1jwM9OeC
h/7sQDmD8835pw31UrAii5vja7EoM2a6ijBgksNvo4Aa+vQZ52wcEf8A+943ViwqMmPp89BcXr6P
oN/RW/70PCajOSKmp+NHlaqBbEwQvT+tn8yKkW7Z8vxpgUEJZBegnCe+h1Gb6b7e1FnTgSwcIsk3
7j2KuwkcyUzg/7buWB0nWEBhLA8nQG6Cu9wVva4jZbZFxhGZTCdzzuyJ8YobWmVR/5Ubu2iqTi23
rPkhO4HzcsTWEQlj+pSQuUp9nV+OLG/XV8imhLJtCUpbBwsA4pxatvhJMh91T8GubybcWwyELYaR
6f8F8nlCV+h0bg1D1z0wx1nl/Mh92O4z8b2Ex/QLLH+G6zJfdIngmvknRCTTpwEN4eIMFa76VWcr
BZINAESKuNWS4T4sWV31TevvVY1E9RNSdeQmWnRh96LJHycDXOUFY2if6hfO+5J5UvFguNf21yXG
2N3rsV9o9w+dPgN+8jGGtqJ/2HZMbI5CE03b7O7JitNjkTjsAmftIYT4s0TT6ofmZrntET/1S9rr
a9X/qSujmxhTYrri435Hmkg3PRNpMehVpxB23LR+ebjd2sjaS0OdIcYS5s1gGkFhUFefs8PJa1Bo
xEn8u/OgTT3PmkFl3pK+ATynw7WWWrt9hz/reNSD0Ihn24WBAT+Dj2cqkft51m5swGRZ6KoI6IVP
xkZBCDhTcN+uM9S9RxRtj79qo1I12afBi3InMxIaWmZOjvV3Q6AsL4UItEPwIU4r5hUdMgQpPV0c
C4Riq1Ew1dZkwLe4cTaobk4hRNIeokzirvRbzTUnvklUdiVh/4VTEOOFwNLPWHAsudiiTfR+29SB
ulGM63gR655n4YbWCBmG5+f2C1qWKF1oOZLNOeLmvrbJY0XXYJPRJsRuLIrz8ntQ+409YBitDh3m
DXyA/8ObY4+5Dfyr7jZxFMbhCtHTrjGTaLsQlO6U0aVharcPD8yHSqsYoZWjPXXU3gjiXqRG5Ef4
rB1jP6OI7WY0i+CYu3eon578DQJdXd7KGdqpt22JNUghpyRgn60U5+MSsclWgwn1Tc5ZqbK2zJuE
Va3Ps5ay0l4mmgDH8QblxoZA7yMJ2jB9kdLzomBX8Dr0jeifORGhP+MXAaJpsswaS1tj82FM+ECD
rQp9EgrCykKRA6eHGqTKUeq7JgK7iqUCoJu2cI0aiiCj2xttsRmFeQSCHRDa4y1PPRgPzQziL8FB
kddqQeVWO4p30nick9ROHO9ytSXTRWQYz1i7+F328Be6yPnhLzcQArkvvQ+O3g6n635iUsIZyaOi
bDVcZhJmSG8dWmy0JalKnLx9xmILQHv+lf6WI3sGjGFPTVn39vosSdlVxw8oEuEb59mtQ1H0K1mE
rQXhtO4wRtdYxV4WDShJGBTruYIxtxBu7t1q2l+mJZfwjh0bYUi9J+HoZ5dwQ6uJG7HvfxHo1fFg
zCubXvplyZwyD6+Yu6ryfPMLUTSqccuULHepvMNMSykoIyJSyCO8RqFHDeu/JQI/guZdXz2EE1w9
og3K2qRRBosl0OJXZ+YZwSDqXniq+VlMFM/mtMbr4wwl7hDluKCCbyojXhz32CrEXkCdq5U2d9PZ
WAlPVrVBrBq/fzDDwxZoRNi7RAatCAFDEF9k/4dRH237VVgrhQAx8jL3xTdml7iL2F/Lv5NIfkD9
Q5W8RGVoAhZlBIzzrxpSMf7Q36K5vBl4VBml0r17muZpxSRMDpBOc2vrELGy/yrotx6waKyiTmyk
umuQFfx5E/EJ/fv4SdlD5HDoXfTcvyDEpM1T/xwzQi9tpRcnPaaqwx79z+S2gK7faHt0QjkhMK1j
qeMGwZ+M+PhffmQV1q3ysCduvrab8kxjwAwvdt6uKQY0oZ8HzhFitafULE+izz7FbnbZhBvjExJc
vPtOwUES6j7pB2gb6N3s0F7Y/Ye8ZQF+OV9YpnrZFS2uH2RtUi+aY0FFl3WDFYtfP/7bN8gsttzx
iESfrVBCR4XtlG3dumVv75szYAs17XL0NKXyG/gSrdbY5DmmX+d8SSBsJAF2KBPjhMRSxnD19viB
bOuputJ3HOmPzN+nGFHGFs44ye4wcCONWv+4Bb9DBsOTMYScwgHVEDmofTq9/oFmN7rn5EEFRLsG
qLwHG2e735A/CeOcIRgRMm0WQarKHVwu9OM1g8Q49eOqTU0EeYLbjAyH/ZySb0L1cm4rKIvcfelS
O7cRYma81U9e8dd7VV5KxKEs46TrNFNQzVgzvm/04P+joSh1ePSl9ml79GEGufpa5dVYeB7lcT2q
kAAVwYvkqJ0OwvZ7l1Kl4Wt34lXWd4REmaBDry758OBpjk7AP5sulnP6avHhNhOrmFW6vooXEVk+
skYjMCKXhrMHyMO1FkUpxgMvEb1N620uin3XrUYcaz/fhxgulJqDzWzN8QbmHaIz2/1TawYn9vsm
onf3TpweUQvxXxd20U0OcFSSrx+Nyf07TrUdTWNS0Tr1Gub4B73/sb74Ux4FaG5OsBdpkoqypT7c
jIg2s/JqZ+/E52UqKOjyq95kH86tnXR3h01IjEOgT597s5zL8inHcl4pW8fzp0q7lkEnXKqz9rmO
LxUuxF0BFE8fo3U5i0CV1xhF8rQp3dYGudYsbvlI1yDG0aCTRgGcDEAknpxHBxD1JTfLvTFe009L
J16EOAvOZVjgoqvnCgYszIAPVOX8R2c0zxA+/nTSfKN0BPCHVVhnCxjeB8c7ftwmBYBaeSbENYMT
Gke1MvBMcAy8uekBALk9N41/MSkMvmDJHD6IvSJU4jfLzdHs2cDcVEr20cioBlRUJ1XcvwBJHq8y
oILrAgF5XFzj4wxsXtnoKke1qV4/tT5YyNgesp10xh9Z7SDH7ancfm50oXxA3zLeGE+hL9emT7Jj
wFCI3+cidqTuFnfTnYgqPZRJImJtJKHKHyTIJyfafMwB/KRYo8FWsOkfwtvtr+ckn71IINmkWaNT
ibKPrYXpE56Af6fKfMPsy5SUtDU8PTVgDaRfdWRkuMvkEPGXLSDt3pzR7R6V7S+mM+aQsUwT27js
f9fwLqkzWncE5XumgjJN/zIKz0s2aKzfJ6zShTgzZzdRxP0DDlKYf6frTGCaduUjupk0TJimc5/Y
v3Gy1IcA3FqPBWn2YNhMfcC3o69uln8oOIQtkYrsSzwAswA1dSrm+pPW0zSrdw4mKjAtkfPThfcQ
Cb/Eer3cbN5A/s7qHxq+Qcpj2lmJeNrb/l5xCNOsPLTGBq9axuADtW7uxNNEZEM7QIxz/yMGuYeZ
G9dR7iHW4/kXe7N/rKgG5JuM6APbMx5cBp1UTanIs3lEWY77W+hJgD9lwmaXg5S+JiPub2RIbr8c
lbvsOiZZDx+HkErq0o3Va1bYyeG+tnTkFbrdEFiYKTW/0d5VB2GdY8UkrIvj3zSjiFzQMNEmDD6d
d5BkiulAk33/ZBJsG51JZqMq68m6+XplJjqAJPg1w8k1H8IK2ikCpEi8rP935+EqJOCO63PFZjYk
zd4VtPAodXeO4kaBRoIVjwx9lTDPyeyFK7FXMzApKp88w6FyhvtCw8e2jL9r+LC5ncVR55U13nsI
oeK9qBXPIjUIBpK4MQqdYsnut/YfLS+yCnDqyHDLYPvFz2HzmLBjZOR24zswpj3XcdmV8RD4ZK0h
7QVzwowU25Tm10tMUHrUDamE1sZrKiadc1/TpfsEAzHSUpXYFdZyTXmZULhgv99Y7cbf77iKUtwb
iTkJWbsnenc/bSf/xeu1bcCHjP4CIRGHx9rKG6R4nGGH9PUzjDzy33SRIcwHNGm70SpjH6SURqgj
vAkkCL1gX+0TLbss6MipeVNqAP3zfF2E3r/YOqp4WWIikKqJagB3sbopHGhbiuZaofEB1NXazPH9
TXZUd42G8kTIPopJhcH32j3O8C8/fgaRLLosWKMu43rJW0qRKkU3Z3DcqVtqsq9urKkWXVbEpLet
YkQu0D1DppVIx4hQkpMvjLLXb0wzwFzyWIvQJ9TxLlVAkR3c8fRxRtgRTCAkLZUMBISJQ0bQk6IT
cVS1UlghBlTlymgFio/1Ykbh1Lpovvftc9o/YJ0PFfeQKa8TnczvC720BrbBTroUuIACDCvG8yKB
wEThRlaFbVr0PrN0+A7FZJ0peVKkfPSwlIsdTw2PHkINbaoEXfIFKlR7b7PhSkfRWTiqBWpSFRnt
+t+mctB7N1WOozLIglXU8Te/FOeMlNsDCdlRMkl1IUPnVTcIdACW9WaI9k9MlbpVdqGEXH1HgLD+
H/FPAKbreCsJi/LC12dZ26NZmFS6wpoZoU4yWYI7asbVcOftP4rjumDgLYsxEsHEGTz9Sn9xo6L7
WZeXSTSTraP6qVjwZsLTME4tXqrGq3to/Itr1iisaZFwICsF6wedn6Kssyc4fQ4mMvl8Y4JT2Xx9
zuWeAOFbfeCG4ImTiQ7otrcd8y7M0BFoiYzWN4WdiWIbHUw/G72hkAhgI9WHSfwoNAcXYVeDPYG5
mEk2zzZj4qlZXjmCwbZeZne6SYPqFCocU/UahZcoiwF9VXbBPDVsDGx7KJK/ROfxOZQh4tIlJfkF
PjBd2Ai8YbFfcfhFp50819ldiPCG0uUXq+AcRkzk8khv/59QR47n0eUIfIt/zQzFytDz3UInmbXt
xlt4oAsYD62E0HrtOH2VDL61TtlXLh83LpY2cnBSmTieIwCezVF/uzFBBj5rAeGvu0s6HKD/Zcad
Kh2VRTeSjpIHu1TrZ5EfFBzICtBKWj2iM3tL4U6SJdPkHYooqmvyXE2savfwX442ya3yX+aauian
1Tq/MPbBPT8Z158XxNsegEM5BWdGX40HS8lnncvrN4cP4S2cgQT+m2H9ph1RZuL8XOrU/ZpUhK9U
/yMX1HPx2sWM5lnodfb//93r/TaV00NSxw9oL07USKabS3UOKVh/biTvj77D7p2W9R1EIG8enmR4
KyToT5+sbAHX2Y8p6JlHXeIAH9QHTTAndv5aegH5DGUCpOEa1GvsVyPpnwCuYQyqKpLuanAW/7I5
1Y/WTo5v7172FzzF3+acumC2KavWsdJN4jxE/ULbANtkAb3ciDEhZOByLIGjdi74wPeDhcIWE+8w
resIUpBR6a6k2iYls30jF77lx9MFwDtr1wdQPFJ9pJ8E1oQTfC1R2VRAvC5LnQ5cKH5PKoWqON1w
608tRxuy3bErTyiKtAwkrBXV+TMEhLUm7s6/l+J0o6U8KHuN0X8jSj/vxOS1ifwArY78wgSn5Zmv
F6jg7AnTipbYzdWVf1mvF4NL4RaA77Z60wV9zqa1T3cWntHtz3dWod21yrnsjRc9lh+OTS1gn90q
3NFOoumpW0V5ibmNDNFE+/RTPyU2+j56Ae8oLR+kYZh3UpTX3FoOjwbRZm6MGDQlKp8/ygtVTYlu
fDajf+mBJgk60H6oqi9Abmh6XpuYqxnZpNdnloF5S/bJTU7cuCxL7+Oytybck9k2eJ8tPcOhChd+
C4oI8lfTinayH8lq9YeYtsvy40ned2kB5DeUqlmHVjRvF7OdbBm2ZaBHR2QoaJHKrYQeyantZDk8
mCgyBizVgpMtYOnuV3mnk75/82ZXr3LIT8M2yrHMqN+Izt2v23XcKHpjlhYY3MgUZnKYkxHgyqLO
RvPWnTgMvHrvHNUVLPEtxE6hDrtn0L2S0Z782cfSZhCPHYLw5HfQCEk8lCBMHk2Y18HCEllrbxSp
YhGqBB3MW1Kp+/vU0ME4mP846PD9Kk43SkcOqMQRByzGroF21x0G5TpJncfG+68E0DhJdfosOrQI
1jJXS9BZ5UBItUoe48A1pgWfg7g0axKdEnMbYpaeSpNjl3ExtQsJcnjPGkLybT4xcULdMXC+D+s7
XoAUwqrwziQBsPICHS4utEVx7bfUcmxDtJJ+RwZlbmSyN98UCP94Z2++r99KqRFog/b/uofd3jwV
3BuXRzVVgORFxTHds9PLmbfCqcVAhw5jbm/0YCnukymQtVnfbd0/mlhmgsdsGDW5SyuYQBvhiQPV
hf6V/3OsUnRCrxYbjsz9n5qmm/9juknCeqaZM1ZwFiS+jA7jIiJxu6pwwyeOgi0r+xuVgoUUDi0l
EIo/ZuzOhiMns3xekQfL43UWLJcareOIyiUgDAQXQ5GWZYL/vhlyOp1yrGOT5Ubz5rlMa6dWXkEc
eWmP7mwYT5KI/7Ae/PqYp4YpoyLWjiMfCjsx8JqW6lOajv5buvRpMbGtuJNkF5MifgUMiof6T35k
rBses5L3NqGFXp/vDacYbPXaIa+SffQ0hMUojmk4mMJ3TIwe0rZnFGL4UVWZQx7OyLt84nQWr4HE
hu8HakfPG29H29JFyYa7In3SD84/3jP/2YWuDTH4iw3DBpI1q/4XR+YacsXE/1vBOoI87atS6nX9
CG7kto0Gyguq5v0OvqMq7LjzhkU9TDC/7c3qbxzyOrXKBA2ZlFnaOkFIdpqgCJw1t0EMUX/9o5kg
VU18pkSLbrYh56iWfeEF07Qk9PVOj04RT3WwaZv3ZxHgvXwHa8gE4WjYDDc4A+9zguBndZUy8Gmn
noRAKUNhGjuolWitTqAzxZ9Pd0FxW9CjnMpZDmWxIKt7YQq1Y53pLcHWKQAwrtp1wS7n/c+g1neX
d+7XombnX+JBujkPFRxjnmeu2A+KpKjfMGH7+LLEe8NUoVg7bgGVBk9FRG/R2E3c+AFHb3vkuLq5
SudRmCcJaVzKtKe/QN+OE1erGVW2toQRWCTAHXhaeidz76YLMwuQbdnL6NQ74Oprf9MOUR1yrNmY
/IOZBJ3hl63WirrLZrWl76reDBCO3CPl0mfJVKF9WH7VdMLanNGejpxAKbOE7XZ/6NpynNY0k0fW
86bfK9sMe39WgFDTiwWqHVrx2oNvyWW8CYlYPlGp1jeQjpsR5kFkc6xAu9ImHSoo4cn/hlISELKS
gPBkR8xF/rFjRhd1ibUxoywbfLsG7jBwIJToTSFmLsQ7ylWV9xqKjHmct8vWU99C2mxPY0djd6H9
akCIYS/wx1zsoGKh2mo0+k2W2pfo/NAgNd0HcKf06NkkDv1256Ub/KMlnzfp58F0s7vBWCjrBVVL
sXSSlKJmK7LvT67tNWg/VSONFkS9o+EkdU/1iyYigY9WzeBq9+XjJj255cj6z7fmyFhpjy5kgaDr
iU1sAqAGOnSTCXyQ8bZ+ax+9PQfMzLinYqjlAaqcL4elsc+1WOolf1a9tZNAQUlPSgol3cKMWijJ
7Fzmzrpj3wcnATM0o5T1bFsibcQ5ODvhv9OkBQIZY5t/NSLwo0XiFkTIHmrD+7v8u9DUPFeLsAk/
udLN3TRuq5DojzhduAksmWv+cPYZrq0dLRaYn53lYcHEaeofTMcxHWwdqnWPeVhzGF04wNSqirvr
B3o0CHCkNMJLE6Mt887XZqLD4zAXmcLUJbDW4pD0w0mye39sOajcnvpVZ7oemWeoGZ84JsISfgCo
zdIPsGk+i9zZnUGU8W24o3KEoQ11njaC+4lDId50L1WfNbiFmjRadVD0i4WVpH5D81CIwxV4TBFH
ugHPSLISTCYSOojhqVn+UFze2Qvuj4Q9ZmBUV0vk/UD628DwW1m+xDB1YwudG6cunqrOmLfmgX/q
M3DlnyJc2gbm54oMAHnsQjMq6Uj7ksoq5wQ1o+YU03S8hONKqas+BfFBlXMKq2ler9ITC2KNrkBz
EFgBX6C0Klr2VJ/wTQZ22tkiJkUOMg24M4QXGSP+q6erzrLvj76dbHsngH4zXhboDqlP19JSgVdV
HXDuLKbr/ihkqPwnbvh5BJW3QGTHpQRoNfbbmNVMZ3XeRWa0ab1oSjjyRmwjP22DZf0Orxl7WTcq
35DJhwYFZytD7+cb7QKfqz0R5yfDMMgMFH0TeAfjTdP68LII1HgpcQv4PqApSlVFk2e1tmaFGfVV
0a1Cp7wjR4yqwqo4J2OIHMAQomY8+e9x4cQF6eS4BYS2kyW+a98doEEaVWGgF3H/4odRPh+vI1OW
VD80xtC+d1CF73GwZPQ+68LOTtOwpiYEhCzjPQ1wmIrXz8+iqw8OPt5pzsSuP+90fCO00hpVfKhF
CvqISTA4pz8/+G646hTypo4qVDQontnkOssWbWMiINgiCNBz6mSUSEVELBTtjGluJIphr++rP5Oo
jdm7V85PFW/tmdEGQ/TIoKmvyju6AF1l4hoKmrV0jE63n+dnEMvfpICf3vMOqXSwERLQMxHdGq5u
ZvPBEp/kJeQ5jFXL35Pet5VQ/8vTkbgkWd1fGH0esbfTht6bH8XQdCTvia6T26l+Bt7dUA4YIOgL
/VhIqEOO83HAb7b8HwmpG3IMn2eLCkjBrPadqIb2i6sIDf/flneNLmxc7pi3qGkQnfKXiLaTkJw6
HAuMDCw3Wp4fUWHZ27W9ixaKyB/TTEzd+SoyyFI6JZSwhuzE1tZBkD2o0WsIGlhaHooDk05zOBUd
zWU6YDCXbcGay5xNf0T02+xtEA7YhYx3oohTOz2G8Vm02cW/HhSSiXiTfDhMs9jJFahOpTa/Y2Hi
Yw4VQNRFTw+0ApHXUPQx12hFL353B0hDm46Kn5vGvSEYG/JesW1kgZZChDk1kTClPc2IlMbJkkK7
q+7fWa03U8U/bqyBe/eQJ/GFQ+/nJoDNb+g7NopcCxm4gWoIIy9sjSsCnY7xZ+CwNDhaGADXkMJY
2guvwwOLAFbZf22uAbHwQT6CUy3UlS+IrgMDmJ0e+znYEIh1isXlhCOZPc9rhtxJdSjSZlcpN/vZ
IJTlGAc7/THVqBuQl6KR46Y/ZzUuBsqRz7eWoYiJ4shZeOsWzgiryj5F091xMmP70Xi3Zic1o0q1
YIzQ05oFinsOiytjcG9tdxOcSOY+dXzg4Jr+jH6aSyZdPkwHZ3DtuRP4oeknxAoCwu1DHYl+rib6
PkjDlw3a7wL6z8z5Z6wKLEi8mNkknznhn5tHz+dj21KreiSISfoSKTtLvffMHFNWXjcAfM9dJafs
shqCNge0A28/4o3WhBeBKsaJrBQrR4kToDlEBMINkEtPyfsrDQhFXi+BMF59ZvJsG/zmUt5wGg/u
9hgl9t/EaXjTPGE+Xj5vGuUEGtdHIg4SXDanoBaGSmErcnVTe7eJRP1o/v3KdRwMD/lMSUN1c8jX
A0FtRAUdiHt1Aqn4/QHQxYBHyC7CqUk64+FUfiXTtDxs9dQOX7lQI5sFc5gcjGZEFifHx2v07Loh
BBdEkRcFNvqGrdCOPbNQv0LKTswBqaRDHiVMA65TZbvTcNGlhH0jZja+q4C/8VAUUfBEQpgpGS4j
q0ALNlf2Og2K3A3qbyX62lIxwk9MCOZZud5G04Bx2HGZjGFH9x0OFibUDiHPYzuGNbyt5TH22yct
1y4FUEHeDNbCRvImW6pTtLb/nlRKcBR8Ix3L3SK3v3fO6KhO3bFUo1vQSPGa672IqwM4kkSYVbhd
bQ/o1xT0PKXfbda5RK40s/r3snzHL0JxDzM7sVD0kFuXBWexAWoJBbhr769uJscLojD9eOwMHcN/
oneIXK84J9uiobE0i/XkUBLic2wA5mNlUfeOjgctJ/HlkgetkfliClnmMthRIUpOb85v4p8tfYwP
B+boLG1LW6SXNljVHgkVknby4km9kws1h/ydy5boPoXJeXh37lddQ43TS+aKCjK/zYlDfujak3Hh
m9T/uv+bIcZ5HK6VszPrYJbIB1IJ1brl6S/uuDEgSkBOrCuSuOk2kQ4j6oI87koTIb0FCOPH649o
6noTmc8nM9yacX89hf8af8jOJs7uIqBocDm9L+VkgSF4PuPwrsQVNwBYEcbvpz2noDJvp77VEunD
raz56d8mddbW+LYK0onTzX4S2ftHwKWkRmUXEFzo/7hjn0nHpuK7PGXQ0+2GD6qM7G/pBctCB6ww
UXuZkOACE0VqakXCNk7Z+n5SpGldZiKfnCVuQ0oQSG0P8783dKYtcstLnd6rAbOLqElLbw8uoRTp
dmSA1Xh6PmLAJeFj5a00T5bVCw3VT/xQceE7qV0Qc+GrB9tqzAp+aHaOfCeajH2KpW5GGaysF2In
jO5w3kxn5IXJgm9GpSycQM+5Y4VZojoQPROBDd8mtdQ/YoO1hXcLUKH/jLZJSlSZuEfoOKpSITF7
U2CIeMljFO0Z3eaBU98r+BibYkfsEifuMRPFP23tJrrrZDDXy4fPJElonumHbVdacPT6FTgUBpTV
C6nfsZE/hlDV/sn2f2DWf6OeaZRS108/0aD76a5vbZSZXV3qafxQAn9XxhPDnhsV53EdJFI4Vs8T
AiQDVFfQDtz1p5ud5DOLEdQIUSrNMFmaTDDkbl3TOln9SDJaIAzTiZneJK7/LJv4vJBUPfEF6/ZU
s7Sl6/lt5uUW2Dhu2aIrnH5LpAREQ/FJ647HxvB52hX2/ot4wORG9ytMwBE0/kWxfLZx8O5rSbmc
oE1UQB28njLdm72KulLKWFpmB8SBBb26fw375h6Dto5YSvQddjLgJhvHReKJxW5eLk1TMG8pVQjI
LC7GKBUUmMGUSCMzQ1uH1adUOAYrUYPwSQLFcim6/HtTzJQZkhuy1Mh0P1xbhu9XVKTvgNezNBbX
XcSSxsAeiu6AxsiudtBIea778rUVidU1N7g/lXvJuhwqkheXl7W/U4gs5N9XSg0XQ1W8p21A/HF9
PXjrBnJb6/HIjmo+r0+lhrYkkE2rZWLSkPJvowgO/B2T/w+2jHPxEFCZwaUTX96GAys7ehYeWz49
QkABRlyPB55eSiMkrr5QGy0uuzSFF/TT9+1Jf4o0zQUapEVnicY0BXPrJ9XgF4sYvJnf2NZ2l2aI
kp3TAffFHRvesBtXC51j6AjM4MZrfUKnR2Z8oTC6bcVxfFVeuDcv05WYkE/vTel5V7KM+/t03+Xd
//qEzCQseVeF5Qjsw3NrnaaOQ4vz0SRi0+JxkGTDTWw1FsRkQ4rmjdjViiiMbzylolnOHLOtgcTu
4U8YCJJL79fpY+ieBL+VNgnKHzYVJuVuBtwhryllHiThu2cUNohJNtdP2vCKhMw08Zgq6wcdZFJ5
OoZ2/b9TzVTcYeJnGRQ4DfGTW83rYAolEwW6+Tz9hTjQVPiLdhLdusrH0RugaAAsbTmLYywBfzUJ
MyCuMSAqidsKKRzTA3SvxHA8HVpPHCMHlYv4k1tANm38LTq+1JzspJJmj5lKRppSBfkuXhnHJEP7
NRmyOHLv/oM4UYUjC08CBNOoljA4BMXnc5zsSVocF4tdCxlUWofLuUq8Ykhw/uIQ+jWqr7PU5dLh
78g13ASNC6V2DZkxa3kINp55tQmdcFbqbPygps8u0A+E9CvUle86OKHfTeHKHF2h3Qva6uJ+TMZN
kqObV9/2tLHQMJo7YLq33p4onhsk5A5CYiyschlfsjeCF4WhPB2BTCW+hJbqC8IOQT0+XG+ovaO3
6/t3oATI0wc9/BoraqHoxAp/JTIJvfyGX2bLSMT4Zj6KHAl090IN7YOCWoJ/BFkOOuAKuxNxf+Jj
SYMLOhCew/p9wi8KBVllarsweyMRNy2kywvsqcn2KuAGY/AtuZRyJFE/Pt0akwFBBr1t0ybC1t2z
YXO4tWoMfV+0pX/8mhkpNcup5g6oyp3Ma9KTsH2oHNNsowAWt1GUvvR2WR1/szPCPJsLH5dnbIca
bkO6h+tWieuA89B3fgZrhXw4nbm55O0qJgHYuXFU1UysyBU+4Od2sBZEJAj0qG+WWlQfoRXyhM5e
Cq/7SiVd72/bwzuUgzFFNWB7GYadm/3mOefGTDffO/c1N4Y3GlhXyTFurVyV4fPE+NRdqIIrBCl1
pcjyquz35K4hHe8Wna8DCqFN7axXp3HCDP2/FxyQy9OJXusJ+ID9V16uKKVR2KP/x1kosCR2GcvH
WjOYzlM/t0Own7YMpya6WQJv/RaorKRsDll2i0q8QJ4lP6PgxiiXDoLBj3k47W9qBBYQO98N58EQ
YJuQGkkZ3H/CUA9rLBMbnKmt5zgBUSejvTXL3SvWXOTDdJhEtQCrlQTgLBfUv4XpyzZ2yavR1w3C
Qo+JfnXY7M6+l9DxZWq6qX/clL+GvE2NeBGtzSWVOvQtwdUQzk2+Ya5w7aYSwzSOA8Gxw+DOeXjt
zBFVxSByhM2H+vatC3qURJWMEsKJSOdhbqP4/74F7BWyOsa84qUl4BQXvGBZf/edtz8PvC9ZDYQK
4OfL6XVUbw6TvcmvYRMZQjwrLQJHWjfeFF0kFewFPo8nKmxoCBOhXzzfTKc/8hKNofkgkI+s852q
iK+8caL+RXiU2vm8oihR0mmWDCPfFIzTfSPyMxiD/P1Ix4zo1x+C+ibMjAoIPkZLSHX0/HfduHyq
0H+/l4EkLHxXPJyMnDsc8uttCbwzirkrRZ6vKthej96FCnSC3Ff44dlroksdxAP7rtCs6NdwPLjl
upDVh00/syzjcj99Wrf+Pxk2ui3wfYd26g+gG0YhpsnUriy5iGUSDTyyc0KbpYM35wKQMUrHVEYJ
JPBukneUZtRsH8xf9U/8gOJYygh8cAbrEg+ajrFOrUaRH0dvlYN+OByEOI34RjEAJtbpgf1agqXb
0pAvtw6zD7HW6+eTCZe6ZTz43r+znJxu+nqdyDMP//RGjEqm2cNqMXhuIkbHEdlraDjmd/R7y0Zp
moAMfXQyz+119NuGDIRyjIvs8uQTedW3HmWgVZV7K+3EwaOeVpv5M2KUSUGdxzLf/bqxJIgF1TkO
Z5K0yWVC1KJKiKkO5vDvZXr5NAh93Ax8/+6dDP0P4Z1iL6xVc6RpkRTVwylurhuLMGTIrzNkOjfj
eK0k/BIgXCq/e/SL8N4Z0ubIgKhNA0VpF51N7GDDoLMWDWotX/NwMFXzOX2UwFwX7e/nsIwoISkv
LBBAG7vetkTiFoMImuMuow0G5lv3ZFDowTyjq6wWIJoU7BLwYng0ftoXZ+fJrRi7s2c+aXL2c1Mi
RvP9+j2AQmIBdMTxEbzobNRP5QFSVATyV8PFgf+nmGBdC/bWHA9eD8eElXYXhrRM2mCd007q9MaA
t+F2rCwLhjkvws5np5+HoqTyOifnGdXLCKh76G2F004M0JLoJnSQyoeymNKOZPyB+vWV5/Lz7pr7
4On+4UHrs0WcqnhBe7HRZGCMbfpOkRRvFQxX3MuqetNRjwBC71E8W1PwC5tsSaWQ+sfR/Yfw1ls6
KzYpktV4MVHaOhFc0r/pyRz4hs2/GUwDvB9rcijl7jbTUaE3lqFv8FJW7KUSYBnL0tJVCVnclwhL
gC3BvDV6upu7f0mwTVBtup/y0XtmFpF9S1h8EoBST4vmB8TVjQwRWpjdfR/eUzIrqLLuXvsD4fNq
pw0Vw5BZDAGDv2UlvYt6BdQ+mlEpes1sRWO0ETC+Gk+ziuNrl+lCGm+tkAMeLDZ1eQNgq4XS00t1
1H6Y/yX6KPF8MClJvDgouBmZU5EJycYAu3IvztL5YO9ygiLnTvYQdRI7rdojlfxk1gZ4JU82cRwP
Byd9NVyKdRL6w0lxG69rmOIkpHYfvJD9jzWSPXr26ROyJbNJw5eRJddTyfB7g0+fJk5ZTPzgWWT5
u4szHK7itWllcRbn2Kd8A5b8Sb/3u111ulSqyoyctNN+SLrPqxDy31vpx07+2ViNkPkKwnsTzxO9
pQbAs+13RUcId4cQfKS8rEhbs2DpBlzEasGpRpWJ0+7/VbKB8KDzDFUIVommWxL6DvTau6IWVQL2
Rdu+Nl/XDk5ZS/MekzUNC+ASP1jiF//4lPd6icBHtoikumc251rmYT/SgFDTfRArO4+WfUgeZ0PF
Dij/JGB2ZrDKyLT6sqXJ78YlmWgMMW6jWdA6MHda+zX9FANrY53WRSA3IMsx55kHz12Q+wQTYiSG
d/3kNOOHVtCfRvv8JiFuGEEghbUrx2Y6O0iHXN8st8mY91jaqx2oSKqxS5WD/fy6So6YfC+vPXRN
3+P8h9YPbz3hgCF/wv2Wf+tMhgpF+c5nulMyG8K+gei4DgU+vmwFE22T9bmTxJAfa3DUyFFYnmz/
yvCzzlcBaeLbcvgz5Gj2Z+SAJ91KBklXYcEWyh355QVcCCVixGe7+RkMt9dLZKzh20E0MmYHJhjZ
DqInFFPgHTMpJxnrIb6L8upL6GLoICbPdn04hVPqF4SmGCzqrT0iniUKs3OG1lH8ayqKufq1/8Fh
b9mVrW2u3QjAxCI1lXHXvBvpWGy+LD/EaLdeupjI7BkhAHq7BTvOX2NaFmGBJeRHkC+wdv7KA1S/
pWu1eEjKpYYUtbO+3/nt4Wu4XnVk6aTOfAB5AhJdp7Zpmr1kDhZMhaiY+3JjywgQrfiPNT73P2a7
VhZi0jZZFCitHvRAKd3iAzg/HAGNdUx4VO+uwxFbopso8KpbOEl7TrDE0WEknlnLEZ4pOBtaQ7kx
R20i2j41EyhZ9mxTTzZgkpIz2e7x8XeVPHd/pZKgjl23ovVqLKUM/rMQ0ynD3i+vCwAnr8k3Om/M
pkUgFeTtwbWOBAGTmn8/MvvVJT9cLwGeJRoXwdtuC4gHeuk+/J1aXpD6lMnMjT5NfunuJF4mZiQ9
YNUHmhrq3D1X+EB81ETQZwb9PIAg9HqSoD8vjnp0gnteh5qJ2qt1pxYAgjliy7SjjLkurZvh9pcB
4efgonAvNZ1DulIdr0rnxHcjNL2oZ7L2nM+Y7YIMGkDL/99bLUQ6dgPbsEMONsjrt3jIwaDIum3w
ze+v59XJT7esHKP825xeSGHO1RaQb8E+pzJKh3aLBx2pC9t4aHlesN6WnbouFEfZpl5wHkapVmdK
uuBX5TDblsE9oltWCWffObCstdAwiXu/+RfatSAiKCuoeMhwUIXKHuHfNq0HWn7WRAf/ra6bZi0k
STOZgKxRxK1Nl5Rxylkr1rsRJGfsdSkk9b21tpK1aui2KbZbOvEy9fM6GMQSu6Tpsis7vv7mLDiy
tleuWzim9fEOvj0RKGS+mEwwYYl6K+wlBMN2TKXOTioyK5dJaq9Sl0DRdcxPjsWCJJ3LYTofidWl
gUlBVAdyVVlQ9vkfVPUPBYQOsj406NXq8vvmO8YrBAZg54ru4nC3ni9c7QzKaSKpitWq4qElrxaL
gn5a95D4SpVx/kNLKw3p+aVXpCSYjNDKcgXjdwLcN6WinGm5znERQD2k2Lc6+xHqE4DQUi07GTG+
sZRhon1+Ws9yswVohekNAuBzzvmB+EkljH1qNzzJwiPdC6Jf5HaXZwIMRJ371oag0H5PuDOYYygt
edx8nACjG+eBH2JYUI38/tgpfX1dalKY/R4iiYuPC4zjH0n9Z4m4YxIxqGP5IXxcF1mZS1ioHCxa
YFqyb65OeeWypnz99BQWaCbgOGwclB0vBXeEcCCGDhqNe+DiShZJP/JESUWpZLHMwDFayTXSKvjR
petLyiKRFMajHuoXVIZq4samluZUdbgJ+SbzewYM5LJALt4FfRYAsseCer3z/cnOLZJ7TbCEcrWa
j6AkPw5wISrfG+VxDY9+t6Zqvm1XcclQzGRVyKMk1FxmSDJJHm/L6VxK1QKaiWq685FBU2k6odLk
Htg8m2xjNqw+KG7nKCh4BOkASIP7bxkjjpJ2qtaFP0gmcRhwmqYqxnaPlMvxOqqL33pXLopTbh+6
Insdid8ud8H5/sKeoWfOzzRq9jbumSn4ZXsdDTmNcLqtTQ/zw9ZQdEXWXVU71pW0Io2chDySOb1f
l1h0pOEBMKNpsnpXzgIzHuWMi1rfZEBeZ3HbotoJWFjrQKVi4FtHqkcp2qbTDSPHTvWgmQ8auQsy
DQXbxZFDhLDfkMFzAE5NexIBfh+PUJxYEipPiBerFEP9Z6XqyDuCvtpYfFMpkk0A8Twb0f1C917t
LFm3PSU6uK9sVUeI7c3YiAIRRGHpNWOyJWpz9Pqsa1PS4DVkz8Cn5g+3yvJHgUfufmv3qeCiXPsJ
lMK8VSDmimr32FJYvSrvO3nn9F+gfiioL54MpWsRcOhY+Z5NznLrc40xE0EAUkwu4UfTh0GDsSag
qza4NLgeqkNoEoOegmk1U9jozszSco5184Y9UFq35NcwlZhTXCW4CQu4Pnv5QZPKxAIGGH4oeVuq
RRj96Dd4w+zXRWI72nYThEJ1Ct+aw2rRD7r/k357A/jJtI/ik02EW5NXXrEaFE7Pf0Ji7eN7WkzE
OAZNjFCeL0rUEs8AQj2srsMshrZU2e/u4Cgdlwx/s4MVPlwTfm/23i8aiqECGFmaGmTojejAX+l8
65SeM25rzUGaCyI7cPAL+7fkWzWob5Sgt8ykJKKq4fVUa4VdBj5vzncPDfVs6W8lbaSc6dxH5Bk/
76Gec5MfsfduTDn3Nh/Q3YYAFF1Zzd/iqfbkjYGp/QzaGx9BpmOgbBqE2D45t9oLbuz9SQgGQ78S
kmFiJSgaUrVKeJQHiAHE1kZa9jYeyNemXkUqS8SYsNehd6Eq1JT0IerstOkK9NCDchaU8a8Fu+Gs
Xl3YxpGH1lY+kSBiCKUiIGQD+xMI0/DrsAgD4JuAYhLqWlWTzMoO5p8blp1R4HNGNOB5rAi6+Mv1
zz2TaqdfsCBsR1iQYLhkwzY1LU8xsPwr+2RgJi9pvh+3qGFrqgV3qOyTQIGNeSaHhMGWeuIs39Od
FZ/4CfszuoxlhbB74sTvmgmI1BjPjQkCKawuB+oxXvbMJGFjrgjLn5V1yLPxMLOvItKTgz9SgxUu
RMBjVt+DfVi548MC/kUU/K2kCgechULdIWYxV7NzKyR5MfRo58+4Ib9jEas4oUiwLsjfnKU8yTLC
UXONanVQmmy0iyJuRa3sxtL7zdFJL2UA2krQzmStvUoMF9BGZqrgO+aTsaLpGOCR73ZpnfmgMR/V
kRQdpiLpV3xLui0Vri0xx4whq00+YS2F/a4U6DvkAYSNV6N2oKrPWo1PKg+64tJu9JiFmB9Cs7+d
I3D56KBnXNam8bzN9Cg4GO1OiTLi/0ucmKAWNhSTszuOOSMAkkdxULm0kUjZ2TwE1O4WortKuZNk
DkgX0iGeUBDSrM4DWGRB85/xVbtdEXA97njUcwlB6fodaf/s14vGXM4DJYRLtp5LV9z2BssDfLAr
OwiXLtYml1+//WNeFVVOtBK8Pb1u+ZPYSMhAVUmUyuYZFTAjpMeDIHbnMXoFuQJpTA5yrG8/tld6
Vl0WgkMZZCigPk+WvciENCKJssVNU5g+R3bs4pVkimrspWKvTMoeeDpKDb8+1Df+Y0ymANZpLdD4
l69ctZOwTsnqZhDQ3uGmhC/poUXcDTaIhCRYvbrSR/MNTs52LXvRv2WL6/OYWUT/QEeUbTj43ejB
BlHz6Wu4mFz48h/YDWfxir2ewxsG8KjDpy1Rdbi6U0XLsKuiE6gZSbks9MzTkQ5YV5IcTVm8Swio
1faqsWW5MOcIr64Ih3TalPER+t3SW+6Glha3CZ08RSoxN9UL/Rb8oDCBuBydgp8UUmMXH+BRP1wS
LEXK7TxbLXOg8SpDT1ngPc/YA55RlD3n8Gy9zgmMhck1GDBOalap+4IDFs1JTp7KMxKE4IBTJfFU
zvDfPbLdEc3oDQlYhn63Es/TPTtGrXrVilYjuwbJkf058PldnToSzif6+puB0SzQwdS3TwusJ9YU
gbHRecTl2SYrZJ2Ts5IpEE6QitNoNgCvlZ301Vh2UZyxQK40X2RdBxd3CyrRlVzTwqSJ1rGUpqBG
Z3+ddkLOnAoUr/Pv+Y7rRWIlYs4W2I4R7TDGgxl93I709/UELxxbZzHKlc/ksipypdvupL+dK6h9
pmMwJI3xg8UKRQPgcLPL0KUBFYPfJ6v9E5iEemgRq9Fmny5YMtsL18F4Mae9sQiCly7YG253o5NV
FEVB4pQdJqGugQlkLm/A3f91jl8G+tP2QScVc1pqLUz+AZrZlHMm2Qh1HaiVmTvx2/nZRQxywjiZ
HZeFWTkHmP1AjqEphUq9ESCpMMEAaflHxrFJF0jxJ+dGh5erMB6RQj2Q8qi6lyxOjeLt4Rsd5zTU
x4HUVts7tlmqy7qpeUTi0WV03ky5W7jh9R6736W0iQeWl7aBmZKsBG98iubMJgrsWYgfoKm8gA7l
B+9GE7AY63LRjSN8LQlgBUl5INF1xmmbvR/CKCrPNK2DnlHrU9XsH0jdjWtpw1QUev9UBgxvAjmI
sWwBHXkpIco773WRVr+gjlG7/yYbUcLUAsHWjwsPvZM0Eajnhr84xeEeQ1lzqlf9AfoTskwtrT1z
4u+NG+1pUEn+2dAYr+CVWvg1eR5t2wSzKaPlVuh492zFYOkIlojvveR2qaric7cHMAf3txXfYLu0
udRiQn4d6ZOxXvYzxEs1foDWiCVTSrpBYwY2GupUnYDwIEQuxFrhzWd2SkhPXsEkvjGp6Ny9XYBG
BUdV2bd/q3HtmUQz1F6onoZ/9lSUDzDB/0vI0iBJGFDM1lz+Z0uek/s1ovMjdKfzlskMrEOKg5GH
w9E6EkcoMaqAX0AFl3oj9vPWiAZo1uR6ESruTAkUV7pmBTJsgdm3Axoa0SmbhymUWTlyUBhbX1xA
clQnhhLsDp1aJHH9T/+VSIIHey8faWIfeyScM1vCnXnRCXIDzJHszXBOjDxmaYOTL1iUrXkjdQiu
trLD4fapf04z6viGgHCAJfK6Mvi7ke5QjDqsQmEXBhO1Kh1FIjYaPNxi6KzOZuBVxLesZpqnbCbC
wo1ZjAadxAIkxSUT+xkG5ZKyJHX9lOsxwMTViWMwnRAph1qeuSsM83/Xp6eVcumjVS+uARqxj7Ii
2MRIStCpgOUZGTBQc+WbPGqeCsxZdQcHAkLRP2CCCE91ebBybTE0UqIt7IBj7cNgS/XqhUgLYHWW
mPsHEFj4p/mzUsqELRiXB40Z++YwAu/LNq8Bm/eK+bdL8Er4sRqET1LY+ED7MGf6ZXlxMDpdg0MB
Za+9lMIhXf43hJB2a78qe5fyIbfuEscxIK2CRuBIW30nPwm8A35TEN6FnqfEkyw5vXp2hqGcc0M2
9mlQ11v+3DUiozGgn9dbajLsv8y9O+F4uZCm2T8c17nCO7SD0hk2e3hwKtzhn9Khwes2LWAmJU0i
H6N0wwVtkm98AQPeVuJVVe+7YNM5+cREeLCyjv60cI31pFXtDsfMNjrPS07G4DvtUucqp7XwuMWP
kpuUvEau2Kqc6oTjskSUaj2rMcbVoE9PUTgckhNad0TSssrWg4of4yFJTR8e2WqNMHy4RDCWg1q0
T8QlBJ70Zm9Ryb9Ni2Sb/HZj9VpeixXkTwpfoUGz6yVOkxohZKOGiP3Ev7UDizcXy3SF03JcPi4t
lsV2jVBymGq2FdqWNcBSW8y67UDlQyFTiGWxJhLdAmXvkh0z1IFVJTSqvp/Ay1kB41H/+ZOkKchH
h5P57Pls1yWJ7GwiTuRbI9CXpaDH55zWmRrGx9A24iNpYaKiDCxsrPaOLMjYr7vCvTGfiKnxrVO2
gIE+J0B1ZCyMmj+vpFsRV+KyTCRvWCnx+VtEa75tXhQCNNK/jzK+vXEkSS6TDZIg2vcWSchPLSrH
o9KiNainHIzPd2ThUseOmVI/mzQyVa/+EjbvnGmDlzi7DExoSKtr7dArtMxYw7oBxYP289b9V9MF
39qYoLrA+PFBBr5QNo4ILqW5zGLW/1+p81KVsBNN76+UMUkA0mA1HdGdgjYrQPmxGJdXUPtGUVyV
OJUluX6c0dkKOWb2XZAXx0MQgdJhcUggMvqARkaf7DOjRmiIh7KcsxejWdSIh/8tZSjYfzmjm6Vj
K4tbJ3cN12HOIRTPMSBQwTeKv07yQ3L5KRdNLYWNImq4JC8PRVoNBHymRsz9VKY8NpV4ugXFXTk5
oih8q7xS/7vnjQnPsznwReI6Sktjjbd/i3LFMhVZoZRhbZEN7gVnA+wnY6ftGGW/AlJU38am8Y8+
gSDt0k/EtL8TWEu8OcbZ60A+WGqQFC8zQfJNzS2JiVmwMYIB3TbNF2+z55aQ2eiiZpO5qtI1JlTZ
tM9nTzDCnXJKRxe1c2/K6nyJDEPuiK4InyoMPfBbCLnVu6NBl8232ZjsW0WI5H1w/K3RfpYzm34A
wUkzZOIp7P59L9TtNtSgihaHMWUrVChap5DNqLwa/4mxm7Skre5AXSqK5PcDGC6yoVZz4/RA3efj
UEggipCEfr+fHmxIe9Jgzwd62ldD/tOHBiadyCAFGOTOrbfuqwG8w2Jv7xKs3xLOinr6RpykXt/y
kEWl36wmQ4Nse3LmBJARwzt4K69s/kruDbxqa5hSmzk6236DVRo0K7GlvPZiCbNsRp5o9eP676lM
CjI0FlLP4Fmy+daZI0GcUeTNskIwNHuD8ZmefpofXUQCDtH1HHJv1JY75RMFQ4G7QiN6qZkRq3e/
x1RJDP0TzGphud+Yg0ZX8Sjg3sU+9IS21E7esMbsnt1nKlyuB+NBb3x/walM02Wclb70zSil+6nr
vcspmBJxGhamU79PHj7PSOmcU+Ah0ZdNgaV2xeZXSTADCzzEy0HMnDMNGZOGF8DwwtCSnQLfFfy6
GisTfQmrqRn023eWLPYwf/8BU8Z/Kgz3iTZ5DUc4qQ+clM40d141JwFYUrbQEepnwEKoGRu52g7h
ZvFLrud9xRSmFtCM/ga7Mue94jyzHZtWOYPZLgoFFyQlGZWayVX5fMrULTxk2y7JM39JtIBGAdad
Y2ltm7DP4koLnpbqG6SiB4CuB+b2ZiTMIAHSfdlu9R1RF5aAFppr5B6imTg1o3uXuDCMWQDWmWU+
uNncBY4cIKKTTO4AEdHoXzURI8/Fkjno0riVtp0+fHYXIU8241UEVlmWaUwAprdQjeny/lnrjzKB
qsTZCAAqw9gaeBIY2OVgAKAzcZKl6oD/R28SBjQL+gzYxBuxAa7QUSF5wTqQfLKy7MoItdImJaPC
3X+7VB6kWaWRPAZiwfOBJvi9B2GSaFH9PtvlYlYwmoz41ZIdct7hYYpU9nkvlilupNjYT5Z0WeZ8
zRo+lMqyxHm3tgrgjasWBDVTanTEuixwYmZxHBw+1xBn0ByHXX36G8gFN7WWuarDn0PJlqHgOjAw
dj+lUPtLcaqnYmNPexSzmI5ZFliK8hrxbW1WLU/Ys0Nu0nvfmct9/4ERSrifHmR7bvj9P+wUyY2r
3GHai/fW6zqEogQBJZtgm6JfEdlUW0lKYK5CL9GwCoynVDiGErP6BzEpSqiKvmpno4tdG5nrd2IG
+EEN/rX5j8XVI+w+T1JGxPq2DjD5/j4A1HKxCJLOvdk4G8U/oAXfzOOikPv5H/gn6xMj3/1AmZLg
JwNcemA6PcVLHQZZBHHlpM+3J+KRZ4EOgVsjWMDBlaXRc0MEV6EezVEqSSvZrvJ4nFi+jmc+izlg
4Wvowk/x5nJOoLRhq5pkchSKcvofsdiUCTiBStYO4EsoQG+s39KQgcs1OyxyEzIxpHaqtwffUy4p
Ng9tsGuHl1V9YU/ZkqhGsGXYPfLLHDeql5URjU5UkKLH+KNLTNcWkH6j9BHRXSa7z715Dvxj92Zg
1c8v76i+8zPmGl9zPwgIibrohB3ON/3+19FzDG8B9fkxt18gSQZUI8eR7k+404gIsWxqXLbqvZJS
ZPZXkumKrFlgAl0mVHS9e7fykaoQ7AgeVWh7ZsHnKolun+Mot0pnWA9xvME/6D7aU49OM9Odn675
K4uPupQfHui1uqQx55xNi8VSGbJBafT4uc5CKiuzHGAUUFvfhiXpvuD1+EiBhHthRJqcwB2RirZ3
zeUTkJbDRaiRSfcyI9A7YUnYn2uz55WKDBjTtBkPUUSf2LRCcLEdd1WSEhrNuey++XWMY05ZksHi
P/a0eo6pqKgBaAy5Ls5hThHS3N+WoHxA3GSpzQfQnjPP0NlhoVw0MOzXQJDHItVbGeXWm+0XGi6j
tzexYU8e11kLMmvxG7xbMU98MhhshnjObqkqOs2qLSaLRiZQ/oCipzWz0cFWlKG4qutux4tM0yLY
XFm42q9nMT4P6x59j7u5OSkNIOG1pzJOH73wNG9Zlkvku9ZPYuJzs4r2ZfV42q2PDyOaVf8cGkDW
JLM2tDzWrFdshHzDVUGDB9Vyz3N5xlzDF31/oeT+82pBc+yMEWiH6wDgLEh4HDWWYpXBcx/mm3jg
hpBaMErL530rzqVuEQ9y4gblauRWAyLEqnwDFXkS82qX0WVAkUz57ciR2AtUqE0VMu8W/s7SyHau
EvyS6djbPv76kvUpEjOmahQQ1c/WnwlC4vBfstdy53JI196emh0CHdo4UfVnc4xGSHAR0NLx5h42
nFYZw977HRb2yYxf5GYs4Y1Brd8OH6B2YWjYHmWEccY0yZFD0z5t0pWM1l7nR32MLupA1yGtzQA3
5GrvMp7LNEF2Y+ZEDHjgK14+OQ5Of2n2Mm0zjCPbEinPYCoq9Z0MCIZxry54GHOKNU8IK0UJ7Ggo
KupZ6TL1XHvehvGIo8RYqJ/zPfXOEm+3LnBYeTG9QhmGA8MlNtgdBO/Nt8nWtesl+qi6XPm2sLJ6
L32M/TMfN4ed9IGUZaND+mc2KeAdKZ0b7G0dOINtMPcZOutoOAn2YxJYjGVXBAiXg/wCTVM4RbPU
LHSacBvIFuxHWt+pIjJcTykMf3RkFp2ab3/mxI13C8RmnHFqvGq15KU9y/HjJnA4fDnWY9M08Bwb
XJy+nj4sa7kfpxXWq8No1GS3DR2OgHaYGb9e+tzC2pbRWZDGAMtOV58JuYeWNO6F3wRm94vrjwBy
ovaxFGzRB4VNU5kIrnBqYu5VSnHvKkFXfrKGsqV2qTarV/3RCKpe9nL9e9cMYYwLQstiYj3m9w0Q
XKDzNQTWz3fy4HXHdiNIlYzKgnyBiqGRrEMwbLiU3Z4gS7tkftsnuXnGQ+KDUze543wNdjj0wyC+
VQfCb7tj4JaDfG07luMNhQM7rOpbgI0spyYVK6vsiAofoa95wzGuNnjHUOFAsei/UgCLmNHcaAbv
5OAD6nzu3b7vqzVz/eMUDVuWBRU5Zrjubk+VkrrLF0aKevmpi1X86VrNpRXdCKKyw/R8ZIDI8gGY
hKyj2xWL/qppEQz1Aih20d9cgim9h1zfvYHDH5Q/pOsR+f9lK/OlR6B8UNcBb7+fmEm1QkSuEU2O
qD4i7Zo3oq6OK+OhI5/EZv9Tz6eKmaBXqCqMElaW8+7GSr1/C8MVHft07MQ7gCwzqFnoztRkVDbD
bx9RjQDA1x+nRwPf3ythoQdLibuzpd8GoWSw110mvf/8I+TdoBb36YoyW7nz6YT7zWlP39yJ2ax3
r0RSYuNoN5/vsK4Ar18m/O9kpvwJQfGdM6NLlHRFh/sG6SQP2xfu7jrY3tKIctNEmwKylMCi9e1j
Mq4LlR9jqLICF3WYBcWeCSronNfc72fHLGn1ohaFPhxXJJIuYsILHWIRvB1/d93ixBBdpduYCqB9
t3sph9yk0bsD1LlN8XERZ4suoifeF+TkzVVCsOqNS8QPiJQ9SOBitLYcxU5yyA6BbNqSUGi+vna+
xkS6ugUymwUjLM20CLKsvqX/NkaNRLsHmB36FwFuOBGs8ZUUun7dhY8VI5C9Uvicm1nilFZmqhff
gUuajKAjqZTuTL9nxOsgjgufSnEBM0vL8Sxtq8AuzfC3SrVvKIH61sVQHiK8jZR2V0fbNmDVhr3I
uyyVbhQS6HXn00lH251XGDOJ+XnWycphAb9SSKNdM1BGlIwOsfaGmoGDdOHY0W8MKhsj7mNuiCst
7AyPhBLB3zcDf/XkOOx0h6OSSw+q2GcYPQwbus+YFKrVisZWeBa1UZF3dZUrU0I4xOPd25a+K0lt
2fqYMsP83c12GH00OuO4nGP8YNIzHzBlfa4SlBJkawDBCyvaWhomkowlvA0Cu+UjFB7GZWrg2VaK
fneyHKYbB4MA1CHgKz371Yx/xpRnErPjnCWfmXfif+95NzFTjaBMhUZA3rqKft9zBmNB5qCiRQDj
S5gd+a0dzcfcVwaT+nkyQ7EB+MP6Xv8GNzKVnU8ZpsqBSvgqihJqe5+4Y0E98tyzGckjyDVtjiqe
e8mYMF9khHbUCQxEBqxJur3NDNd/sOX73/r1iiyOYGvMW3V0KANLdpbGxVwRB3tbYj3t3gXQbVNL
LQNAeZ8JRl3l9tFDQIKJX3BFzlh2aSMwG+8uqJn/vxuGpYqlqovMppdc98pKl3RM6eDwzXijAcEg
LXW4GJVf1l7EWCvcuTmHpLA+WKj47B+nH58btEls1eq4R3jLTJ5crHzfN8f0hGXiRZZMfEP87bNS
zS5YN1tpCwwnSj6Jag1uUH7y0T/ix0CDbJr4TG5JfKy9n0GrJcOhM9JwHfjeoOsj+sy1wWubqalF
z7+/oG0SyLkGe79gdv3wF9HUvTpmlIa+P0gnEI0o/qRjWlXFS/qFtek5n4OchVoaWdSpqJDij7Xk
RB9gRjnUH5/I/KDcglE0imyRtuy2LtLlBfjxh8r4T8+vYc/G0/UeoGl57LwgB1u00cvJXMEubWtC
hpousUHy8iWhLWoCs8hTCQWnjgxpU/5WpF5eKHI/YiNTbGBbx8UR9AGtBUTrnwyUB+TbJHIsU1iG
PuT0wQ9d1fneXd7NsrCNdv3IuaJRCYZgVadGDHS7cKiJmaPCAGdQZRJmxLy+xn68ClTD4r7YVOgz
o3HyoPc6R2F0uHA8tq9fMrM1lAnkmMSLAPT/TIQ9umT6pTr1ecdv/3LcxqfjBgi/Ccve3iHUa8ED
SMx85JJOAc1BqgAyY3az1dmW4rEzJADZq9tuUxPY3Hd1t0YlkShWI+syhrP2+MhUtpYG3V7hppky
unQHFsPKM4LGWCWXHQk6c07t/5jMNdy+PmC6Sj/iU9Br0X9HQ8LN7ESK5nqvKh3j7sJhvheUm7kN
79WfqAPEG5FNWDdDj1+/YQCKcVYrIox3D8+2KlMX3SRmHRF3pAJIDwE+jrICj3SmXWkV4SX9m+rA
2NgkTYUxsYcOkixRMWKMS3TaZFtsintkrRX2TyMce1fuyH2R2OtvlIBFbNfQxsYsfB6tjURMyq6c
pu2KkxR3bh7/xSumqsfjRXQi6F1YclROQNvtGO3BaT4CmuIgXWoTTdqPMieao/hmlYKAa+1NFggJ
Y24MoN35tcBZwKRi0gZVCcNwmCf8L4UTsWLOHSVjC9Z7wLVw4uqhQLpndo1zK+3uqwunqCAEwwxR
lzUyL68NZAsSUitu+14a7cuWIOc2da4A3Sm6aw2IjrVcW6L1g/toWft28AvFMx4xVShF/4qkyl6S
OZcJj94nihwl8DVyf1yoiZ0Wsk4pqLJWLlXLb9jUo0HW1B5VULCR5NnmBT7MBBbhF6bfTaR/fztb
PFj2w6vBoCGJzdT8PuQBBfVX1lRZYmYicjPIc2WVyPY9zEhr1nZDD8N2ObUqdLUs5QqjG9fFssnP
MX3djOyFSHjSCvwKIPpTIYkoBjqhzAork77bc3+15lvQhPwuxV/TF6nO+wSI9bK7Rfdv01DvLpcY
fAt0xClUEPcSKNaE2MpRxxvhT+3oKJtkmY9hhJWrish7uLY3vgtVdzUATG3OVssmLNEvKp4jNJjp
JcRCtUCVCTEdgYTwwCfNAQgFevwHYDULkzhF+2PdDB30jhQBZFIF0kMyk6jESyF6dhvS/RTAosvP
oUDwRMMnEgwc0jZ0phO4lW9W0KAqTxANFrJKzx8mcH1xUniOGdeD3p/oBcusGcgAuRKnnYrgeCWf
VKW76WXjQ/JICOClA9pSjENX5rxThiG9RZ6fKBIZZ+aIdoPkZ92yCkAYkKeA049wgArgwbho+trn
W+4Qvmb/7rU4e1qjz1zGMLcfXldhWOAhVLQUDt9Tue6vvUj+JeFsod3ITsaki8q/keGD0tPtANsh
uAbq+gYHA19JPrg3VCXrF8AtDq1D0p1TPJNedyx7RwKWhIIXUF67UqpIaqDkG739eDER0q8FX9XU
WN8gGslj4EiFkihuerkYmXrZ/MjyDXYSzO2qwv9MkcdNhyfQ1dsqaZ9nMmuZVk1f/6AFwgH+QObv
1QU7J2InNiESNzi2CoeNqZ3+/MX2DTWeduMLZqIX6lJlNhQG0amDTblaX2MkD67NcTDBZWxqfnc+
d40cgMij/DE2nctRcmLp/Ium8OmsjtzONkg0Jw2t/pI7K3ZTuLZPm0TsQKlb00noxLH6PerV2ITd
gSYPebQp0RDOzGPn9J4TlCkBemNaHMDsLH12z427hGRqCcZBye9fHP1FTKXb47+hL6CrtXRbN7lY
xfOqlQUjJvFViGFVSbCST8Cdhxi2C7zBtf+rmeOBjMTWI8S0AWAMpNRwUdC26vpEtvcuqqihYzmS
B91OM7xp6e5FL4/nRPX/HTbb0WgdoU0aqEUXWiUrBgTLx4qx7aP5tEJV8K+RvpHbKHR5FVIlCLXg
KUMU+aDIprWGdkn8mpMo+CH2UKpZbvqT4b/CgP7q97kIqHL9PDniK3vaAaD0jFweq2mris6eqBay
z++KO1YK3+XMMnH9V5kB600al1h98hoWZ4WZ9qUAzzn1AgKbl7spSsCuf1vPnhVG6ZlFdfAum18t
Rel4EirzaLV3acXGAqmzS0kLBKQBJi87gSuzkV6rqV0phGwf+83FFst7aBG9sgRVYco8HcKvJFMJ
PAIeSrt+ExdIf/L4VVZM652vIn5EuSFslecZeUTuF5CgaHaxMOf/EUsjDrjUtHhfA7/OXQikLESr
mkX0JBNwn/+MSUTq7WXie0uJ7FuiiuxoZfNAj8FAu/zQbHrQVl/W3b19N5lAxJP8a+13whI7okxr
TdEPS1wMtKtt0cKYnAnVZOHgk1YQ0BaeqnQo2BvL14wdBYItTJ4KQmyBG7wnspTZFPd0EMe0Kurw
3h7F0Ip1FMxI2Gs+/0Xobn3ZvJcN6MhBqnDrdWuZ5YEix0TVMjALvuhqb+WWv8MLnAd2scsZ6Hvo
c9auF8LbLKWV1agvR+2qL73sLYc6bm6GPHhx8N2U8mhHxVhhZzS5a2w4IGiDqRUaSwTExJzRMH9/
HJKYEmx3cvt4R41ZugkRiga0jzPNXEl2jIyTYZxXttQytfRrpRZwY56pUEAXxgyGfoGNmiXYvmKd
677hRhkocs750wWJ+d1AxS3RU61HWoEQ/vMi/bD2PZQLc211PR08y39EbQoUkCoL3HKlPIKmfZNA
Ozu7JuH8a4aTQFeUnZQHv36BJzlB8S7D78Ux5jCCYAT917EfFQfTt+mHpSX8Qflqomn8/ZbWX+Tw
5VWdSvxBJJjEe6H8F4oYhLa8LwfX0lNo6PyJEq83hoSjURO/BpDxqZSTFMtE1GgtBRmLLRXnp4Qr
eN8m+yuKlL/3IcBFwp5GyCAkmtLQF7TctHoh0Hubz+2oOQUc60eHz56VdKzdVz09AfJWZzPAoRPF
JFNJkF3BbIIygXzE52y/1pmMuWFNmJck0o+5FbWoXR2XtgUwodeAhIJUQpETYD6FCth1Pfji4uCB
WlMhS8/IuMiYB18W9z3gDN6Fk+ShMUypX+Psj8l1tK9Pa1KyBjhSz71cYoO2ac69+fb/7JAj1rin
mTc+Ho8oe4smiNOg388IcP+pabJK4JfSawKyCqStUBwbxRMdHE3uCWWssJIaMTg+WmkZMZbcXU6V
OYMvYYeRwBG+vAcKtALXuM3m0vjYxKddrEnd8JKugX8Mz4hw+ImkTwzI90YPmvL9gKkSLmVJNbiW
iEO0XYvVwj0PtO0qkDPS9IEx18K1HqXJ/ZdYqPisEJSfL/WAo7zNEnju0JshVCQh0xDPZSldMug7
Kq19SykFjunu/ZgTXna7jxA0FF5dW+4tnTo4rLsN1O6bgzl0aOnekwmd19zJWAKz53T4vPydSwwj
n8EX8/3uROTnsLv6IZJ08Sm1fqo1oKze3y4sjKm9fhFCIroJbphq4gWm+RDP0v6Ji7lnca+dtKjB
OUzS0bqTPn0WkXOGz3Cd83qY/3r+aOZ9az0zWNho6OIMJ16iXm6UDPM+JqNRdzNpJQHs69tNMe2g
NbuGrrGPbcoPQiGbFAsiEWDehsw/lImkcC/XbsZmz/1WXQ541qpASY8mGljKkHlBlL707/nGGs4/
yqK5fuD5P85k256SvkAdSHRnW1vHlRMFNl2OhUHeOYYx3DxTpBkHMHKn5IOcT8pGX5UcWX0N6q6c
qz/I5B2DnuFU3aWBv4Ua8jJEOR+UyhMHV3x1whSANNzokUUWVXtAGec7lblGEOenLzFuzk2NyFnx
P+KLe8ZLvyMGDCDdny20vcT7ObwJDm6OjwpXhN5hoRougojz779wexkD9SonQvfaWwljrqAk08r8
sdGp/rMG9fFHcvZGzXO0DBldYdEaYFmkVEWYpLFPbpOEo78UnM+qABaei2hpvYnYNtgWv53seLYc
4vIqtD63UZ5u0sdG4cWBl62/HE198yIS1znBqeMB4q++ywdEaVsctZUzsROszPO78m2OuPmPoarI
PnuQtzIAw11r5fb0s0wZATgc39o0jDcvK5v5wFToVNeeet4g9UNre0u+C1DHRq7WixPhxEVml4/a
cqzSl1nz+nfY7TFuQHRXPCyYXFeNFOuLnQsTWHhkb1yv6FXjwNjFDzHRw4ay5eh5Z4oyv7kjl5Gw
xTwRMdwUt9WBZtHEnUzEdjbKCd0LW4KP9gMzSn12AJSs/klfIXsnjW7rVbq0QPJckpMIBgo+P5c1
18bFs9XUv7DGKS5xE05/iAaAOwbJ9zL15Mc+akh6ZaMcEgMhAluyIxFKO/fr3Xx2NIHhlkyz/D52
b3YZm9eIcKwXzBCBAdsb2Kl7VpIqL+pEYqimGLhWUq3yJeaq30W8UatabO1iu0H9BkGgzybLQh1a
DPdHRSLVV9L+yc1pghrL9z90JlTm9o860EAEKXU/LjAlbxwELDOchGJHfZ3H9frXPAdYpC2sMtau
gKJGb8iXKS7P3VXK3KsRvuelB+n/amXVQCaa+AYoPtk2BNgwzVN7ihsLG7gY03x6n/L6pIgsjmE9
HsAcxvxEgtCCK+8beGqbkycNnkxrojpKYtR7hkXpK1ek5O/x2n0VsBdZMAdOfSnUGKlGo5f57pgx
C7Ca8Tg0us33/aSvVgwS2o7JyvXPovUlgpwH65jq1H557jHXWRktKQWDBGUvUpVFKaApEbo5QA9h
uy3o7Nov6llhhlCgsb9914R/j2FyfDDDi0eUV1X7og6r+cFRg6XWr29dPrf5yDktu/GTkOMLy2qn
j+4JAxryNGqNWXRVckQOIwod8ZH+hh/y5CMiLIumJbPqalNxldp4pWAerbFFc5QwlpFELUuxqh8+
KAcOC222JZtC3M9xMx33PEz+4gFYK2Et12BcX6I+lvaueI1t1z3CpbvSS83usehHADk6lJKYcQh0
EttWynfbdHWdfcZRujyZn4pt2ItjeTvEIERrL6fUiwCnaT29DgKhWWx3UnYR6uThEX4zwFe0q+ye
CHuZA44e9l2Q87ab+Uds4jflhi0JLRHaiEKtqBNDvN4SP+8CWNrlpJMlvFq4XRikd5QLdr5yMtZU
QhGzDy0Az6VoSaf8MHAFVNSkUqmEanemV/Oijj+R12IWozjP1BM5q+aDKP/QW5Fc39RFrkTbAga+
D8zhzW6AnGy47sxHVhYpa/FBihhZ5DJFsv+hiKTOo6yVokQWBphwFpZVzbgmjlHjuLWKxW26i7Zt
O2ZYPeB8i1/UsDNGC6mF5vj0AEyE+Vg7u0dh4BXsZWn8YCIEjP/PVpJ3cIhvf/cuvwSQ6+hrdsX7
lbz0Fr3TEjOwjcWnPI3AVFIoW9MDyITfbKdUGaj3iUyHP36ADsEbzhRsK1sB4Sou0qbKRhFsq9lQ
dzM7d1Pdq4BbKT1FwJvIgBoIKglXNx4Dnm5+BMIxiNfje3/Kt+XhIwadiqiO7gmvCRwg3DX8Nh17
jmyPUMp9veFGZsV2XSbmikjIyO1l2iZTaJLXbjps/fgD5jjicwYasTuPYzdvGNzF0U0OwWXYlMtF
QKQmiO87psdTamZbSfbRMH5c+aURByCbcObB1II9JtlULRszhbiTRHgsz1xpAuPLExC00WMt0+3G
72CJzK/e5bvMhJeRmpOjhxpiWpPcUjacu8lqESQHjpkLiwOv5lTstsewL3nJtAGcXQIk4qjpgzbH
UGRZgV0iOs0muV6dQMRSzngXI2lBIDIf7YsdQ1xlJlHtc4iBcUxBRJhOCdNBkzYjLBBpqz7k/+Yr
s7YnuyNuHl4v8ySIS2tUJmHInnr+O52nhV0FHyA9aOqI/6qdJjtZfO9oVhvzxyKUML4uyjbUlEJG
wcNRhXOGRU8T4z2Unihvip1EY8v3Was0qWGPeS6iPAsIe5+D5PuuEISw1sry7za7rKs7GeYAl9c7
80eM/dg6Kr6ce2TdcuenkhXU7nK0Fd1rBx3NAg5Gx8qGUG8gJgqOOED4xMRecbuTUyQTNtni3LkF
zqCDkDkiABRj7ZQLpR/DNZHYftcxZJL5Vf8p3h7ylR6llB3CJj6tNHIQEnRPpMHEICI9LOHiCqRv
kcjahRchdke+O/1dge8h+eXIKlhXUb/oB6EGjznzHxzDr9QMoHzA9TEQU+D5GVdU6MR04LbbCi5T
uU9eQ77Nj9wtYiH+5dHThNBRfUGfw2APGF5Piz1YRGBj2Eho9UG+FiMbd4JB/bFCowbgiTSAYxuF
hCFmQ0BL2ZEpCx3Y20EBzXNqxPXzXPwbx/6edwdJRhD+LT9Y4CKOWwNu9w8q0ldWZZVPjrqexmbh
qRELrTOY4jBcz5rPnQPZZJ5xQKo/EYiKaMnZsUWBz6GwQhGfRD+3jJEK4xQwFWZ3AlGTpnluAZd7
8qZHb64IRuMVbmuMCmf7Ypsl4eVzHhsD34impWKFdOFaras8O+o001xMHcQQ/4UgUbgrohriRVPX
yl5ZepzYxwVnIP+1Vx+ETtWfObHP6f1eJAUxfS863kkF3+CkpEm96t18C11YhY/eI5Moo8kwaEwl
HTf7lifaFMMN2eO3MTEdRgcnIn9W8e5L2a4VC+j8Ris0OpxHPUkeSLOH9BUv5KhVdkbIZ0YhQfAm
ANQyI0qyMNHjeBaNqQaSmxBTA1ItQjsh4glQZsfI0wUDv7nb1O2EWJIT4f92FuZmAGSm1H/iHozj
jzqoxzTwGBqojf7s4pT2BxZJJbTFvfRp2fZ8ygS8yStUNn5nCHWUSqOLIyH9GYRZ6yn3jymBwIY/
qfb7pEYTK6cSu91d01mnn6mKqlol3QxQi6mAJhz1dXxAghNp3zoqtx8Ic3MFSy7k0xODLJS7pm+K
TxHGomos1hgUHuBPujjdiOG8MvpHHtciyLZnVlFWkJlG3SoLcqgbRhcnw/odIXDvo6Y/zNUGS7fy
Vtjle5dWXAfRr/JsQvTsiV1nRS6EBq8BqpWtzx5jRqAf+Z8tMSByZa4g42AxGUmHth8UiEXhl7Rq
BMVF4QvYmJiX09IqFTe5kGJZUWbVL/osvdLiohJCGKimx/DpJz+pjbhNZ7fHJ8MROFTV79OH+9mj
qAx+Oj3dMyi9zjvdkZ7yEPESbJtBxeLK2UV6O2S7ZK/PP11YQkEEwBGuZlUKBC+9IAmeFd+OAko6
2bZ03L3JZRxoLTLRY7E3ZXqhwP7JTIceBBynidvIkDhq3z9vsRv3oj382S35oUqvNd1kh44okqxR
Eyp++kOolHIi0yESB7cfxZxbUD/g4nx5eWpUeC34a5GrOgbfLTOjy5z2A44JTQnTikZ+5ClRHC0W
QETcg6plKBjqDE///ke+Z07hT7bbtkQLKpJ4CVJDEO6uTwiA2mapl8VgektEFdiUQWijAwXTkiVX
7XF8OgXadiK6q7HIYoFBoBgd3IdBfFYYbEHr9xWltOVVQQC3sI39OGyG/aIxss43t0rwjOsYBwd6
QxD+dQReJ95H+x59L2PfJT0LpdcJ9WqspuCKBXT+eZ5Lp4KGX61hO4SXW4/I5VCDTJll9WgJS3BU
m3zlpRxM7AU/LIVDXxOaB+eE+CYxLHyb8Q10YZRm9nWzJGpW8GDEQWKa1VvZO6SiX3C1QnTkhPBj
0Uhd28Gc5T4+p6Ee7kxr7FksDj+ObY6NYPYqGyy0tBjW3itSxnN3vEcNhE1PcmHJfhwdYw5oRVkx
aalJ0+IuwYRf7iWgJ64rkHktmEr874be57I4KUp2L9hw/Tsayirm+Aifafujxql1kSFKwY5CUkCB
pPqVMTNP69E4B6kt9HnyH4guBlKDsQ4IL88VxGoCOIZIpd5ELZ7VXiyb3KYRDxYzVjvfN5x//KBa
fek1DtrAISHjAm8ZZoFrCn/v61tK6gOiNzEwMq77Tfm2DGKzdxRuUqov90CPMNmV1ssw0wXOXjxg
Re+SCgxz2P+LRSyqmoeG0Rqs4ZukhBADMq+mJOGq9wS0j5nO2vQkX/mDcxu2Ejr0YneBLPsAySKP
VshGAsXrDLTe4pi9fIJ6E2cMx/F1F5Qfkp3LrJZpmf04eRoISOSt4wakS2d6shB5IMB7ng73BDwn
hxXTL7R8abRHSLGBHH4Nyp9svIsyDFB9WISdDFcFI04f2f9tfX5YwnwWb8+aABw36hbOT2pJyslE
K8azr7e/0ev966Q8RhJjkt5GDwlorzFLlZsAFBQ86SWhEbC8labmBtMJn1YWS8/V0tJym1PnhfzO
wvq6Hb+i946tYYCWjPv8vBuc2+rfh+38MD4pS67J/bEN4kvhMWz3CsNJSPe96Hk9UA+r5LfdEpvl
UOf06SIx/k4rYukuV+xQyDVA7WeON5YoccSlQmexhygu99NhN1KgAzbK+J/2yxY7Oyod5drrvUKH
+flx6Vkz21NwDl53SNgT6rNTiDDH1WZ8ZsnHajwCrcuc0kh2PBATFewy+Adp82iRegIUueeicHdy
21p3n7jCPtXIgrxww48+lu2LRWEDCIZ22cpJz97pNbHKdoHVGCD0RjgjCrgXyH/8VtxdqPOOn37I
hbQCQrmuLys2fM8Q/rB4gSdrT38B9lZ+2kTDrX+1hFF479XzYcZNdwg8JsIO2s+1N17p6sxvktLc
oI8UAgKaUO0k0/tNJrvhM9qICVRDaQXMTXuBtu2fHel/JYrDKC4dV6AeuTh8Q221H/eXbZJx1gj1
qbcsNV857zrAWxISMxhIvzUHj3nnSRXGWm5mqb2RK3XW8U1wQPJf0kF+fY0pZISUV1LC2iM7/0SV
nvmM104S3Xhaw6C5X/DKT8BIaIGgycC08IUgeTH/2lWMr51ze8rcMhX+2yPk12FXe+Wl2eH9a9lQ
ZJgwtufd7BGX8Rte1LU2f+Z3DxCLdZMLEalarbRiWQwa35d3wJnXZ7QxPp7cI1wEkPSFLHLAb/4i
Rnm3AmET528CXDrMbJJSmOdsJCrwgzz1doKKrAgJDjiGTQt+R2x9k6KKOqpwftAJgOyO+lB/DWBt
FHO6y6GjplEoh6g4Z8nEoPz/PvlFHpzEZ/1EZCFlfWZGnfnIipkZGBPJyi1HfpzN8RqUGBx72enI
sR2PvRzOuvKcrFUcxXlcOjxhPNOwpxDZFgEzH9YTFJLpKo0Iqd4s2rgJFyv0cun6YTjs7xpGJcE/
49w+DL4vRRlb1YDzOSLc1ZJ/WmQFH8m2oKlG3I+KfMAjf5IkJGVMHKrqzI9Ty5ylWk55K80jzPRX
PbjincL5KfRU4JOclZH70r9sBzWYTOKWvwsLbDYgbMNoqhtHtd4stSEulWyQVgqG7d3pz56mGqD1
gSvQnfoLteOQjuym2hc19X7ZTjfN8qwZeyGlW5pJODTpKtLKrojIxkFkciV9uq5vBL0E5K1e1gJF
YFbtwr5oFpOLrr53G+i41ktI5sVx6mbDq7EIEnSVYTa3/XYhAjwNxY1Dl8RTHfcdYSyIz+xuUAcM
3EgBBpkWTkx9xdnLNc1xKc0dS+r1OYPauX1ubrNcddknc+pFcKaO+Vva6OWYqB6xDgp5m+U1oKg9
Xm/bWHaK/KjbOoPY8to+0PxJLqKsV8Rqs5WXWpcOd211dBJLMM4sBjhc5v8TzFOZKRXOcGoZqNsL
9WFZ7p0iPiHfNyIu2w2EBVkHxML4Its9DVOf3lVot67frzawrZR3uNvWpwmNOXy7h/qKuL8d8kVo
w+YbsUdhcC34dEMBUuBy6ZfR6s877kOq/TOybvkJLfoousuu3/7isWxaE1fk6uBBFKJ31D8yZcDi
nmm9YzKwWwTX5JiaL2US0kQgF+DlrJuwtWB20IkTyQzxiHrMdDZyfNHzkVLeQvxnN4m72Q5jWMsW
ixgwAOxFWJEOdzs0sk5Gh0q7pkno6SGm2hJ8pVxSkldJs5YcNxn9YQryTP5rKazpP42LuQIJnh9j
H8j7e/1sc0MkLHBJfnAE7UdOS0HSdrielQFfBMttXYuIcyCgBhHePztS8HyunZgmRTMj/ABdhm9P
0ZIoeMm3wqXsOoViawzRkxAySnVgGUVrgILTl+HL5I8f/QZat+mZ0yUjH7tqCxj3Z+4csNvwXH8a
2Ta87YWiKhWeBykLcMjFHwczEARz5uE2vF4uBS+fUJuP7Snu7YCGP14ZBXZs6xXXBc582o+oPoOs
GWRoh5Ge3d6FI0QqmqJCCVhlqXhMuxc+OXkmHALsjdXo088VKL0pTVaa/E0zY0Ns9q+SiJ+F1/uM
m7RHjq2pC4vkbuwi0e9vwLHcYwJQcvmma3WArziTy0mIBbGtxk4UMd+ZJJMdWqFz15MRegK0To/d
7Qve4bqxuOKroapnDL9ZOJWMfgbRtxQs0E4XjrJbWcEidtmW1Tnn/8pPniKlMYlYIFtmbVhYXkdI
SV8WqZVAM10Tj5nFacgHOl9oiV6WE53tdcBLFFSsWs6umRzBt/Pngu5oKj4eXV4f/BTMTytDtJse
sFHHPz9dDydGhlg9Pvs8Ybn2qVGO79dvMB4G/KywJJrHDKqmZFefVZeCdtqwQrSeqvluFhbR3KID
dB6fZdUWrSlsMucp/3U9nCm1cPdzA2l2uv1gKv4n9iGh4LLpFId5lqgB03t78xKKU5pEhpe6hVfw
kSKUmmO6otMrLWubtYIfABlbQMg2unz3OMvpGex1vOhvp3CVAb94JMci4ZIx0o224ziEpf++VKGl
yf5CPJALRiH053F3ij2zPl8LJxBkfKHf8Cc8bK8eeFY75jiHO8Stz9ha+2bvHWr8luPDHXS7Kex1
EgKS5GhmGbsVyxVYh5x8t3KyJksOTevslRlwe+AyHOWbW3EgnGPCImmjWLTKk4bZmxeWf3NTdDZN
w5AroX6mwL37+t39giA0v1pNn0xoKmr/vdoXACdU0vtfYu0d267O1/w06hTkVvwOwAViIVy+BQn+
yqUq9R0YpSlUxaVuDM0AlG+oaDGOU5A6Bvew0B+JTMwYgWqfryl/31B6vmHkUGrKxdS1OvhBNNuv
ILsQc4quL7MvCtn488fRSEGTPHl3obzV2luY8rr7svYE+LvPNZzvJgCntn6tNZdCXZHA+/Eql+0r
UKoyTssd49kBP0EgSraOZb7jvso7/ek4/NdPrg0Wf16O00RFY8pMpiLTKAGvnGyBzVcV3K5iaDUr
uztBkEhg0m+1BNghU4jvevmtdL5mNMtyYaxcQ0TqRgJWohZq06ojpzewlSFRN710WxECV7Sja1qF
Vb0524iSebiaGqTgXYO4qmqPwv+uT97r1KyEG2biPWmBrtqdfKNi+jXlkUcF+3fbp6OTcB4B4gxx
Ams9HCA1/z1SSe68ZCT8YLNb4Mqnl7+G0/e/VbDXPPz+KnWwl5qPYRMAgu9jiMYJ0bHgv1CHxxsl
y5T/MF0D368xkdVEyVch8zzmYI3Ro7DEQdtTnUNqOyoM+N5K1bpBQtdP00dwCa9MFiEfz1+aMnYd
3/0r7Mgsh/cgOqawV2c3Y8HkJSFKrYZbMI+s8CJ/dP/N+2jnTjbCyO6UhWZrsXAxtLPzBQQsFEoH
hqQs7sJdY+PBmzzU7iJ2vwCYFeiUu8ZazxUiPUqokrpB+UZHSA2j3Xja0oN2u3eA/hGB16gKULIv
HOkWbXlzOL/XiO0ZI0q9sd1h2lecLuw7enEyigdpFYZhM3bjj+OkB8O0UoSrODZ/su6XuIvmK7Id
9/MsFiwnWDWiZ9DQEQrwDbc8pj508ImbTqIJ55YqAHb6D14XCQxdcBmcayiuUh9a2jVUcPbU3KFG
Jhpcd6Hcmy6cAxPKHwJtqPXeIk44V53fgI5DjNrZRboaSrCgldqO8UAHgQXa5/iQF9MVDhsMCsRQ
t1qz2peggTaFoLHqlnh2WPFAra3XuB9qucE5Htw4P2dcWR/iGGHxKQRtX+93Ense2pYu/VCf7ddx
8M6Ar56GE6QI4dkc3RThq4M3AYqM+36YyXq0lEzNT2TrwJ9XfmXUE2Vy9LfzjDDYdW2v5kmzUx8a
qzf5Y0cxnyvmm6SyMDp8DzC+2m8V/gNonzvR7VLC8/3A2J/xZLAS06qV2QnwWt0h2Gxoh6iFeko9
O54otmBfZ9mpAjIvVwI1DLjPhlzQH6aS2PY6mMSqdEhgN8253q7Sa7rzYEjYhPUcAtcjCjt96Hnp
/PQb76ey/pvbgqfuuhzSve9ZqZMrBm/RTF6cczv/yU8CUP636bFuz5DeHrj0BOc/QY2EeozWTMhn
q1JL9vtSR8L6kZJEgRAKTpozg4cPWk8a7i+0TrJDcXIF3BWXNNYZCB9lt+KumC6ezibCxCxkGhuz
XbFb3tfhgfPou7iHPHQkewZ0cl1Q8D8lKbijQcSsERVsqUYV2ppca/tu4xXeBUgO7g8DB5YNcu7S
KoVBV0uNJkYWV71L5soSYpLagxmjUsusDM1Mf3ZhChY5OCo2mGE1MlLFgt3SPEF7ScZ8QpeldKc/
U4h9EfD2Y6dlshLOzBQNktd4j6d5AeTIIMaQgFhJMxmkCoMcKxbtF4OXe31h4IMexV8foctTkwfQ
c+Ruk/lO8l5ZJzRuraGTbRP8/zbr7ORP4BDj171+PK0UOTsaztZeKgPOTHhiee57AxE6scYwk8Lf
YFGBafk7PLbNLAaTsfDhfQZ6WNA+ItLfbitoEc1J7t4YgFm7TWhhz0oCjUMANLRvZjgtyVMEZRL9
tUzpp3VH9knn+7OY2FRBPksJyHlGGKJiYS/6o8DsemWgcA11RNi7YgZ5ig0+W8rbRsOdiGr/h5Za
zHmu2cKTwD8lI3VBbW5rEQhbuA1hyYKBjGWr5w3qC0neZjtJJrU/ZFzOguHCbkA/uFJNc8VVyGd8
y1lTU7qyRdMI5egFfPNeNZNVF1OtV3RvKcRNuzT1mtqA52pW3MtXVkPodM3A4045y3V5QVatWYtq
AESZBBsts/QBr/kj6hkc/I4LHfIKZOcHHt/MQNlw3WJoBkJEFWetjIEqaqszDXsa+h7dVaabDCtr
ORm3dYt4OhrdhJcotPgKs5vMVF92R64bKR1XRPgJ901T7VhZARFjOl+Il8udOrlHD5AkX6gcDwOP
FMTh+3I89ZtnDZKhtPfE5mMXp8mEqqyBUofZF9xeG1b52dWFdJpGo4ex1FtoIiNRUOOtdfieNsKG
5GqQiTqRxfp1wrQyWPsslwW2SuootBOlcH2XkgIOwlnHxJ3mEndiuRU07PKBed8HV9595rRHcU2D
E7INoWBvqSLbcpx2TM2czKr4SZ9ce4T9SyWYeGSxGQfBVmWOjbK3kwQ7Y8WzXBH58roiSSLRq2XZ
XmoVrylwO3Sxd2OQat5hl0V0Fn85g/7mUr+jGQZA4ubp3rwRe3DAYPQgHKgikTZzCJKSh+2FkmQF
JtPgKG8DDJUfARlYfphoiRKR0lXk9vToA0Itxsl1yuxZqf/oeDlvTZXHuwCYMdwarG6I1aQbmNOl
2GdlRN5+h+LtVQYm0HFnYbvUEDCqGcqg0+1y4SPvwNGciEVtPhpshfX51+fn6pxLY7mc63KPwP6W
2UYTQPKedlMU2Fd5BIfF1S5O1xjn2Q1jwMu2dQTO4Vka71huRANdxqt3gVsM118aq40g+/aPxwGI
YGhviLlrx9Dv3taw0cquJ6C4ZTOUeLGjTm/Khk1BPmikVUWMaZ1Kr1c8yt0HM2U+GCeN6kFbCWLG
LgmI+HxQ61m981+7xZe+NBLlFQDNQ+kL0PooBs4t001KMwGAfJwczHxlhrFnCNjGJkf7iuG8RAR/
5VvzqJLSNkW7rNful+uGEev+XrU2+s667OXE62mG2WDzRfLWTocUfuoNHQS65Ds1WCUrLGL1XN7W
AGnOh1Qx5fw3kkiaz87ptLJeCtKzEVCL6KxGkcHuGwC7VPeiSrgYB7pVwIKTYm9UPP79M9QGpZBb
r0vXpXyzwCk7mZygBK3bFrpvzwCFgBh0h6gU8vdHyVssMv7mcndKyX12YO0dQq9XIsBAo/xtK0T8
+7UarlvxYeucUytNseWDgz6ngl3dbYKRnsE4HKh7SBl/S+mrScr/NHFqWxxMruQClK7j0VbmnejA
4/Bz2Endts4+i5jtlYW7tvVqYeLPeeT8CYrrdRfVhCGLXVATfIV297WvmyLf1CM/4TvDze69nc5T
hmMTEecAOq5r+yrqzf3GOe9RePM14hi42s56UOvofDnnNaDqjEgejCGy/ovR9idSs04oyy8R2qhu
+ZDWZUQasC1+EagsVE1WTnrGVkhOD0Vzv9LmLgKcOSPS5Q2nerw2fRceJKfkxs6RLvLRv1VZJRl4
OGrD5hY/Fr18IMBOmo7lBZd56Ka2DMQc7F9Us8A/0xcItBscO/qmwS6J+6uYnxS8FfvlVT+Dvt4O
DnlSDjgGusv/Vi1maIXpeQNnFFXuMnEPndFK+7eECBceLPewluXXY6yD+bmzTXhyDmWjFE6FXy0s
sbBZBGLhKvVFRJMKK7Vd3e3sxS91BME0QT/O1hKnqKIR1y8WEPOVnAn31QNUXklZoGTRX6WNL3Bt
Evme7LF6iFqxehBksKKzLXyEXZgJoC5i+V/velSeb01QZc/GafuABXuT/+2bUrPEOyL0fWch2Hih
Wdkqn10gnXN9nou/9p5fM4nULyKnfGv//Y4mGDc9xjE2/2GvaauO8PHqfnHr2sr9HmQz8pAtJPbw
i1BpTVFEiXAFPhb4vtRPrf2zaQun/3n3RXzFfWqXVOLky0noCP95nmaUiA7mGfQZIhBsozCtgVMd
XDZowT8LQtHBQToSOsWk8wCtS5uEVL/SG2NZWMLKad8Vtm8VCpOSdfr9wWWvEQR/3fAdcOFc5TPp
k4nqKN9wqOyq3wAJesiDexpddY+jN9IbVqgYd9trtL+nDxlhVKWB048w4aybvHJtrQbOGFf8T0GB
IjBNiXLTh6a999id5efWPKp+Cd0lZ/cvICOQ3DdIxegY0oafFfgwryxSBDQ936ESU0Re2r2sEoTF
4RzcillaspiddhpiQ6zD/WOopVKEeDc6W5pvV0F4jQD9PXThR3wbgBsqc+D+u3YK24vfoD+OAwdH
6y43dV3DirSyw1TQ5wHHP08y+eXHtzRBj34kthghtVRg2F9jwv3mUTzShW+ZWM3Icqus84h0bYG7
XhBn8/oviVS7M52Dm7U/oqDyH9D5rBNVT2ih6or6c6b+eqwQi9B2b0jKHkdMnIAmVROx4La9S5f1
ATwRKbuFO7lE4Pqk5tuOkDhwxQoNKuqydKrB74GB4Sqs9Dn/6F7gxVkdXbATtCzqsysu4/kp5c60
wuoNkmGf3ioGe9daORwK6z30+gVGhi9PVUIENjYdDPTSfs0K3XVFwkmAScsTSTUb+OXy866G+O4L
XwVLMGohxsYN0EVxrOHcwNqmJNfrXIRdJrTftXEJlyKKQASzwy6B+BS1x2PGRR1KBqRaKaQpIhoz
7SL8AfqkpuQhGnE1zARtpHlQ/f6u8vjLkRdUx5UezWoMhZzqfXQyff9NQRIlBJk0MEnCB60hRPLf
3wvBezVuj3HfcYyX82cgLYfpyPyrcvswrXHaxIW/jm56NZgzFtA6LcCP+xLR9v7az5QdqHBr1EKd
q/HRjDTeKLvDB3En6hBsPcVlAEPrqEYFLR0MObYOWrsN8BHm7fk/+x3PnfvvOaXVX7yV+wPXs3lF
FQWq6F6G4FdqF7dKqhy0JJnj1IqTbIidw3yIBTJn87XG3acM1KJjucN7xB6yqN29MGnz5gtPczLw
uHgfM//z79tgcq0+HfIcCkShvU54CyHpPE5tCPT+56iTt3MR4sp4wj7XSl6RghDBYGNkMxFiY9Qw
Pjdd7klpkYJUw/f8J71BQo7cOmPCKfLsVq0gucCNMKv/dIuCrXdx7NHjVQQ0fuKbZ9oj3boqzcU+
1tbLF0HrbdX/Wij5HfO2R070hxUb0BnQYKsUTLeEiZgSR7j8/iWSd/b7N6eb/WizW85Ls6iW6ehm
pewE4UcdNE5p/7UBTTCp99DCx54ek825iKWGZwK240at2dxUWY3xYeh8yXuLqX32cCPJfC6TbAX/
U1hMIxok+Wfvc3q9M7xMSWmWG7N3d7PrxaiYQwwwXbpNrEBUEOPcsAq3N1QNiSA4/F8IDiFNodUW
OzBIMamBtU71EAbNWimN3hcOTyt6PqILnREePqNRe5dWU6IZ6azl1G6KNFN9qViCDaGKLTv8SVtW
n/CA9uCS3fgp8fJQA/7+HJvhzrJkClPAPHeHeTRl/vIKYkWV1/W877hi1qrpXGZNeGHQ1To5m/9d
+Mrb+UFEMeqiIqUrQd/pCpynGwGmKq3ATEkPcQWmJaeUrM9bCb7YfuOC6T3kiegfF2/Uwq1GPWQk
rjS1Fh6tzYmIv7tmsiSO7Gv5rGXliUlCS/4oTUjqaZ5Gdv1De1h0fcz7JZ5wz3g9KkAcya7r8ey3
FoGTnH/ASjKBjyjYIbWMtLnqA0sVoD/hnd2Fq3CTwOGS7aPHDdxBvsRhxRLGGlhJZrMOa37gbb0k
jBz7Ftrlm0spUvsNvnQspXW0hlufIjZkeNWaaSTLJP3syKKC2lN87/sEVO3ZyjcTLblOCVUNU/pj
Sc5qGOFxqZMZbu5LWLdBHr+Ew+wk82pPEMokzYc5mnRNpECSvy5aicBmcdDSJyZ2iZ7gE2Vmbmd3
eGrYiaPg8DpShm08ybkPwbTvgj/vAmgL+nRMdh8S8x3AglU7B9mAFQ9GrwFaCeLSg68ccfZkh/ZO
fmYt/a0fBMIQK1xB5ojYW9PWFnRM8xeo6+/qzIS8v0gBNo/yHV5HRw2/yVccEOqq7V0HNxB2jZjW
cLfoTsdkkLdv0nfa0Tr7oTAzGu4YlMwRdvG2C+pziERefgWAUA0J+Qf+3Ww5jU4zTdODAx8eljiw
+FbYKzK+nAT0bvZnMJU/6p/HwYoAHaKIt8nbsC4Eexvw3hzzDAqE7zweju+kaG7ozUdDl2YE4wSk
6hHjy0sBAgsI628hVU1JsmCaamNRS00Fde1//LJTD4JWD65nNAy8yHXSEUc99RxOxKQcRmta0wJ8
3HOooX6j1y2klhNdds2x73M+z6vlHsMa2dWahRqyyVYAYtL5JO9mxqctdrLMuLqP9VDeeWg82TC2
52TAW7Cbv2rN3RTTBV1VcByo8Gi2f3NiiFWmrgedciCbmzi/oXzG4l0JlMMf2RpXi78g0TXevxFL
pAHetYm87svktJUmBmiz2JNY/i4wyWRPeE+hzWSmWgHz1FRAakpjXDMhhqacxi6y9gp8pYGhCCzI
yP9yrO14U+eJXCmjSa79963z3YexRRMsc+RMaoLfwNmemV01fBuoN317jjwnyXqQ8T7TU2SgFy6L
2+vn+yl06j1yN6PidF0Q+xyLuc+MNHN5WJRKhGQWlIfVqwPXhD6p4GeuEodpwJigqMZxe3Pf9B2S
xavEJtElU9VUI6lmcXq668Qgu1KAOHdf+Cp5xth3LQ1Lb/hpY2LOn/qdsyTOkbU7FvwndJQsTs1Q
bUcIBUqzAQcZKEAE5McNvDm580k+QnCUbsJFylCpes8eaSHYpd2PCfhggCgtbXNWhFKSLzaxB1Sy
gtNU8m05KX104Yj6mkPw2JY/mr+wfb/y03AlEqudIFh4W8zTgsjOpAQs8kdXnOxcopi2hvSrDYgA
P4DVChk8c9LLV2TdxaZmB7LncxTM1Qs15EXd1v9H3BKcrHRVlfbUm4S4vh/9DZIRxSzk3aXJ6EF/
9i5TSLxzzjbpHgvVbwXu0miMUrgRYdiVr4CuzD9qxDs4h330ggBOVUDMz2CBRFJUrPjbNeZaRini
uO6Cn18waP14cylGzppSqmH27nGaWpI63dCP2XihGZJz4EEwHsIZ5Bv5gpCSHMavrmx0zHTRd3lz
788QizmeW0AxCYoxRuwsKk9dpO7u6ELK9XFRnV7Vqdo7jztnuHIF6dE1cYyJcxAIpyVmrAIdtnWa
SvYW4Zxw3aLg0OLjwNIt3AyIYRtwIn1plXPqEIbwsXvCHOTqkTf4x6YVhCTcrVdxHlhDGXIxKh9v
SYdidDA+8QhktV8Alg4045rovmPWK/xncV0shuqU5i5qFvLTXzWUn0+yDZxzDuyB6xGxNH+2++pc
K5Bwje6JJOhF8tj8q0RB8wc+mEeBY2v2yiAFO8hCGkZ5XG/9quTiDe02rx3aY+hbLjD0LyZb3UcF
OIeZjW9aIVbXH98G50lgoWK9Ikn3fTV9nJr6W3ijreCzFivyRpdD5QszB3ImNc/WNGLUcovGmjRS
mlqESkmxPxrzpOB6NWIctzWyct6h7TtwSi2A4ERhs8laIXazFmE/mAW7rXokE1rn+4TfjmWDou/U
2GaZgCsk+rH6/OzGnxLTtbXusQtTl9vTxAi2VVTgAZsgKIFkGTIKjNl2b79b0JacdmEBtUBYS38O
KSfUyXsaG3LbYRjyp7J29rKcjwJ0242i9rGdZvdu2VvelpiVJUE94QquvLllOl0d2vk1OEPUpSbe
2Sn3k704MG76SmRgKcxfw0guypZy1vnZgB1OmtflUX3vFgSlTO4pSh7b3IQly/RT9BXzJR2Z4iGp
7LU2sZ6WSggN9Cx5fxWF9EoPKy2skhB4XBfzpWh0qCVDARH6/ByMlsbHTk0DmBgMZig2T/hhYuzR
INo3AXyM4qjXm0LCzZVKdLs69PKMZdb6iTEY9IuEEUorQgXQdgCK2XWVrVb4ORmEAeJAi9CHtrw1
coFBoLZiLy4cVD54iFL1t1MFq9vjL7g3JdXWxHvvFxgKbaWgrQtjw4Eg3NHpfWZ4yDvsEFClAPwq
PD9CgMq9OzQhzgXnM8gXGNYnOn5rUXNqlVkDGUaXNGWDVTYouz778Tsu69Y5SBoB9e5dt1l8A1PY
T63ICmcoqGbYI4+QgGwASq+UnIEeid4GoUAtaRLdhy6+UtDnFl3n30R3k/trkaQb7y2xeyiVH3OS
4CR4Im2D6cY0O6tJOmmWZNRRZP1ZjwdDeQbcvCM0Mjn834f2UXB8S2jLQgm7tnLUR+5ZiKYkq6AH
iIjpdbEHoyPtk7TRgpD79/9pyL54k3PKBAVgv8Kh2ZndrRCn3DFtl4hZ/5dJgyhbvC5OJo45UG9a
uMFXlus+0JGLVMbvGKzo8KBC7Ul7sJArQR6nfoKzZPj8aJvnJfz0/yH9ue05a9KjMNmGMknEl7eC
XkJCCqZbnSP5yreVZnTIBoIqMqrJGglDskl0nb9BVldRiLAzslq4iDiX+xXPD69ocpiI9JfdGKHN
gm8D3aafnPtfgJcH7/fHoq3HZNovxNTtp5E1wyMqWMFPNpeY4n2Qh/sJDFChNh6vRd1NX4lfn8dX
qzarvDmGJLgdCJmKdiTW3W2yOBOHBRkdjR3TDn/hCwhXUD6y8ypRBnNoHZmPguA5+TvoKECxHbU+
cRSGOOGV4QYLbZDyihOyKu0MPnrQERaGO8KBX78UwzEB/joNcAzPAtPXz36glGZu2KZn2vawtzZ1
sP1rY9Ht+QL+09CUUSj3eTZOxlSRrRT4/DZrUIENfFGUmNeXrQwnJG4kgseO9f8nAcU7ZPtSXuZb
Qq/INxM6aIqdMJ+ReR/P5u2czJh3IOIc9JRHpegdIfu8uFaO4g1ICJmJTlDk23GqkNvqnnhNZNhN
peryMESrDQckHW11ok89GwPVCmO+6wFCatykZzuXy4XaAJFTHaIzGf1EFAhWQFkFWmddv3ZraTwx
xJ75OOSks7u0hApKFUYHdpFiafMjU/Ns2DhA3vGdyIvckt4R/TKz8zYswJPrw6PTQivzCHdLiCJj
rKdqxh+IlPRGqDhJGeNHXLjf70TcQmy51xZOdSUnYWCXD6LAmAWSiYZayqdPIOnC+Oc8LB/M15TB
HyhuR7skMJ7WTVfsRjDwOTlbyLmhrZCKY6sGeMO1cVcC5v0SUzpssPVLfRIJRihcXfOcqEPVlszV
4EgwKFeGG7mKdsUSFP1onR1rVx+yFZ28pgYT0QWKDFCf2Dp2R+v4gKiKzg4TidI8y3Eb35J80+iU
/u4oIGQT6k9MdK4FjYnqIVaZ/j7mtauWhTMgg1glrow33sjSHDBZNncivQUPnfaJfPO7FgZ2sEvQ
0Ge3TCS4TTuZpUZ4YYoZa7QbfzATkpsAWJAj6//C3xVlZmrugTt6lKN9NxJP6n1rKtY8ckeZ3lTd
Rpjqy75RHNfDUTHEPw1bk9mtsW6CjkhaIdZaZhtT441crPR07F2oiDV5Chle6Fg6QTZfqsoygE5j
321FsaNjcUbS++fRB88+LAQ+vdc8Td6W1wO+hhZJ0mHvnO4MwTHgSEgJq7uKBqSVIJnv6DK2P3o1
qa7EEhAEf5zM7Hu+hoxrobuybtySLgFDnqYpA5xRjmZ64s2catyiTTVnHRTQHGPxBC94oR5po5/+
wQGvUG/zl6bqVt7V0t2LOjZH/ugebRXrKT7QhXhypviHCABSlubqVpGycDj2J2wQCcvWeX1UoY3c
DlkesZa+eA8sqye/RO45fR3TZ67OnkRQmEptxL3bUIponEPzkIXgYXFOJMVjJNsh5tro3Sr6UPTu
oRNI6CwumilVHNNSRtFOWNm/+5iI4YGwUFEwzHZuEttqV4DlngSNSuTu3RxeiArCPQ+UpwauJoWa
dq9OQX4gLvOuKkvgfD8V62+D/e+RlfHr9IvpGDdusJIQ0hahaMXu0nD7e9TOC0Z8XbgbEEx7FpIM
Kb5dOylq/q9Y5choBK5GQZCB6EmXZoglUCyYlcU9PhogbA0d9Q3iJXC/92tVPcjE2u4vPz6OjYwE
M4SPVl6yxB11UtTujH7Taybb77R7M+l7YxFQQDxdyQY7ot53hkr0W6nJ06psW2+RybHmGcPCaIkM
d6+UqzfINL3OScqa0vPnTS9QlUfJ+3pLK7kmZ+ATlUAXc1+uOI59fDE4oWytJaOlebSXkqHd0xq0
6fEZCbSf+xZmgklI/I6xymtHOE5EcIA0Y04LzI4iqJhFQs1LbUI2y06nHdYXGtpJ0YIO1wrLEKJ5
A027ryDK40zwSiDNyIacZBGb0Alfj/d4ySwsssZeBz7HKqtxPG2klI/Jfh7w6nUgCh1YBNdbPAMt
DTNLfaUSriPUA+HeJKZRktF2lu42e8ClpKb6pmR/qrhbC/w1PIeShJ8Vn2AvMT8dYi2pBteb8GTk
CY7pxPCwTe5lX3yjBzI7y6wdZYBz6tR2ntp5j0kNDDozpNepANdpPkD2Ra5tzB+NXlS/35F6YJep
3Iz+xuPaIGz7scH1z5x9V8Jv5tgoTz6akJOle/1DxUjGKqtE5p228iatQC16gQAeMNjfC7IkR+GE
VIAeCNEGbZ7aEbN8M5pJm4UPac8M3gL9h6NCRrutqBmncEcoX7+vHub6g8Htqmc3ImBjXku3l/nq
w0RVbS5I3kO96jJKqeIJNiLs8+aCWzYmz3sOGeRVcv3lY4aG2nnXosp52tayFVVwQQtv28FTZy7V
V6MdB2/p/GaaP9Ppi0ZIO0dJdxWbdclXSIJCIxVXlDMLAq1cZp/Xbv3j5KNZAcL2t4vMsyuzcLHJ
YbqDC7GUqi5hsLK9/6MfZlnpGyLHQqgJx8uQlWuR2E4mgkWPGiFIMnj7Vp68pPnY4/IOuPpp18qg
AIn2kD3iwfZZUzaWzRipkd+YR2KppNm6Unq/AmPYlivhYyBZWmwphfgT3SE6kZfLVmIJK0ij/fH1
2g843+AxsurNLdYnXITTVQMFp/t1KNZXnATfyzXfuXbUhT5hrZLFtUfBH+ou71ZDZonhMN0ZLdQp
3GMZgDd0/2ovndr0YLacOR8/V4qao4xURau1xVQPXogWwGJa95WQrw4+wymFwTGuKo6p1/DKtjLX
hYZZ7xHgaEgEZcv6MiDoqI9Lrc7vEJ+tX2nwVIybq5vplF4WhZAGtOXMYGKW6t0eaHzaOaN517EJ
XuwoIeoYjqTu6CWdEISrSpoPerS3I308+Pi9vN/b3y8Wx8O1bav+QwaOQaWh0o8vOH42fbixvKhi
gMZS49JEs0YH98/I8VXD8Cp0MI1tQaGVzD+AYNEyI/2SwDMxEBnG2IWJKDMH5hzW6jO7YYneaEpM
+pAjVCfMOeP6naS/zccL5fX0Kd9Aulsnj7drzS/hA836oiwvSr1hOLt1A/U2VIuVt+Sg7GMNaikY
/lzuUns+h2/cTrZi4x5er44VhleNH1+8tOrzhy3beZy9batSDQKqBHrT8BlZqIaSzzjvN9Zis/7O
rz4qMHNeMWcakzuRZCbvuzkEGt+fVjV8t1mHEGCSbHyTNeuyoGicrNRH7bzZ5kTcG/T6TottCUIC
O5M0hwYFdC2+tXFqphZK8cCMpi0V1xWYZU2r9zGKCjwjGxVNWfzcxFTpBGg3JaV6FrNr+/nXE3GW
Fs9yoiY4wdxuZcLxWJ3pMSMc6Stpp5mNGzuty1ajaiuqZmLSDGSMlyfevwZ3MiOu+4Oz+Oa1A5rm
wOtz0cbC5P9Wh12+4j0XTJt+DgSFizPRW+5D2l5QIxUEDXnLyBtgE3Ho7c9XgusVykohMJtZeWJE
SFyZE0soqTrdMYlTUR/Se/Wd0nNPJAbFFi/3UpB8KgLmBsUA/XuJ6kA6KfTu+pVOH6zHaSfqbES1
neqC0C5+087kr65l9PqLk7xefmxuN1j/N+K7fDkaXkL/t6rh05Ps/1agDYlpsaqBaXDdiuQwSez5
KOT6qEjzN0qS7ezSZuad+8Ep+8pxR3BF5D6QZfoHjUoDYmE6l2VkNHPNn+2V/f00ZqgVZOxJ/N+R
48o1+rJrlFd3JM/0SiDhuVfL5QQsy58oCCdvdBAegfT4Y321sKNV/zKUiPfy4iIB3P6Tz1JZr+ht
ZYfJZuDeB9MEcPiMooHru0w8ahUPvo4X7ZvwYS/mNb7xP2VuZuNpdjLuzP8XiXo4V/UanIOspafK
FuJRVjU87Zrdf4bQs+/nV91NmIdCVW5mLABIn5SLjE3EKaCJeKooUv5HzlQ+3JJpG+fEZONvErRR
Fee9c/YYSshEvnP2lPecBGfc2ATj+AoRCJBF1pK/CQn7U/4Kx3SaowZaO/hO3dFrs1Ec4yIL2iKz
EBSMQsI9InwqCIlN4HdNd5OjHxl1/ewCFP2si33TLZLpFhJaEqfCJ8Ja5aQHHvtxsxbWetS5jHUd
Bh1YxO7K6i7X09xDLaGv3R5UgOfdv8D0BImIH6fmji+nNL1vIrDtVSMs5QF8WxUMrUYo17wILuZo
6e0lwiUHWnxIUya+MGaXI+D9AT1eoNfPxpTInU4ZPZyzRCG8b2dVNM6EF0aQZyJZLgTc7iQ3trMG
LojsSarFHnx+SngiQUqL2BnfjAKJaYRZV0YSQkg9201NuhDP/1RNQANLKK2GjtZAVcSAQXJAr6WA
9Wqe6dOgi8U8LcWdwPedk9zxr0bblQ8zb/KJzOtRDc+G2BioiHulJwdm8l65GNfIJLOULP6QxYa1
vkVDLdLKwDiI7Ibzb935MFyPVWvdfS/uGJddqpcf5pJ2UNaVa8wXJTp/6rRsXlGAX6x4UKae6hNv
7JHRET+/fqhvGy4jZZZtx2lo24NYbvYKXkdxLh0q4hDLZahppNP7pMqfv403V/fjlMH4gsqXa86/
Vf+2PDDj97u0s8sT1Q03PG3UEW8XSacSUCFYSlX2sA+asQpj2mdyyh24C/2hadezyQ9xUD6lnK/n
oj/IW9/ZcUxNS/sncr4H9ePM28pAd9CCnsVPIvVyNeQLlWiRl9TuHdx68V+Bp6+9vAGE4k65SKAS
KrLBS0h77+I9SB9zqiWpiAvwpva09uqa+QOn53TByut6SGQXOvx+W4ltu8yLWh22fJwtjGl8yv7B
bu6TOS/ydwvH5zkdG/34+WQbvFImtslufKdLuD3lY5UNGuUpCu59u7z6QXcqieMUXvFfy/gYntXx
WrzOHBhIYx9gUGRSpMhux5hxzKSsfa8xBXsl9Ih4CnG34AK8Pn+LVwUigIalXjKPtVOpqXy8E0zZ
6nJuS6eE045mXet/S8wrqSQN8tdNPWO0I2Mjj/CHSM+HFNbM02Rh8JpFZyLHPO3ftCkGC3vodlXa
zN+J/s/mtVm02ftSWPEOgwEKptO0IlA2WVNdWG3uMJiGC5E0YGdxVldIgUHdWd3/vOh/E1M46ZeA
7XcX/kDFT/ZYqtM/Hrl8ZVFaQuPJa+yqtkv9voRY4x5gR16XiPXDB2VhOtmzHz7pQCAHd1ARiShU
bQQduP6tU+zt6FYv7vTpELsONSYaANj7eH17wYV3cBv3TsCzlkF5/xGHndf1GMe4O/79/Q4g90tO
dAOtIU64RGVJKNcqGF+gvUgvqoedoGAk2gOUwYo2obZehhFgUy5NnVnrxkyXOIhuON1iHYdMbHYr
CjqUxns3mQaU93Ds5WoNL7HNJidGm/mA3LvsPKlzaJkyShJlO5VCocWgNunWeciKqFzK6h3pzIbq
NC+gKOauL/83GLXfPO4qgBoujPDEOF0CFTWo2iaErxXI/qp17HmajRMafqsGpYFU+Xtcxr3fXuO9
QMJ03RqrDUMSZVAhCnG0/6cjQvcPYxugmpVsy2y7INQOcwjK97ejlOB4jpnAWWmAzMeEohF0w7wQ
69LfBuHJloIX7/jl6Mw1aH5q0Kd68oMxULHnKhkLP/3isew/EEY2YjmyOontNj7QSJ60Oow0NXoY
mzniBQsPvUNZSK9s5FOI24fPFk/5G+VEPL6I6R13vihetDCVfgT3DBfN3uC0BXAWH0yVJVMmlJtb
HUg4pq5QbDHtjlN7ET/AtRNm1Iv7XeizKZifvTcWAeBpg7hRKbRRyTm2jaWHe7qQKQOuYWBeFabz
j+l/I6P+jUuwFHVACQARlPWbh83in9VIsgVLElMnZPvLV7KyjmcNkqsKpvVoT3uuPhg5Adyo3gZr
1qLynnN219NfRib7yzBmgcxj6XIbV/46zlCDs31sCk2puoih5h/ZaiGM1WN+nuqSoNbPMKhSMnx4
5ORJICfiNdz/gMJB6XAMRHfwGBTtsLsy5IujOLBRQItNgzFqp06grOfex8r+jMtcINFGmLFk1ULH
AphIbsLy/7jfncqBMD1vvW7iw7SacBkDjtk8Gwmkg2PaSnhEwAXv2hDX/1VFuRB0TZic1Re7f7ie
67CB41+A+Q4EsLAFGW5TqQ7Qr7yLNQDpVG272HZ5nqnMcSbLrgzRHFEoy/5HFwmwmig3N4ShDfyP
Rxyz6IS6eGMfQlGYV/ibPsxKYczpEMQijJb+Pv043LrJHSZgZdPBtMVgisyWnY4PpiZK3ZFrnfR8
60WYcorKdmnOkRyBYfbL/+2V6FhcLi0ultI6w+zf3RABBo5DyHzfiqTbpEWTA26nA3Nmi0Jspsdt
L0n0iMmKyf3YyYNayViqTA9ULjl5xrPj7qxcjy3nIXHVos4K0g9jnGARSqnM5umUX3e+IkqAQiLf
PZGL7fe4BuQbjUw/BJB0DW2GMPVUB5YJMZDTj+ifaAhbRqeQIXxbXATwFHpp/ebmnuyBiXjnZ8+B
L2BAc5v0/kgeFRBf6Dswruq3f7gl2H2k0DxTMoly2xPnclr7Yp7JiNi/ABGjwQqblsmRsN5k0hRX
7wSZ56L7+WnYBL0RAu2CoFi4qPub46LPgNqv635DGlTBODogZNHoQnVcUbtLFKBftUO7a5yJyv+2
9dGhMNa0C+CfkeRX5lyhr35f5jikfufZjVmPPi7Rg9v8u4nFb2AswhXQrh3FFZ3VGrkZuIK9t9cv
gBUVlr5dXjgqbvDmnZZ2/b8TFASSacvH7XHxv52g2ZUJWCEcKSQbC+lMTBbzh6coJV4FYsKVXEyw
w4lj5EwT1EnnPBkc6Af0Ju8mDhnLSYTyM/FAk9CJZAJBThOEFihm1ygGowc6A3BAaqHGjtBGoHzy
Hd1tE3hhSFvYDLmejOPLum+l6ok3Py1wN332jea7fIQ7biEkvrtcIeOmLXU8UVj1z6YSibjTlddk
8wpzUjncJo5jvRNF+wFnmA4Oljh85bzIrJutj3TyJsDwE7sN6M1yPHv3LP8mAqGvraWW5ACDr1jZ
+F0jqmnlGQa96jkH5nXTIrfvJ/i8c9bftpBwOR0i02BGtXwaagtVp3PX6fztRfYB+e+NImQ30S0x
yYsuUTZLFGmEq1WP3UqGzwnA1R1B/25bS26AwNzmsd3uQ6dRqGtNLe39GKpFyj/3Sy5+R4WYDl9g
QkdH1DNDoGlYKipe1k6u2gdxwZ3nFAqhZrAzjCjntQQ367KYK6PtX6Oqrb8LaUmkSVRAMxFXMr6P
QMbSJ60tcyMGlU4bBIhvUwePrt5V4SPRh86kcHIpDwmQfz1BanPH3lshv8T5KpbDXRoDI2GOnHRI
O/CJ2GnH1m9rd/gj55m4ZylK0Owd7Nkl2IhWTTOAdoHM6KBPs2lHeprnv4kc2+e043BLbSj4Enl9
5BUi/MLJD+vjBMa2AD5Yqe13gW38F0IScFCWEmwKKn3+DG9axIcpFkhtzF/mpsvyKiN4F6ckbxUI
BQ+BRN/GL6USZCYJ6M5e6QZNRtP0aylXKq055rzJn9tqPwds7hQ15GztRAyR3WXhaCPtj4x6GiJZ
Sz9vE66ssQie8jZCsOa0jOV6FcLw6ZtM59/cIi86eiO+hSBWJMr3XlYHBQrQreeCFSQiNmYLKTDi
Cq2F36s0PL2afH2aKhcI5jrAEuVJ4e1OHgHRNx86XYF/4F/GWqkVDfCLvajKTDyh8kAT8DAjmglU
qvFwi+m6iGJinwcmJLFxWCAig2P1QY4naJg6zIu+5QK7k7PXJmTMzksv0H9pYLKvSFZIUTzlz16O
crs+gvyE0hAWJ7NAuSacnYpnkTTPATdI849AkpoQQ7mSW/D3ooQPjpZhK4oVKsdzDc5eKVafD4tp
oEhFf8ia9x0XALSITKkcBoeoawPHgH7+Yo6sIj/hWe9wqvnDIeQ7I2X9eMb3o2xGZHR7oFL/RJR8
xSBq5QWg6yQdBPs1JFEhNBy1ty1NCqh3FQHxYcrAsJ3lmx3djCl2L+YY1/ntr/Ol7KKY5shFmiDW
zHaqVHTnCTuLnp68fwx7a0Kzsv1AxgW+/TdcOqiYaepFIW7Va3cT1V7Bvi2S+ot+TsvjuQv5SVRY
T0FW5Oho/3zoIHt4X696Oy/MQGaAM2B7Eeb0qHv7jpR5aoOZoMLpXcCPDm0Y0FpR/NzdEdidW7Nd
jvAHSv0ScF6WuOPsLPZbsclKf/Y38FSQhn3Cyc2mLdwXYrS2UCd+lrmGZar2zxChNn3IH9POHMsd
RrKk2U8FbZkM4gN11IteBLLv2sFDrX/at/GiK/tFvju/IywBhp7tyBaX/bybrZ2JvDwNsghJJV03
wINHrK/T32ssX4jB1qQEXShEZyyoRGTraU+xA2c4smUbLEKhlgEvsGQCQBXw2JNZdff1tnXqtAZH
giV1mCFJDWrvuBYQN35B1oTw0VzkFoAmbEcF+hpkapGvojwHRYeZR8F3iy6wlc9zh/ZhtKeV1nDN
P8YUL9a9irYCZmhDzJSLabkdoElTt18grqrM5gz7MIz9hfdar25zbG6sE1hnyg/jjYGZyO9SOE3w
M7/4z0IOsredwQvIciZhxYzyrx+AoboICG/lCPheNx/cA7yWkNY6X1b27ZUPQR5snzsrJjxIKSTC
rY1+8FDDjWmZkqYpST8LJYL3PIYnCZayfNrCniRr8k/EY9nrEeNaSOm6Bdf2k/Y0twIJgmtF9/dN
9k6riHDbeRttezpZ39z3neya2I/BpvimwmGt/fGUFbdbcib9PLttwnBFlUtZTD12YZtPVzi2jm6c
fHeGHIKwBJ/UtmiU5AGShj+uAuJKk0nS3vzwO0FkbqBxAhsIzvsG0liIRuXBWK2bzGGQTx80hFMl
rJQW53MeRutxuNtNV9VuH2M/a/OBzK47vAUAG8Ix8yBix5FikUAgMMxmZdCps2excK0MUX/oEX3v
Roj4lK55Dg98vaD2be39hsCCG97AXzp4QE05+dLHYPekKZj53bPwuLHjVFzS06pc/3latv7hL5Mb
wZqhdtX4QjUDhyQTUx4cBhjXep7JAElEEbKTtGUTpjjnRjT3dFAaRZFvfHminj7gUUQoIJbg4EhU
xRut+NocbgFpsg7BWJIyZ4VNvFh6DbZj2cm9TUi/YJp4dUF3c4Roi2iLJuYaw60qj8EI8eQgLQBK
GOOKGnQIhehOZ+igzdP3w2GH7Evui1gt/+bDdWJv1asOa4zK/2dOEN0jBOLU1oMb7hq+rURketgc
FH3Cwb5T/qHgMQQueoLftqHTMOdw7EKUfUskk/cbInxbKaeKNySNzZ8ZTiHQ23b8NdCxEqHYFOf2
K9LSvGHL40+igo4ZMIMAndg4mtVq6wsOItukcgMd5gvmqxXQJH2j3ZdfUCPvqFIAaPRRi+xJv/mi
EajmGJ2i5VnPu/3rS2LpZp+zHbxpA9lJtiiPI+T+a32umn0Sg2EiWm6bra9NLzKloODcDIjyOyIq
jeAn1/9WXmw3S1oLArTcLRcUi1dwThLiImTq9+CadjdrkWr5i4TVlm0507TUxR6UjeQWx0vdnOdG
QpJmokFbZT0XbHETOF1LTXKDSkY2+rzK7BkhFNrSNYz8dDUe2oV8FeX/FqmOAm2UkRprMyyQiCJW
8/VQqFVqn8ms6L6L2biBdWnNZtMCkyP1lDKDDE1aQKaHGS5+i2uD6u+5jNqRtqVfY+g2gDbwOKW5
qOIrKg45PBfkTP3hynR1tqtq5wGjTLx+MKXFaATjCB5ciKoTj0cwUxmLPkh/NvLymheqPneFk8sg
akjBBFQPbQe0vAoKUoyp26nVf7sCjVnuISQ2BeJSrobseNEqm5GdCDBl5MmVvxH+Oc+31h6oSMd6
DmyXVQA11PaG1Vs3tlP8eosfDRbZRAe+MAyQLCjq2VcFLSONqlM3LHt/0osG+Y1DgmQqllXrwwZK
/WQ7N6o79wTmO7zRwOldsLrj+PL3IxC/teV+AZrpW/Qu+p3S/XvkQ+CEefkHUxxbUA2giir4BZZF
ATnfbBq8+v0/+lWEjyA4/0nJ3Y3Nc0IelJBXg2C39hdtzbaEExaUhEVV187uh504z54t9sMF8w/D
4cKiAdd8csRaqdUoX2y8hpXqym+eoeBsUuRfOj4wZv6k8PTtCTV1ZlYWR9E7BpjNShl6clIo+5X8
1D9atT8G77VVQf5x9pqio5EmfH8gLyXohaV4Cvkh4hRyQDsjj+JULH4xq66PTYIEb93/oJHJSK2j
JpXEZh+5m6PPAu42ekIy3B65AJiUTHvxOa34eVAr/Dmlw6owYFC5svD5GCQlolQAljeBnzcDj6Fe
KpYf2OL1S/zOhPO+V1X8odqP3YIxUe8YnOV+O5DbKnHO78TZs2hK+bbOXcO5zFe4sqZ9ChV9UDnn
sLeYoYYEM++sjnJ6fxDs8RvX837dxQyD0BCBpOg1V85sJy0s3e2qQ+d7ARMsxIe+6/4///tupCyJ
tpbowWCg52yLUJrfU9aTIbXzkmNCfjgtVyyl7DWZiAvZGadkzPZAlLTQsdMsjoa4lbURYzljEyFc
8VMwiGrdgSbeIj9qPDOUKClTDAS/IcCZ7UMY+3uh7TtxNycsEwXH8EBJW2ecBb9bPeg9sAMN3vXD
p5DShsRsqrY8gmKu12oEaiIUxUnN0nKLHnqNGz5L5hrz7p75n7ioNM4/asMVMqh+j8hTVDoQINME
6NIkUEogARPBrguMu6PZsQsZpdiH+qKxFSrJHurxuDh4bGLzoLfNBiw5YwMqZNQpMMFhi+AfRdir
K4U/YBTYphexQHEX6ZvZZ8O3Frv32LJaGsCD8xNbp8b3hr0LNwNYvyFGbOhNbFTvMI6myOEBcV6M
nP8AMjFM/JoAyoY1f1otTUkECzHo6iO7JVwn7drk+wH2vzZxzEiwJZECedYdT9z79J598Qj/zeyX
+fuHAI6w0CG4kuawjXiDtvY34AT8AHjShpfid7MPvVdn4b2SOX2SMBaARV/P6kKVC0sdnZmltUTj
N5u8Rzi+s56TYbBvCBYosDXA7VGAIs3lEI5mrkJTO83YZTKtL7cFLMuUYjhXzRu9Go84Dp+ihjoA
PrCUfUESws+h2csH1v2/kVixtE2RXPZbNdbYSlQCb/rXp4tOiybizWNSW76WX9gv6rBjdbemU6qS
+HQsfHmervD7VIViLF/R43OQ5+WeSf0Cz4pUGUy2O8zmTB+U0uLu0xmzL1yD1faDjju6QsyA3rtI
28Hto3sPuhBpTsAA4hw37vWxQcikTd4QNlhnmD1fGyrVSckuGyh6x8UHGDqrHP/BEK3577gl9OeG
1Ncyo/Xf5xCN/smU/AfetGeTVX2FgkwLflaq0sEo1AqYCEakqDJtEqoesmVtLcfLt0/p0rXIwVlp
ZJLgyhEQSWBEps4MkYsbigaldfH6805aeTAjUSrq34BgnVSfADPu3zp/jmKO+fua1fWD5G6U/gNz
2SDv3cEFVVfghzcZ/ijaMv/12Jo4ti/T1Sy4aec1CcvlM9U9M2jxUNJqQA4TCH2rWImvjFg+bOfB
tfWSPuTTgwXnH8Ap0LpAQQI30ygt4bTDdYnCcOfwl/dLTBeQ67d5V49NAdCT03n5K6OPlkrlZWyx
PL8+z3XgQ/lwG8ATYk9O2qXbptGb7xZ9iYVV2O10sBvQx6EFGP2vxas6HvFftSfRoZEianm0LHIJ
5VUigNj53rzK9px27icXfnynntMYDhYWMIt29JWjIPpcnazKcSSgaIFwT1PcqBtGegaGt1W6+Bws
/9XuL0ZJ5DdojeFq1DMqLXxEsgpdc+LesL3NcRETg/dOnpd/0W/eHGRGPy5SQ0SyCJw1olJyFn3B
eqAPrnArcVJNhqAs36WFxBnlhjZZ/T0SdY0zDVpiaD5jHdPfcXU2NuXpkD8hNTtUcY/qIEZqo074
TJRoV16XF5k+aDhMEBT7rOQ49mGudXhhFvqEHCTbBpM/ErvAzAv/XtmMA+U2o5sXtOZDGmBswy5U
LjWVrqnD1+7yHj2XCM2Zm8A8qapiXgy6A06sLpWJYRjkm2HIWVtGFBXQpMV3G1Or5F7Zx025tOLg
LVeU1OCkgq8MAdqOnCEu2Hr9dXPzCTuP4CY9ZbAUUrESrmxZ3iY0aVg9n50PkK8hrU2AzIozKVaV
0U/zQjqiO0bXB2zlTWqjyxBF4K7ufNu0JyJGvOE6w0KB/D6SGmsSNpqgGQB+VKZ+wqt/A5Kn7BMo
0MRCtGCLBqdRQNAhp6AqvEH1MPQTDiSUOOwv/TIbWqoRE15WaFAIeST0jIUlyH2kOTUvqfbf8324
zS1WQGSFZSruN6a5ELWFuNBx+AfY5PvXP+7x7cN0GZkQnHUK9jkle6MBheaAqVcd9v5NAuOGG8dt
+npmeLUSVLNhquow1GJxQYzDjv4rPILguE7y0qCLdogXLLBKF+ilQK698SH0pR7HnjdmJO6rh9a1
fXLCY8AeF4a6ivy1TxVbyMMAwxKbThB7LoMOQ0ifGXrKJr7s5zVpRePe3V5GJtqDbw+e/SVgfxnR
IZ4EBPanbihOF+if+iTGi8AP832YS42ROIXBG7DLPV25mdCHr0S31w3w47i56MYIr1N891kNtYiZ
L6FukrUbIjNGZhCW+KzeQ4ZgP9lte9JfLbeMYogqTudzpdFS7uoh8iX4JazJBpJLG+zIOFeXQt3w
p3azHWI7sRR7HhJBUMf8tyHH+Xber0Z7u4O1tJtJ93JIL2GV0cT7IIM83TN5V0j7lZgxYzPpIbBP
5UhpOFK0id7WLYLpXMN7aQVNs8pyWjOOyrlTRh50v3x9aHm9zGC0Iw1F2yUCKD7upZg+lPIEDPTL
rkZmgS+8wSEfs6WRyeiYnAI5P9fBi6hOH08GWfjBZNYaokeSdm3CIyEnImB46tUFQqnmAtyj0jVW
wo5+8KYaraOnQ+9+GvTlG0UAlJsciFOaKYwit76GlwXinpLYZqcsFrkVpBjnY2y7fJRzd1Ondx0g
8vNRoFsKhuUiwKr1Uz5b1w6xqaCea9uKvz63BAcgJWkXq2I0XvjxDg1ATa09z2zQ3ECoFHTbWAWG
iNzgoWt78WTDPGirk9PTQPMpk+Dpuo8MkTxnCDGCb1ELcl1Pa0RYSTkBsNk8LScAZLTTWR7myk9t
sxpZR0rWjMNVCnSppM3IJJFqpGrqk/ftTnPuMI/oWNatLUsHRLPRuplXCIsVYWgD6vWPSTT4cMIf
nHMqlrC2sRJ21NTk8My7ZsyiSw4WK35Ze1GtXqvYs6JCgYPSvYPbIiTzgNqOrcg+rPMdEnCnR+tZ
hAgjeA+Yidnk5qJG8rr2EI7Fpqz2rihPb5JZ220NT1aX4M7x7KSpm0iYhWZl4mgl/zoGjuXYzWY4
sO7nK1TeBvAwjakj1SGs1poDqrhOloVYUbQE6zlnRs44r9e+KAWLTs1n2hBlBl/WPr7XVS+A2GNN
DkHASCLbiNY4+y2+XlkdnSd88/1GEbHhY/IVDwb/PxpMnjJS1h4ewrx8fLlGcX88LitRY8e14obh
fFyRTbW2y7IjiFVOx58f9yvPlCiAM2IAlcLgDlF4fWj1KUkRKuaHggSXPm4cMeyNuKsYmOpGIVOx
U2AL+TQPlA/eXfvOm/Itt7qnlNedHfrkiBsBLRmXzpVJ4/cNgvRpTUQHcNAt1hB6/1obxqEL4SP2
i/9WVrFFw7X/nFbKWMxn8CZaRTKdaDiMVzLQu4WwmDKVAx5yTsDwbmvGqYCixrWdNwZbRMkYRNKd
dJIA3rR/hfgdwHYUH5NmS36lTiSFSRqnAAHpQOy1GOOnkqEh36MXLcPOct1zAPYttJKfdGll4sFn
U4+pMu9D9sioQ8ba3IducrwQPLrotZYg6xQ9gnXD/NDujiVL2k7DB9bgwEMhPVzFMPj5E+Xg/T/b
sC7r7atb0TjyiFY3Hl3liBlLGO3LH3i7z2dULA36zpZsyoB133nl/oDxbEM1Out5pSPdlevnKAok
15o1vottYqlKixlJTHKopfWuGPiFNpQqqNW7en8o6Cq15nTRvNUdFZ7eiseTNJi8JHKVaZl8uDKF
+MK1mminsIJRn7hDmEwD3Zn9J5ZpatQ3pHXFFnylR5D38f9yy2/kWmH2oDJXyEDzh2OX72VqB8vq
Wlub4rGY0m+FtHDXSzyl9dnLc0PvYzitWNyOyX+k3wcNGpMOSkw0TUhp1kfYMgJEY7+5ZOIka5FG
Zal8gjsBVKCWNNhUPC09RuTo46g0KX7jhgg1SGfKMG2yhNi9MmqD4xt7xE2Da7FHQJ2qhPgCxshn
gYvazwwFn90zM4KeyiHZ6b8ooGWT7t4mXEsJmDMoBdtVgo8ekMgJ9jH8fQ8NuH8eTBCv5m+nbGrs
awdbie2use/2tZhoPcAPvXG2v7Yn3547czltghNeETQtutKdtK+Hx0oIJR4+RRAW6Ex3KhivZuiT
vk1k7ppS53b/2+cYkpLhN3YeMSMfD9dFChq3WfuFIhl8dvJ0s8U0Ez38AZokp+6w9TNXwcPoMnU3
XJ2HQC1j5Xfl4abTUtwz5Ywg4fA6mPgZ6ow35MD/Px397KIamdtpOXXw1YMpGFifHnylwVAVx5Y6
FdVYdbdL/Yl62phjy7vkbejHVrtoTkmAESIJ8j4cv8g72o6bws3CsqktZtA2kuRt//OwJA26lsHn
ytGdnnBnS4UMdxLlIXC+LjySOteTZV1A4wa+xZDknBKbRpPqnVvFJrStpQZADIlF5RdRzuiF5/yu
JeQOlaFgs3UPfEyZFNEW5AorgPccJV1RgiLBUe1c2HxsmOdZ6Pqh9fiKPNXLEuOon94N7A8FLGm1
5nZZvdAxKu0YC+S+x5KcvppH3GOrNgqXRenHIecF6JZItR1x8hXJuSmSZZMVfKVuUvc0/zpGNBEe
r8NPYwFWKmBXmr+hx/SjMVKjup9Eaf/985VenDY1gKRsa0plzYVPS1DQTkJgMim+RLGRr8oRwY/o
DPwf2aj284qLiw8NXbXpkLy6L4VpPb1JLYIU3J1SvJ8VcxyUJdKud8L5l5+EF1zs+NW9Au//XeoK
3VbjeS+VzAJORlo2C1RhQHJO9UUrTThfONp83PkW4B/gt2Vx0zFcRpE7TYjZhR5nfcdGIocIROdd
YCxwjFhkgzSniS93AR7+LVjoFyQzdZrAhS6wxMBuhEVzM+cUswYmMiEDRJsqfeZyb1/2K/TVFATf
+Mp1T9ymBJRbFW/uGSRJSc3llzeqpET+UsWOtVP6N51mc9OIpzGfHPbwuLA1cMgP4ExPMWjQwLAl
/hwwB4cfUgC0E8ufjKeFjjYpNTu4Z+xIG1OD+Fjc5Dfdp4+zBYp5qudXKGEgNJjjI8OMXlcKqUvC
9Fi9p5on0KIYQHPpHeE3870YDr8sPK1P4VMSFB4RoPi7LSOCZP1884FKH7AtyFGZJ9SPFor35TK0
J26h49p6CdeyisUOwSEJ50I5j/z1J0Fh30jVyG3mmOR26OBwXjMT5KvWB1/0YZvq/n6+hGtcZYeY
wZWqsOEkTP+vpP+m+FU+spVcNlGxLTM6EBchWs5bjPchJaDoEApasidphWaYv+EnyGcEO3IDZTVy
TADHHJ6tNvCi7MaDP2C+3pzq1OnBCCiAwy6lzSBuDY0SL7UcG48EEVmZYbTOIaBZqCZmPArTxE0Z
hjjYKibXmOlWljfJPVLLBC3Yi1eODYKDO66uEj9cW+/MeOQBU3OFyq9SS4o2ZArmwjJMu0FHtWft
Wc0Vmma2I+lwO/i4tz7UmEIPVMJ0dEf8IzFMQqv1bJQeVqgmojPbiM6Uet53+Ohjb0Esce2l8aE3
YDUxbb5ELlRBUHXmCRyKusCjPX0ESnhEo9EutHkfn2mmXBC4flxVEDdvF3VpZcDTghU/wvvZ1Rkb
UustBv6OJNSHR/06/mwscppTqiGzLa+yzeVB04zUIauijV2WokwRmwNqXyzbGfcVQZtrZbfr9W8w
6SxnDm1VbyrE8Y7ijR1f7MgmCwa1uFLDRgiS4uT8cCtOAIT6m73DtIA3cqsO3ptKWbTs0dcHqLkJ
nWekOxa6KcHomfwX5I7p+47hePUM0jDExKZYIKCta5TzD0mzqm7xGZq0hSPFUtflT9WoWLyzUvgv
nIFKVtDcLTml+E/3rVb3j8k8YwCsqWdVkVKvIHtYFu4QSlWABioC7PvFdneIWFFB6zv49whLg3Oe
cqHNf+A6vZIkxIlNmWDcLMh7Y+Jw8zKALZPCXrIjwOLT3KJePCfJ2TPrw3VB9V93h8cgJPhdyKQA
fHK8Dzv2UzzNDDuRu3ZDVwj6HiieXjg+iflrGFiENdqMXEzBWsjjWEdtwcmGN06yCzZeB1DTSfrP
gNtjzd4KRZGTT5LwY55xkVciCHYPckwxQ/WUZROou6JvK+U4KaQ7gSvYCCZwg2M6+uOMaBJs6buW
udqqQBDpt9N9at6LJNekslN0FhOfVuTJlEex2laYwPBjPAlsDVQxV1YkEvJ3Ej5FPa5vg4/wL28b
CNN344eURttbOt3DrhXikxNqxAg9GgAiJTyFXo+DvC+wRzfH6RdOLbbEEfYbt/A5YS/AafzTDo5V
9Y/gAS58YK39PMkwEmvQqE0ZkxnoaSOa6DTpfYtbnapS272JhjvUCOiY7Spz/zQPnq+jwuZgAxKj
2Vz6gp7QZzPcDJPvxAjrIvYgl26MUn7ANGL4Y+Qfibbjw4GyLS5MddHqcWGNmM28XT9dRe/oZtH7
aol+RpledBKD2G4QEcLVfhcNeR5MxFtJg9BT9JczD++t7wAGOM1Oz+QlNKp7SY2kF0zZK7doF+y8
uqssxt90As9dRk0+Ehrb40OF6Tl5AJDR2BMvCcaHeyCuv2W0pE0EfNO7e5fVR4DvM/2UNASuehCI
ftF5C9KS6kS0wzraatM5mvARFY78eOYU/3d+fp64NcAsftBU0VlvkPL5lbkSfShLUTXcAPn0A+cm
o/reRRFb33lWKffC3CExiUcSt0VYF4ebyHN+sfcCLSbxMS5ITJT68jUS5gH91ru2Yie5LLhNZSeA
YskoLHBzc9aC6aWEF5wba1r6VzS7sf3iMD0xHYSj+R7eevjGPtUHEy+HoWGKreSMi7tMkNDGiroJ
y+qfuvYNGWzl8Hht+8hv73adWF97Y64VxVjVuinLy9Jz4pxWmmvAF9ZeNZ8CEI++nD+RgI4GnQMe
wgQUrP0cYeZok+NcbwwrFD0Wn/PgqVRnl5zZXNwaKksfLO8D2k0Sv4/YEJ/yKjS+Ailb4Z2nmP0s
uD+P+IqzwzrWmAC956Gw5v0DTyExdjz9QTgt39ivwhVm0Lu17bnbpG0HLuZweMFgA2vf1rfg6j24
loTLuI0ErvPGrZ9mEK041xeptHNXUYtV+NXxOJ2IEv2Xj/bRcyCPzY/O/BIiZG08OrC+04BM3kab
tLryIU/ie6TUz4lg03dT6iI2brMJh0lSySO4CxQgrzdagqU5QDM1pzemHItuzNHf4X7Bdc0oC8uw
zJ987XfK/FtvurM6PSLO/zMcVLdB6Uxy+SixHcjrFT2Uv+qkjFkiUy7VJ+2uwTh8CDIfNm+GXAGG
MSAvF3ZjWXDi7DCI1658E2EoPTHPML2b1iF41QnnO6jv9L4LKswmFjZU0z4+DVOqmLhsiIIW4DdU
3nzXN/JxFCkzYeDwIpnlpqsqF+FIY8EXtyCp05SF6+txnCuRT0UlDV6DK5Zw6Z5f8oIqXWf/ITuX
6jBCQeUeL23HVLyipH7cqMKJK/znlLoD0kh5wnsrUDsjmZMGps3oS+j+F33SeRq6MfLXql/F5e9A
g6Pgt3thXk/eO5Xt4a+JzF0JwueZYk22tyckGezws/uq7etm9oxUNPQVKgXGegFqX42437O+1F4q
zRIDHHZ9SekAC8wCnmrIgUw68r1TQnZXiLjXJacCUJRXltS0vDkig1HYNzpZQqH7PCL/ZuSjYvzs
gqdIfqGdHd+rNYBSCPELh95AF8dYY4pGzRF6TojdSyvfnBsCxrLndEAGPIlW/av5yzpdbxolcVW3
ccOrmBoLAIjxXExImiHtceSg+YAoua+vUO0oM6+eGGWemddQqmdg1adKgetbRa4r+2Z5nQCK68ew
jOMRmsLo+vqYX49SEWqpJ9DgJU5p4UVJxoW/GVsQ2el1ksx2JzmqmNzz59hxdt2UWVsb4hoxHr8a
JNMahZKWVhR+er7V03MEDS44gUQ1x3Ie4yeOoOHJxmE6PDErvFphgMjs8kOmHvR9IlixZYGjuWZU
EECGjHUDDb3AE8Y++dVCcLz77WP6v1xVP0WWRz9lBbz4eSDG8cEKy8hUUN1GyVcmKVkwQln0JgBE
WauSP2SIxXaJ/Npkbh1JZ/QmdRoBGtzu/QRemiYRSRrDLiV4HqErWjjXYr8Gd0KOXZnO/Gkdiv3h
5hCqXAljCNM5AbmZvqqy7rgQ+KIAI1NceANtn/3+aEkFV7ExWu2RErU7XHmEvd4n2dL+pE8eH+L3
+dOaMO10qKwmWXyDxA77ErLplWho20yqt5UX/WbAFF4xnrdP7YYNWbZ5GyCxxmjEVl7aSwMxZUpF
3GlZLC6ibcFIExKlshM6250/Qu6CrvZag5ctif4glBIbU7XHijOUHYCfA4hdfRsppHyRQ8tAvTHb
FMcBUmKS0cYqFhnX6NzzPSc2CtIfs/O4zenCRFou0+18jSMKoDwV+L/6pEFDrV3nOXCPBeSK/3KC
pESB5Bv92wDssJbu9pLid/q2mQFF2VS7VmQqr+stKDrrcbyUuuXSwXqTs6cxrSjbS1HLE+8foG3g
Cev+lsVLQmdEr+dZ2nI5ScRLtMSHdIoHjtyUzhSDwc1Qym2w+IyBa7OWOttpVnt6BxztTsUUrOeh
304uTL17VWzZLRkMAgAyrqecokPbtLXa3IZK0ewSRCqGas2UcLp9l+9Z5rWD0SL0rvTqHEXhVlew
p3bvFp4fN3v3Q3n7Z6m0hRfQB5HYdSZ8H1y0cgGQuQf0ayqeNC+SiwWl3KwiDZLc5abR7GU1deAG
e/zuNq87KRgmArnwoeDO9h/I640I3XAZaKlJHVby7afgd36n79RnlF3LIQPWMVz4wjSLDBlgbVhY
XU9mm8KRCVGUZx/CmjlPyP9YN25Z66cQxD9nIQ1qRwcTmxO1P6EQjviAtfg3FWqK4FUkQfianXm/
VUDE69PU/XfjpU/yf1EroJWRERaXM8GeBThrNkqwOIHnFNfBDnXqK2xw7NwjlPw48gRW/O/be6xd
93vCLd6KNd91sTtLqujf9WWTEmxcXlKGzoamklNIZzA/74YYGJazjTRyxUIyRPhlS7rMo2bjtZv+
AtE8VX8L4lwT4/LIQqBfdDpmUHhSnsJt13gkbUkGqU1lu288pIxC969tkSv3bfRbRLNWA109MMaC
Qr0mZ/yOtoS62etvgwkMlW9LGU0XrhUXO8vCBz5K8u0T2X4DndTagB1S4J8LTsvp1SMd5RSA8evu
661HsJJh5t0+A3F8PQEFpqCIoemqAyxVam4DTFF6PwABS8JPFbCVjXZ7/VcMEr7bYRedjI3v2nTE
6sxhocw5yUaxy7gfparPkslzW+LM5t6pV2I89yr2tNPyEL+H+gunGbb1d4VczIBi2/jvNVcqFkv+
Ath0A1u3dXpk/Th4JcNCcGy4vFmckqlEgZRxQ6i4/OYJGPPE0ZfViuENkmfz2NcUvhMlBlhMn9DY
vAM9bh0JnZ/mntHtt8rhwXjDl2yHdSLWeC38tjwRQtAoUCzC6iDuMTfhq3AN6wqYl2yUslwJycld
lGr1KmnhFpek0fiK9CtWSCHR7by6woFPKIrmwmMOSd1i0c2QfkfAD9xPqGMfFEZGnmbpxLp6kftF
BIwbxHo+p9WNjXO8lMWpFJ8WyZ6cziRVXDekNmPeV0JUJj5gnShv4xWISrQWAAZSnKfNfDtBas1L
ik8JJGdVwQElsOK9m6OMA5QEwcb+nvd1AZlVog2ki4r2+RRaRZUkHRyfK7bqEI80lpGzhSE4hR41
xLh2ETugx40D10+cTr6Unk9xIRBrelLWwYuO8nlG81sVMP1U6e3Z2pq1LfK6xB1DR2nOaervyybE
OCwSWtHKslVhu2NpEI+RFbHbJ9R4C1WriJsEn6Za5m5Rd8EZJOBwxQ4sS/t0GVdSSyYPuAb5Fwjp
ejN2cZW+M4Rp+1N8nnEQsrgWBABOAIkl4RAo/ULCora2ll6OOLKBTQo33lSGIXF5JK3QQ6ctfXGf
Y2nz6H05gGHiv2dMOoxFrVooCe7Ur3kxOc1xvW5YXBzjH8SqpsPTgxcHTy74Yiw2RiAjQ1YJOi0I
iNAtRBMB6rVz6OWlSPKooMO/m+tYKEMg1dAk8NeltcZo5gsiQUANzytmR5Kpzgq4k3iw5ealHDzP
Y8N7xsDo1n9ccztp3Zj7fBP6cqGB3ZHZDFuv6a2s8xN0FXnP9svq2INhj59j1CVwdHwbvW18a5MD
NH6Xwubjk5K9A7/gDxmZm6GmfbTv3ZWkn09C4+BQCCmnXnTQnfhQo6SWwGCUbRMW4RTHlzRct7jN
cBsErUqKwEIfjtmRdViF+8w5utNoRuSCM0zfF58DIS40QuqwOgc+oXBT3DUqkVwpch0KVErtewtB
jvTuWspwgDEKx7giv/qwQyRUqSrZMjYiS6Z2mrBoiu+OHvLy6kVUe5qwxpWFIty9+aFBaBQnjIGT
QNsSm9LKgXW4JYizFP/kvd5uDYBGJyT7cJZeFbLAzw68OusqBYaQEmEQqzxVx3RR+rEG1N1Hn4NR
VjLbz0+SK25BI9jbJB4pYC7rRqYhscDx8fL9mOSCn62lXVvTxIU9KqQuHjDYSC4xwhfXyv9UxgkF
/il9uv4kw2P893Bb5kNFUfkrLWMU5jzc8TO0NN0wtby4gYokptMtrkLDU8T4ghJYuMJ0wSXxce0p
hYorxaA6VPWmg0gPQgze/cCXN9P4+zG3EmauTrmac6VsPzein8aZoS71UcqB379sPCoVY/VgLE+W
bBChT9BOvZEi1PTt+94ONd5pLd4ub3mBEM4aZ9Ri+tQ24ipM+fOgASVMKVgBu7/vnkdnAiTNqPAN
8qq23gYuIt4eCkhWsDBn7XO3Adx0Z67hDRfrdLMBCCOAObgX1puzUzgCeHoRQqiaP7T8oG/dJ0jM
0O+cPxNIJQbIhDuaR8HKrNqTP0Cd9/8qUDk0Y6VH3Ws1lhsGQxFRJU7GKhyMFVQCNb7VjKycaXM2
wHNom8oVAXHsVJxllQgpMJdVZpvMl5JKr8LgYcn5ACU4XuymHmA4oaqpkxY4s+CCvUG0fNTjZ3Ug
tUSh98vWh9fwnc1+E4Ktq2EFX8O4uYKxkYCMfCFuK5FGgb0ZZGC1QFY4sCBbwiiZKtucXQFhbxP1
FIlEUTC9vzknlGjdhdb9/oT6/P+hCNwouQV4OJ9k68KSLSgOGe+qZ65CQIXMtttH49OoqGZ0dR7s
IB+ScTtPxacqVLgVNSA+ahbH50u6QMC8cjf0HRYXCW7X92dh0rbp8R7rOEC/pEoXFvwcyzcmtFRu
KeyH9aoH2bxpCGQlxJyv5g/+UDYLBt4XzDVqQKIIyNv7t3fNHNY78ZiUHb2PHDm0cXSu6J5UVHEv
0kuVYjZbwg1ClNWu09r3sxNTxYIM1TeSXamqmxAbuddYKq2oV4JVUdquoZH2RBM0A+H4SkKq59rg
J+dEbuwwOItaS+nKJueN3/g4QOBuLBbzlSAsrfzxtTUcwLU1k4l/RFU9qzbeeL4CF+6Wh32z6VY0
WEDeGPtfRLM1zF6d/XOTWVpFc6TBvAfFvRHwkpRnh9e5EIlzcsIDfG4/8iEmgnKl6BggeVu6vBAr
yLeTH8ktp2eFrL+V/JZzjOl6DzdqcL7zA2ZKDDzPg6W7QlIcHq875C50nbs6PiAEI79w09rwNI7V
WLrCuR1bBO/LGiDFehYrpaxGlBzcmghOts6vqXpKSKGClTrZXdI37b8Bf6ieyX1mR1VyDkRxdA4m
mbttnjNDj92CJOe2kaQbseZ0+ZVy+gcVZ9BfCiwPWUN7vLrkVXmpeyMYyUdNDfJmwh3hpIJRbA7a
HcHRwr89q0rcxoepoWVUQ5c6GApxxVLRdpmP1MZKoiHD1OQ6q53UJeX4USdhixnhvNOT0Oy5qihx
BgrdSA7Aun0b9E7KQtt2KLDAum0g9hgkaTI1HDcwwAx96Sp8haSox0sNP6sHbSg8jSgQeLXew3+k
frF67a+hnGh2foE0S1fLSp++D5gL7Pa+RVSVly59yG7sFK+FtlQJz7D3Ad7hjQ+i0IJr+BK9C72I
yukY+8ekLakGXNrk8YccBC3W4+PwaT8RfGFdq4n4YoRBe56ELedk1XT9zsfQgf4LtVyuLQAa4MPc
pSH1WQUdn+diN0OitQqZn/QvBQkmWeAzQ4ZcJ3S/UJkohDz6JsFtYf5S5ahCqkKmAeK9hlDD0ztl
cQJEuR76DbGqm0r4iz5ny4nT2Pa/5l7v9l6GZjh/JxQDmXh4SJ+owZJpEa5X7bLiyXZMAMdrq1Q1
9NRPnBi7Q1ss9du793jS7XcpKpwVJ0j7p/dEk5m909yF7TFAYbcMbE0kf3MumP36Se36mePMJgaK
vNONCNxZ3KfTrZA9E/7Gk0841meWsenX2GBWFATUE2RGTB+77ODLwPD4QmiXJC6spY/XTFpieOWb
rwmwCrMGU5MrdpRAMsyoUJokhJk7vWRpEAaNlCz30cyrKFZQgcPccqRYZnZEsHp4W9Vnq7jMhhSM
2o8BAsVKKCE3VFRpjnHJluav0sTMxAJdUkM2vfl9KGdonvKNDnMKqJwdhiud3beCaKlrYVxw90If
xreW2kHsQoLMg/ULkuirdBiwZFP2coGF7clHVieSATuvBYng63XcUgSTWEZzmPvdIAYpk5lyzrAE
L594IuyStNbgApzZVBOMSjoVWoBB49CKrBa2uGwD0EpgcNZIREhIlpCKunSisHL9GcEHp02e5KtS
pbKeDp4zkd05dgpiIXHlz5eIi4ix1fjMNhTrsGhg0eYBcyShvOODQ/vvrld3onvGqIX12Cu67Fcg
IZNfHx7jZ3dyUWdjAp+R562yu2DGGtmzYbodsk8eIpUsFoGzxKKq084OcxY3IBraY8LOkI8OlJg5
3UCHzrLlr/IeEKfXqZzJS9g0ttiAdXA39nEusxqZk1n/dbYxI5NmT76bOLZ+TgsM3TUN4gYZnsAX
Om4M0Az9P9OIRZREiwTlev98/hcGt52+s/41Mi9/QJHrXYsC7tqKD8KQCM5v1Fh+NplyLDR4uoLF
M5sja4ZuOEjSg8bzMup4TILdVNE8brtb+MColtiMhFiqna7CzMa1Xv/eFNxTJ0DGsMQB+Gyq3zUy
/bN5xj7VsB9m/H62mK0rXrGgSk4k4jY1GqNEwhxu5+PU2rYhc+zVRYua/U2fwrgtJewQcZna4tpe
CHtKcHpkwURyIbge9uUWn2q511eb8r5b4JufgqKqH/X7+LQqrikBZ0W/ah1oLYPtEt3niA4UJQuQ
sedYz2IhD6/7OqOCuNK9LpRz1bb1qlQunzm2/vzbiEc9RfcKr64xoIXyKiLzweTB7hlgmcJbc9dv
IwULHv/u7xRaEgs9xzhwYQw2ROlE0oDGso5TB4QwlijrGw0RDjMq+UyumySoLgVSnC3QdLq5+Faq
FI8cPvWZzIqNTwvgrBfXeeIZLfHfpZIR5k96NKjUN5+wnpffDaJbbeWju4oyyKdExtnYf8PeKJEA
/95Ve8vUHXRQYKchV7bpJxQQu8Dk3ON4iHRaV/jJT6x/mvXLZwfuT5dCchcO7w8OF1l5jQbdjnxJ
mJ8I/EgG7zmY3KZ93t3mR/DyEsabqIeGvUT+/kOVGHiiqKnxhZfkVQXWRlvxZ+vKBLTcr3kwSu0h
or1erDz1b+A3kRykSvNIgMyM8znzcc97J8GpUGisf0e2HYFBShnMkuWThoq6z1tgjCiXLR+OZBRT
k0VtTpQWDB/KT4/PLel1D+qcLRy1wAKXD3rYlvV78e0dmtCJuz3QHV7nypyT07pGizoJsAljWNkF
iyD9Ka+IVBcSvWQjLtPnpyW+vscA7lGZ8Y7AiNYLD4WVQGu7dY5gNQ+YXtD1gCimiI2SPaB+tTVO
/YsOKiYk03W6tQ5VASoaxflUYW891mETRnK8JLebco931mr0e2pdjPBQyuabMgMab9hKg8I0Mkno
XxtJSf9clBuqoL9uOEShLu33Mjmx9yat1bn2AmB+K+mFQmlGWgd21zSPI6HSQS5l1OAu96P/mUgK
9rCkz+wwJqcV6IoEhh9kGpk9OGfShCKL2OUtxbt1UoU6e9c42U4xHBeJxAgB+JUoVPjg2dCyjVqD
u3Cn02gY9TuuX0FrKeeHB2R0JSZ5m4qIZXYqinLa1NFwYqd/zDVj6i10kNLCFb86oKsHnshR7Nh6
ZCH3hiozPrvvCLPHG1nPNIzmbjO/eaQ8+ToUzS3ejCodRbBSyMW0y5xYN7e/4UYJE4L0JqrWXw2S
1yl+oDaMuI7i9F9vdkVIagdvEunVTZMU8433e+fAfp/ZPifyxk6INadyMGqdxO+gDUbxgX5cvEuh
C/q04ruZpMdpKuPJxJ4KmGrVk1Vdx/6f0zQ35DcQr6a61o78z7ioMA4UlEG88yhqk8+a3iEFSz7H
pLy2y0+rm2yU9U0SzJN3UlV21K2lLoSWHczauj9r4aaR92X2sOv5nCV3fV+zqE8gDNX7KdJZzntG
GmcWJ1SdNMmsS2ZZWCyx1G0FJgRSsdQ3YSbErZDAt6GyX0HC8iCHrTtybFHonaKNuGNO5zbbgzvt
60sfyoXNId8qrF5blnm8tNyyeyJvp9qqUkqMgGLMhVitgOd23Ji89BedoZ8Gc2I9CaxCmq3U50GO
mYHbon9bwk+PFIZIDkvl3gSv5bYl+a4KSlYY22YhdCsMOOH+pUR6+d/bx/DbvOA3xqfdN0kltbQh
Vf9ZJjV7kNJXshIOIkvRT9Ky0LdmgzYGMIprSCX3FlscOTT5xXY5hOgYVWPTB+l/dnTUKX47TDfk
WHWNX1VxR+u6wn4ezrDsMVkxjothX0w6eD1kdeY5znStD487Gr3OsLijvOHAkTvGic3CvpB0dWGt
jbOEQObPVz2x8tNhGxxQ+nntHLJumZX+14j9bDl5LCuodK2bWDtLePIL4tdLl23v5Nc2Mdx+mSKF
+Uu3EsVN3IMZp+PIGvegIg3daQU9WDJRDh0XktQ+cLEMF/E8mjXcbc52o3oCa/FtZRulVyUHRaig
txXLC7U5fPOCRk6wnSBj5mrscjui51aouGRxEh3oH2lvSgHRgPZqjX94Haa4IVQS//9cJyUdp3SZ
U1bC8jNr3r/GupmGt4Qnst2WEQqWqfxJnQWM+v9RrfdDMPbsbvHJeSIE28l+pGgxN8VE0uwIcAXa
Vz8IsK7dtcy/AVT0BmAzbAWlCmDrUEfjD9Gocpx80n6+gPQ09kOG9yVDeYjiyfqqXCbmfrsKnDwQ
X1GWwQ2rnKOgr8FnxTcwaSVWV8JbrPZjp+hu5ZbXyjvnD3KbhBP6DfqCyfhXFJzxnNwoZovr561c
hCCexewCZLlweYFDIg+NovvK3CCpY+1qJ3AcgQ0KCpjqsOYy5qUeEctbUqa4Cqfl9v5vzh+fJtfe
I4xToifynJvh27hBEiBjlv9T+MXRgyzD5oK1bM7aoBg4rFfE7GWHcPkGtRxRkeSoMHfd+F21byA3
YT6jCUCmsJAPfwJUhDv45qn/NTZPTFW3ku6plSWJyfbN7NohF4a0NZX6Z51JhPDzLqBQxRD1pun1
5vYjvGaU6ZWv+oRqKgngV4XJmtf7vt6RPVWbdb1aQXMMBb6rcg9ueghbwtf8xcQQNJpjjisGGXvg
nltXS7Jqm70o8xXiRB6XLmV+NU/0lxDX963HXNAwl2RaOngWUeWYcplb0x8Dg6T2M2a6gLh7LGn7
TzcNj79w2qwd9d9sO3QEhdXwqe1fLJtjYNsKJ8EWhE5xOx+6qs2C/lq53Z1ep80N1IV2taCoMq5i
bzBdH9RN1gZxUEz+q+6AiC7gT+Fn+pAeL1ONjf8RzhBEwk+GhBgW7a8C/znCvSF/ZfhddIRxMUsg
4LPCaUFNG2z6z3PJLzzHf8PSgSMr3dsZBILQLhAAAct58mAbLSUy2kGhQOvSTHzVcvnf3LTJ4KEu
6C3ClL5SRFAZMDEygPgHjocKPEtSUjZrtxHBrye0+GbIPcfzvQjTT8emmqR0ZOA3aODGiumTeHOF
ARz43FG0XHollODwhawPmsCHS5qGDiyspIJwX+6c+AysR4Hwhay64V0v+0cDUMBbLGaOzH6mAl49
JInwt6An3/b/4kPG0EvIrR50QZHetFUfb8W85MdIf1yBFIt9CF4jzRgD2p9kQHlT6WaK8DAHRj1v
WCQeusZV6Mmg9UjW9FnGzKFAbh8LrsyK9G/UjjqI1gvZ/JufwpoGrF01PzLidaiolCRSlEQulD6L
sYhLjZgINLFfy01wNviNnIk6ynQOvV6ZPrVXtGWNGylri3UGI58jAASoiaHEHdmJPK/oL3kz3l1b
M8n7KFraDoDVP3ezCc5Pqr5Tez71IM7mLmAzyJjVS2cbPYQtzjQzXU2niYwrtgtaPimMFyCN3Jm/
izil+ZNZlqhFpK2+dwqopkkJBdkcJ/HZDFlEdSZt9Zr1Utqkvf6I/IdwpMtZpdCjp+E2a4pBF29a
yjjqsyl0mp3JHjySQwWcmbWsKdk6Allb/xecPR3ydHHDjuSSb0ZsCT7QM9/Xi3XOzspt+poa9yns
jz9G0DGwRDZ8Ej4+57cEoV2LKWnxwZoqsDkUJ0JHa2Bfel/jDQjH61siwiGje1dl374FSHXF6ft/
tTEe1Vp3/0WyRV/1OJ7UzyuoMm7VfFuh3GcuBNF13pyiFJSdowl9UmA6Ym6+YZpGIpAHfhL/MCif
TWKAn3+qbylQejHU7b/mSyBe4QoyvhBZNAX2D/0Eswp461LC2jqAm6R8q3hEsQLvlXRkRshrZas2
zO1REJ3HaDn4Jj/uMSvaBDdLZOChugCkrR4wxpZN8bmmDHEXw4wndN6B7p7cpNgTaxPerLHPjCU2
38Glu4ZscqPYz7fobgkifTbS2ptwujBmFhEeSDScrUBcH4a+Bj0LKPYbHQVe6Cs52zs2D/9QI9ZM
ua//OyMNIzpQx/47EmK8au47R3RzGkyk0/ljDNEIC4lesyS8THQS/QzGDHWBYjekGkIZcsvhXnCk
0kdENKOxQzUBsuF7//i/CCrx+spNhLU3dr3XabGIErUeTvu+Pzs+A/bGa9P5Elk2pzQfHgC4NRhc
9TounCFwxlp6+3rqsa1pnt1fhxcovzfHLsof/tpzERa+ZP2ziy+UHUvCtDabRMB4LrcLoxm9YbK0
6ZtPftzH6MSswaRbYxgzIdGBn7WtkyLkhJI1aifRg3QVJbkjq/YzW4ypBlMEH7FUjM/WC+w3p4xJ
tJykBxB/pY0mJEk6AK62sAB8Qt9DoyHF+rLNKMSVzhUMLbChLV1VMTD/flWZcjfTePFU/8R4ejob
TcnKQm8jwFXz/Uxjy+ruzADIgjLVzB2j+CO9iD7LOw4937Hxh/EhFEOjbl2UKbUOntBd4uhsFoU3
Al8Q2RmBp5J2uCKtKQcJOeMP9cpOTx1uduwfCSjqM406cLj6UT7Qyb6EF/lTMzpB7wqYMnIUuaWw
JrDrGtq7N76qPmL3a5Ay2pcd5vlYQsZKyl+aMMiiSmqCTfC5gz1eVc578UALlz5GyG/B/6vuNPjK
lUhGJrDphJvpIs9GAvRW1qZSO1hiR9/XF39c28aeB5yD5uND84IyJuqsmNBVUlYT0OYTOD/MBSvc
eXD42Gk4Mla/sPE4nac+774T9ufJRP9Led2+WYiKMRyvdbeUmHFJ+M0wDVrGnYMs9c22q58CD21J
vRJgLDi5/U1bNypa0ii0GjssPE9gFmrbenpyhz8DTDF3j0yacfeTW1neoeqDNqnNAB/gc9r3Pbtp
pA6b1raWqS0PDHbEFXvO9VTl4qdv1PtazaQindvJJCLb3M+O8DaW1Ga8MFIbntcJw2X/2nF9TVLG
5ba/yfK+fwFn27CTrU44NBD5Kj8PbP6X3EzCmN65fDCQvslNTl3JiSwY2P9TVhzAXkDCUM/gp17d
enRGtITw9lGUESstBbxxh88mVce3rwquyF1C1FZe2ldGn4EOAomEjRqnLzEmza7Nxk9/Ow8LWXpI
RtA176PHkz4FooxmJQtSmS8OgJ8/iCbrRHG8xfOI1r22L8fP7WX0jUBFXwtRMIpQr7irtjPIO8Z2
9u6EvubmmpAmDdcD4snJIRs0oL7dFtVBpRoP08elY1NORl3r+G96ITnepfUHerv50INo9Brd8N0I
4aj44GpuJUkWyMojWpRqFL6Gw7nlnL395pcLdH3LlZ3Nyt01doWofCyMzVDm41JY0oYxHf04xApd
Q2hOC3z4TNOnyRbD09Gx41/fiRifx9jsmWc9bPn9HV/psHxT6lffpWoMAHn9yZiwEGs1tvINyEmL
Eig1hObhBVpwLZ7mFURUpmhlLZp1L33lxvQ89q+ckrHTsoGJ+socl41gVpL7UwXz8sB2Bz5TAnwl
IHjClX+2kgki9PVItihSdmn8jAT4v7oxvmrPUGHD9KSdsyj2UuhyDSMUdBnF4cssZB2WjTTARjqW
biL3NMbdwQVw9H6bJhQMi6pKXYiPjg0ZiKf+nqtYAZNjYXpJ9QF/71pb8wRS8wF9FihOn0x7+l/r
1dI9ul3kNbA4nB4AWpLTR6J91mro6jW1tlk6X16W79typgzBsiUv3f/c+a93692VcRdRJCCcybBv
Z8Ua/6crHukP8CqwKoXcmwEijbM8V/s+7ebgw724W80Fv1fjiBsGBRusvyfkVURCTk4uzydJcbi4
uJ+fWXhsfa5ODfG6pSi+LVXsUDnnPWq3FH9S9XMLO6iP1kAfdamvPRnJZEcRUQpYoXFb8ST3eZYk
WBElywYv8qme/M+v1URQDwksC/SogIuWvUycPdP3Q8Fnw8fIePB0OiMevT8CqXeFoqY5psNdm7Kp
L3JcX3zCkwCLTVk2JJYIXoF9It6HKNUzX3NC180n9YOXbKqkQXsw7C+cZKy/aseDu4ySkqLdHNLH
OXOxV2/xZ15xy1xAMEkQgUYtsgRL4uYJVZCVmqEYLwbHwWD+gYZnISb0dRBO8y9S+ma4hJkh3eMZ
3q2dVaxacam5ZwHTmbzDEJvvTonpKGqTSn70lzWEs+4bMbIuhEfziV/MKkFs/q65eLQ+IBu3vItz
yv5JkPNGRQWElvQsb6ttFOIsGzMfFeHrqFvC/JfcFl7q/ABgk07J/0ZmZpjHuMEND3AYUR2tw0ZM
3jSA3KtE597KGWgibtIT5B1Qd3oWyVaGE9zSn1ISvyW/bE0sdGPNZMqR5/VABTrOy4wdwxg/iUcS
b6a2lpRpVHxFTjC1n9J4cBWO4GO3Mce6TfnCPFa9JOYUcSRmDClRmlU7E1L5J61DO9UI7jbcCrAU
ajR+tLbpXyv69MbBY+zUllQm4LnmJeYsm/WyG01GqIZb8XxZreev6hPc6yyiuf2E+0xCzrpnvcVn
o4jyUGGBAHghjKfhNlw1VWdBO9yVowp6Wk4qMV2Oui3DncfPKljMjt0AoQr6sz7Qo8C6ga/JUoOZ
EuJmwYjELP7Z5soiip8bhmaU1bknHuo2MRMJJ4dMkKvkQOD6zqbn3arfiOEs4JzOgbmdHaTWX8mo
QZZ6W8zfkUJ1o0cxUWzZZf8wVE2WZi+BVwTW8qqgNANi3aRlsJ26wCPQbN6+RKFOAsURHOVOVrhi
4BzpWmewKtigrHmTlSvyguTpCcwq2U9L8KeMz80oFLzWqhydCXL+SmwIKJViBNrDIVXp5Iwu2zZt
Ew9de7Hd8aTTfSrQnBJA1qP7H9QMi+Z0Y8eprlZvqxG1qMXpmug/pTjgt34a1+kv9OiVm22EvJIC
97Sb6M2ESBO7sOusgnbfXQrnrQtr4LCTnZES5db2SGlQHOJ9PjmzcLzAnrExJ5purbeFkSeNMEUm
7a1JT6TsxzW9KItWmuLs8n0xCwACFK6yDxqX4gA4eZp267v0chCRLmPfIGx5CydyizXK08Ps2xlG
pbXM3KgdCMvsqEp/N9B8Rr8bgk49XGTTR9GS2YGQjsuntnI0F3sEWvqr/FkzhtoASYCjggOznyXo
9tHrrcm/vsfFQ+diXO5UhxESKCGJn7NtG7sPAFnK3cXvMs5HqcRm0qizY1WNKL+faJhAYlCFn0qC
tc15k+MBsaNE84L/xPn61MssbeC3w0rvdEoFB7yDzAmpnMMlIq5IFW89u1pxfXghYv3f9eZ8fipk
cgNZqZUDjjgVmzElrkUCQAqzrvSDHM9e5FQu5fIBIRAJnnKw4fEa06EHOTVZeVl9biGgHmp4Rcc6
LFK9pVscZF/+RYKgrOmxYkruQ0i1B+vDZek76dDJh6LRrfMFjJyOG/OdaRxvgi+1t21I/s8K+Par
QvTkR5g9FLRGpLtPAYOCIs6WpP7Eflt0ZbeWEiWKYNVUzj9TzbF1DDCFy2u1w/sKlfIc86oP+2YO
zM6EUOMxk7/ERf6KCJMtE24hhejzT9sZJH6ymHKb6aIx0Qc0/0zzXeKwtG0fySYROpprn+tUmYJV
Z6R0hE5VwzowHuIYx/kmjzBHolBVZSXXrNXQbu/GerlCD4R9/sllS3QSolols15XQ/PcyR0YpIbx
NkE+JJ3pfJfjI7EBsHDMqtEibqic/e2nf5v+Cm+x3XROYwAtDv9f5qQqykUoIeT7miyEPWg2fWXk
iLO23vyg8mgzxvntKXdaoehp9LF07z82LmHVZ4sciPG1qli1mtJk854lrwGJ6EYbe2Oa05jaRSgo
2KXi+UbtIpXx7znYtp/JWeBwg9oM5bEZePB5sw0KPyzvzCn47Fi4vWDSG800SqpPNXpPgAbVIzT3
Jbr02lXXSoigzlHagLt8mLROqSq2f9U5X2aHvNYE+QT2dchJinjxHpS+9j09Rx2vw7JrrM4lPBhE
CWpkn+ebTWiJ1zHpdPc3paf7HLjb3jJL6CJTe5Ta2ZVrNgx9vV1sBs4KLPoWSgO6ByQoHRl2E94C
LIZIMModRWXQp1R3X5ItDnwE3UdfVxrfuDO9uYbw8I9bCb/lYTY4IWRQ8HlspAX0EfXh67m0wowu
ibOpXNki9q0giOzK2HHrz/hdFITrJUwRAZzCKYKCw7bDkZAZ5duWQdiFhzSwAuZJQ0UsVRFwquPC
S2aw22PXan+UNP7JUGR5XZkqDv6xslYg+y3L9jNtcoH/mB31WoiXVvZMF+DkiioyIju3Nfzzsvca
DmFU+hjSFBhahk9bOMMpuF1MDPrEWb4dS/9o4lWpwPjXWwYXpxu1T5ZZWTCCx28erpRTtjJkw9QE
cguM5IDrwUpMU1oTL3obqGXI4xckzkSVQYPbYg0H/krPEoF4bTOeW3qLBOf+PQmkJ35NFspcppje
fjXejRFPzg6oMhEzcFaCj2mS4Fr6P+FThtRUWQXVlW4chFv2dVMYRX9ZiBP9j656IlchE+Yg2kjj
0t5SNeCQ9aLkrlpT1vp2NAJabdNk6a0Sythg1xuHiK3dSuaJiI3UiEMqSWINCfezNiRzhEs6AVOM
yUgfw0pTj8A5yzJAC2fQ72FVNMjiCYsRAr5TigmMsDWKMIIXP86ORLkKrXtUhlSLwDRNZzobL+YE
Dwg3yEIWcjnOlBvF3LUoarVIhpscUkPxQkEKOw9VPT84ssx9q7d4N7pnBkMSaHeKZuiDT/x57ShI
G+GhpoN2Xv1qp7LTQ/Qt6OnAn79kA40288rf5/ekW1pUpvq06AX3nfjZW31az9rbIkYxMaTzlP1I
BJUartuNR6s73Hhc5XHfo+6e+sauyvM2JTo2zu05BiYgF36BB4B1T0o80XF6uU7SPARzCOvUSQoi
iQeniBkZG7kcGMBRHixalJiB+2tiUH2vqRpiVsuD6a2mHhgh6pkXGalcus2726PtRyCYAoqPcfH8
C/CQNSOFVu5kA6gV9yRqG0FmvHQheis52AB5HNmsazBjJqv4HM3VVYin8kO9IP9bVDwEEpYxGRNs
R/0r6OwtRH//uimWWwo44HpKmRP9Bgo8z9ANGxLgRdMuJ1Di4w52lZ7DTSqROyUT3KUfBhxYQU71
jLtsXjIY5TgnHsx4iDLfnGTdD11j3qWUhBqQ6jtppccT26TPv/BxQUCuscCFEeYPkE2t+E9zZZPh
MdikRrqot2pd2lk5h+Yr5YGH2QElJoDhcHTpoWxP4FmlCOrAjktKtvKlwlsuGIoyby1mSyyWvvjZ
tcwZUAn10JhfScVJ0dFaX+tooscJA1YNYar3SSACH0Uwqv5+z/GiWyyfnJ3MwsUmoN9k+4NOmeGb
dpPFVkSn/Ke+sy1rx/NYwFmcDavcT6S92zA5QYSJCLzWBIq9NF3zAiBPLlwkzClEVfVpajTRnkp0
vWo6zU9K68pPyvynUCX60iFCmrpvOQvvOdtszy/8xK/CT0lamSqGE1E3LE4PpVlzXbMrm2aiSrXj
/4HzicanjT36xR74+UUm26Cf2bIw05ragTfV4IjAhZD8o6ELUeJrhQMy1TaoiJCbvtBMrGw/kL3S
+EdiHUBWP9fWWnwoRSCvVrHpXFJgKdKWwTb3Z33U2D320dlmKM4Xl4o4wtQkBZSKFMH3UmQ/AUL2
WhkqaJtQB0eTWWcjgGtjyBooC2MyM0hFRQX4qKcThODI/AYZR2gvbxo0/qRKNi1ucAvhuJkh1kH3
rfIr27opQwmVT8s9D7pKGsoreMXL/ekXNNggXWHuoBaRcG+ItCVkDIHNuvCXxXNcIlTnKLdU0xVs
SCEi+N2dK5AgHCzEFeollM0i3mRIkn3jBA2ZBCmLflqLqkWI2yakQz/EYSOiEElWjmtvT/2VWFK/
PfloGhg2Tj9pjr8HZnJsx+BzhrcfzQ4tGVhf8Afgvhy/aqxaY9LHd7/blGgBJnPGqXnVdApVftKf
te9M8IayFtFxzYehpPkEPpGfzYlGy9uknrVzAs7xwAyD3kJks2O+vIlOAxcyea1p2X1eCCVXq0hG
bquk1n9K60K59krSSxxDsSqrO8g+WUpdIQz+ht3HxSWLr6SyT6twBfxcOD5vcL9aBrqcFSdnDdKo
KBtsDcTyb52x6imAuumg3zOD8E40ip86w0Ob9cIkuujWaOdyjBoscnQIIIFQ7yt5kIF9br9cbslG
jmjREECJazicxZ0LQM7TrVqGbbWcWtqh8xX5r5tvLad0xakqfzPKgiJK9JgsTmwZ6s3Pkk0FQTps
0xIQriNmchX60NJDa04YCk0vBBZI5rXzPAZBNNklV4IuNlUTM9TOHcJNXkfK7q1klhiV2D+z+5h1
/J8nVl424QR2sUvQ7/aSpCItNQtRztxY40wxfEx3MqZUz5jEDDarcG0k7xS3/jcC0GNzJqLCxkpz
FQW6Ff8SAI8eAcWntvyUdNHjX1KNa2eHjYJnpfb8a0U50ze8Yj6jEYSvsat4D/lUwLvHGjG92rSq
hsxvt0xVWlOOPlVxt1DODy9wpuGG2/RsLWFASVA/N/1YmDyxtPgKjpGjfvDXBzihcYirnsIR1+XU
94huY3F3PQtVgeIOHSJZBlEuFthk7DufnW9CV294+HTUUUrwDlN+PaUt6mV+Ly30iXmOgHzRQIRj
+nsqIB8BTjAwifwk9Y4KJt1mARY19YgbEFje9eHyfzfnWNdVIf6AozZy0FzXvjr6pQVEWqnmn2rT
awub+fM05FWx7Si7TVlzn0cks1doMTUjduQ+9YR35CYfhw1hYYww2s+VhuRCXwGq9ar8Bwoxsksh
DSzAOyD+UCb4ZBrnS+VENZ/V2UnCfDP4ex26LzNYpEQUX6vNT2tF0NgWpKIjdJS9J0wOVVAYEvHz
BhhlUoUPF6jiMfpjQuYhRjHH74m3+D5RGb0HdV+FIcmHhH2aVFAqtqq4DRrbDtpVEa/fvxK2pobb
cWwHmuV118vB/WPXCpU1ccFA0JofyCKcSTDp5eTtFB/0gcuCO9cZ1CeUaZ1tanSgpm9Sy9Ck+tgi
NBnbQRTn2QsoMq5Upc2UC1J/CbAVEmtYmoMSIILJvS7ZG1LoorcIOPP/irJ4Q18qOkmDDLTlqsvy
gs9VMDqq+Sqy5Her+5JyF8CYt8U1cr6s4ix2uzyr10pO4+qL5nC+P1f4ziKgOn//jTpXROVq6XNR
/qUE/F3qZpY0wgFDkjMrHzWgIclXHnql3/2VguXFZBli6Ly07Mon+nK5duozEEUK684u6QC67tRN
v5yO0MFmbIWXYSTlaTwjuM0utPG16JpNBU++l4qqHUaBsHZPnz7kWwRKWCciF6WJ8Ff5J0CbwQRk
4lsmPiS1DCIW/ZgDl854OejvXq8UNADUM+y3IiqRvxh5oy/VJqpcJ0M+d7Fw59dj7Q2U5r/i2NUn
VDLLrAMBkhLWUjlXhgRoUjEwc/9PKNLrE25ewQpgeKX9kHvTyUuYm51hg/6gAihXC6DxTX7NoM2r
KnXDG1kxBfzSCh+/49siDaRextukbBxcwdU6yWDwlf3O3KypZY8QY3AW9GJf6QIWNjVlMaRw20JV
57GJMfJdMvdgYNfTX5KHyjXxEyDH0EFZ5n6u7l/rt93NI5YRLjbeGEDvsFhQKjzwQeupn76wB8Mx
P0f/4w3jLG8YkP5k286MgrUHsI/ecG7ofDRXzQyEvWhEu5Pc+5TwdKmK9nIpJLbB6B29tTGjCCro
hZX7A9N681HmIGe9cyBQqekdIP4N0NDYypFwchjIy7+5LgO8teed4+q4nQownVxwqqg173fMB9a9
Xgf4tBhGRZ2G2WS8e1ewaknozP+O0hXnGgxBvwjsZDJMX7mbReRRJxqS0jor69eFzWU416AfeXr0
X0b5C0SZP3fuezg7P41o4m+KZKOz695cVbwTk42Fv257WCln2H+r/hljCPBlxMD4cVPpH4K0uW/O
sbMFl1rta3ilZxpn+t4zIUhH9rE1/Oa9VxnyFJaritHkEnhWavq4gCXbQoSBZwtkg7vsaj595FB8
2z/dnsnrs0BQz14B12Ka9Bo4/wDKWuOc1cHo5idjL41mvpd4GkkspEhbMpsEiImDnZx/yfF+jc1I
kfxZTT2lj4dh6AIbSunN5jHkCacD9f0oCxvgAOXmu/CKWTDxDDDVlDOpV1Ly9ByhxW12cBuHRWFU
Fj+IBEcoHW3BSdFx+Y7+F7qPgk5sWoNpUZr+tpDnhJqCK48YARt0w43G9RE0qr0W+8Am+v9QI/I1
v7ND5YMHbPLwXiZvr3jW5ZPzPXgYN7B4+RE1NSTFNxMo3qOU5+wK260lpYIppcjknOrmS0Ze9QEG
qZKnl5NI8DvaJyy/HQndxGDqsl5Aba3VYeOCciX5yLCQHH+mAS31S04JZ1GGj8nrgV0H5kC+gdSY
oGj7riDryNSNqAuTHsSfOEbXHhRKau0sIon7Cdb+22Jt5bFiq5nIh8C4VQgj+Jm+48wrxtDjLXQP
vNdGsGJ8vocPIr73hLS3f21jzX5A9Lr0bKWE86w6pKCPd0lx+2gog7hZEqKIqNglrax6r5kNXuwh
3GhShnUPOjlMJRtTcO03DuAKvaBriMEG4yTgcN3wloRqJI7dr7Bca8prqYVQqmDBNd69jv5O8hSH
oSaBU6mw3kYW3j/rlb5JrrlZ6YbIlJ83LB+VUeC7ixgbVfWB0ge1epLDxo8B4T+0ZJXv52YTe/lb
p1Low3LzSf9I6+vnSf3kfBnu5yhXGpoa7rj5YGd96gi4vcB+Omy8fCC1FWgcIgvL/LzS1ilqczdl
nOcw5RobvZCxJqgEOqDVf5km9rkQbeMisNO2xA8ppu9uxMIPMbwOv4ZQ9FFT57xFTBBwyjkTTSUk
E/IFOMbZLxPIF3NCQILFzUnbtpK1h+88yNjdYj86BuG+iVU8VBhGobRgoYoM59MMd5L6+8Zkzim4
PWq24G/yg/+GyMGfIzfhqJSxuJWzsHKsqoV50qJ3HhlCpR5l1NhoccOMrpu9B2n7KVFWSqRZodmo
ZJ53ZUs7KvFcjeOv8pPuLdGNCu1iSVNmliHVF/0pFp02yZCaIqcfs7KhrNezz36kJJ78k1kk2vZ7
c6l4nlS2YKRLF81CN2dPmI2L+5DlHiNrgEGsrSFvQzSzXZAnv0Yr5xAt4KXtNFv+BVqK9iM2MoPM
AlhFbwc+/mEn/njB3XRwNTkbaP4oAfLIRDvXd1Pzh2YDGygVPa57Qy/sS5Cfuje6EGALPzpLaJ6R
KRUBwe7UyIr7D851/7yMOV1DL4KsvEv3TeCQ6dG0mAiwFipdP5na8cQHEvjzSLNupagT/A3g99yg
ymOALtEkCQQO32JQqTtyZk5xrVLEwh7/DEWPxuPj5TiXtigQ1XgpqqClnSI5z0d6BV7hKbsT90Xk
yam0I5jouEbVRNrhBrp2gnsOVH7Nh5m6gKhqrZJx0YEe3Rt/R3hwAlOiXf3FoIf30nqlPKYDXHje
J4fX8qzW5RZNHJjBXnoGHX7m3bjOYWOUs5oqOtqDre8SRkRWk+BJLhVEY5+3MQefqyZDF4unhLAi
kwUsI2qveBRbVDywL4qRkNPBLGgHfqAAXcfgybX5c1cy7ZY97vyN9lQUlIEZLBSySxYDTLXsRV7L
io8IfzpF5ghwFAz58TYtV8wNENnKPeBdk6VzXy2NBnl1U0J23+JsRA364soA5t7sdApjgIRXP2il
1n95d/gmydJ/lxTJQKCLQ8C/ALmlFjyS2cYfIuyB+h2Z2TXDaHeUnW1z5tyMdCMRNaR62/FRQ+n4
ox+RaLZHFpyqhSIJr2Hq8977LTpO2aXj3u/HOWBjMjsbZvSwKqw4ac4yP2gLkvRk3MGn28N7mV1W
HKaWPwczY5qjDTmByxmq+6djyUA9is972y+m0nLRGq/iyQxCPLIjK71ctrpEd/Zt84qdu2u7SUgA
c8qliWQy5CCjOWimMM2z4jyVWHI3YJGap8NYFQ+hkVE8hc2r4B13YfQoaQYKI4jJ7TYTgfHp7tqA
wS7wDgT+XcEm8FsqJvor2dsYBipyxrt4M2X1SI1gIuMTp+V3MvD/Nchl6yOCMkL02tLq8+HHJSgi
j2SKlBNQAptsmoST0R31fEqI+0Gn3NcByBpq2Lu9hlTnRZC9grARqebYkTOyKROPHI/PSWykfcgI
8bW5QUi9c2Ha2the/PZxuCOXteuzuuncmbNfBVrUHhJopWfiuOgoSbC5CqGD5iZrpZo6DsZFCGka
P24PUoWrtaWjDjDIp2v+5dtKNd81Xwt4BwOwxqV/IZtNZvltkrqo3ktltYmoe+U4UBAY/H75WNCi
wKKRJOpMvtHcTzHrnC9fDpW0JG5vJ/l3BOOqwG3NdYmVkvRDDixMPCvRf5FRk/vOxc6fyyDIOkeY
VLUGphC4wZqSvBzIbYXK/Tsk57LV4oTTh4t2k5aJzYgD7wo3f8KyMluUtgJ+mqmYHMu7fiBHt0xj
/Hff2wmVQfWm6cTFvpna3baj+blzUOwpjb+GTgPz9iax54YZlVcwMRnbPJ9kC3EIa+cxPyDzOHou
iPfM10QUNHH1MRLWl1VLyMSFKNiRrnqVFV/GS0G+k+wTWUICT2pr9IZhTUOIHKYpXZCAIIjezoLU
GBGoaV+JcHuoWSKlbDBQkegtI1pBGpqEwjvp6/dFr3e2k7q0SOPpDoYJM+nNTjC8IgRMgyJVhaF1
cD7FCIi9Up8PJDow2rjN7pxUe82a5Za/hl09d7BDmrSu+fQOB5pwsRL4wshcHokyYiGf4qp9Ipc0
lE1gJVkAglFDC/zQILKRAG1bPM14g7z6L/7nbFRlzocUZ0zqTiuQYo37zM6sewcQSJowRWp+Nfpf
446eR/+9yUs29Nw3AMdgHpwtBoAmJ6cX0cuDdcNkusaBIPCCKYkQRlFOgC+/15lWgz3/11KYS77W
pQsUYtkI4N8CvH6r+XQbcy1szQRL9K/+EjsnqqecOOgKoOQ/sNhlx24K1IgVfISnIBH1pMnj4upp
JxFqaWDXYaIAGgsKCtMkHfz6IaUfeYYKXb7BOevz7KOklz2KBsAxP+JjYWUBLH5UPQDDieo3Onn+
2jVGLfN5w0QXQk8eLVLHxACy01CqbxiQTgTSJgXEOlJM40i3A6KnIktsBcgubetTo077f0POIODR
k7BWnq1eYaa8jd9O2Nzgxv6RIVoZKqan98wKpHCLi/bRLtoUfOaO8qiwDgG5HJbDIhdJSnFGwn3s
pR6/LX6Rp8ah2nYp5VZnX/xQcXj5MOtBR1tARDvYBuufMT6fgEey2ATSkavpqprxsSxebBjcz5vo
HB8x5ARJ2EenKqSPBCCLdftTVlDQYGuXjNwjJfyKQKsLe+CcTGysi06fRTb6KmAG9JpZCJqQ3wZI
Yl5MJ9w7yAQNrkJvgGoXjpNhky5OVBnrhsZ0r9S0w4+e6d3FqTXrwoxGsMPO8LIUz54F6pQbD/vQ
OIPIYLnbyiw7e2ZyvbhoGpxAXCOA24EgAwWAwc+hohr3fiO3VruI2iU4zo4trkQTWrxLK8BIFzHv
+cT/Dutz11BT7jt47E0kedgbEfKUIFTLUOK/PFLN3pGrSoND08iLns032WFi1Pa2OHxggmUFMxJ6
bc3yhsi8uU7FeLc1VhKBOFiwRV142LFqiQEizzeWn+bOETUEr7Xiacc4d9GjqfQOpYycG4OmyvMm
0seO3xjAmML0zod7z4DUrP1wd8WujFCNzVb1nRfrQ//vSpDWd2lCtzv/hxagrXsn+9Tm2IHngZPS
/DdyPWbPl3xzAwPdiZpXUXLiRPVlO1R+K+w7FdHKpO9xdNibKu47zwtDeQ9Gc2RqyckuO2+c+OX8
laikcjZGVD7Zr0LLqN9u2PcQbe2SARsnjNbKITA75Qov/6Z82E2Cin6ccTdg5e7CDBn3jg9dAgJ0
is0mBXUHbHOgNO1zabroEPRuT5t5Sx7St6JdViv4l7VzF/0M8Dg5qwuwN8azhZNZV7kwVQYGEBGr
4y9ftdUBADNStgg/ybgqY3sTfbp1Spqs3uupbE358tNXwGrehvlWJMLXA9RKtRZC8QHApiQWFu2j
qvdSqPUv365KxYq1DasOXeiX5/E94GqxeOiWIq30ZO3NfT+fyT4Ek57j6exJvLFTWIL1rhLcc4th
xSrowify9AeelOgIv5wVNCeMbDF558YetZJzbZttqELQLffXLAtCfpkOZ88qIk+7lfAx8M57Cq/j
h7xFb17fPNqr9cuhlRhck7cyJxZkDPQ2Tmf3XWVBwU700wd/zwV1dljzx7P9JIvfkT4UWYgF2aPT
34vQhZAsbrUbBZf2BsDMxtpaQea22i0P/YlDKmBVfEWLPHGTnz6Oq5Lh38FiG0HG894wuhLf56m2
Zje4753842sk+EilM2XFWoLFv084MX5geObc2jD3dKdCZbOK6lYohakDIpECChkLZ2NXLaPJ14mL
GZX1xMT15OodP1DV5cQZEt4S2g3E64I946YLrDiTyrMg58Rr3NGEje1yLoDAZ7fuoVYycQ/FIO5W
czoQk+r/ESu1Quuyoaw3zW329UGb7ZHc+oyNrkKtU2JLkPytiDpTh/N0oiBx+mOUgWwY9kCOLdV2
YlE88x7yb+xGErdHQQ4+q8tN9FYTa3UnP8L7l+zSP2ONBoqQlBmHlPBo9hmLL8VDGqut28RrHaJy
GoxMSP1e+4cz3nyCb8CtH21YlTCW/18WeDL479F8z1XGvSbEoJf1Pjgrzf8dgqtexpZDKjSwH8XX
y8Qn5gVxTvCjNvj/FhCj8wska3u1z9Qq/7eeXuj6Ylwh8hl4BwuRu5fmJgCaBBvE+rTD3JiNBUVh
BXSWECOeXQ+sPtS9NpgoKYcQA6Ks1TWuP0utIcYA5OVhCD/zPL3Ngnth7j9g+FIqs8DyofA1gz+R
n4YHKpJWJdMizO3vd16VasWtKCkpPWe1WpsSjP8/Yaw9JsJK9MgnVZz9a+zxcb97BtldC2xX+y/a
VDoaeaqQqMO53I0YCRHlgrTQhWSa/ieENJfSMLU++HOVFrWIiAQKn8IIlhg9Y447xqdiBU8+Clap
r+zffYn6bR7mypVtpG1gYcrzwJVroMyeH9CFudfiL9jmzcrcdrbCAHBWRSdSeLs3audfhmWQyRdN
ke4tPcn1gPfuhTEHbmTyWqoMvRlInpzJFaNUwJOOg5SC5c7zOjpOFVCQuiTXZK8edyp8fVr84Nfi
XsNBmBuEgxWAYOlmFy1qUwF0ntJcjviln9k9ixrRRp9KWZtde+8YtgOBFV+k1iQWNj9Nf7IvG5RT
5e4cRA6fN55v80NmBVc1SKFmuqYDpIPtdGeE9Ksg4d1DoBRhYjAa9p6ZriMXKAqF00TbB9EO6tjC
E1QxPi6bnEN3gIMfPudI/ZWlUStTuw6Ynbrv37JTo0pWNaTu8B2JAynOphP0Qaibk9GqFxUcC53m
c/PJalwRYJfJAq+hbDwnt5lFn69jdDkONDh51NdPBARy70+/td4MUXGSX00ZjvcqVKUIJkxd78uv
9COxrS9xY9XK3NrRT0WlR05ho2zfzTOt3UScw3gX5J9bakWMTrndSgKJxqKCe3U1qrqMidb/h1IM
5iOE9nLI2LEFpPAc6g6KtWoRVcu4oTc9X+L1fSwrTBO7RrRRDO/H1P3GitzCSSEmVOEocJZU/Q9h
iRSddoFKrdtlAJhIFEaYuwt3v3znPTPesaOJBgYoQmyj/VtJWgQWkgIxxpNjkA7dKSP/xAn0BVMD
F+6JcrK+sPoax8Sdn0u3fDtM5HOynHmygQVL3I1lS+t/n3dVIXbyXvrFoGTNuqdRK+PWaLAoq5Rn
BowiRD/nAGnbt0pN5eV7m/+a9AqVe70yVgRumjVk+MlvldfyHZdnFG4aroUNAAOvOqfGO9GGtfOM
WJUhfF6aC6sH2M25Gc3T89lNIz35oPeMk+foa7nckjfQxg01xp4PhxRVmDnPJ0rPXmuiQwjVSJ3D
zwBO2DBN/S//ZtJT9HPYr+30kTk6v9I+bnfHZkiGm2Wcukno03Lpi8FEEl9gbx0DfyyYzzOL9Jh4
taetL2wMy5r50HXQ9qRVxW75AHYfQlqQlAm8lthkKnncP9cPmthWA9i/XZyh8c+WOrSX98kYN6Lq
ZsIez/lwhuKmu/H1ZzzRQ3BZddUD2W5yFrW9yG1Zg2JSynw0Y8UguRJW3rkvbblI0tvHzVaUF193
xlTQgT8ec5Y7adcY2eszKYskryLWbCNyqymPpOhqxoWG7KCwL88NeK5u8UzLlseM8PcvRtSqSn/R
SW+lnfHb3Fki2k7jqkWvjJGTJVROPQpvezctxOn+Va5FJ9xpGyNd2k7t8H9EYtG5tL3O/sfUOKDJ
YltEi1gm03sp3foZoslp6bNmFvYhzXWoIq9Ip8cxajJA/mkqChybEP9ZGmuonH1ZXqDT4C6nrUjU
p+8WncaPBXF3jFIs1AxE8QMs6RsbETWGwLKj4bUA7W5ORiG2XrTmhlq3pMOl9pQgFur23H5ASCmT
wIOvPuCzZgy9LfnRo4NO/tlRxKnrdh35DcqUhIaZok1jUu9b8+ns519Gfnfmwt8YEid1EZbK5JEj
4qOfbv10QRbgjY+peZDbQX99CRoP4xL6Qx7+AEd2hN0eYFTlZYd3v+C4evs+WwHow1G/wQYhyZVD
9Dlku6rmYy1mem5L6AofZDmdrZP1rcmmKUDi89qP30srksYvjZDsCuYz8U4P2legh8Xy6+WVVxAk
z6Q2mudaq2+YUxfWaKD5USkW54iowWTDitzoqdrWOUAg5/aML0ZUEcscb+AdDjVPkmm7yBOLFuGN
HAu7X4lX3Nn7GNZ+hVWvFbMpOwThsfMQD2ADrZB5ANbtjl86G8bZSZckoMZL8vhq/Y4m7E6oqTuR
CCReFC+BVslvC9ehMSevV847RoqijnsigIS8cgfDSk0OiiHPhJXNY9qQoOUQ1RjySHLGEUZyyuzf
mgaVvZHF50seW+yKr0bE41ePB6RB+QPDdrJp9kO+O+wVZOmcWmMAUzK+3/pFYASayL84SgInlK2h
OMpjh4q2NrdcV1/DibHO12NFuq46LSCE8zCwYc3FuoH/IWnBwySJ68XS6knApsPJzPR0VptxcNHo
jMKnIDvlD55hO7A1h42ThujYibWAy7Xi0sQdeSCB+bs9bNjsx0qxIqkwCMg6XtSGqmvImvrRm8HE
Uw3DVqP5lZokAqiarjGgQGC4TKtyqiTFm8GLuFKh/3EXOgFvAylagJbJmRKOwC/a/LBrz880AEyV
IX4HtltiFhsU+wwKaMWbMZwnz7fWKH7I77w8NxtfTQTFoNFv1ubBF6+kj+sD/myq/YPFLVsdVSa0
DDyYhpNsOt77dxWFHpuSVmuKf6tQJna8CLKLMX2rOa8131IBO7sqwn3ULEpZpG10aLMen+TAUVUC
bl4c7J7bEF50oqLGQqbJPf7kJZq1IbbIgGRgG64h9TF+p4pQlA7GlfFCi+0mBH90O2El6tjMuNhj
6Mqs/TIBAH3Iy0p68TjQ0/BVebW9zdOBqPf1dS5ADRwP8VoSyMnOvTLZLZzm8je5g9KzoUaa3sJP
sTaxE3M+YP82yotQih3jsPXDkaHe/9E2OQFE3USVFVFLiHeGQEq2WwV2O7x6isd1NVkESy+E7onV
nh4Yb4SZORbjDqfP7CVDjuZdjsrIZ1No0IM2S+i7mwKUKaOgCie85WsLfBqYTO7LICLiQJfQh4df
wVrQcrHJ4W5b0waT8QxvqVOKA5BhbtvXiC0m0tYdWkL2Pj+2Z4hiiEwEItyrrFI5HfmQbu+MMmFy
XBstcUUpa72Lh+imMQXvXo+a1YW2ovVztmCoCFAHNY06rMqLyuYwqnEeEIEDHEMT3ePuY/33r0s3
v3x97o86wJxy1W8gAEpRgGlQc1m36cuyCprStDStErNPldLHvUtiv4g9QMrLAwZ1Q2GU9audwknQ
/lzofccbB+7CR5rVF0/vOblGk247VBkKV53L1yMcfEbXBgOHlyhqRJ6xH2oGVSpmqRZGi+XSKhuI
mYciTXCPA/71dYjRhEZlpEtIMgN1+429X3WQJ/7IE7RywHZq/ON4r5o3S3hw+4ZhaptaBFVw0zeg
/Pc9EndZmvS/eCaE/DyTnVWho+Cw30eieFGwuebXL3RraChfxq4zbjOAqubjCNTgfHkp1v2AXp4b
oo7/UsQFGzrFdQDPvUWuNub4Sl7ChhjUUYvWfL1ZXWrmhWyarD/fku+g4b8UELya8+lmGFfAnqtJ
OMUbWolpWYvG5Dstb8h006gTVCYdcQ/tgKj6aVVJgrrKCPZ75IJv49sdbiBoK9UmT/OG4Mx3kw37
XknKXyiM6xsQ1cP4L5/oW0NyU0Tz+960o9XpR+oFcBSFa7mGxb0ZvK2jDAFeh2WMYCo00kZq6sGE
eLAnhsrL9UTKWHeNqCeC6pSC+RtAsGbjuZxlijv/wMzo6QeshY6SqeYEnsvaM8WyTMtXAaMGnzZs
u3JGTENOPa7R3oK/hwG/MIj91cUKtuuj+3APE5c/1RI9SGQ7/BujBprT2OR28vHZAJ4N/UF/CVj/
+CHg/dp2C49x9JI3r6Ik/XPdesvffSdQMJg4rwcWjkJQaFjyI6qcZCCwi4YitfajGvls84nWz7rh
V8IAvoOqePbjBBgjNTX5w6Y5Ce5WoCpmLfiivLYDtrckC1vwJlIlNZQ7/+BsGTg788p/2RFm61JH
hZAGd+xWkJnwf4oPxHIciieUOjpP4SFNPCgT6y8rJ/fCvTyQKbyEbeIrjVI8uR3jVDnIbrPb9wxH
SbBR7Fl8N6ahCwGhJx1yu+RnECDjTUtUt6+SomhSq3KlxU+nyyfVkfWHJ1O8Vy0F9RvKbKuBmAt4
gJ3ObH49bFGLkVGvxad/LaTjQVjxG/4C2Tibxt+BuUJh9XSPAOkWnQ6IdKi65CFxi2swNlcg/G0z
Qjmlx91IRGy85CzV0dxwJnlN6euL74he34SPWpQ+rG7QPArumwlLjOohc0bcEy/81bhf+0eR0Qyv
XAmkFapd+/opCRH+SEfDRsVu+oHeQ6OzRgX5TptNDzSZIIhSxTV5+KTTENdlofkTU/nEq4vG2L7h
x6PhOK6DzZV7q682fPurZJ8MU1Jsqn0clcpC4/Y2vzACp75nlSeHXF8Noq67vkQexVSBrhpNy19X
k9+DZj/Xp2qJ6gbSr7DoGPuuoDZhEb7Q+TS+PhgjLKrKuiljegsyjRGKTZp6ZZz3ascoEiyWZ/SH
qTlEwM6F/1IC/EGoTFD4odmxRa4r1ZrUCjqKOJhdpbbaZmFO4UXr4D+DWNhv0Zg0Utnbva4v0O8b
bdPwMyii2vxHmmhakbSL5zB80yscE9+pl1qPYCcDwPqgjP+Zv0UBWCzxJhnyEItpRG11sQ9yQU4G
km65ZXsOOfIxCdX1KJYbSyvXHz+lCLSlo1gNsf0uVn4xmUAho3UvaLp8DpBXvmpOS4YSnOeVi/hQ
QWD3ij31X6zX/e/IZGN9UPhYpgxvsL8fKj3L9sRSlMsmszGXWSJ4P9Gisxb93DsIs6EIs45qTNCj
RWvcLMYIA81bOEWlZv95L8ZWOIC3nq7XsvakQRDpq0hRVBLvfwb9/Y8WuuAn+ctmKdPlGhYq6M50
qHLdko52taBnirk0ULvTHN/Ljc359NnUHyha8i43cCyIzuzCATeJUuBqWOkioQnKSehT9QfZ1nsN
HLUbPMQNglmk1DrRjUNxpdmdmTpcFPmpvm40lVmhIUMX6ICpjIQXTBgOUadjbjOMgUDTHibknm/2
Pt3ZOdvQSaCRSevm4TyfsLumgHQbWHO8+EjKOMNCCunRv4H2ueBUVY99w+brjEfBT8BjC7Z/NNH/
KzvjU/plyn1gkiEtU3FdlKs1BNrwdZ8KdnOk89HsSAeoaun1i0MhYXKJY38BeYRSuAnl/VbQlx7m
dvKxFp7vy00+5VwLdniqQy5WgD6gO9zN4hnMkOvD7czvTDOba189ulRevoBS+rRDpXdeab8+Zxn+
eoihObTYhvIDzG80269uf6dC6+5byFeQIrHWeRdS9WGFYSOwk3irTSBjB+tSKg0fHjn9qdkZtllo
+GE51Ys07UK/pR99dA7I2UW9Arw9H6OCkdDn5mRxg7aXdtHmIW5z0ZOzoP+vgpOfgKiHbAqzsVRI
HkJYJYgJKqNH7rQTwyP43NUM8ttzkKmF8yTMMQ5rva1faiKYj7oX7EIA0ZNse9Ij5U1f4lvVzfZz
e3mGSB9mkhZrJePvYVkItKJA98qpfHBPGnH9C4dWVdYf+45OoHJ29R8z5O+4Nv6Pdeix2fKgroGy
Sd3HoQ85HKorC38G/UzvV8oDE0pXqZW/rGnAqhTzioI5c0KAXe/OhHhhk+ciMYOYC3bAD0hYxCoB
SmJrNycqDGQanxQm1HMSACQg+kKaPV4gSfKZGGEbmTX+2ZLvUD1bbrjU0FHToJ07rMoXPciHWURc
hdmcRXgz+q4QvLKDK8EKulpPyWw1T8sbP5ccV/DXpJH1oM64t8VgdZ3fgFFk7uuGnXeDAAw+ipet
GJuGG2uEqxkgl/2wYhnhJsFpVMPZgPFxY9qAMaLKnwsMp7PMv4fttt1le4rjcb+egoorrsmvFIYV
MGv/Lf9CGxgmWtfbW6DI9Sb8cqkgfBdLFztaNrhfpsuHsxSKGvnscLfDuOk4Qeyb0ApDcl1IX0zR
2W+5BPsaDKeaOD3ARx8eLDg9ayOCNYsRFVSipDdZrKleU+cnDSs70mvhU7ZWBbsDOjSDF9GRHQXo
kzYVQE+3aURr3yWv1m4m0fFuSIlb+Eyp77FwkTrgSZkVVIa8gP+RagvSb1MRdhvosCLuyyGu4yRN
rg0VYoSIJmFsQC1SRoMoiS2u+AVRZmSKpWYqiqCddvMJNxQ/QEsH31UZtSNlubcYMCJPbDj5TPgo
22DjqDclcGO30txefd7FAV2+9JSk9uikRZt9aAgGFR7EuGIRNW08VkAYVGh7HowCirEcCzZ+kQon
qkdNYR23Cc9YJmwSVZbkpRTRNd/Zwu0Ynqt/fenihzaByV5g99HI1Cl9oGdpmHQSt7kx3X0eCgsb
gt2QU9T8D8JN0A5qz57nE5w7W7JjSGfXgZ4B/lWU4OHuEeslOjXOEGQkS3zMk/nBNjD2BvwA8lA9
+dA2ATmjH96GHgQTL0+o+bi1C8noQk1SOS9ZkLN51+Q+04XOHv3AEdI+sycoE0Q/AvmItWU/UXlJ
p8DStf/ZuKJn7I84iZjBdQUZlDyv2ewgdXU9ep6/R+oDRDQF9mv/JcSHU9peqrWQ+d6k426E5EPb
87Fj5ClN2A8Oo2LvY2mU2P908cppzrFWFcevCJ6X4JZiIqDHlFASmI2FQDeFnQIDp4hFbIEvBttY
qLv52TseOAtTggzywEmdXDG9xMUxjUes3WThCaUrraXmK+fs4gAonXU2emSAa4jcgNXeTqGnS36c
bK55kqDJLCpxmM4cEzkHnpu/atdgfBjjt/ya92CXBTiWspdemXHAueJw3oifbktTXfS2d29hwMVj
TXIWbZkmrwh9MgAOz89aS5j9BpDwfdCsAQBieUJvSY1OrgP+AZBy+H5zcA+p8EIzi9OQKsMv/BQB
Lnowb20ttqE1zBcsZeMy4CJCgPnhM4g+Ijq6JfZkxPHplTA2DgGSDwkR4CEwmrEkzfJauXAIj5eM
Tq7Fc79aiimKgEpi5YCBFp47HtIKBrqLvqDVefAeW74h/A/3FqQc3L/ZeGTWQTx3SWU7jn6K2ltU
zmTnI8AF7NyAcHMh4YlwOI6ZRQuKq9Xo/DLGQ84xDPJkjhiPAOsqnzvt6/0aDkxrrNx7co8ABVQC
zZvd/FPLUDTeN6sBga/Wd9OeE/pckhNQJGrfEmCjGP7VrodDqfar2y98voEjaLabwTQh6DWT68rD
1nCgdqD/CC7ohRzjQpkXFdPATcFc0WTyEJwWbCVEu0wVOLUjmspjHE6UgdgpWUytKcuHgdzeHPmb
920TuULd5uwQ9KXeexuK9m+FUfxY1jJ/FzNMZ3JmB2D1Pci1xY//GbtXiU71JX+KSmpFuHmOZT9W
EMISpsdcrsxqKm3QUgrevDuijRe71LjK5Da06GqAAbt97F3f98HlgGykx4A2M9nPfHrFBndF+H72
DMA5e2X2p2QVfRqqwfdYp0a+Els6wlx5I/98Q1CqFU0ud91Wf35DNB2gUMrvsI9lMkvpQz1ObAs0
fZV5MYNluHDMvjMnR8cRht+n66ZGDd8wU9gPrXUpffahtGmiX03PehkENAnUuVMTVtlM8EYaoy7Q
z7/bg5Nl70BVpsz8/Qvu6yn6vMCb7XNMr9Uql8HG9sa8l2nLvGH8Fe/pr4C+398MhEy2EZe9nTBB
kR/mMqULwME7XH4vfpt+srtdZxUDYOHld2K5Gjz4x93K5hd2j/7nRMvl/xOr9zCNvV2Qg1xsgEYU
13/znfkUfLrG0W5GPjCIY0Okf1+taqs4BN3y/QoDFqz98osRDzWJ9OcgvQT+f6PnT7kXbzOQNbQ0
Raf6HJd/PZZG2PBAuFH91trHkWr9Z9dhz8D2p8nPArfYqr7+5ArgTsc53fgkx2j2v7BmxFZFO+7L
EneShbDbN7j1zuRkJ0kaWCghDQ/tBHKRFyPHhjDOsxC6SPoo8FdWsDIMa/LZwdK49fvFb6flddHj
9y1+aXUHvYGoij1rYGm8mS8r/Ti1Li4h+2YOhQg4Xy6Thfk0bNRX++nBYNEzhG1qZkG7jpOJnkDD
BPvJzpP4yw9S6Sooe0dvbVDxGiKTCY91+b/zIKVT+0fKaRTbf2uJ6UnCw0VWq0LVFmB06QhvcXNH
7kbWPkclLOAB8MIm59AKGCwxQQ4vLwm6RUJSqQmqT9aT63Qzoyn0mpeXGR0tuVBkwE5myvY7coTp
qF/ZLVGjaqVmZQhC3z79ipdNfPyStrm8d7wAd8OJijeodZ36S4Nc9BKDYyPBqKMU5K2qCg7xPg1a
bJGN9EaWwK5okYMCz0KSNs0Kpsz1Iv9CYjW6BplGWMR9vWtNFDcYi5X3cJDraDiNJUchYtmViKJT
I3SrgoMmsHR6QOP0QAWi1Ufby2w2cj2aBJVFkgJpMh07KM/fxL5p7zqZalFpwPBd5mUWwdNVD47L
dJrIvpfkRmv3gDJdh66ndSAdycZyWIt2mKlzQKx/TjdKW0oF0LufQRk0XL8Yd6JUIkalnCaloq75
zNQ2AUBZisscs9QmGwROe/tV1JwFjqzR8Nk1ZujEt30ZaY6c+X7Porb66b/sYmi+JyYir7z8heUq
NU51O76f9GsT2use8tUUdPRSVc15LEywNb4+kaPqwKa62iNAtVP6Y+8/mtNyehpI6AN+wXl+Uox2
dtR3ir8rzz3Xd9ew4ba8m9jTmzngQmH2Eerhg4mNp+ex0L56Fu9aw538YAQQauyUGEuUza1lnUBs
F7s8+kDu1/cqJoWqPO0y3fkvMc3i8kvVNqdvpCxlEsvG0hbIIQ+4/qi2+G1aE9OOVmQ0CRULiLEk
VNMEJEbOyWfXz/RPYnLquWT4Gfl/XSe0CduLrs6ns9twqup54SGGEdVa2fYG6liPX9+kxDA4y7LR
t+dOjl2E596OwjzzsUSyyW3vhk96M5KP7gwzI5yGJXIPp2SeUiWXiYXZKkf+3ozFz+Q6ScufVxbA
tdfM8DTVlmoc08BhfxQu+1XGC2FPI6MQrltpXxaffW5aMQ5AtYFCViIzFq4BLp39qSBwCZktnP/W
BGd4KLVeHfXO9GBh1GPJc50t3mj1Ua0jPeb8blTv6tOjI/jOARloT6a5Y0NzyFjZYJzKVwzcCael
/INy9BpjHT2vTzQN4uCN8u52VZXXWW6LzDJW7DaEQ+iCwvPMvsOVJsSupifalwVA7khJ7U1RSgsR
y75hDZB6do/lNYLpg9IyYDrcJn5KoZN6CJMu/SRVY6jIHCnvvHekAheqmZGlmUPh4+5J2pmOxguz
FxusVV15xzhfbnh6kjWYxsLEkqMJ+zXbwPgBhn4utzji4Hs44weg7+gMzE7rCQqF0xBWyHdXB9i+
3253uQ+7JOHgMhHF7UrRYc9gxx7b67x3mGAkhnkg8nGMeXZqYZ5HdM5m9vEqb3ywGc6JeOuyW/Q+
n1yu2rgi7WTisxzhgSBaI7TQAGsyFtksb5Jo4BgFOIAEj132owMzrYVRkDaDeW46biWMjxUwlfBt
0X+6ZD8oOXmCH4Xi2Z/vjjf36tvMH1/4sghOUVVjeiRTj5Tla1qOvnkGNX9jx9INyUHlzjbmvfV0
anb40NtsWA9Lth4s0LZ6OyxJuz/jpT0QC+fT8ApiKNKtEuO1N4uMVP3ek5xJZ89CHFCpYvpy9ijM
vZh80he7BO5YNrqyXWeGyff/OK2RAxJvgkqmi+NoflTx6xjbUIyk+N7Rp4rNj7/38zH0Y98NrI9b
Lf9wnHML/aEjuJ8f+51Pz4If1WfJRLNfhGK3aTq5dFSRUgZIfqNX6LKacttnsjTCXhT3L7//U3T/
0wLagX0i+rSE5uO3G5pD8GYhKDXu20BoQm1rssTAVIFNHSiesno35pVcvjHs79iwypVUDjcYp9cs
BjXfB50wD6yM4p1IM6DyhsGDcfrvN3BwKSYFt+iCm+D4TwZPsHZ4UK3FzDxwsV3Dkdhg8zCIYoMd
Ex0p6PO1/tsbcXsMJjm/e0hVEj9ZCYiWQ634Mk5dIC4dVPK1d9o4ygVqT1GFZmgMC2kE7Al94mJp
mjZaVmRLyN79LMf5D7aRIuzkraHQo2BmQeyLo8vLMhr6pqOT0JMcDv7SYAtSM58Oh3Ib/vvHc0Fi
uaMOz487LGurTttmcAjFrys7mtV35Sy92htyEGkd087CfSYE5hagNtqUeimWIHNVom7pOwFj+9Jk
AnV3Ru3ShBNs8gRB8IQ8cqgNgFZdHRnSrdZZtIFaKUFhDWCz/7Ky6hlrLXxJD3UMppXN+rbWDxaK
JUd1kfZMZBQSm2N8UJjqGmAuXGFWMO8X6QGg2ue5pJF/ZfCrI97mDx9+UgwxoSD//dDHNDcJ2VNz
UirVqw8a64xZpm0n740RK7iTJH7uRznaWsrN8t2N2NOEvUV7tsQrQGqKOZ/l672OOO9LCco0+WGd
xDOfOMw9JPp6CRxaZ5YXFel0mPJ09MEqBAKTocTtSlInGwHa2NzWYLKou1pR4Y6BnVME2qESsN8G
chrqPoiDiUXIVaWnhZqoQN1zKSoZGLZrQfbphdXBY8mz99D1pxILvTY+g85Si9fnWsPjC149qmQV
pQuKtmW/LS40Ult9QD1H1t/MuNJSyTu0qdb/fEXg5/0XtyP5HKBB/W0xtqH4zgf5zNMnSvIVH/B6
c78YDbIpcSckIecVzt6IPtGnhkoLp+c0SbleJlWBXeGRocJkKn0PfyUJgFUuEEzTHW96yrCUQHDZ
e6zc3JpGg/X1bQHIaIfigbznJVcxHQMr0Gad9zhdvsaT7GXZgPVbJMUeFNsuWp2xGPc1D6Bpo7Pk
RToU1ZVi+ErtCeiDIPxw3K/OvWqSwQvW/l9/PJc3PwA0oClmkTsnGOZDuypHBHetDwwpG5ogBuVW
jGbkgeEHtjx9mrIgV+EkiMVVlSMDCpliN5ybXI4ucoCaTp7H7OdplhJQZm8Uik6J6BPf0QNCQ8LU
hPe0dRqLqmQAPNc0gFx5L25t0bNug7sqn/dlG6PdbObf9UFugH3gBWCwBguMDjP/NKy9E01C7BPV
WHLtV77jTUpPoZyuml5m5G0NCC+/cqluM8gQZhXzEWHGqWJjOe9LZIJj0Al/lOssk9tDRcZRmarW
ViqflLwxGHUpU5vEHzoy3AGAsoLEWOhfUQXIkQid9WzKvIOyy0ubV9cKDYq8FfDLjqpGgdFG5sBc
ZiRWZ/mjaq6UT9AGkneHEWi/B5uVldjGNhQfYL/Z9PhS4OWq8wBvCqrpxeSjwgUSX1HgcK2oEUaa
OeTF2vW44nnx5Rbsri70OOMkjaesGzukXPEczxeyIIh//5ZF9dHLf+gKMnje6cYcd2QfbHSqGhNO
jbJ7mqrahf0utdFzdkNYZBmZid5cbKoKTnmNPZoREQG+nZhYidX7fqtz2gCTCUXm7sc5M5FvWqLw
LhZESlpJMnQ3wgRliVkGdsLHZI0fLThTYSBPV1TtTkxra34VlI/CJ1BDIydXowDW+9e/1Nki2Jsk
OyFCoJvBHtN0rOZEj11HSsuBlWEhy7oRaVzU5NP/FXXAzovvSbSRS1MrKS1WVTsSRGLdOijiAzWP
nPDTQaVSWaFX5dUPuXKmdivZFyQ/nu3OPiFq8H/Are4dwGkn7B6xjyszetKq1gPiPQrHDtvL1sMS
rfEykCzqzeNpYyDflzz0j2LiXlccPTnsXy45S68FX0raP2PB7urpMulEpzI2sSSWR6veiBVdDIkx
0CupyQnhzp1WuM2/GsBkMBwh6k69AzyMi9azuXnfnM7zzOT+3KjUupRmSsJF9msCDkX6xUTGnOP1
Z2F/N0QDNjlqYXNobMqzuIQpa30RlacsvN/9xMW8mRXOtGiDSbigePXMWSuop4/iT1S9+kxLP6Ms
hWEUgtDoeXaQnZEqDdQnoHtPNyj3CfDIsWurufwy/jgM+ZXv/h9GG4eqQxsw6H4Xd5ky38GZdnEl
ww7hvKqDSMTMX/+bDxlecGg9jADz81TqRJgm9Cfs4jz8d+yO4JizUOM+YNLjjYMMW8dou64+tS7w
YfCimKgvhKOBPMyRu6jqfekQ32fy7LNHp/OKNkvKfialN4jVclYrLWhMpVugO5pvsZhN/O80vWAf
tC6KyIxPK97NAeMAoD6zSJwRICr7iwh82/R+baMfiIlF9h+yJQF2Dnbh+Jmg0mWxVy5cLIYOa3lV
1Lldgsu79pLkUDPB7pcp2b5VSQbID69+JLC/EU17uf+1PVC6SbJMKRUZgqkZknPhnSd6/LekqM1R
Rt9MyVU+RaSF7zV78jB5a819IKxrrIfrIfjrtXLU1FozhCUbtmGBOi8CikcPu7QWwk/VFwhkQTfJ
wmjAN6OQNT5fEOkDZ3mfCAhz95LOWy5ejz/fo8W3bITZI/zmdCeu5YEaoQOOtnG5CIo9cmu7pZ8u
neGPTm2D0f9a1om+fwmA2a9X/xw6DnIKe3Tb8L305pm3PApbM2VgdY8ukU0XgqduBpqWsBG0DHpo
DGNy21pcimvcheSYC9XryFEwyifpM3q4jlj6nvJJWsXsv9AnJi/OsSvzn1jKFoqQC9penH9TUiT2
WqbiPfyrz2AshHrgYrbEXkRL4Uh7ghS/bqyVr/uAHvKT3Q31o4Dy50LMi3XYLMgAbZz5RCG0OzIc
0As63McdwZKbTBKa34Zw5zm0WiRFtJyAPTuJp6QdVoZBz/5jOl5IJaPKSEHrp8LbITSS4riL63AV
6HP4l5VWQAW+zRoN1ICLJF+JdQBkQeYuFcwR8W6/HPUaR9iTAz9T6m0ql47LZv49zGt6Kq7jidLV
9bGwIDJeQ8j0TzymjR8eESPKiLrAMIqndw8f7bYdbKb3MMFx4+QjjdD8abQ1M2G2TrwVJfMcU9y1
66nupi91A1PBGlI9+7s7Oh7J/0ovoODNzQO7kYdhtym73dns3zKGVQ7TBOtQFInYq/0buafi+1ew
cM3VWXRYuSIEnuzF1S7UxziE3fNGJPxevKtTnRyeY7oo82VPlFmDviHoe5dOhbBO1vKkqIeAm8Lp
Mx0/o6ukYrwnuX0qQpi/PTmqLaXYpuOd+M0mTw/G+/QkyKaSIunt48xsATupJ0NcQmQShpu4nnJw
o6iRk6XcABgqXlCWDzit0jyuUphuaoNEaUnU7brr5bOsozmY1Wg5hde9mzAogc1jduLyUzKVmnIj
yXd/hJvoJOeRFR4sbilACTXlWovCx6/xEdABlBvF90Je5wLX5J7MfQwq9bFAirWRoob/DReXud6B
VSd1YvR/5+E3ZTbgG4gL4dgEraQejh9ICpSUE0DiWlj1Bsby5allrWvTv1HIM1fQVJlb0eoS/p7R
0x0LAC4FfqD8Lovp26HD2HjBQhUEmfE1t0fc4LUJilZX5vCHdp8Phj4fpwSvRMjr3t4oL/NfF6nC
mcqOn9qrMu0Le3JakBYTi2/IAyxviYucnr9b35tQJw9LMU+dNhRZRng4C0qf9GJscVreKO4I5bN3
c0cNPHk4mZ36+9oYg/hkf8veuKn9Ol/iwt2q4b6gDc4SDvI2ccj/6gMXR1y0lekZIoRfuRCVK3nO
yEkyITeZQOJK16fzFSBaz7rEHVEUzaiCAmu+15FMEgv6kVQ+foNckM1dUTptQmaiayi4OGBUNVGS
C6imBJnzzdd6Vpgn/oG/UmFUa1zJTVnHmnxHUlY6GplHxInfI+Fl4FSsG2vYVXfBSmQI46qVVSSR
YS/25JpPElog3STKGxueaMMvacSvNI7vdzvCxw21fcsEiWO5KSIpw0+OD6bMhuGqjVeqVdWkW7SI
rSKuVUaIHbtbFTAAH6xbzLbhdDRGsk3ZrJgViHt9oopXNy6mJHdjA9fSyEcARsmSNinhrtCMOVB4
cZr2pNk2c+cn6qVmY9tLLp+EzEuWz2OLfeecaqChYK3AxCdpMqZaB5vGv7KV0F3QMNAG4gQjnW/q
Y/f5nkuSOrFK9yEV2yR1ujUIJRrkN4D/U09Z8ASk/NITYIPPivKJWFMvrfggjm6t2pnlxrfPgDo1
oxGlJZnFcYLkyA/Jzn3Kgjrqpz+P/G6hEmy7ZyaWVUk3te1GHxC9hHShgS0b5/yoUSrhQJJiLvyT
OsXUOkF7SRT3gBLEpGIEXsEs/KMSKx7XhkSwT8JfCmBUL6EKoHFdph+Gs1vzk7Kp5J4ovvNjJrgC
6zmH3IE+oltUkYlTe2H9rdzG1Yhga+nlUX3K2ACGNYxL7j3LLGMvA60ga5Q0/oTlFVP4Dfsolroi
cxwhFsTGo0q7m4vaEbUo5LJYjv0zJJZ+W/Rmm547mOjGk0my0Vfq8DUjbeVIWFe8tG2wZj24Z39f
xM0HGfASzM9IZFc6YX728qj+QEtXLbbQv03dysj4l4zo92GTWKTSEUcypGOLGdHfeWhJZ8m8lKnm
4t9lt/4NOPjKuYz8duBcjq7Bb2U/dBjp31dgWQEBRnbyqvjumpbswudR7C1aIBqEUDV20QU55bLL
o9oFsrQufWjrswQjBTjPIu+cyHNzofZAFIspRuyJHWyMVrNejqA5SfRt7JqJNl0AwYWYNeWiQJFk
rahnBVn/7XmbIn4EOouEr6dq6k2bTmA0w50HRHr4QMhBiajN8AifD5WKbsIl465i1D4YEjAdYUh2
wqIyvuXb4xHuWNrR70cZongonDUEE6QgqrM9KXSFL/7Kx+l8LRKOq9nyRCV7BCP8oUGT8h/F3OxW
Xj2KgwJIpO9AMeQn4hawDBu092N9Meqy66GonAHSogZexGYYy5NCv4aAfEc+GX3TiDUXi9VHklI1
cEaRtUP606R99SeJUdz/RmKvnUYCaN7mV9X3G30s1VUw+ojqZQ/6bEY2ZKj56BSjC4UflZqU6FGz
8E8hpXUCV5y2ZyYH0u9TRM4X4DsK7hhopIR+lEgraeGt6mtLqLuL+GRRsaQdAYREiO3sT3sih12U
w4qKX4RnWDvlSBf9Kw1V0hi1Rr8yCBQaVI9JaDMEA8XDhqhJWT7cHWh9BW7JsNxndDUl8KtCdd/j
1LmLsObWihqi5cPIfy/gARvYIrz2kXkViQytyVhFJKEeuZMcVlhhaklBeqRzrpuTgarcTh7bvrZ7
eycKw2DbvzbD8di5asLmJ2sexalHFAFpNAn6/sM2kDw+FngnNnxJq7f2c+WtKM6jeKuujamOh0vO
Ou9JJqPwgZCZt7b++ggP/uhWBGa3xkblbD8oqGeu5+b1wMFVO4Cd3rcnLvLSiQ4pTx5g/w57Gue2
gdoDGmOA2topqqb6BvqCKu3CUPwUbUNlHPjB8EDa+DqqyQSnpoS0xVFpE82cQ4Hn6sSWoF4/EmNx
L5GVb1uN2clrWwDBYNiuEH2oskvL5OuH8B861tnn4umeQn3HRBNsEV9xBSpHBJ85N/n4lk69jb3U
Apsv2fzcFXRDzZpMgygmbH9lSrnEzsAP819IY3bWyIiLPGZ8eANkzCz/gW+BNQHbHpIPPlhkmKjt
Xkq5SmUgZaTKUBj0C71sfuCqCKk30KNEsJVll2otpz3nRO7TF2L3K/8q8qsXcCis7Ig6RRD5KMvg
IAMxRO2uEoNR+arZf1UyB/Xh+6TkXyBlHAC42Rfiv9Ia0iaVsRdUglfqZoyP7JVdBkSeXV8pPQFc
kgwaKXsTtZcEY7IGGApZ5n7/TDa2XOEpmhMlvQVmnOQFe4lK17CKxbyjtqahHPnA0RtCgdJnjvoj
xbei11VVfaNq7Ukiyeu26KBF8uIUoCZkCLB8gWnjN0ei4FAC5MhOjYWQbIApUbj26ppXhGcGJn2q
eBQagwTaaqsZ0hcfr50QD5PaeeDVCQEEvq60O9shEamWPXrFIJpSX1ripn1uqKHhSuKtKygTJtdh
XWBIjX3hOLvhI0eGGEmeC2yPLMBFe1UcRgLi9Es8sewp/vNITbbSCVpSDCpI51uARo/VxFpahvrO
cJNULcOpY+R3BCCxF3fnLSzmH4Zloqy8dLmfcuju2U0C1rNlBM32d8Vx/IMpRgF7uIpDfaE+Eq1g
IAvGwBdTcD2HB7Er4ifDuHXypY+3mCq/QLSTb5Jtyl/082ZKAi/LpdXD79QPoNuHVlqSrtJXY58u
hGZRvhlaJ00IsA+KDZL+Jdv+S8i/VZNX4P87DS83rATcCzCm7jcfWgqiSlbY2Ztqb3TNrzV73O7w
/p7KY6yhhAgHysiNAfA8y4L/v46ts/GMpRJqhzdnBGJb3PCajaH63ia2Zlr/P2J7oHuRFTdxa88q
QGIrGIEQhWi7hzHrT5h6RGYbq8T/kS5H6Dm46oCe6YYnWwAVypsDdWsjwf46Rd9MfYV8O4JNAjOo
+2qwCckr5ikFr6X0E5vW5nyFebFwFtcis/C2HU2P183Kzun6TXoNc2I+mrvAhjtE+w/PM+Osu5kE
D4ZVqFdP+K95ItqN/KYfdOtNngua+9OFnnsM++jK6U9RpM/wbjAjE44X3qpvZBsV+vrASNzY85ut
mJWTZnrv7ef9xM9XKd7otsRkbd/+uY0N9ar+digaePjFUgBNpdnZggvpXeG4UBFe6rlplrapOVNd
dkc8OE+ahQnH0W+vuGOrNvD0Lq2MjZZgoAiiWps3aSkgQ44bQG1hXVmlwoZ5NQbiVbgxu1WBk7mV
CmhUwIvfVBpGYLW+q6awg1/Kgv1RzwitzhisXYATTzIors4D6rrfM6LMV5+bpjlywfpgNrTAYB3m
MF4Hu4hh6pYgZQN6BinSKZrMK3N/Jh1FD2Tin/Kd/dIm9Hq5Sk5X85NivfWrZ1dDs0jnWhLR3cvy
DxDRI2yPe4BbquDXtj3f+U4RyETqsbwG/y1CjX51k5rHcI9auw0KjDxZUunckq6qUjKxS8+QRJC2
SD4wQqYafhXawr4fy4+bBQybgEy/erR3iDzhuRY1dQzz/IcfHpK5zhEHp7vlRxEIxCphM8NdiIy+
MbSjbA49zOpMtMuguNpikqm6SdhEpqXeAx96VpEyulLcuxEB+1P7SjSz+D1LSIm/Lw1gurUJDdGW
U5jjtL3npx7+4pgn3F57VzjOX5WpmJTXYSzTYuQSIN2pBh3MayoySpkaMAjovBMnNS55krf2cGnQ
LebfCPR5w3jbK8ig23XvlCGc+TRvEA8zjsET8o7R/zsI5CUsWfCRvmNJsMoRUaYNbOQbTO0brZkb
LkqW7Z3KSJaMd1N0cYeaxQZ90Dus3wxFtjrR2uR+5Rum7aSbkBg3DOC7dbPk9QRxgp3MGcgXcUSV
s5V43/rHyMf6Tub3seNroGV7vAdX4srsoV75goVdfLWy3l99XJUxJMyo6Up5AdVX+YRPzI/IbHcp
jGQJNA7dx8M+CVqES9py0q9nlwONemQTzHf1dcaNJ5VSBTMHJQEq0sW3lr6sq2tJmJ5aDbZeNl4Y
sUNSnjUfE8/wh5pbcbirDhajcuoghtcNPDWWRMeDLOI72rHwxuOKTgORuGbVMYTP9mdkui2GUY7l
dzIogex5HdTw0kdawpAw5mNMHKZ2OoNsdhbOM38+MuMzrSgBpNbp3ftsPocStritaLkKUp8OSgNA
2vkOzIbEgv2hf0RDsYdftrSk4FZK12glRZgM7XZ7+3QKVr5cADSC9LcuC2PnlqSv5smuj2skLCyb
n4M+jpAONBTF0rtLpRBSiC8Y/FpgtQWuPLnDDUISuksc95HnR6+BDglAwsj5keG4EZg2rslUbxV4
8LFQgiTTzuuOawMjPfE6E/Mh4StV56/Y86MsoXllI8vVGgo4wDOobXYSLZZNqaqRK/dyt8KmvfBs
aZYh2f+O0sKOUVVA274EjiD5XhcCIS1xVgytEV79AvWMJqtueDQFuP0NuDu7Vzx0XlSDZCJrOeop
RMDkyIRbivXJm1R/E2f2yNXz+S9sn5G1ksLcBJSmgJrSrV+BH5sMx9W8LANKRi46Ab1PcLROCGRx
tc2AQI8EWNBgO1YoH5XFWdsXi4gIjCV0NNpkhCqsmUsjl1odjfbHKMmLSWsYp4dodUG0aNa4l+or
aBTjGRVmsGcOv8xNWPsfch/cQ2xXB5uK7SRc302AnjzUDbv3T2dmdnOTqwFejvgrVWa183Z8JKfy
24R7MQYN0Vpq+tZIx/1PZNpaQ9aquvYpEU1I7l2x1WAK1qFo+S2LeYcw3IPIgdFqerb6btZjGVtp
DJZbxyJ0vR8IiN/U9SzYyIIZPbcIOnX//kHtQOsQXR3WfJprfYGAqNwF0R/Q0sKoHz6uzEtaeqzA
tFoJR5NO/rwt3LYGwJtM+dSs17FEZE4wHNod0cs6uNtty/FTuCJS0ZXMQkoM6+XEEl4SbPiD5VBr
mt+u/ykSZw+3JTdlhDh1xXEreZw2GwDb+vQ4DAfk5oFHSalEH8mfdTWwIvXhfM6ECbZepyjW00nS
VLSr6bTltzRYGvhnXVMwJ9hJP2qrrrYGJnkwBLY7noE/23jrk33NL5gBBhKDh0DaO5xXhfO8VG/b
+JTACyyGdOSl3+cS0woPiarbYXRIRFgJiNQKOErDezHiEubVjZf8w0MHTgDttWzXamjnggBqCJ77
6xM91VsxJdBwJTRrdRx0jROctH/nmc49Ri3uDMVYE3RrjLKqT/Yk/7pCXpaN1+vYKwyTurMoe9vj
Fda9ZTaOJK2mCc7v0V+MzQdxl2quNuT2vzs0VdtHxix7z5/gTB9fld54txH1UTEPhuMnNo5b4iRN
V1fcRet0o4CiVPAJ7MMkAfvou28PN2OygKc0ktPspsefSJfkd9zjdDxfoiJQRdeyF1X1YvQvplQi
76iN5x4wJ700yx+q8c2XELYzqGrIu8AlgjSNtyB85rhZ1diU62gPKSqNr6mNHrupo+dBwRDz6V5d
KFQpKjSGQFyysEwLxotjdJgC344F6szae6C0ffC5gWVAUMdny8++ayPNbpLGcrjvTuiZfUHNils/
c2lhj1nvV8iO4RZkKrdzYuoNqrWlUTvf1kJm3sNl8LNSe2VLZp9QoZpuyUugKT0IK1eNP4ukNv3m
H++GRMYI0nf8FQzWbEKhD4Qm0L7tmBmmeI+vjlI2CZwb6wk6yyn1QZvxZGB36KTKt+EbxQJkyzj+
Hsb8IcoIFR0nuaLF3dae6mfpR1n0NgEEDREjsrFzHmPPJE5Y0czlk4ZZGn6/OjW+HGy/SYX7PMgf
CJkXir1djsGAEaX/uG0+TNonGtkSK2FKCb//TzjylB3KiWYIlo37K/an4E5YWrIGHzXv9lNFZoPZ
8rtDDoA7/FjBlfGnpHXaH8n8XOdaHlJOrMzd6JxV+dCEucT5tQKoludXfeHvEGzocIsH8P9x8Tro
PrETeVB+GwnJQjwXdbItyLmvH0At3Z+AUCbvj/coxLoURNtRleQHVvtYlNCFfDo0GWr3yBy9BGap
o5wOhEa+eOXJ2x73cW8iYhw4Zmtb237TZK+wij50w4p3qI0BRfh/Cx7yWkKOLD1VpdXF33lcQDTT
8WLfy5BwAjJb0Ni3gyCx4RzeBos3POhE6KncvHeiLs5j2kph9Fmv2wKhN3425BhfR0/ympQugOOv
z7l9woifn+8q06KAtpqyz8AlOF3jrqWJSX85DWko/EOWscm31gtIuOzZjOT+F5WcRV56EPgIMyeN
rCe1MK5puhEgMrxUEg/ad8K84kmavu8tcDEeGhN9IVOAcEefQR6TGqFVmfWUxDKOWw0su4r7Berr
i3vypBu4u9sKaPzjC7gqjqqJihk1yuglRmDOZiHs3MMkX8v/pXgLK/Yc/jPKUdLJSGIbUeD5Aj4u
bhYvMnH5vB7t2BLwxxmZWLMVE5+B2dlwFvtrdp5tFZ8xEROIPa2Y+iTe6U31CEL0EA5NuBRZSibw
u4ii5e0+XUeVF2T8gy1xugmmCOhypcMxnfHmD/4TZ2Q9lv4+yaxMT1CvzUuBuhct3+sGytZEItU1
u4ipv+4y6Z0x+cLcA2vv6w8IEVJsJXqN/sdnI4aoTqvomaaNpNz4bblHgapTYvTUFAzm+O5isrw6
Ij/FjLt7smDpT4ULc4yLKZJRlEvZRTf1t20/gowgxiLUEDEBDu5m5P1iqoHZKnkMhFJXdwWz9gUT
jreFhx6qoGkE12gK3+bMirY7sXl7O2rgi+QRhX16Af7J0yCySLS+wESTl1u9MZnmtd9RC4ACfioc
2kIw5HzNzmxa9lykAruZMYybpxznPmkSw/2pyVreON0NYvSqbtpJji1zRe9Hdqu1hGt5J5gLRUoa
B2Olhwx/jP5X4eXmapr7/+1Wbfl4/lOz2WphGA3Qp/tVStGV5afFC99dLtSU4QJfLIHLEOKJkwg2
nJeq1hk90vYsPQSXGDPn/bpaf1gQYkQcrgcf0whYbBQWJZS/C0UKvWIVzxzJjRLd/lnVu2gO6zvh
rSCQQm0ieOLc1NphLtao6rEpc5kMW5Gk6F0D2is/wbGkCqbAci+Szz2Caqu5SRi/Ff5pOifF97El
SLDl0YzlVlkmjtOfrHuhscDO6olwNPtYzi5rXpD3LSM4ykfxqdz0NPFeUMsnkkU+CJpXnv09Sf8w
gk1f2yijusw4mTyNIr7wiBzj7EUCuTTtnZNHJc4r8voo3forGc/XczD+qnUiW/v05dAMhwcxh1vn
2WOutkdr7dtCY8A2NLh+Nsw4gmKyVOQaNRGPedUbFTGAhRv4qafmMQy4fWdXBphH+knhlQ5/Dn2B
EgW+DSjh4bpMuLH5cocQBb33UgL/L32Gfu6zJ+MGxixO2K98rRnrhHQIqwRk8w53nhharFx9iyDD
xs0+rvulfJTETN8h9MAiF6cYO0IOmPTFGSaJOhZGFiCQ6MpIC9FhVMWsGtqk2DJOFQlZYNDsozFy
DFkVsmQbKKMet8euL1n06yy95boAHnb6jtJSitbPhmI3TMufI7FW0xidYf0UcD9om+uVtzrRqK9z
6BzWKkdI96B5+/CocW9agz4BVj72BdAxg127m/BVFET0qJ9zkIunEn4GYrqmhhciF6hyf/jlADk+
D8NMhcQZ+Q7NRO2b2JWsmn2HeXhNgjPJuuFRdrrLYvAFQSBmCC+/HglHAc4l3FFRKplr34qXWOLW
ya3bhCgY7JmSyoKPbKEgOpEYg/KGnlaXCVXH8Q4HZ1upl6pAvtuP56FQtJPLMwTtg8L+fzqHkdmV
V/mqfk1i4GkhtvIrxfpIYD3b9b4eqZf0FALMw1TkaddRsCg6C2Lb85HRTKYtLX90aNpVZOYf5651
54nCDldw7jE9tIaGHELVddaMc9dpfZP9oAnpZM/wk1t/SEjB8Kwys1bb2RIfQC875Ygk/afSpNyI
YX2xED+v0L6fvRathandf0xjlq3wxrCjeTiFUZB3MHlN8NaeCj7i/O2K+ZZVKA85nMVkcVvm5mXg
ymbqsqTb2A6S7pNo8H2p66fxEsTwC78rysf5tah+2LIfFExbSOI8/cC5zCDunZtPKGqTqukXkZ0M
LSZQW+u6K3PMEV1E7KfmH0HY8pUF+bTYa6DtezO8Dx0I9iQkX6izH13lR8GQsfaLflv5XKXokfMr
5N+lNA3w9uHBHt3Vistqy7/6FW1nyErqlH5NyvLWxumO0mEjGr/KdIiIIeS69TYuOT3lUerX8aIS
zBoSoIwvrYSmQJLlOASBqeP76ZqMZDcqjMpqvIwyMikkc5rfxwq6d0Xc+4C5MuoktTWoAPNHmuhq
oCI1DH15fIbzRA+c0htImOC5e9hKjepIpNaSez9mpSw01Vh0VA5oPOUYZPlm8MOt9SGDMekOc+WL
w+W9eOdYsFur/HOmYzJYxzDr4EjpyUYSQLmIxNjz6e3V9awF80pSRsD2R9mKosO3oemw4rFe7DSu
iCKreWRkvo8xjnJHhCQi4htuFWAYT/ACWaKURvHXZBsRWqG28wizm0z4Fl5eRWOSK2Q52BLKqW5x
71FMkot7jI5k75IvKOV8fA9JrS9/zjsiL7nNAXvZVZNCBawFBSbUlhGyGsBOykhBCjMUjynmaDie
ajaAbRlRp58M7wmOggB8K0rSc6lVug1gespHmMq/BxYtScqTDl+ya/LKpZ+CjiFhVOzhtDlLQ6RD
UEQxQCqyzz+vnwvXyReONVtN0kTxzA6eiz1VFxEGvdL49tuI5T0IYBKUdZIKDa4lhQJDn/xj9Efm
eQ38Gp0g9cYnQZNeDlTf4sq/x89Vv2yBTewyS6yiH2fMKMxsnB8IO3xWIJqi6XM8QHtaUJ3igz5l
dfldMs2UWjcKHTv9Iolo6ZGfAsXL5GQb84sN/9QCmLV3fvaz55OfVbpBAfLLdaFeoUaJViUbAGoh
JouPgqtC8fmJ7pGp+jB025l0Ci+vwVtR6Gkc6jGXYgH2pL/l90V4TA8Bg0KMaxQy4h5LnnKswidE
k8KN2UuaB1k5fkwHWfN7Yyd8XO5IlszX40ZORYxaOLMCfwOJJj2TMraVSTLO+zcMIsF97hLegjKw
GD610NXU4D6GA135Z5FosGi9HAaxepSVhSqC9gYFn/rVHvUFcsx/HXfi3brRty5aafRXR+AJYue5
0JtX2AsMr7YqSvqNBL8vBnOpbO0RET/inezqWJiTjcJJ+gezS1bvNuFKzuAVzD7ZPBXjgQsHCLFf
heRf7tj8gLgiaF8v6cvQsmWV/sJuTYHSpxXFKPZ/olFwik4olItvHJ99dmovy1+/odWzFV6/lN6x
BsUyPXQkobT/n0HpaW7eK8QMrCGTSodIgQpzkVED850eDLCwLnvKpCP4cEgPkAVwRp9YoXnKrvP7
IPk2Wxqsw8W/GvjuKmbmpfsrBsCjC8iXxEB1pGP84EBOPNYzACzuonsNf1YCDRCpv7eu4wJHO0kf
WmqmfYYN39oRlu5puyxISDuHC7k8/spW7WBJ4OcfcaPVOTTJsucksD11HZLElMqXX0uF2kcYsdGE
q6okMtyncxGAztR5jhq+wo71LST5An5hY4/xRcfLm2CF8FGbOXJ2wLttsT01kuTiElz4BHLByHcc
zVar5oAcL7hdJSkHti6At574QcXTpXjUwxy51L+j9hBHMIroHr1mvWgmM/kbxDqB1ipJTa//bEoI
NNq7RtReC4bzzB/H3IRRH0+7PJsN4XmG7e2dIMmvQ1+7RtwtkcpAYIL9XATEfp5mJQkaVR/Y+bO0
GJzVNXjuNLOyK0NkpemxieYpQ3lL2sUvhPqQ1d9681wDOSlvgaKtIdVuAdUoFkhWjQx1p5eGcwIv
0Zsb0m7pCzWPsxIE/yWUOuzWgbtuYVPVF2hXZhrC9rPedVC5fIvl/+qQrlOv5i7Fk31mm52tBeem
1efo2uVsKZv9jbHTzFHqGXXZWx3PutzBcSVyWu32+97twDhS1ZsaqKcHvHopAcYniZ/2oUY2Cddf
/bmZ3nmFHvvVy9h5j0aF+uHkSgWh/GDgEzPzFeXNNcegjr4NGN12arkWTTa2RFHP9YlgAkJ/7/dv
QuN+ToE1uPdb9BSfYZda2qLzbbqrZOnin9i9xy8d54av/VoQTIpdFjlgnwHpYSgH+JeLQ7545HpI
YLTqXMuNqHns9e7afw1nDr1xATk94AxhzE7OYVO79Wthpk6ocYl/FvjR9Zr0T4kL59ogrKTrH6z2
MnBO5mGpD8tu5S0jfn7BbImm18F4pjhOrachfrL9uJz4IkAHZCP6li8EupwpmRFUUq82/zH9QvM2
vMC89KWZf596yvF5S/Fhp9JUaz4zVX9J5t8NKjYOtIpeOpqzdvqDdzytBOzowHx9p+qp7jZmzQge
2YGUsC3opE6373Qk7d9aqCPHSLI+oTLFu1l5n4XF/cR8Nd32LJOhOLenpR3OvkHpWYtxWtYaUESl
mBx0ZZ9+enG/aBLqGscT2LxjRyT1E5Sc92cjfKlltMOOB426abFTO2vAhQzNy5r6pHUCYeWjExpd
sTPSUdJs6h9o96NZX4sE37kXNO1BD+kHOaWQmL1y90BxrWqxlrm3sgvnpxJXVlHenUNlSP7FD2T/
wPPlXiSq69r0V/LiBoJEpRz70GMEXDk/ua7tak+hbbb3iDSC8TroBc6Ga1CHNn3qfxwfCrAgQxJY
AUNY53x/6iiXMiptyQcwUvVVZ2QHKG+1/hIu+ePtpcju3a1GdhlAA0T04Tcw/KzROvO+2xY2musF
MhbQDUA7m9iFL6eFA7IA8MrAeXWpOgpu95fG+5UWIPxhJxkIJDpHtm5AAVNdhMsWrebI6jmiFX+0
OFRGHUAVUBbieEiPd7L8OjJx70QnwjgPxGx3CCWYCSx6nzjjQNjqLNm1Wz7rMjnxpv5LivRXa+qS
WcPjyrnAJwoBEb2fRGg87Ni4Jnlhyaw5vnj3vxiSxSd6+VvHC6RpmaoC/MuGqARuGxduuxlATwJs
KhFAjdlKvErsYMkBfMJYMxDPLBGDvrdNCmIQamcxQ8TynjmDsNjG77bSng5CA9OIQ6k6/Q+d8DPQ
egJl688Uh4PS4Pdu2zGXvG1y2D3hXzJnPWQctxq29ODkZ+3G6oiX8l0/4UEQovyKrg/fE6B2iV/f
VFQaoQCOcS/1Za2UYd7x4dMUFJrEyfL8h5AExbHSTZJhY5GNgfXdb/j15t7eO2tB3GFfKS6n5Z5w
pTYqEU8KEcx57B2eSCViK68tYNd5GjKuEC3yccctn5LJyjdcgZv8ZsFNRWpOtZoC1pFKFX5z8Q9J
ueNaBxGZ6I1Nj4r1IYbVikEBm9dtSSDxnV8PcpyX3wvAPHDKfpcVGdla11xD9ajOg3gCX/S+cKjz
2UniRoIw72irtOhy90+JtQOmDaGrd+7yBFG4UDu4M+BKIcnk22mvpJmTkpyZhfdHD6p6OzPThG9n
5cD+riSNi2TE43s0W5Gdg0ZRMlGOFee0gW2Ax1NKmYbQ7pmPNPF/ulJAU0RkVVS6iWnIK5Z2bHnV
yVy0hyk6/ferT0GZ5QSlvpx89DpAD5+aXavBIT/LKvY+/GvK5gcg36Q6PtzTIojLHA0fE2BWGpuq
7BMemzi4iFjP0IJyO0A6JP3HYvlmjbqz/tY7pIV9Db+w4worMSU2TYnw2LH747A1w9eKdmc+j0J5
tJxyBPq3uXVvTa0+xpIYLMW9UZTW8moqmRkpk245zbSWZ4jFbNUcjD/vN86QDtNTlkkPybK454gL
VV+QpFVYVmgNDCwx5mIPho/Dy0mY49SJu95WGXhJfDHGkATmFDpHAqLbrsBiYoyIs3YdfsufbIuy
hB3zi9fKhl6rrw85q/rWoAqi++usmgzia7vp5CAvg4jpjRlpRcjlKC9QWpWMDYRouDF4Uv9gwkM6
MZvYzwzajQuCM5YtxYi5YFYBlQEKdcVCAGeksqbYzAWKtpqrzRjkQIskkfXi4opWcWg3M1sotKUQ
3ZFkZfyMHlBCXmqu1cBgPibBeMZ6fODtiJ+PymErUkSNgAB3oTZxfDkU6J7piyJ9sqNzawDCgLmI
1Kc5CzfenjZcS6oQWZeOkpeTyAfKosvZdxLd5O+EG7tdxU0wV6PrjTJvnU8KvJtVsYuDH4aLAh21
RGp5Hut0KXiL9CsHlU5YpDbgMmkaH5oUdJgvEzwz1tSyr40/Kr+pzTOe7YHQZuxPp1JwfNoD4oht
0dStBbw0Rv4TqFv2UmNnNmPqrxIyNM3ShAt854IMRFaFNampXQV2v+kVwLameM/Cq+fc8Mp3J/eM
2XFk25MGQTbQ0ydhqkLhvE5GyqLTu6KJ7bx9v3sB8LEtoPMOUO1BPYKSEWt7tZlejoKauURAzmhV
KfjwB6m2ZedEkMmDbdDfdE74lQYlJFSyI7/DdijpJ/cIMGqA6Mfby4tzWznOZwCFWYD5pPabvdZz
O+nTK6V1UYOxHNKnZ8aUQQlf6AkDgjLPvHa9Ke8Jf+DAMmZ0dvezYWdOdkhOEbKevU1WHr1hs5/z
uehtWmz47vhbwD9Zjp3XIMxHVjGL3qhZQewgax6wgkHDK0veLlD0JHfdzZSR7A5oCkOxd/7Lyazm
Yeg2vCEcnXpXmrRGV2MkEU0PsLTAaYAQ0zBHWH7UpGd93qIEHOvGf2S3g/3PlYuzX0H29HK8A703
Z+/hRqoewgfV+15d4+gFIOor/InuJtJioR/yyFmbTQgVqqppCu0VRDYAhGBYfGovXqBYB+qA0Byo
Njf4L9FXBKRrASAeH9Z1rUann17mt16AMB0ie6Khc2I7OGUfR1hbLUengUl8yO6paqzvUScrKOUW
CCS46NcShcvX3VUOUuukvG5pV9EvOeJshElFURtYsXe0zzkeSMhF0+8spnpNVRGu7SQLgUDKscO/
NRaAW+J9fv9Rlz3x8JKpZAhMMmmBw5Jy9+1IvFU3WBUN78PPbGKfimvWG25S/EGcY4F2h4g76qeG
pQ4TL7/eP7qR1o0ENTlp+YaKNSDlhqUk+gkxJpYOjUerK5Iyt0hJRN1rlGLrEcaRsFGVWyKciM+x
NsJBMzTwYdQaqGr6Lk85oRKFq5M6aMauM+B1bixou6NWNIZooCfBzdSNUNIRn1A+xujln0rMQg1D
oK3jMJFo2lHwAb21S69vDSDs3+yAh9Ykf94HsWiBKls0reVs579SvuOW/WFpkIcRHAHLWUORId1S
Cnml20A85jEffBPFBxPTktJyRyN3SXKIRwmwRsi6EoIGPZuyS+RpZpUDV65CASWsMnqxd7KnZQb8
dNwa6FdjWeTcrUVYyxcihNrxPaTj+QOcu8hdbc7AfOWz8Y5lK8YP4+hxhjf8F1dfp9vPOevH75tM
RSqZtwwFUSgpD7aoi5P3kE5I9Oqg9AGJJm3U0RAqOiQx9CqySl8aJR6VhuM6I6Hmk69bt54k3FVC
gEW0fVdx2lFL/fkDZsQ838sIjlnSqnPMSPsv1owqG+JwDGNnZHTENJOM7phOgkjfY4cyPPTdnKrv
kn4pfldq1nryryjoU4bd+xZbpntaDQpmRpn3kP6NLK8+/2w+0I5pGxBScLISG7DCQHsmcA0vlYtJ
+3DUhbYMJBbPfrzvLj3BBdn4w3+FhRJCsovnQpoPf0jlm7zc5loapB5PzfiADxBjY5j02HuA6AlO
pMfbdD9XwfB4qSm4JK76mJ9Bc7D7qmUCgqKjM5iITcMiQrkt3hJhIIfecTuqNRpYIVqNwQCBzjj3
tHObiwDtOCOFQ6/FKAmQWWURZlnfr6eFcolEsMUuC6I+VpjymhJGHk+kKQ02UDXsVqoHyzZqK1wv
ojPOgcFvGaT177ucA1m4DvaqJs5wyxvAL+AjsAMQNrNw20tjxuSg0b3TnPlCphYEO2H/tGQD9N17
g70eS3z1Q6n+V0E9LQVFxW8VCf1cvtxOqET1/vpu2HvR/d4m9X1uaa9RQybh4ZHjBZNnABGX/ypa
v4uJNgx7oNDh8nAtMeRtxT5+6pLqclYlHF5s661M2vx9UexiDfTg/xbh24ToSy1ycmTx+Ns4eDFt
Hzu7Jqo3HhsmSi4ek2xzk8Eszb1mzizjLnD8mplkuilungv0EFf+Ju9SduX5ob+h7O65yri78pcG
C7bSuKDGAe9xQ1aHAVaFkdrNyWq0l4sFGNd+VHdI5ZG99arGvanQ9oGT2onGllYwsoEjD2ZNTYij
1eUUW1yHX5+JTj9fg6LzoQ0hETiTNArsknd6N04HbN8YMzUCf2KKlQzwIRMKB44gd4cPN5tJ7NiB
3PwNuj9fPKf/wlX5Onthtr9aWQTGaPjQrfduCbvnlYbHFnu3W8iZLy9nFDOaW5KByx935Z/jEwGs
AHnPMJMoQGDVtBAsc+BWerME4Z0VEd2O9acbLA8hSqnfdV3gcPNGn3zKF1CVDcKi4obRmtxZqIGz
PscZFjJ3CkP9sgEAEaUegWgruE9FjuecwoU1OaynF+frqOzig/GgMtN0MWvP/dU4mDwEo+hjxSB1
VQNs92wje6WIiZlTdKmoQh5cOrz75QwhYStjZyrNjJ8Aeh1l5A8cV4Mcm6EsVlklZhrSM6h5QRA5
aqMBwILbetBGwTpsTNMo+A4ywcgnDZvHBGIbgwIlwq/lOpj889dSWCLFqSrXxOMStYoBUORs06us
hHvgaEt9TF/Po1sH0A+f2yxISaIfmywHpeJjS3p0/nKmYXH6KQOIkx96433JIm8pP3qsYGhe2aaa
Sh9+/14sB3zkv0cJeRNKDf8MqM/w2gj99yYyOT89BXw/gAMboNNHVXvCmoilJCizP/cQrIF8ZCAZ
r8ZAEWyjfdUF4jzgAn1W8hPt6hGdZ896X4azUxwyF9iLqFwX5Fp9BHzLt5/m92DRNEVsVHCvVcuf
9yTsBIC7eOVwnChYgOWaiT66Vx0MpSOBM/1722QDVl+K9MTzHoO5SnMeEw88k0CjnN7tn32x5d6G
x2ori/9X+nojeEMGhV8GYNkczRGob3jAtFbRIf9aMT09KSSFHmnWrMSYwCBG+2s6bKdaIEVDmYOl
usnR7oCl7H2joMgEzIz6FP1z4F8lHP4P8iAoI1S7h54puVN41zb45mNwc+clXwZTACCA9vxDoJRx
s5+ls1JvyhyifSxWPLZ9lBuy7I5xt6d0jYyRhkpL2IVZikdqR86zTYE2JlcoknYGxq1+h79MqvDu
NOniAfV1hAHpV/PdA8xFpNAFxiyVHgzdDdVcqbMKmZRCp4jxl3T5q1mkR6uYoHxvXpkKobyb7g21
9QYFB/a0NpMZxgDIWrYU4/Io93kZ60kNr809qwaNtF2lM829/EjEubvmbR0IkeRjMrvSu+excfpg
/fHmSocVNzfgj6Dhx4gzxuIZ4q2xZcEIUUi+miwPTbx4rnQPScZ+lMf6YrkxZ6BmRBGtPfXEyIjh
lvXkk8LUMSnaEy5QFkalc4OxGJDE6yFBODjCLMgoP1AxFYCGMrSJApq4lbDwMnph5ItdHVp6ZRy2
hch7kK/nT1xQPl9PDQP2o9cvkAPpFIkIqMNknjuXeai+eODfVBRk42PvvYJNqfj3mRjAc8bQY/6T
vPgn0LY39/OCzrn5MNr9fOSghRbEQ0x1pvJY8A/6HlThCLSx1YrAa4Owez1f++rg+DOB7fCnSAaK
y0U22A3WWCmTViH6ntQjk5DVDbeQgV9/pJ+WYVaInCuMOs01UsbOujrHhT52NWS3F6vnNkpt4Ynf
EFrgmp8TbQ+GyoW5vdvekS9RlvO/zSZN5kCVQmmsLAJKVL6zzavYGr8ECni68ITKVic0d7ie2wfU
uhZccecJVU99ZwvPNDbLizUtAowhz0oMErIwpzndtlwW9H+BkV8EMEtlX4Z+5Rks+dkTK0h3BNHc
OlUVV51+Cz1PCF5lWjjPti9vz6nit00x/kt3XTnB4dvBrI3e9S+XVr+nYpCKbDkg9QhZhVRAMjfx
4d7JsS8CP7hOFaUQIYlFZoDBTQMNDxhfHZfMp63NdqbqJzGDRvI1HZc54nffWDzoWKbE2hY74YXE
7MfUSjVZkz2tOth2DQTinxsldXYxJcx4vgXWQo82HDa6U/HA8QqzXUNNJMoYBLW2O8j3QS1nkI5Y
wPZTIyT+DGkkcLn7PUR9xkEBIKyCW73411frnVEcvaB1zJYpx99a0HUrzYCNHk2eVEWN3xEnCJ4k
wGhs3meHEVExVVSczQzu4sLRyBrq2UTpA+VtliUBELpJ1zH06AHs2abU/KtOdREC7qIomazfqx+Z
U7bPpYLFl7HSMuk33JObXVw0j3tD7VltIFmHV8eJjr5E+GidWpoyKp2AE4u6SvJ/mAJ/hfcDLpBB
UlzcR0dOWe5qss0P9ZNLe9k86d2qkCuk4stzyPRtgAR/6TLihMGKTvAk4BJEay0vPjwPVkVi70my
OLHB0nvyczgeLBVQ5TJAHnVGJd9nb2l+sjogOVuenGHJVEgHM7IgOhBvxS4Obs/k1/tW2p/xBYim
qAH/RVsd1jg2BSH8SJtWp2zspsgmGdEQL1KmQIIvPTOUHGoDFFC4sTgX1SR/ud0mwXOEXTVuhGAr
9pnoifE2ZcAFNpHsHi6UvYupE6EEH1d0V6kAkJ5tAoseL08rIkO9YUjiJBNnFdSIWRuoQUTaklG5
Fu0c+80A8FIC68lX0vwU82NdlREE5pK+Ecbg/a+fKraBqRygyOWWWRtyvYwbxZHEK2AzemnroZBV
tjbX8HMP8j+TzqFsqImwEL84nUwVHEqrtuvfU9uwl2mKhlQCQkcTUUfN2H3FqdRo/75//BpmwX/f
SnT5yOKp6yTwvlrGQdpTaHYsWfRMI05a6z0t9tMxCzJ7Y1YYLEtESbkR/TzHDyQjbLgUBP/c828q
SgduS9nv/xTOhy1rL1dRVweGVJnJR7lapFh64sp/uZ52hT0A4iloHXMYcmQpue5dU4QquLCv5UXK
tdJNSm/1xm0Q8vyXfYQZZgqPvDf0mpeGNLc1lnvnl6PPwbLSEaHeqza4KnQIlU7NcFlXSPj1NvtU
Gd0xetjtySXaP6+xSc2IsT1zH2xYeBkenB04rqaGyGlPEbCoB+LQjFffnW3V16Hg7D0+PbyfT+Wk
5+qinNxjVa5sipEDuz4OHLDiyUa/nh1miiWuXcBXgZeiYOkK5Rel1wEXinJW4Y2O3EJOMlVVt7Y0
qd9eaZqhLPjzWI7a/368iI7ytldl8dowgFPEvC/psjZP/mjRD2YZ4LA4c+LqnmnR1QQnaeMUPR5E
Av/GJjPF4/0kzi5ALWRBcty0gm6eleK6OmzMx4IOOaU+/KTmwJEk5ONni87BuXi9lRfsrxeJlqKY
K3wkgrvI9a9SSvPuvhaI0CLLFQy71EHzOLtxKBU+wBxA9dA7dGvylsa8lmpa4GXq1TDMN/BpDFDo
OV0xI10gf/HQpYf3hu9GnFy/yMo59HseUVKxnTM9+MtNrZ/TXhHxb01CZs4SDpaTVI3mOuu7EdtI
5tH2XetnIA/NWoWxkqwMLQzV/7igecJ/NWI9G1SSYRudgLtZBqtnhk9lZW5ZCsEdd9aWWUTBB31L
/C12F2bhUMSS81c0BjPpk35jte80PR0XaswpaoeSrNnmKZLZ6fuYrHcMH1tfNIse6DtUvxNJ6xja
E5UBzKgU4svR1gqRX4AmQ+GtxNQlzgDw9S+cDYqEx3G8qPt3DIqz5/t//r2Dv0VIbGoMi+Qd1K17
3d4xoWhvD/Q3kLlNCVaEf3gs58chtjIbiS+ciFFj/o0AxM0w57SMyMlVuLxqcXJy7vLMzolX5Ufl
5m6w7BHi29vn5WJHB8igCjPWOYSA+eGHF126xYbgDtl3mu5VXMuhlY8jcMamPhhKEHObuDgYL6el
RO5YbCPmAQQKjbQIdEOKflkEkKQB4nJfeOmktT/oys7u0txjXjbxX9SENEflygXNflff5+BWZqkF
Z3GbmwYFftimVTkwkG/9GRDJZ4BZAjU9LGYw4iei7PfL9St/IBLiPJRaz12DePVNVf/ofePnckbZ
m5FI9eUq+NxgtH7DJgMU8BkrvlVDMP2VSZY9N55RLJWNqNXwWDn1l+wVhtjMu4477u9T+EE0evMl
ESKXvunb23r4B1Zo1v6HhbZLvQeDEHxe7lEWnWU+6DIR2Rpy9jGMjpeJKHdjTPkXenngLSPFjXLB
ZOrbpNfAaygfD6OAzAO4vwErSacSYIFbikmKH9Gx1ItnWg7lzNYD4Pn8z82Z9iLiK/z6LVcoQo8E
Ew50xYs8DAuR/25+K9yFpWMChA5TuL8c9MhQjopzm3jtXpMc0Jb2UJDLn5qGDbPZpdJjmbdXBkKY
2reg1/DMPOw5bH4El5OpV/WxZXlKDvoGQUu/hbgUNIn5plVLGJHlGJBJmqO+OAUVf+6Ucc4DmsY+
U9sNd0wYCodR1PNsG2YAcaHz36dTkoBJhrxlScigA+wEmfnTdssYTwF+ljnRjBG0NvWk0UDt2+u2
oLyCksckWqZ3z80hU3cttRSS/c5qZ6BnCVBxait+B+Wn8/S81vE+eOS2iEQFt3AVvE8HW9Zxmh6R
M2nnYn3hyp32vuO46qG/MSuuKElFvIg/u3/2rNUkpulXdOpmXlfvwYGIkIv4uz0EtsrIEqIrhdEx
NLK8vTaoAijqZt1M3R5oFtvXmPXx2ffSi/5AO0jic3YDixndqP+Un4RGLr0Q+QNQpaI4g+DJvRAU
SnQk9eB7thqtk0Yirp/RerwkZ41st7vFTOYStbmJ8Zq51oqHg7zfh8rfARHw7IYZ1w0nl6JmVlxK
UihngWHIDTbfpst0RyaBA7t6dBOp6PVp+IItREtIimxJbkY/Pc4FPwcVwxU86IrZ6DFTApuIUBBD
SpxYrZy67OGk+k69IlPaF7OympLKs1c5g95j+YlsbybW+snhtZZpnkovgp2bMie1xKJSPoV47xTf
3FlcJL1dVKKYqD8J6e4zhzlAFm1DKaJS2oTgctlE3W2v+NKgEfqUIL5k3TIAgtanwrufxnUnfUQC
nzVuu3oKlT8ugxGkQsilaW5NA0qEYz7U0++Vc3HFgkJARPBBqBSSyjzh0w0t3zk+xqyWNwR5GN20
SstQX9NIGnhJxikrHbEhlWsNH76r9YLxugmVGCsrssHlfuUOXRBEaECStRw5FBelxFh3IvQ+d6PD
gL4uTrE0xxBAKvge1Z10ZrWzmvJMCBoeAY7m/1f/7JZhfhC+CizjnR+srjm6yuNQFo5qzGz49kph
WBnE8QIwyqZs3lzvrxXKPHP1wRVWxtAU8Awyyf5H9SlR8WCxu7senac7oDU6K4vTFukg4TX43J38
L5ITiQKr5aEGVP5fVLsrwU9kNZHiUr3Jeu0Yc1//LfJ/znqjrouNfIraFK7hG5cYqHuOVmY/vQLe
rkQ426WeTtH6VPcW65FW/FgJ8OdlspGGbVflscF2Le+I8WvWal5px2m8coQHphMKWINBbAMCgUL9
ZxCVLunt+nmQzW4uxsREvMztXIF0CaTUHi//ctO/A9jkcUPd0/XsAib9t872XeV419E3d5/aAXIQ
AITmtbRmF9AsRNaJsq+VGWjdPm3tZXrA5D0QpxXqAU9HNxv+5LsyKdYsB9EVzLS3rmHUsJ+V3yJd
dlPC1SeRVpVtBWFFsKnp2+H7U/8aoIbu6cR6B6iABCqtCvKXPE7S21aFZkhIvTnVgQ4cCKuQDpcU
Oj13aUq7coSqGEhnGloIdFHoLEUcIHSGIvVFszqPn4Eg2e0Bg/YobQRclOXFm471jlT07bFWGBFB
2VLtRYbCFqgFoYccn9+snY4fkmukgWHBPdQoR1rKwCxicwKKHaGM8vNF6kAMKvVd4/sSQH6Krpix
cBZPJOVzFqJEAhEYnwUipJ/LFFjuLqRyJ8UpACmnaFhNFZYd0RkcU0AhgUDCSMyy8g+spsVcEL2r
4MFdp7xJifl3dcNSHkzzrjudQeDPOAWV1Hhhgt8OsJGwdmckUwRcpiPJzVPFNpmIpX7o/UlXbsIX
JCyI2AodNyQ0B0APWptrtvQLtunb67Pd07FO4NOgwwg9y7StZQldcm4lP7WwyBMQ+3vv13ReRwQu
9YK+DU/wUW68phoN9i1aBr610cJVrZmcuC0PtnPsOktdVTCXhszTpt/UUy9eCih1XX/SY018+Irb
nfKNAgjmLa5XRZiggq2SGyLDP7TCedLzPWmymRAQh+wxZz1n88N3D/x2Bk84bstPzsT9S6ju0E6l
3uQTWbo71WwYLvzBTtS7Hkbo0XQxNrK3F8lzb8cpxr2o9932KMNEMCICSl5rFO9mmYpQQyVLUgJ9
/YNk0GVUuOq7cE7DFy7zY0Usxus9drwS2IseTzaEsCDBPSw8nhRt3/tb1Wz8SvctME9gsxkUpWb3
zHMWzLqVpK8DthnfLCqooQDrFJKRa7SjW4TWJJCX7nkt+Hrm9fi8bp+7k8eBR5AEh4iOFtnJxdGp
qetCBd8PRwRBr0MIjoMfZiLyzLKtt1TQyF/9GDfczXXdI5qC4BBXfltcFqP51ngzvoNNFg//YZ2G
YbSJVG2SogvMLPf4zzM57o/pzH/QC2sXq+5qQPfpVzs6/KEvj17exuVDfS81B8mK/C8PygZ/Nszr
sCgn5nZLB0TQNtOV0ozr5XdMOpVR4IIsJgXRXAqxXQ6zxHWDhgdIEtbBGUrscI1y2v502FEv9r0v
e5Z3fDLS8r1Z5AjIGpxCz1Twt1fRq/K53NYCLHnY0Ftsxq1XVly/98U5o413uJG7Rh1yu/aTpmFK
OF8bzzKJ1Ru75D3j5LgUQMBbFNEXonpPtFun7YtREVEX6G+i8m3VBGKddD3f7n4gcqiXyHCE/KlH
CjG0nHetSepkOauj6VBMZZFsHmApseN79QilDe7nhGvhpVx3zmRgZLYIUL+A1v1U6EDOKe66abv7
9ZvVk4w9rFgDngzHaiv3PgPRX+jELEGBru2fCrWF+5TgXRRnOhhnr6ZPxoHak1871vzDT1MI22oh
xovfpEheKH/pazBKwlHAFVzhQG8D33FFiMf6LWzdPdruyW2p2wtNbLUgQmxe7ykCR+F8vKi6vRPw
TE+wm8D36t7SURK7c5GUOUhFeNk5sEjNpDzVXDwLK90oXVetQogsXQhJAKqd1X6o1lGqwd2NkGcY
GxSU9TrF81dheaF+qLtgspkx5SRF40/tJfbwPWaFG7UFe43PMQMDhiUFtS2opQnfPAtO2gGKsXAf
8B9lvNRvI/r12nq7Vp/RD4Qzju1eXeIcBz3cnwcO2Nd3B8uCNrwEHdQUV0jS7QcMkTwOmCot7i/n
j4gPzvkYtN7T94ci5Y2LAyd3rIvFGJU+/pmpdFfAozXX97ma2N/029XrsXaKm3+XG3owdxGuxr+Q
On8EPEuKDZgWxGSRWVNs6SFmwg6CkZ0TdXW4vqb+k9Q7PrcCQNCfuZACPkoWxyjUJjceD4UH3lzD
KG275DoNYAgLzwRu8WipULz88rbp4/ZwovrVQKQX+mPA3jOqQaujlVKhsxlyemeKaMIY4D5Pysbk
qksbjI8YRTwmnSo8TImIRTzEadER9IHX98VpxXxxwxK55sFoRegvTnezPx6eimVYZ03rF3eQq3kE
NoRyvXozaV3Y61ZArw198+21VGtcGkXq/x0W0csyqqfpA7O6MPHMv+6Uc+jrHsc9JuQn69OFSFso
G8UtMeqOvtRvueUDUk2b+KSbDVmNfP7tlqVUOY1fcNgaMNnSXXQ8uHR5V4c+jTVdlZ6yDiGDtMEu
Q/kDp6FBYnP+HIlx06tuBv+eIPcal38cEXYIcYDn5EbkvHzbOvgSg9rKpR8pylXuDF0zlXVDjnlE
/CQR48syXwI/OuWzhbs/LySNP90GUmA9Dpyb2ELrC6NGzTM5OFgIxuDvJ14uQaLZmyW9PIm5OP5u
jS6wpLU7A5EZwQpDm9EBA7EMqmjXLPpqtSYJi8LWiqsYj2aMwWPIZa5oxIRMyXJr+kWhPWTG0+us
lmc8ZY3q4aGz22PmMcGM4OZB9wn07Ff8qqu8axDCVWI6TbU/uvYE8n/z/5sXCBn2SCgp67ssq5th
7bXJmyJ3jYsfGynytOc6+wSDrd32PXyD+4BeZE/rAiv5xO9bz/sXvYncncn/dwU4n8C7ew9MGayf
JjQYkA339Q3jyO020Oh1NwjI5THPYCjeVqM998lQpkyEQEge6aBsCr9Ai2sQB4hJLvafc7RbXf0K
MIOW2J7xWtw8rWUNCNyjTuVRCOIozeA+v5jy+huCZvatw0b/fA3lw0EC2U8WBASdsxaYm786nUwX
E8q8V18aVPs0/SGZw0VS0ZILCHqpkgab6RdilD61iEAW6/FSM4/Dmayp03DYYROjrMTofcf4lXBP
tOuxK9y5Fc69MckZ+tj/X83ywZXdOjk/bMnbRfhuOClB1aNuYC6jJAPcgWqYBy7i2zvVd0e8F0dD
Lga8ThTC8Sw05uFL9WaXC4l38uALAX7lGZ1mfdEWrTH6ShOCJbTPTcPwBp0gXFytylWbP8a3jX88
dhHwmAWhEk2+6pa2tneAG+peiGcHuDUWX0OPG4AX20rAYToD40nDUaJeZOhb4dteHN5Vz9Bd6HiM
SmTaGq03haS0Rq//dS/WxvME/hGx30DUHqYWyAWhcF1Fo9NQInG+1qlKfwY4hTdse/nuRc85wPFs
lenUCKhRDOZSFuJ4N1Z2RN+5rufEbi3K+kb8kwQ+LDtDFXHuXA5wsJavyrpwjZAnP1vFByfd2ZwB
Tn8KKzbig/iq49Of2MyJvijllY6KJUn8ylScQf3NgmivuR5aWuqxI0T/utmYOB7wf5PYHoWKlGKm
kSrrVoYSjHmxG+bdIGS0R976y7/k31JS/cBL/gMdzMmX3aNN0OIrSt7JPv3AsPpP8+LWHxDTsYTV
xX/VGFHcZEqkw1F20gmEhpZQPCTM36uHB1hJJD/UgW0xfOzKuDPA78GBHPbCcBQ4rRiuOjnOpmXr
rl8ZaoexLovnK2sjKQnOitFm1NiVM8nGmJPuY1YyOg8rYz/mpEfKp6qEq4BPsgmOxvhv9r2jB5ib
U3eRAXZZgrfPqifSeShhvYRafxF9uVYofAWDNnRXEb/gYKvOUmwsj6grLItBmqZkKkxnKNZ+l5pe
/+tPbO6slqNOvzejRensvygLVuAQIS8QMbzjGeWWkZIM6APtZ6YSZHN4CFjMX1+3l2bxETNy94kU
t5sNLcBf3ywAOH0EjOzgem9rcOIrRPev8tPnhVMJ6gYa5UxlrhnK88jy2NuC0li7d72qDtJ4LL32
+/OfVSaHu5tVcR/cJ/T/cxbX0nQEGWMQErQstWkjECetG7jiOYRFHL312aV3LXlUcJV34XVPrOXF
LfMzc3QQThMBzWNjCkY4V6lVwLpADYDwTVmaE5fVAcN4eqwMa7CH9MmRxk8kCv6d+t0LXd2Ui8r/
PNTfKPwKKxPhsMJ3xQgVYCRRySEp+TYYbyasLeRr29CJ4rEc4dqW2KGpy4f+hSSw2HGKvAnSr9F2
GuFfO/ANAcHupdHX6kpy1OrCElGvZbWgi0kb/vTmkcSvvoEGv/lVMXxoxWQ66lVNy2W/z9Ij4hbl
+arL3KsS5ynZfzXdhVty7nhN+BFikf5bL/2kQwjuynVBRZn12MvjbkGONRfzNv//jiqCqHroRslY
hrVB6GctbneGJlbWNr0arLtYP9Xxyo3WQmXxi//JcTMHvKFjrIv+jShJc/PyYzMMAAuAkX1OJY3Z
9AdCgWF0RyXTtSS0xGk3ffjszDQFgWF6SaHR/rT7Zj5NJUrfkPmsL9MTHwAT/q8cw9Z9SK6epil1
fEwV9EKnmKMjTq3CMMIQJj4XHnpiBZshnBbNYFvZzz39xuncWpEV3hfEo5m4m6IPn7XI1S8F/68G
JtbFL+yxOlxOQqHNyJqo5ZQ9ITY/QQOctI96r0irWVs1XdaRlXlPZt5eIqC/TvZcrES4COTSDQZk
r0wgh0Dc0FMVTfIdFd64btbHCXrcSxyTJVpfFZqLELfRw1iSCJdRO6fqc5buxizmma2LRhMw3/Xo
57Lh0eTgfMdhCzQw0i5ZFYrjiECY7ytAwFv3tNCFY1riuKTiUHHKzWJQiTdwUhgi4SAOGmXjSZoM
v1+qsc/v+xC0i/L4bbUn6WDow9yYHysXBZR2CB6aogLLxcMpldSk1sJcGgOaN/CG4P9RNLyZq3j7
rXfVUaufM6lUqwCGNU0YLf+iZ24JXZeYnvVuCXVNsTuml1zkNuoQQhv3+UDuTCNtZYCf/Oc8OeAv
HPrwzoaZGyLabDP1IRaVlykAYQr3DA7evsgpHWht/shOo3SHLaPj5YdjVZ7Zk3Dhoe3peFY5ZQoA
koQzvI39W/dcgYwzP4aQHVoaLyJUgERKvq1R9QaXZVcE3uKzGzgA9iVg0MJ8tXQDjajtbamGC/oc
P22ft65ZgSaex8j/H72sRm2Ljy6TtPSCkx4C9snDKyFT+iI4PwQM3bubX/YDxSZKqT3Ol7BLf4UD
rn2SLRMEa6ZEb2AYogUTVwxZ6CVkMUZ7lQa97VtOVc7sotYq2nqGsyg1kKG0ngjIfh1/MYm54ADf
fNXKcICrHmdeZxWkAEv2oDbAuvW4w8pa6gjZttwDXakLiJ7F/vfIfFe+xXXor2ZH0bupO6mZtTzv
KTIfD4hv+kmy7d4b6FpKySrKjYGmB3fpxf/S45rdZi3CEBPaCAXgguyg8825tNNVA7pEJJNsd196
gcHEdfm8eltqybQRZB6XDfB4ye1br26Nxo87lwRcmLyaAeHVdYEiHr3m3AbNWVd0zDYllSvyNSn9
acBot79rvHCZpa/hwFnTPXswXm4BgdS9P7c7rcq30a3aQL+dsBxcKJAVRXSr5EXPBWcVIJ6bIKz2
DhsmiYGRIJT1gcnLxOifcJn4yGbUD6r5aI1RSW9gk+6tZWquq8R98qK0Csf2CBSwV1z4Q+kx5Vkr
JhqBOLKFwMtrY20ntm9ikOzLMvBnhEmLuT71RwoAZtd70XvDXDSmURzXqKoNQLdi9NmqS+ntfMnX
X3GnILuojcYj6P6rIV0xLdo1WpQ9DC1tlqsmHdm996WWEy4jdObvzKvSnS8eGsYzCRss6OVQmxkC
oyXQTeN7enl41BLvAIm4sRol90SWB28efx2xRfA3ZZbcm156CuxmZ1CCjXUX6jgY7E8zUMpmcWDm
Hcgm7la0NttoelIOqTXRWIPBWnFAthk8lN0S2WSMyUcdMg0/67/Jz/RurEmYAavWR4p8ArYp82h9
s0PZ0c67I6NhxZ9tCMDZFUIVYSPdygX22j4iWIMjozZm7NfoezFrZtiWbH9vmIzJIfd5aiMjX73W
+/czW2/qFje/Qbj4ZiPHCQU5QFVqTGNkyncqAQLaLeb7XWXxAZQ85nV5U4lIDjhmEbnj+QDV8Hio
lOFnYBkUE+q+ts/MpZ7SZh3cIIx3rY4GP5uU4+7J7pa7QahuT1YOfiAf0fPO8xJLmWD0Rpb2WVCi
KIas3RgH7wNarZP3WWjIf3LbHiUCoHAdtM9UzyAXzv3RdKhSQtlJ84wcHfh1HHU/HPZDdvMJhFwz
d5FQVd1lzscR9nIM4Xl6Zv1wwv/M0Dz3k8rIjfCjamXtKQlg52pgT9cwRKAsLQypE66FuZB1HGQL
i3pajqAgXACDn7APOP+J5NtUWRRuOOwE9/ZTRxl5o9+Tv/kIhwqvyS6oMphCoab86lnpTp7IIyp+
5JdWctba8P2AVoDwc2lSORBgtTHGKeG1KSzG5ag4fGRF1niPefNfFbH67ka9vYB65UceimWQKrkV
5+BeQvpYZ9x6FWI3CjDP8Il3Ht6Er44kUMvMdv3AvN819gAGuwj8jGMvQ8Y1NEYzGTuRLE/keeTn
Nt/1cqBNoh34UzGJyFJJGOahaUS8Q2gm4G/MknsEpnOG2ryiiNMAcO7DmeznbVWcHo3haYaFlMBq
bdaR9RgCl00EC/dWsjZeLvEsHo36JrrmjKjnEN8/g+FepJXbvOwiTViy54FDxBgxwB3RzLpSyaZE
26bpPCUlfAqsP9ME8UyAtBTKy1cBxG/CTVYKWAvUe5/6zKh3PM4QGwhHL57w8eSY01dGfqeLnVhv
QcScQJIKDxMnDoig8ZcMxkARYtVV8G3EoWlsWCDXo7TB+AsBWNpilJcg6qdBRbPEyW9xWgTn87uK
z9F+5EPf2RiyWN+Gbw0T/YshmRWbr7cUoNTKjli++1OiAELAVdj3p44/062fMC66a4FWIiV5oj7m
Al5m41cORMO8jd7GLDzeDO5TcePo1cragCoum622e+u6VplRIYKg2K3VfS6Izcb9WnHcg+Fw5n9Q
0IufL6bQJSAYEtg2A0p6ZFop56+diwQ9aBDJlnS/JtmYIFaQUheY93R5+oPQVPcNSIcuhIHXpA0P
1hcPAK0/LY9MbhffaCQmQF9OQBiXzzMkyXlI5nFjGWt8cpd66K9/CsUjqbU/wcv/lad7C8TrW+rb
+G0i27pYhjBHzRoV/jYun5TnIkH6YMf76QqbopY4AHvjrUMVvE0zyWrIwzJAwBog/TPNkWdVtjsp
eVePock+lvh8SMfRb08qJloCeveS8HZ9r5YJylDIhmOLzjoCYzqoKIYp5J2RI6YiX6+NWt9i6Zj1
N+AxSpwsZywS7eMdjO4DJ5yrL/siQ1+WkPeK4t3zRlslU0Mc3g5ZfMYmhUXmLLiev0g0XCQtuu+m
dNGaAJHVcoqCGiPyKVevxAInQuNki7FbNEH36LJBekeA0vr//VCZxTGxb/Mi+l1aHpwOuy5Lj0Ox
cCfeq1KP/o7VNyPaQlR80A74l7TzuV7Zlvjqs0HQhIMn9xJFo81nJoXrXh3EjUzyKC2gWBGdD5aT
YrO0m/6BmsCHTNtE2zQHpuNtSBcpNzdtWZad53boioN4wahaGVY0w2U7hNr735+y9hJZhUTMLcnd
SOE4RY+l99Ozbp8A8WB6bIuBqnj/YNTzLSL0iXguwy5xW1aTypBJICWiasW7+k10YOPomiXKSIRr
FOf1P2IOjy1hPVsDavYHf3hivOfy/ajL2gfa7Tae980E4JGU6JrLcC2kEjPJ4WnAA3+S7sgsdOTa
7b2zNmwuFLBfTBrck7Orp+P10Mvr2XN4xoyFfW9diq6jgcfzlPjl6n/PUcVYsGSiRi7MmnU7TXlp
Z9TdEF9XSmdQu2AU+cNzLQve+9cK5zeDnwGr5dp7LcFgeKtOuFQg6jMuubhprYnMrvf4Sc60DDkG
9lvGFeBZZZXCKB0RUaT9DHC3Gkp9yYy6EuT4GoaiyGwDgmahHA9iYY8Oai3Yn8n6ej42S6dqcS8b
Pl/4OFb7BmiWkk8FlKytx/fRLE9Ip6oQuia6XWjSvEN0hZ3wDkMp5xHuzRc7XGXT0UxudbAUv6V/
2JB6qMBCHGdFiZVGTPQSMXwGuuyFKc1kp4Ed8ZMroJeDxp8qMkErlYD1mkvtyFX8KhowbDYaRmrX
KGkBw2Xwva5zFMED7kmQWWjLqZW87whYgVNSHAN+tycg0wvoJXH2g+fx9wwCqrLtFJZlos0HYqP/
lmEx4/qWnDRxUYcFUBrZtiMkvUoSVbLoBLcK7oWUHjDFb26SC+jGoTUeS06EabI2IEgrv5zJZ9Pg
uuJp+pttHhyc24eyn573LVvK17LUcYk5WdGQi/16TzTEUA9Z2royAvyqiKvqA7bpA/pkWUUyHx1n
7N0PUeE/XbgSEFzruX5hD/H2a16GdzLNGsl5q/1d45loRlApTwXHTObXACxCq4oCviQg023I+IGs
PWX9Z2IDCNon3RzqMtLt1B4ocL1qzNKaA4FOsGEXyCA0nLtvHubbdaJ4kPLpUpRW/DLAeVFet1vn
/CkBzSpN+APe5PwiC2oTRSzpybHR0o/YmyWB/PDxsq2JiIh4M4qp7iVvzXG8z9z22syxvSHDxi0c
t4uDAbEH3f2R922jRSHsXjQlUoDeuXDpdhgxaNoC6wJWbxsmzEZfDah1btLW491Vg/ZmsYChokwf
dqHeTB4xOJvvofmqjzRpQkU3ocT5clF0RbzZRhNj2ntDV/wDXxnW4qmSFQOxRbx/eRK84owrCTfv
OTJEzU7GgZUek1mCyQ0z12hBPqKj7sdY/trSSQiSHaNACH7iKzt2QCN/mWpDSYxOZH2BIyUt1rwv
yIlUvFby12FWYDGD+x2blYzNmCRYNP8r75WaSbfPK8yJ0hrENvjdnGngZ7zbCPBnfGyim3wdBtkB
oPy9X231nFN+YPcipvakhjFhyONa9TKuLR4UmUAbmGD9lsYVBVGba6SsCN3BIYIHRk1OuCpAURbO
zxO7+fsvAm2SNtXB4wa9Cnq56YNWSe8r2XAGH+msjcWCqVBFo+YUwJlkXQgIaulXqWVazL+8Zwpi
ZFpogudW3E+qCEoM5+JCKdK/mSrRTLmxvb02mDgGwG/wg/+oAG4Iw1PLpgv1qNEE0BC7ea5qL5Ef
qQkUDUVJN7cSPqWuqblCLAjZhXI0jEy+oRJrdnQnPPngkIVpPdJDPn8HZg/yvVzqRaiq6N1u5zWF
Mgfql1YCrwnUqpN38qKAe+Mf/vVfWSON0KuURRM3JAVhJDbwdt5qwMWtluWfD2NIFr6APYUnSRJZ
Gtd99eSS/+lVkejpVxbbfx9eUP9zOVw0SsDv8dzHKnpKeSPdEPCWZP7DCWIwlxAVdUBY2v8hbcta
TGPLrGTZMxFizJstFAMX8I0ogiXbhgTJKE7YgQiHAgqb+FIIX4UVrn9QzagoHx3PjaVoxP74BB1Z
OSt8sOmGExgiK3uZsHLBUGzMo0pBYngwgGERJP2SGxtVNhab2Cpd4yHbqoUxRLnXXoI9qEuFHrKP
lQMnUiWVBF2mJApT0dlveLpBqzCWO7BGYW2XKv9ESbDsoAm4jlf3ernD9ezemMG+vQLSwZH6bE9s
ZXLVk4sfYkbhc+YJox0Uw6e/GY2dvVaiF2AI/xu23IG7gA4XjHZleoHJrTiuUkFZVnnoljREQQub
5jXBq0XqQtlmt8N00Uo+SSUewhKQwGdkAfvnZIrxtKh4xMRRmW5BuFgTFeYMsn2hW+l3vkdsq77f
jFmp/gJR8r0WtzkZC+xHs7bFUJcnRnEXHfCT7u0dKYof26pXDavBvvpBH07ZXQ3n0GAS4LrW0GmG
koZFzV2Bdn4EV55u7xUAT+t3xCmd0BnEfPxcEt5/r1aXcJcSbPlClnV5yQeht0I7L7wNe/grDiFg
Lr39j0q+wpezAS4Ve3WF+WzI+sxjFEl9gPtyxNlzrQm9EzXwl9cNLXSOQozKTbHMFXMIjeWJjWMF
R2hlg7S4I7H6ABOP8r/OeZgoHOSxOeqACYduCxWjaIiT4I2fVN6rOdGjMpqToez1zLUnooCKNMcF
/UUIrJp6iJlvehhEYuGs02v2Igna49RMxZN5NjH1YzaD40zyp97RB8MUB7EJn/wuu7BojJxkrJFO
IQkeGVY15yGiFIHwOBnMBqcMl3yM0plCTah80vQ4aDqoG7tKvpLk1Wm0i6lKkgINLdo1HsYc+/Lu
FBmyJ6DHJIPyElKZAeYhQR9oc+x+BDdOk/qmm+62HOf0E2CCmufsLAus5kTg1BSawjq/LGGpk1NH
7UckVdklTn4OsIHzZb7kg50AsUd+mERCo2QEraagQumvfgCmKVEDffxGYOiyft3a5D/AlPvs6Xjr
GfZh+pEoZCI3k5CzFkAMQcdOCWJ8N0m9kubgyHI8A16+yTi5lthcO7dmlnDEKqhuAVw3IZaaDvLX
UtykVTgEr5Plnh4eFXoOI3f7dL5l5GJdDpy9WKPZWSB4GYKNuTVwHy71SsXmCImRyT29UCAqFjO3
sGn0eU6TczuOWJafH5Oxaxuaq4kDlEj6InyG/axgDC+kewlFp6uoPC0HpDSsfhrGKbygbs1pnpNk
yWW7vhhM7KQl2UlO/jYL4k9didlJ05TxajdZlt1vMXL+tE/I0c814s8c41sLdvwGUbow9bJVDGoz
+K1uHZhPffiE6c5Il/bF9Uwmf94Sb7gF2OXkFH8TymT9SeEv6YryS542wE04eFHeXNWXHwwjXdcj
htXZgaJG8uzOY8JqEklc54aeDppMwfE8k9Ogy8rPYNV9YWqNEuKMK62WcT+eLMUYF8smZLiR32Jp
CzT8hzA47XJ1T25MpIQ4v2btXmiu53EvAvXVCm1XvP1hcGJRZzZhymagYs+JrccpieqBPGYi0lwo
tpxAW1fZkHXWCNXjYvWpyt8q/ER4vMkI2IU58U/lfc7PMfgufigaWa9y8GiiE3CQvXhTqkSgjlDj
JeeUyFVLR1uExDx3xtMEz4EIF/rfhdl6jSfACcBHgRC8ylodL+4ghWdeOvN8NdD1D0MXjTeT0GHP
qc0SA+NImM7AXLg2hSSsCaQ4gON3+7Hn43JTta6PNs+nkfJP+VQedQqC8M/X3x0KRxwrF/EpeLk3
qyFXcDoqE8Lxu1/fogLpz2uEqSsP/qB+YJHyB0DzO5Dd+0gjSzkuzh3mI+kPjGBKDqy5EdWNw/7f
MfyBkCL0/cB5/VXvwX3u37m2hvFxtuwePQ/fQNedR+0UaqqA7eZWLKV8H3Ks6FsbinlamTjKGkDE
PGx6tUV21KLJvCw5Na0LmLiYkfAdmQVl3X/m3gOawMiFRWOwGyeypYGJIsK1CC8dfySN3JlvDemZ
c5bZx9EGRr+o0jiNh2DLq/3dkAkxt/2/sL/KM+AXVWfuihzy68pcSN1Hxi+H8pT21TVsfGwH47j3
jqfogK0h82bsIMu7zcVrAOIbBJZp8QdI0JOVMhy8WAMzkTJjT4YT1e1E3aFViOJAifGjpjmaYXYe
4f91nxELv8ZAxHN8zDLnZqXMl/l4FhoMz2xH9XTmxgf6MPmdr4Ysse+yWKvYtynEfPOHCoZpyeAp
Go///Qp00pXQA96GAFMMMOojZW3Sw635PAZcJdrqSMH9BuGYsc5ltvvN+g4R0qfpr727b6cLrNiA
NuvMqTZ6jXCcuQMBAzeqiff3+SPqSICjVDYc6zmL9avPpolDGjv8Jjf6CZ0AElMPUk7fJUMKD1IF
29DGSozO3bwuMqA5cGKGqL9ca8Xh+YM1+xVvjtCPBl7drTcQ2S0vHueDpI5FGqPWU0zz5oW5Jzod
JKbbKEOJ+1xx62tf1qRH3EGvMMKzvthSlzoYqw+45derW5ahQjI8dZthachaklBbd/Mi8UlVL9mI
mUngIiTqSb4RFYOHwxa2VTkghtu6zOG8ZaPQfzQO7z2NIluEMGRxAnzv1q/NPXfCBwTEd+aeD7TZ
swDj5lqoxMemCrsemTxBMjgI7ablFxLhfUaieK8d4UHJMXr5R3tBeMSqGvzhxVPBvldDsBmJiQoJ
1QQ1xasNpNPPqwQ4EWyoEP87XJV060QuAEiLd0l/gUObJ6ATDuVDC/3T6manFG8I/Ta62W/xm0wX
Dbqq+eThdCz4kamkEqBXVUo4DdVfE1kudovG5HM0cxe6LlWBq8V36XZABTdXd2HFizY0FCitAq9u
FojiVXKLekmz0v9VWqZtqATL4QVkJ8x4VuiOV4A//X/ys63M90DIJMS23KHYpXweZrR3exCL9aD+
yuJKeR8EsgZvdF4MQOItHMsQjPPKa021CWnXTEjC6AsTzdmlEgN22/yyupsJprHTHe5BtVzRw0/V
L2PixsQwgzYMMwNKWJ+X+J4qWKfnX5Ph1X8lDjJEFP+AiMEzhof3pcfi5rEX2n6ogoM7Xf0SrLCz
As8BWKlYSgYgAnB1ZEj6kMKYZCgOWhnZ2pf+qow0OqplmjckgW9QA44DzGjYxgY0+yCxyfUeeBE4
9VPaZ0TYmhSQvIP30+rozG91MV9wLbL+REzfWJFFr1YxkJ/B+wmlN1iEMD0fc4ylCfnV/wKDxwaF
lfN7vK+ITBy7Fh64i6FduazlgUMJw9o8ITBsHP38tf3U/T4fqrbavS4qimNZRlGpDSx38/f5tgzq
0OQOOWc/x7mTUlbD4v1zw1zYSg+9w3M+19oYjEbZaINL3tVERArb5KiDnrGCmUZ0rEAuIONAj1hR
fMQSMaOK4WcAvl1MIVULMvNKoAH6qyybbUvGOGgzlohLA3Aga/GFN+bxrq/36U7LedUf9w+BtQ+1
Yq8+Wi/dvaN012XQlKAUHElM9VamkZJ0D1+sR9QYFxS0BPdR9x12qtPpLUdW1+ESBIvjPKp1PGo2
2olsucYd930O7PeFVnrnuW7Po4qtHktM2F4/boVwaO422OrGhTMphdMqTzW7ncDOruThl+r6mDZW
aAFn8facQyfK36leMU3hMl/GMwGls3Cs40xc4mQDSHaFMsvXq/hTa19Sje3ZJZbDiOzFM54Q6sG6
rEwG3+6rVuuelkAW/TP+kXQACJmFMq7+fBt9gDrg3WcMTIodm1LI3wzN60qU6zOq4Snl5RX+p2SD
o4rEM4NST9DRqZzuz+ENhOka1iYtfbrv57LH2BsE+2BGZpzSlyzCG5RYgNQYMkkM2DxaRQUKLqRh
y/SzSSarX1IaF/SKveN4pVEYyZVz5riP5nnV9GRDLMG6InTwCg+kZIf7qZNPg0k5W7aG4eB/u3H0
eezXOTHfwsIisIg3YLhC3ikJMp4ndCl3lh6cz42kJdaAURxn5H2SEEGxV2mJuPMx3r6Qd4Nn8gf/
TGi/xYidLXf45oLCzez+Sc0wHo1oLqeMWbdi1O1WmBEsaVhaobsorTn4afWpVLmJin4LCTLUav05
vQTpLnMjQSl3pwSWWxsT6aSkOUBbOR8hSOr/CCuhnpDGZ7rZDkYQORCtPfDSJehBroCKhePE9oS3
Zmdz1vNO+yKyrxpwBmo2IGTJseex3ipchaWninPcGwwDXqGh1S+encJZ1OeJCOVzFQ3TLnlwjOmD
yh0PqPb8OjpcImFtjl9FeRIBoNIhgTrvpYfbTLh8zYhcZK+ZlCollItz3yfTUI8rKz/d0VmBSRyB
79KDc6ZTGu+Fq6/cHWBZhxj9FsZztuio16B3N3f7O/CEFmLVEJzsWkCQJZzy1bqlZxh1EYOdlEbW
osTQK+W+ZelFDpknePF2rrzPCgWrFirWyPNeLHCok1HZ9KO9pPcf2Fs3PJfbTNsNb8T4+dI7Qo0j
t7v94t99UxAKWQ1Eio9sK/i0HA3Nbi7lv+qe53UOuDCSfs4HS2fh14+Hs2LtbQmYCZT/irYdgcXJ
SGdyCye2ktb27PSbdwzi68dmZHLCeIB4xKCi0+DexOJVEDc9vfEO6Bf1ckPps9favce11qqdRoXQ
xT92VV64mbrsvvsN+P7oYtWIP8Rw+2+3Mzn6TNfxiZUvvx1v1X7llrGfZLT0otYzj4UHj0WYef61
zAjxlSK4cgfGCysYqkstzZSoLLuJjPBmZQZu5DWxT/SbSsj+E8yFOZUwGAyHAXoEu6F7Kbtm6kFT
MwwhMxQbyZp4mkMN/TCx8zJdgkfWijDSeY+jTql3n0lbkwneMz+hcEQEHm+8OBxSxxAq4iafY33e
fGaC3nEv6BPqAuAoYFXkQNAkLUV+F1jdi306v+c7WrSU0RvK8iMWbiZhj6av6olceKXl1G7GNN6i
TMQ9+QbcEponIYed1VN6dSWaebrFUt12CQVOUf9FZRZKj2kwCxynUbXE6QzKrl2830apxK1kGxMk
HLnMDKR/r+vfhksfJk/2fwlDBFteEJaTvG0E7A6U/v8UjGV2rXQbsYP83loiPDq7GxbhriTprDAA
/5MQMG6wPUNNm4zA8x7nEbV/AyLnUfndYXSPw33NbEg/eJcUeihbwePOTGB+W4vFd4rGv67CRUWo
woUeRSTnV2X3iGoIldB4JqszAsszrCPcie6iRoQXD82sdFz3VMAdYMtE4jiY5Vg8dSBs/eQojt+t
yh4cckRNtIGTxidUd/FbCxyXMqDOhqf9NpScOf69TdC5Y1uZyhN1hL7h8jOpizRyNOKJj95JozRN
6c8PSEpNTi1hLTINjJ62KsS10yAQrxvZWwBODiV4aXRJYKkzPzUbKwUZgMbwTIFX/UjzB21bm1bS
jbWCrinyZQx/xvuuCtfry/BmDYf+6eu7JRiyrWS7d9lTy38Gqbaog10PesBWijJqmQ9ng2Q7o8WF
enW+76Ae8exdgzIbKM+L7BmWn9BRALo7nNDS6qq0n5jI6OD3dd2Hct/ZaiqhUMmGXmbHuxB56OPo
guXeB5L3ovC6j1W2Q3Lf+oBknyRBLVq4HIaRHiZ/B/1o7Tg8kFrtlA1v0j0RngrTOPiZJ6Zs4V1o
Y5y3l1PrPCyhpyNR7zHWM6YdnwmWcjGbhOmeBeqEQitfmxeYYVcrptTJs4vKWIw02MQD/ZrCO4At
QAvsB8d5iOCDPogmVZFO2W7sqBIo+LdTqK2m0IXlNyTbkrZG9BbwrClh1tGG049BKN+y4xfL4lHk
Y8Mdg/mkFxvJDLImobCeEnW1CwvvepmmJD71xKKl06LOyyziIy/eeZMMhNxY8wd1JLZwKJ5zZL+N
5paWwrd3RdmRQa1EV9OFoY7bjhbs7dOsoU6Vouj4fbdazicR9EZSvuBsgkVkqm4TyqCzEK7OhRGl
em6jybmL3qriWnVl9bsFJ5Cf46t+KJr8V8QkfPw9QqVkrT+6hfihzJVxkTr9M9S/PdJV7FW1Fjsk
WehvrPvjSBVxBogxuKjiP6+LslYnWAmDJiB9CkN0jujB4TOAVZAd/0rvCgOeLxTK+/+u+yb9Pqdj
iVIDIkbQU7SJM02kztJiWFHjg3ufym4Y0ZuUHC+p38xaf5K+jcvXoehZABOyeHGn2D2LZxcPW2Hi
VK7lcSdkSo+MvZXs/3tw4gO2Ajbbjp/qFnhCqTGOQo53/nHJaM8uycQWfo2yoLUGRsifwZBboaOR
SOoiX9qjF/i3fP5+qNSdT7TSaZuA1wDJAmi8tMfiep4XCQYttxqXiXi9FHWUzxFR+E1Lh+0/gOdK
hvEku7yG30ckAo+HyorQWHYxZcyzoiYz6u1PEZP/R9CFxZLbcthMw1FAvdxYxbo7FPGmHlNURkWD
wqFwpM1rbiEP0gHASz+k8VcL20+6lRztmZKnFG0Ew/cIDcG8tssMG0mK8Et3YS08AQPIUrsEXR8Y
qIpxWFtk2LKbZVUM/MM9+p4VmAw+niaqH7wRaseLNGpbtTSCrC5fJTx1VneQ8Po1sJPAIDdboMfY
snft4qtNgqEhw6JV3QGtFNKzJtH2fuhi4R3GdMhS9JnO7m8N0iyxptOQQCDguGBWCE6wmI73MBqK
BlvV8CnEPq2JU3TgeabSyW7JeA3IL2+M63mxHiSPGXwHtNTUWrAAELmU4B0UkwMcyowC1IwO97LB
b6kWwEblIjrNGMPaS4gfx+i+SG7LsQppQTd/xOfhKT/tQcdbO7rGaMnNS/o5+JPf2QJuJPtrksXH
Xsq8rIOvVQpGHBMmp2/fEnJWNM8BR8ZHvej6/8m54Rvl3Pc32+UzCs0k5TQaV7kdfih/EEKxv5Yc
rEj+X9yhh3kY+5MVk/VMh5TLV7/lRFhib1nSYklujJlYL1uhvZuMyXX10ef4R6Z+AAr2yU9w6Jr/
cYsg3K3zHkjlLteSUgK+tNGKXDHaTe8m0QYCfxJD8nlynFuOXrREg+votjlexQEA6uTk3okk2M1w
CAlSbEMHAChCxfXK8YiTFIRLqtswu9h2nEMgzebDCZ9lz613WLaAKEUoa5nPMlkyxvF/CPKMjyw0
siKPlOTWRsmIr9SNgK0aQlxyYfggCVqnTsdDi/b8A++5sRXh9WkqmPTpyVJ7rccrAUKbVQN+iGWZ
CRUA5cCcYMPopm+NdSHfgDL120TBIFMjB1pGPrOI65CioUlsaaJ1S3Sy2lAHMtlGgopgWwvrgnY2
ejQVM6gsPleV92UlgtSnsh7znnw2oG94RS1x+sUUQPp3MB565XtdM4E8Bl1A6utDDy7Zaed/rX9A
kVP8C+PS2hcnjBOUQ7jgQf256e0wtz6lcd1y7oeiDrZcov490PkuypDlMHVjROLCtyliEifGPLo9
AWEUNDTxnNZIL8phcIaQ6zly9xg0mOMNk+mRLnQfu9+1xadzF9STiISlvBirRtw3aUCNm2uIanUG
w2aknyf6/9PT+wh8a0RpL6NQIW5S5Q6PtuhPmCL/tX4pBBWx090MsUgwg6qw6/I2UADSxfDQ3+P/
Bm6rnT+OJBVAac5HlAN5V1rEncs5kogZQQnJSIDsGLHfb9kJMnPaKtd6XktJBLPRatDRn0Y9BWvs
/B41N2WEGs3bWQkMvpczr1boCbfpjd9QNGjEoMGJKuje/htNSckqVsmcU+ogO7U56o0rL9VBdEvS
I4fUG8Z072M6bJcB3Jl4L7sl3hSW7u0j+b6xjauWb9QiQRl1yab0AF03ZDzRMkvmDinmkQx1cTUF
Mtqw4NmT9sWqFVe8+6d5hgZBs+Vn5uyaLvtj8ZcOLhmj8nZRUshVGXRJ6aV9DGzqQCbMR12zRakg
z28oweEp1XY5Kz9N/AriMVy+6k4g/uCDWIDRTyHATBmtFCUqoo7TkF+Kur81BP8VXx9+1lRI2bZS
6c6C2+P0IQ5CyoEOr8cMKfJVxYX08zmV6Xx6H569KSLyUpznsNatJ0XMPdtqcpnckrNTnBL2vj3F
25Gi4lYFMVTnh34OEOON2u2CUujhlJI8zknYy7K04EQypsGfTgjiJX5Es7h4rNKPiJ34NNyCl072
IO2D7xXTv7bkYkgOB+vuMPtZc/f6UYVXXrjARgZUZ7rYmG+OlcVXAzYBy4apEWJcO3JfxvqyFBTX
TidNEVplZNfx20aBXOiDLoe4gIcO7+R+ijFk8rPYPutWKS9r2abNYaS1wVgvigqfDF3SEApR+52Y
TR8hYE9S8yvffRZEC6NaoATfDvkeDatpC6bJrhjlG4gl+Fx+57c2tMvs6+enkfAd3bLb4iJ5VKMF
DRmWxJ0tOrxcEICT9sUQrsTd78HQdAtJMruBSO8fYdpIMc5sg5z/BfgaWqCYHsgLFH63yRlcbmC7
GESIBKL65ZKxjm0avhH6xQzCG/uXBTOd8B6sUYZar6VXx78+AnQzTYZbhFqv9PZII75WwlsqCAQu
D7I/MopJ4c9VIVPMCHdBf1rDfsBao2qus3QiA/WNhMItmRtw28PtVwkN4FlFDjaV05Dp8e9opkGL
urGO60Hvh507y0hKmA6GNulQO85nHAkgQDRiLJQZbIpWAFjh6BHjgHXDsFtpTp2nli72CPflhXOR
jtwuuwBrM8qtQLd61O23GM600fRarLxUGIIDLojH5Zl1C+Yvu+UCwB5iY0BOQNPGG9+K02yqfCJl
buoh7T+9CrZ2uy5Kwet5n8qQcVucLw7DenHdnflEnrY/rkaH2/ptjXGHq+fYBCjiQOKJck6Xn0+v
chCdtqgRsYVFc8S/26IVyInyezW4swAbcD3dMx15hpxOc1+9IPUjbXbPHpddpS2dMd/AHEInb6G8
cK1v712GPcO5Lh5khdgWcGakoHNkIrAWfxL1yi89D22ZNgvo2fBU3L+fJHMkMq0+zGLemeR4Bqkq
x8lJ4A69kbeIaOpYutoUGZFZ/r8EMlI65O7SIYMeVxkQ/15Medvmtj4miVcYRGDmh+bJg6Sh++Pf
uur9P5GjRowAlElZVJTKgtVHWAesnJLhKDqGxNBat7UcVCDcQtgyBJ0UQeKIBtNZHmfHLJyBwfSu
3QKwwZ3OVtY9qxFBwiCzQIR2tngWKU9elZyUhBG4GS4e/9YrvnBQc5mb7gqK0DJAIBFoZj4SZPE5
DQ0sYUoLYUGylWeM5WikMu52IXtBQwnB5WWDMzDH0lBFUL5SfRExXacgJuSTCTxNqZTxQ5FGNX6B
fQrlhZ3AsEfrqeEAgjxKArNgl2eDNjQmqgv/pRTfJMPcF2kGUfqGtBgjrzb0XOW/z04I3q9uCkf6
JimX2uAuf0uGP8VHDMjKU6aTGgRmONyzN93sEm3NEXhb0Y4+ZY40lqN42Zs53bwUE0rcNBcZS59E
EBA1obGdrndyILRHxviAIxQGm2RUNgyN1aDRwE2g+U+ScloYJ3wPjMYBNuaPTiWeG/60CSHBWp6F
3CkXyQ7icQ0ZrHFsoZ86d/bzgmDjgfkg5FAVzcjD+nyHlj5zrktYyobRZh6Gla4iO+9wubdlrqun
JKBWkLYfoXM/ynNxLWXGcu+JlZs8oQxiV1A6oBmPmmVLecFmoPq5Rb/VvnS9UoD9k0W/Q95hXJIq
yJgPU66rfor9sq0VIVoy/18ij7hGT8EnrbE4GsGOONOrfycTPZaDFTzZgPkBay5vfFzFZnbATggV
BEMMkLjtyZ30fvTDG9j7qxb+iP9ZgfrWAOYukEWlc9yUlgg9q3X6mTrdO0qMEOSTy13DzO3HbeXz
u4w3XnwRGEWvm6uZjXXyLTFnlgJLoRqMhTn+r4sgYNjAcFoYEemviEqSwhrl0zab7C1u8IxUb/BI
3skRAQZPo6QouI7xZff3EvhNqiyJe0AeMaAsAF0e8TIhMdM6H/47Ee8Ud5IaKCPgafN29LKMp1MS
4pO9kPqPpfzOPlYoc1SCCh7x6WJFgUmZdfGZpmmvcrWwRwJBqsp8p1JPTIN7sz9VfP9fz3O5DHyN
b32UsqakaFu+0u4C1RBanXG2Of3r1A/YpSifnK55iRZQW8+4fsrvDyal1PnccxYf60NvBiggioTT
PTJswpB/jpS9Wk5ly0to71ayGFIQYLN6272TBGakcPFsTxXJi3Y5MeEA3Xo5pc0o1wwcvV4cvHs8
t1PCK/iFp5g1kHoSFB8i0u2xLHWdflV1Dj2ImvR/ahAaL/9sUTu62CxWUeaaz16c29dhBPaYzpKw
hI/gOlrF4NUzfngR8sYXkf8MJozSywCVCla0TTX9rS4bvOUc8dJPkY3PcXqbRKUpSLioTxF4hOIl
l4W1PBzeCBHB3vRUrlTZPgqaAIooMB+a5ar6MoSFs5t7zlzcXUSuGae1VVVnJrk/KeGUV2kSJ+NG
nXMuWkA1pinJaxC1wTpqKj5PbSIfJbK37JXbcqTbcJ19CvsxPYCD5Bw9QiAmMaMsPV3Hmu9sZbyf
2GW8hAazWdC+4sxU2PUe/dGbaj/E7eyf86r5IyE1M6Qb6NoFRvaae7riFoeLJ9Wty12yLb8Un6yr
8BqOTeF6DjiePct4eTu2n5k4pZE/WpqHLAp2bbG8x48isj1abCRT9OpL2ooT3F4cJ3qOvnj3iqC7
yS7CecYJ0wV40jsxBYiJ1DceHNM/q2vkklOM2Cf/HIb6N5SXn9e/LwpAjGhLrQ8D+r2X0xl9AM5Z
xMuSKNaH3FDG+krxd0ZeJNRvdHpiNNouHOe8FX36ijdKvatHp6dmz0F+h+UDLLXsK3k0YV7PDupV
05odw+iEr2U2Y6TVTLqt8E/ZFu532oMP9VqxIOOqy1GEhTvqt5TpUmcId4GsLM0hU0BwfyDvCS/j
YY2CmETCIiWn+GOXzl3I41YOxnklgWuCLC9kBZS8Xs4kEByMHwYBjpTA8DYlrvy76wpr8lMmvaHx
B1UvN+jJ1FdQjvQcfoyF9c4Cu12zA16MSMUK9VxCHs3u6hkQOlAaSnfe5gd2ts4QhL9koIrRBHKN
F32eJPAxKvxJs1WBpBwT/su4SLAEOnbwD/et2lsXGqyhl4ZP4TQ6jVwJxZ7YN/SV7y/JALZj6FHx
mHVf0j5z/xQCNd0R1C5Z1IP/QcSfPDqZcaUKnFnwAznNSwl0Pqt3EKw3ivUzPVlEPUnsC+eODGYG
vLKX2ERetpvbujY92BHHRKc+ngeGo44PS7M90DlKxq6Yv8L1RTOTfPqWwIY7R55G05olT6pfL59K
U0m094eb+ZcuBBu7ZJ+u2FYdb6pfW3k2ECAxdrKm/Ao7L4detzBuDxSnOSy6/Sjfuj7PoGHH2doi
8IczHt0q3Kva0LQ1XTzoOVJGrWMHbHT+lrSfLbliC7qSqACCemlTEn+HjSqPvkwcgsFvqD8E6pbq
gr3lqLM3BvZgGrGeC0EvbrJf0mMBWSFcScxsi/w+nx0hX/TQQ0WX5fAaJ97R2JuRsZh1FToiC5u1
jQzIYSkNJqiucFqs61aeEr0XevSqIhipoHxz3E3triVxZOL2J9iY+Y/9uthWOVk6/XIqGZLeKeoC
7g6Z1awVUImpB0eACKE3Y/1WsCsl8GcUYC7QkUbr/oLxNSujDmsYEME4i23POTGl4ZcSKEWa8/fJ
DlK1dZhEhNC5cMjkH0BzctBy39BS1t/OBse0qE2KlleOSJW4T6G3gTgCKjD6dhzBEXdlo31ItK8u
/Vd1NeUGCmOfc0ETuvTAuHPpKxlFyX4afmOj4S1FWV2ulTQIUPIS/P5u/1Mvp8iGSsiltSHwsWrq
DATHfam//xWQlsxKFTqzR8LbZ0OHUQXP7saEe8qa9z1g/XMowSTVKOg5I53AIvOeY4HN2ZxqNsDP
+LOCDFUFTH1PGWUK5E/3wwOTd3D1pgi+qj40srVtBxdIcB7qlhJg/i0mgObNf7RtofrpsH5jSh+e
wFUil2MQsN9REjpBvwyUPT+HTJ4e7NW1j3sN0zXAbfKVnqxygGcK3tQuvl5yYrwo3i2u2onYSikj
ZeWNV76PiWNWOG4B7xFu8HvHvOHZhfb8f1IpdSZ1/18KZYTrb7Hp5U8WMEfP7tY7e/rr5GFKVghP
9mdja99HVPQdG1GZFYBKVeplTzjfEEOlq8AwPsZxV3H1lc0XH2LP9mECt66EICwgLZqGdto0O8Ju
+ZHGqzSqANcPQnOgEAwG7JwPARTo/NaEuqXvV9npWmKSDCnYQd9+AHXd9lHBZsZt4b6/tJgL6+9Z
Hs2wJhsS0A7pTT/vyo9f04d4odk1lkm06em3F1OzVYvMX01KUd7bx9RFnD7cZvSGM3bpo0UGB7Mf
AM8QUOfRYuzvBw6z+8dFg0UeBgv25yUGu9T9xFDQN3yam36NHODlQaxwbIru7ygXPCVZIEtDO9u2
QiXgRCHGAezLhhCK8nmj/H2kPSnQp/dJIgZb6NXE7rLEYNsy8rbIf41k87orQijKxFP+R7OjaD1i
Lbctz4tO2lnpcuaIuLWF34jU/vjDPOEfyrJsVEt89b8/vzyiAam3qTRD+VVwWh4ai7wl21kXtwjZ
YUX0DJYT3woUtzUkLlhjUiCLSRAQljpEfstSGPrnd2xjT66YH67M+XAXuQPUYfZs8gipFhXfT1PL
y7+LBOud+D101FQ3Ckm1nn8FRTXkMc0FJ6pja8frCB3DYpcEW8yzGa40z7st8W99W92VqWVKEiXd
Cw78kBkwOstFbXVzaBVrpc9Ztzbj6felFEPG3PYy8Cy0z59QlKQJiH8a8wh3Y9nL5h44IqPpL1wj
7v9BkPkyCwBnJDFCzR4MX98YjraY/WgwvR9/+syfLWgK2hTvrx5HhBfuwzlTf4ogNsidMP5jbBUA
8+MXCWV30JCoW8GtHkejk8WJ0tTTYqktiUKIj78myNSH9JFObwDLEZ21GMYCBsP3bGhycbREy+8s
cs0XB88AFzFJDD+iUyK7FGtAqYnC/M/5jL0OLBSSRAKsb7Duru0n9xUUaXRQlNQ1bb4VtVaRqEKD
IHqA5AvJO+aekDLQUgiGMoqyxDFC1koEFJggpda76la8WADjE2NbABimzFv0L1n26Fie8mjKuEbB
gAnkxUo7dQlUmPw1vCXpwwxFBRIpmc7eekeQQtSsCul9v30PfgjB2owZSxy/mHbZ/UuetQ4Ujhar
IyrcB79rU6htvS01ewTEyoMyhUDTn5dRkV/tNRuFX+KtBzZnKRISi9OP0b1/YlBXEemT1HWPPk46
Hf78N2u079YFhTRIpJSXizirIgewX7t3szSzcpxUPtJ+astPDJsvKFO2EGhMLYHknBe2CnxdKrXJ
kaz6l5TdZ/QNWLKXT1Gy4Hhg9OISA8yoxCk5QO0y2YsF/dCEQFHD6lk+E/Or/3EtW+1Bf0AZ4DNR
KG4VaTOV58Ed/F65pGGM8kpOr5FNuZ1Yf7phPo6kPua3hCvWvPLsVN/B7zkiCTlyNj79oGuD+Pqf
37T+BoO3ayzrorRrqvweIzRreEBb9OnVM3/qoX+SvSjs9nxLYT42mIccTqqZueidwZtRzfN9c3sW
MsrlMw7SRyzfuM2DZRYJ72FVhxnRTReKMy/D/GhktoCpQHA7PEro8A/+nFEJb9vE+5vgDiO/GxYL
LTrYmWtJIw5xwToFwzWvhwsu8vT7AXueoFTZ/uuszlRJUKp4SRVGE8tvTzwR3jIaKArLMc8WenIt
EPqYC1/gryaima9EyGcEUr/PGI/V3v0fYuslaA2qXDAdYM9MyhtAa1bhRUejrmSTQNPbv7k6wj89
wURgf6KQiYdVeH0DCisXh7YFzOuhBhEIQg2twDerrbpw9MtbskKhb3lWVCJOFzuwNtDbucOuWZQt
jQNTzZN/OAfRlk18s/T71fMX3hnG9M0QuvaugBmvPRs0URc+nw1mbam3Y6BKjFdqT/hk5Z+9AKnG
iiw6HxVuLd1MWrmF1H+mncmKOniIsBGhviJgcnWNjWaXc6pILQXG/WTMgPbLt0pLn02TPjvF7817
IV0b8IYPrFjLAXnB2cN1buEY2DmZSPJClf4S27dnB7pgxo/nRRVACuFFUOa1zALXqepePD4P2EyS
wP5t9jnn4S1frnCtPSv9F3AEF1iJUXwxsHZbp2dIZlox5dgiq5mnAGeh3pbsY/K8A4gb6YFzxZog
plsEMYehlxNj6fSNYSk+Ee3H3OOmDIKDWJYUv3llVu7AR7Sq+NG/FPrRpeVyGczre0zIdaujYygr
mtik9vYdBYXTlwlQkL+3174IjTAsLrWvg6C+dwAE1aUuPhSWEnXdgM+Ji5PBeFfIS3p/TT8LSwr3
zgV3EFqe/ggAd/tZpS2eanh4yLlbUGCg4J4ND9M00ifTCSpeMgaK5Wx3ht5Cgf7N69+riK7iW21k
w8MUQ+Ihv+62gBtlOcYWVNSFaqRyx8uLkbX/fUvXZwcYNkzxvbIkIslBY00kqoRp7zJzxmNcG6g1
olTtsT3fS2f+BeaMEOpuZ9bdsrrnC4IOIkQD3kKyGbSdYOCpJ7vzlz27TTb1Mm8V68/IPXau97s8
mBICp+LNoIot67noSXKywUxJWsk5mbhKYNHCoToAJiNDvQt0R45CNXz7uAuqs77CcxBJd0rTjSL8
Pyl8dSoOLF89vicbe/G4JM7XOBYQnI1OeuAnqZ7wbs6ILglCqFknd3I08Q6OeL12tG1HLU8QXUQC
4cVTOJtbz6apdBktARQPyVAhW5Gcb7veU0Pg9o2UNGm/nIUZBDvpXl5IaKo+yIqDgoXOlQfWqrri
/1gliSugUckvgD3cplgsRUxMfpK2x+9/YpOkCnfEjmrjjKWDSEBLvOHdDijaSqh71tQGAM+D63AN
2cL3+32qz4IhxZKm/z50s9XfC1CS3E4KCB3/8dRsIvtsxWmDF8NAiiRc5KfYjnm2csG4AFQcUjQF
0ELXAogyJzKnI/Pv89Dpj4qrnrCVYiUBjxNVeLzYaEEprxxmPQNkbToECXTf8R8lDTFOs+9FxLMs
bVG0LgM3Zp5Wc02el47fg1FkZ1t4dwH+bLsxxUz01+Ez7qqPh7fuSjpeado6W8txjbWYfOdsnElp
0vv91XysfpfAifn4ajILGn3BSsymec8jV9CpdAxKmncdtUf3qU0KjRcm2WpMe+GEG1yUZgnjBdqR
BZEznXR6pUQdsOB+/5M3z8HvOMGbK4Y4nLmeLMD7yXby7Usas5He9zoQB2Vr1mNrAzfCB3NZqMGR
I3AMf7Fqm0N4gGGfrbtEzYyw0kaiXUcgN0xSdjlQrtm7G4mcmNij7Mr7L6qCuM78kE2GYxXlc5R3
T3JIxhtinrhscCYJJ0EZ78MZN808OV1e5RtLiKEEGveFgR+1g8ecWayjK5chJnUYhfIs/zy0ki+5
AZjg3cgZuTDSjvFR60puyn+mpics5GcDdJFCx440ya7Rj48D49d1CQ8Zp+UYG/jB4+st0M6PpLKo
zj10B2HAxapLCUSPGes4wKz+lJJhBBVA5n+OU8WK6bEUn018keunNiGWg9AXafPY+HrgtX/nGXiM
42l9Jp9bz69nrZVkeOEc0vzST2OG8Vdt+hDNPTob3A2XNAsY6XbyOnfM9boZweGAFwMwKviYmc6w
mRPI3ZbeSns88sTK5v4cbzp36C5b/hvRAuc3VgUHa2SnvJFG9UqN7BO1vUG2gC2xXMj4UzRXnoc9
hCzNbUcJMpkP6Uhig7uxaj4cEZNpTxPo0iDldcf8UtXdNIeaS2mpHN1RLhHTRlAJWHxkDoIQTjzY
ubjcqjJhyl4XT1TMhO6mQ3sGgpJgqJjg9MmaHF92g2BVtnnpSnUZU6aysTAHcCtmfhF30QI3qHlL
oReKCOMpVSpantPbCpSGtGAJfT/pp/mKrJkc2p0tRZ5KUHkDMFUar7UfhK1IxQ+WFv+eJXHCgFjI
DXHTadeb7II29pYCxvPME8yh6ism52iOZmXokHcj2Hy5LEhH8OOByiMAR85EJvoow7S1CB4EpA5P
YrDrPP/uupH6J0J3U+qDBaoz9YlEjq0VW9dZ2rkdu2zpQ0mJPxeixF1MtlIhhmxtqQP8ot/uFYi9
NjfF0hyLdesqPJWQ/AHC6/e3PJ1AYI54L/e2HxAyTUvlzsPzXb9HL+Vh3Zdm8nGjt4s+gFCRzThQ
ztqC8rq55a1v5M8hqpEDawidJpfptNNeW8vCCbC0TaqyFKYWNNsyIa2Y+jIGnhJkTVSF+1loGoe8
ozJWDt21+GpMA53i1ynpiiMCrQqICCePXZd+icrLf01FJ1p7dtLkPqNRDs/nwiN7nP/NNVkrWztk
qwypBZImjq9Kavzhrd/MIlKF1p0RDWAwUVTpU3iXY3ccLKZOZkP66Yfc0nP4OgN3xAK9tj/z5h8V
YFL+FB5pZAfGh/NkWSOHbh6MUJoeehFX9OQid0wSoL49SU1hXxn5ln6lZ6m7I5+4NfxFEWxWuWU9
wYgb+svKLCHdiuzED4pGIMJfj3IcwnkroTwRCyoWeeay/uCkNRcvZqm7aC5EZDbD9Y0I7ihR/ZMx
4GPMSqOQlBhB+H17G03EXJAjKblXocfb1Y8sse4Z+jWQIe5p9ej8YNW0a3aSPNPeSU4kyt56KXGP
XdqeyEgTNByQbhNNHLvJmXHgd/9SIdnPeG76tPuiyJFKYXq9syhW60cBA1ZPURYgx0Ki8YvAsDf4
z9f0xmNstxHXFo/Se/hwDWyLASls6r1OI8cByZkHcRg5P/f7oBt3O97Ipo/MegaAElDmDx8W0SL5
q8jNThStAE1+e15BFDFL6Cjziq5ajchNdusmi5swIN+xJlYC5sWa2HQ2zc7Qht7Uuuynbj5Whudl
nkW9g9VQLsQCkUhTcZY35OffLlo8IGh2OrR2dWud6/cXt6A43NTVvHR/7JxNTdksDHt0Hir21eIL
6hh+DhYKq0CoHuFTWoh42saRcCvwXfAZv4/enQUUbIO9tYEdraNhr1+jLPS17fga6hi6x5+DlSH2
wptOv2wZKW5jZgriIcNKFCukvv5d9I7R8qd7chnJerEtRMZr/1VWQtmYqbzCCMQRuqY8K3FKMA/h
Hs+213P/0Lzi9t047oD49lEn65/b2xySREqbLBoWbAY3HJLshlwqygG0HjKQGlGsNfbShHUPmbn/
Fi3YXlHxhpEQBJmDxsgnsbuQFhb/H/113XihRz8cS1kzikzkdoQ3ti0uPiFnxEpui+WdY+O+Twcc
jIGO5Avd/+DAi+xxwklXqPlSUXvMAr8HUs/65TmybWlK0UBrX/y3gUy1gBEr1IvasKIwkEbeHKuS
fcNKVWFvyQYOBYka+wx2QAtbd71J7kJ9HX55MJFJ5T8ZFHAIHRlf47Xs+KVl7yR3wVNUawNJjIum
pR0xTfAiMbRzkiebRUibF4wF1IHeZ+rdpH7//GG+3wgxU0XhcQJ99lO/Jh2JrzWi64denQ+1PyV9
nf2KJE1dmYEsLyZs7nBUaJtUvrXtv4NhYXPKub9nQkT9J4InI7wVBqGQLUeTaYbKfrJLNgx6ug27
Vdh4RZj79+wGq7Bx1pOmXWYUScHtO0dpucpSTukBhqP+JHEHEu1hdYgyNuFlOrVNpjlm8gsa+LFl
VfZRZodR5sOR2BazDK2LL6EFkgcU7emKulDKNE7MSW2cm+FFawbDYH5G+PrtffhT85rEqtK+zZYm
sDS6ASz+AIpJ8oihDRJWke1hwfJCKpNRHzO8N/7gtdY/dexEfkunXLdE7ZArfZ32cZDn5SOUbo8c
xw0/XJzMuDQVg+d2mSjawJ0q3rEkf/I/aiuGLMOmiatxdoKMW1TGlcEAdk/6HoT+ot1tuH85wXbW
CZw9xYNOQB1rJNxMxhKRKxChmkv24oiq38LdIEfwltD8RJnhm6m4rW7kvq7VmLHpVO8VEtKy4rwH
qcZ93Wf0jjDcLJVhGuFnJratnnL7LttOfAdgjXSUeLdCPCs9PlKB+kzeiuvfRzkJSoCrTKP0AGAL
NsBLVz3YulGO77nCiLNEMzyqLEZgdk+QNoog9lDbYyvalG4F+WXSUuKWjPSzqdz2N0PjQxU0C3TW
PRQ3UHm3SEkh9l7vzgpYHno8KATUaIZXurOkefnDR6ALrXfjxDJeh+w9TCxmG4kChffYSpl5XkdY
T+ztHtlfrp+aOYCYrGPieRMRYTGgiLWswFvgJNikDDjQP2z5FS4vWbDCEw3sfN+ewEFB0lRc9OqK
qH3be/YAThoE/Y7xkqwVVVyTv4btAfJdqk0UJ3D9Tq1mYH/4z1zRao6IN4xhVCzW7EaCJeMNDky6
wYcNJuM+mwBxZwLcPWJ8fQX3F5GEc7PN+AN+R4oZCK94WzUFoZytOfCTKgnAKY6JL2/wnLCWDdDX
ICFFcmByd83vbBWL9UD3DqG15jsoin2RuSUSsZexNXe15v3sRFRQ2POiZa3yJxbcRVxDckcOQEbA
LtXVXIopXzP0DqSW4YjuhKGwuGJRYiXAjmbXngC8LlpNur+vHIU/nYrKWyHUbSvo/WnJdz4SwuUE
g2wQYB/9y3cywyOcJf+YaBVVZHuBTgfaJYnQfmk3qgRgIva5FPPx3krHgYu1abD727amHzbfNeEJ
5Wut1Hyh2YXQxzqlo2HRHI8ua21t8/OR50M84VDR7ngJXXqvBJeL0uIE/BMsD9DK+2RuFZWr8b5E
tDK/AIYXVN0gp3ead3EihVQpIZnW/WR3ycXvhJuFLuJUIUJdMB+9dN0gZ6sBIOr6M/O8oNLBZJva
+TtOS1xSvTr/k/M/eKVoAmRHkfU+KT+j74nqAi7LfgLjJi0Ycxz/DCa5IWdL7NhAde9D+2ToZQ/K
ob3HGaq6kUFlznIPUeXbZ7OgeeBpeFs/uaGGpFxsb47D5lQpeq8Emv9wda33ij5puCrZ5p6ABV2q
jPYtKanUdtRPWJXizF2uJ2fZ4o0ClMMyuAsQE+ELoX8DvMKBC3h48V1WY+mjFo3EtAkEhYcJrGuu
lultZKp3NtMrDi5GKMKGJTN86/4e0WMM0L+XsOmUdf9Jka5yRgcY6/CQpGHcFQ4shWoO+0yV8UBV
OZAe5fhGzJvjXXnYXdLSwli+GPDJUuiLt9HCPIqodJejUbE4H24bcg3PLfX0WAtkkn6fE2J+j0nh
Cde70VXEA/QqMXmTHwrbkbRc1W8zcOrg8vRGZsveHbdF0ZU/jQOidASdPiF0ocqtPvySJD/VHtxm
mbeZoC1vVSe5seLnhDJ5etP1gDSr3uOqdHCNuSuCacmLZwrlRdCkX8iz6sfsWrsfAlh2AwDCNU3y
S9bLJXmmniVvjFlgq4yvSJWXUh2oZdG80hEzWTUm2aLJblP4BFLIEFNaV8fEyvOUKCdR2WLJ5SBC
LDFwu/qTYULtn9NQ8Dotq5wttd/l9bd0qwyS1kE5paZR0bQtOChbcxmHPd2dD0QjOadYbHNZlRoK
54TPndTRuYdd1LfDZvz9a55P1Kp8fe0U07JcdtiuwBgF+3R8zAJiqFsgPPyXN548NKd+YGvjUAy4
o8p6YomgpzUOdqI22V9/4gegzVAVIkv+F9GSx/mm+ntp8PKwpBzsqu3lBaRBVbF84VloES/DeMp1
2p6yLTzh2Ar1LeGkrazTg0COBmOb71cUiECBoko5AKZXKPHi+buUuFB6O+OHZEliKH1RuVT8aM7m
F+2mtdS2/q/VBDs7K4i0KvQERqY/o5V60z75pSj2zHK7XWPr/cQtCc66dfXmfXg+K9q2Oi3Jof16
JhQRtFi7UDxo1g3cHdhr6IJNVBto3Iesj6/zv3bhlhSMqfMZ4qkJtmzFtWoiZ+5BnfyEnZMYm0+w
5w7UrMqg7lMOoZeJdUL8kAmAEYm8i5+Dc/cKZrpP8VUhkPo99MOYA87t62GewkG5qHPeRlPODrPu
4KGyJhsoVmuKZGjvVAYjMROCiLC1IvmixW87Fygw2l9H9LtlguhPXB/29nuQaEjrit0U9p80DA+X
BzwwRgeDTqltYLm+1saNAsuj9OVvT7Hj7DGNFhUj9D55KeSOyYFgM151WSJuo9FWBijtbVqFcJbs
LHPp6eijPtGHz4w4dpAblz9KA865kV+YRfuKA01xgn2rPEzNoMTev4bqihjPujuckmjsbkpOffS9
BQr6kCnfL9psg8T/uPO55Xw7upZSn+Mf4wk3mNgkh7SvY9wXZ2ipR5TFM2Msq0OGFeaU7GY+e0bc
qLBs37YOcUpXOQ8z0ddXtYp+K+2QbzItUsDg0uEeK9MMtUetOM9hLEO1zAFTUMzyJ14/NzNYuHV3
y0HM4Y522tSqAN/ebxEVV0Ro5KGzmMgPv2E739FVwz3ug0aMqw0dyuDnMhca7V2DI98xPbS90OWC
PzZMSiwT/VozLqSwvDOLqaR83VseiTJXQGYWO7YRgmPRPGwIK4S58Kx0hqv1q/zRTX9pPtpxijqb
8sWUhU7B6dh2JnzyL5Cd55y+lCWL2xxy7iJo6op+vUPh3SCcyrxYOISfeet8mAxwvNRFNpj2FTd4
SJoBP4jfRrt/5Y3tfqNzJGTwP3CbMb8XaTm6EB+h50QPNQHSL4K997DNG3ICPxtXfsM3TxOIdBTx
krJqWfeLCl5YdYG7qjE6LohWWUYGw1cCofmnYoQacDtjLpHJMK4aOm/PgbUGb0MRyxlunWONZGc0
DavfzMgCOP8nvVD6V0hhDELmj3hwi7sVGX1sWYBgOHb8IbJLLIauJbPs6S5lTYc8Rh+Xr6ZDUlC/
8DjaG8mKB8ezVH1ui0/4N+9tM4GhvHsq2wDzTBfW0ARmzdb39UMZ3qXH4nr0OamwWhRWjP3oY/3C
RBovVFgad0mJVp+NB5jlZau+k+9dyRnLkLI+orodXxWky9Y71ceGaaq+8UriA0FjC7p1KhR5qXnq
ri5YIROBOWpPSW6+KNnIXwLHP90rXYlZmSLd0XjyTmeM6+rMmXHki4vN5lUYLIfnWoAIRaZBc5ek
Grv8pkkPHl02e+YTCz5sCzjb3vv3xTj4LqMQKf8YL+qcL+e+bxCGbC3l5kOsy0rh+3wnM42+UI1B
61s0dya0xJgZPj+Zav0dNGvVrxwDdl+bddPptyRd/p2sqhdUfFrYcMeYVCy6XX9hCqvIk/MpcK4c
ua05/aYFXGnz6/ea4tn4uduT6PxYPVSKwjWiZYiquRgaU4zmKkSp2NPPjnmS+4B5qPwp/2F40dHi
AyWqI0SCrwYB/2Xi97rtgGI3zAH2e8a6BsAfoP/3cIzbcLde4dWV1vimIbT1MGMF/6USIUu0KPx9
ddV7RX2dS6wgNFHvBFpO1t+y4s4VoTV9p8udmj9eKLARURpKTJt6bd9IIDvE1uCTGb8LUxANA9cX
LnxwnoXnNGCb2Y9uahHUvA1O1szvITcMdxVQQ65ZA46tT32uCdb6TIejaBc1IlgGWUllj2VxA8iU
N/2LC1s8V3hVncWRtlgbK2SNwUA0joDS/2bvl9ckNayWaXQb4hiaA67KXBf/RXf7Hijhdajh1+Vf
KvA7+sfDZCn2ZCA2OMatzwDvT/QXDI0iMIWMxK3iHwkBRrogVYpnkWGXbisCxsX4/oOAKqpSFKJ9
dhvscjxbkvGZSL1QhJsNLt+lQn38wk95S+GrE307ZJpZkpAjZ8agz2hIPWVgxD/Dbz0k8vyQfDO2
geWFawBlUG+A5eWykuN3s1yO47axgjT0j9PobKfNLcxuSV2tjM9NSAHR+Sy42lal80gKbfCWP2bF
BDUV0yK4rvGGepUQ4D5ChLMzkeF0aqvxO72AkzA2Fxr6ahoIGWVY/oC1RVv8t8lQy4RpGrjYe3s4
bea+KXVtwBMTuFaNDn5Qn55FBvekUqGK8yVv2yMXjqJprG7tgZHLlSZISuNahqubCjrQl2abVvn0
uQOZkXU7vp/zKVA89tWioioNgyJiKF28AEBBA9HUDSi79DvYMTvhxnTuXTirIL9P1NnB53FB9wzn
cIyxzBmhttEZetW9yNp4o6FTUlPa3slJjb2uArPCv5YYXFeBFSHDKbuVAy0DNG1cRdZom6MiNY7U
xK7Sn3cr9L9ibenJXuE+yBC+u5W4GCeXqJNHyWSuic3yh3HFex4xBoS7/L48n8nKFi1VKVT3x/+g
qN7Y7wUZeEEhGyF2WqRcmKMPfit9bCNVkQldWNDKGV3sdnWBKRRBEuI6rZaZT+JrmbLC5FLx+o19
ycTENm0jAp3am77DVw82+jdn137Jx7MIl+kGKBkKtdmyl4rnItNm0bJskiqAS94p8PGBfTtFSRAD
XTdo1mLiWXHcEeoIQHKNKCgVU04mm+LkhmL4I5rbDETpzGe8QkrdffgE+aMxPGhCeq9OaZBMMJ8B
WZeoMe6/+j9ucDWLfGIcIdE29GmTHVi2AXWKqlePdclXm0jsH9LYPAgIQlG5dtMKRqUg3yicjun6
Z1RsxcwgirYdH6Fyz2iA3yosznNHCfkwnapsFscPs8UTGSzrdxFOQ5vfAT/8Jq/ty/G9T7cfdk+P
ztQNfTzUO66ieiT8T4IlM7pawIfWZzOzSPXGmtUDjL60lA0zF0Iyi00bp5WQPHzaWQKydaSa7Ooq
r2ijhRJiIK2s7JTDmGXsdIwvcHDebsM9cCXLBvsZwkNfAzWUGGiFYt9nzuSgPOM6iodJGRR8ApRE
XPIxLJFALslZtQqi4s4QqhSpeyiPJvOprYhZthb9NnxVPyA24XB54XzjFiYpAp6uJV508zVmnvrc
Ke9nI8wz5Ii3sWa//LVXrB1f1T9gXrL2IHVStkuNY4pdcZtQrxAUxhIylaLWZcNzHIQu+uOFObTB
shitwFiKSZmquVnQzywjCpLwtohWGajp/U1xPXLXSFmYabmNuD9fGspkpdMuKz7QxV0mTuegy5DM
XYg4qO/ArWInuNxTmb5hrLUxfFyvik/RjvgTJ6CwRCw9OuPEhLGS0y/FBdh74DlSfFAdHFkZofNm
FoUxPcNh0oJHYJ484PgWG+yrNWgEZ4ed7oSHov/vlNzoBoeGIEJHyPJ4XYtUmRhc8r7j8Einq/YZ
BsTaw6AoD8TSWVV8e5VNTIRS6GJtqklGBxDZasQqrv2HW6Ipn9yPOKuJ0nE/gvpsWdrRct6bEAAJ
ICWImT6LwQ1fxxZwdMc1EU7+R+w+I34ty2mpa3M/OFk3F/HCexnFZSEvC4zmBqoy3E4u/Nx2JXP3
5qMrXhJhnR1OiJZ0YdZ36Sm5jJetpPLaInkLUwtR1037uyfv9WP9UG6h6XToHSdbB/t1VjSICAPU
eXOr7dOesKS2RuHSACX45KcF5nWs8zYU9D4ePa/81cZ2ZpQSXb/bUcf6Y7NdYb+ZzPlf4jhslisn
EUJPEVqNdj1vhUZq8py5qy9KDlHaL9vm/UnSz2VPC9jWRnGgGzR0nCcZWI0T2Hh65C/MNzpI1s5o
H+aB6XiAnp7nETeFCrdYSPKONbiwbsbqQ1OgsEBAw+rTfnQoqVqf+k87tWmCL2LztOkY9ouAp9D2
VtqppN2q8vipur8w7Z39G48BfZSxWN5XidOIYm3JeUYlr7gETeu+1+HP29PCFLY35Q4DCsrakCV/
9sa3COp9olv0oRNpsvP2ORnHluP/FbKmKZpM2bucU9PKJnVBwndHtLWfcUCHGOLGLsVWzH5FUY4u
/M6ChV3cgHz+qG7Nv6mt2/h0gzyZO/Yb00VQ9q/Et+LqGtpcc5bPM+PKSSIoBq/AyBBjkdCzwqdB
FsojDpdAKTBHtmNC/4sTtT91KPqqFL6f+A85j2R56WkfrPSONLjsN1RDSZqD/g1Zw+Fk+nEt5e4G
QQs7GT9NHydPHjCpZAz5LyUZNIQtWcXkDgO+wi4a/9GhDb7WSlWt1IlYDvoCkljhdFw1cR1T5sKj
yLVz7tJ+9tMxcIalWi3Kq1b9zl133JyZpAbmNZFpHLz84TRLrimjTKB/4pHi/ew3+YR8puwCo0io
bDrRV84Bwz1nfdGUgChRdHjcuViuIkxfTTnSjHR7o/F/UQWBeAm2Ri0U9FLiar/dCpvw8JfkKxAS
1aeLFYUqBbZaYKd/xZbeLJgq9Zi5rO7uwOl6vX6kB6E9vjBGirPjUGB3qst0PLXMrzHds9Pk4KGD
F9VBMrBYfMFRQ0seHyi3yhUcNgrcfT2Eyb6+nPKiOLNqPDzQVCoWs0VgrT8wLNkn8yabYW77gmAh
ngCxiwmY27MEkrcC9ODipHoLBtVbiTmwzyGVAZ+E5OtXdqvOJTQHQhO8Og5DEAbPfjMV042QXpu8
+BYF2EFhHwM9lFP6it+inPEGwcjXIGVIaARioo3RpRNRNTGlgXNShZdVoW2iP7/d9hIuRJTW5doa
NmBvyw8VSXfInqXVQRtH/8e1Ty1+5EZ+l+YDxnwNJ73LCmJj2a/qOzK9LBfGEse+64r2tyCJbbmw
M2uItPq7/V/a4lMKVX7r4KgCm6NxxJyC2HtGITDv9xbdGkOiLmN1u8jI5RTUPaLqqSlnUxwWIw9z
1Al39YuC3z1Z2b5UJNcj67poqrgu+OfPNLhGbCF4fhzYlXY2HbxXnBn8Y5ctaa+4RfsW/4SBJ4Sj
loQ873Wxcz8e42dA+wewp8b/0e3GcMGUs+zo4YRAsADjgDtipA1+GXvcNyZRHFeXbsTdNjcNOlw4
z9YVHjEvkEtVlx9QFSuE++vW/TcZ51AzI1fZ8dWel1YuoxUBW5IXZ5YEyfqbJ5biTOXxB6mE60y/
Gj6iajLy0iEwF6x7w6SLkLhs9F5n8NqyNjRoMw5YEFmg2EGUOct9BTcBDsHmYJxlC7rS0c3XtDIx
PRUE2LC1vVSnm1g+ra/4VE8UR0FRs1bCRroDuob0r9gReSZCtwRM2MJhs5SI5CqJlzKhPIDqEBL/
Ex9fdiBY9+Jd4if5Wn5yopf7CCfUdkPYnltizEHB+6XppWz6UhRnA4Bzgf9/TFA1DXlxcs2eEAp3
uHp70D7LSR5wl+H/CeZ37q+EEyNsCj9vvS4ibp3RZZWWr/9oGQxnGA7nMFz8u3RcsYKCmc8eWM4j
AUMMWmwcrYsdnVUDbrt9X9X55+9RD7OZqVirnKWJkFlrN3B4YvthQSEbfy5sESveQSgA1CB6xc3o
4sZ0prN3ZSUg/g03GN3nWQ/hPbgkaRKcwAUo7AmwZDAv6Gv//3qwi/lCBNXC4kZ3RaULfu6073JF
+cfsqiYtUxQaf5opkdLo9vdURYf6kN/O9tp7ua+Bb0QeGwNQ88E2RqaGisOwiv+z2qT6ycENi0PW
B1zrHwMcWukMgSxECtYgS8qNZ9QHfNn5oI06X6+4TqKQHzLQG65VdTwgknfUcG4/ojp5sng+tEEM
tR64nNTvSMQuobCfVFpESOQWCfKW1i3F04pISk6Lilz1Y5sMm64L7b/yGOQadu20Lqb0eYD1jUur
nH9KgF34TBimlAq77DsxxRxpbUtJfui9hVsZxsbsd8LHYijq/S+uR8FadQJVnVb3Kbu/6f07uTnf
lyCRcWpkpzK0tpGQnwiFE0yGv/rPMY1OiGFzldaAhTOOghezzI4+/EEVrpnSdSdSKTlish3t4MU2
caZeDrZrbFNeGNiWgVajcIsrbyEFzq3tX8Vy0icncmXuJE7ctUGE+G6T1Gkk+53kqrf5jSBTqdO2
fW6/DTYHp6teBdvrc0iKk/VT7t/WEhg5ivjI7xNF3tUHkfjyyTpH/vcHkyFMbaP/o9K89LjR59HG
BZuZUSgRBx7y8wLMO7m8w9hHyETGCts+BQygu1DOAr7unqai9xR8DCnvO8E/o0qxNDySWCUTz0Mc
1tp8ZpBtqo/X7LV7LRPiSNQJbmsAyKxCettFfC9Mc/SivYdqto8jscglh+/oXpl10goCooQkiKQr
MUmow5OWUNs/mnnWuWh+BmOH0zsOn/TFnCOzNzemgVRKixR3HbC9nFm13u3GzvAtVM6q/1fPaVk7
VWXJ+vLNRK3CzLlshVOMrBTbgtD0OR8f5AflnE/oKGMR+nc7I2Dg9vwvJJsaXu9k4kax+jJq6rNL
Dn2/ysEy6jXtt8ryVzPeojdo9b3R951UJDvMCAuLWDZGa3jp9p6qTzpAs77DL52UtuucnXUF1t9J
9a4LkpdEtwXvXtQhbo20MTxD3DhinoCSRuUmpFg2AzAhEVWuS/oj/Mq+i4mTFCupdfadUgr9/5Pv
anE2aQI3QjndKaaMOK6Zsjc4XGtas41742qhr86OMlWLnQRRadxchShsb7aykaBDdiEu8KpkplUf
9RsLQmeKuXkmkhOnpGx3FDLx+Zwa/+S+N2DzM0WngcOnuwNq2U5ScFTvaaGAwhMHgT6fOyaX8llU
ZBN/qACO0s/jGw8ZByOO3LQPrEA1IDFiNaLt5T18mcCIjQLhhjSpNuLONX/n3noyAE7Eexp1gpRF
j5V6bra5qCX3R5wAYk2zW3AbSDdbCffWFvYeo/K4GkJ80rJmBRFSv8BaJtdfzGubbTDILk1Uh8aJ
patzYOMqhnUnNMAYWZQj7Yi9+RhwZmUx5zGukEDtJ5u3646OZOuA0Sz45hIjeTJNBTvxwLRV/oPd
fwV6btS4SnrJvQY9uuwZe/cryH4bsTQQsRPBz+hR+kpRbvpNHe3PutkrrKbfqQzvXGCQpUfMgBUz
/TlomseKrLQra/PQPx1sBryHBT1T8fGVR1DUzGfCnEDF3WQmPoPzPJ9QXvm0ew9VYNa/NBos5zI3
f5FogEd1jKyMT20bArMOVix3aevHzUn7PtZ/5woje66xwm7knJAhI8nd/O4m17egr4L0DUn15xlD
u8GmAt1as0bwMJBauDtwJ0ocnEpH92SOK2IuY+tzbkux7AMREcDfy9IScdEguHJCTdNqcOvBQOnV
nyoFGmURByI1Deh4B+r9+8SThjgPPFMJXSXakqyZAjVunPV5iEGB2Q5xf21NgaihqlDwf/f21Z4J
VbJY6cK5RM53C0xopRMMw++e23JqXIfjuDOiFM+aw5K8av73FIxINJRilLvAnuCs9YWur3MneqOq
miRXeljzI4m6ZalfaYv1+xGRoSEdCUKwB90KpFNjYGOOeLFOmx67FsWoFwyM9pXYxhre1u4Axvu5
jgQMeMFR1WffYYNZg2oJ4Nf3jHF725dJn03lBaI9tToaDkyo3XDhg29hdlnPvJfYbOyL3qwoX9oe
ELVWxVXFVQjznHjIxMT0FGeFL707ii0rIi4ksicOQ0LmiJ9fsvV0cGTxyOFZGMqKDNZtXXzDAc4s
dAm+iso35IkVpG1G3zgPd2qlusI8CXCuV7NcoZpzYMFoQN65piNDPT8E0+SPzXaKKFy+Fu1DO9t3
M92D4dxVr0A3uGmzuA5gUK+BTj/5+2vabXMrFnZLrXGgwh9Q3nE9h2A71LVYSX10WZ2PTwmGIRPB
8t8tnmNrqUXeJRaDH0mthT0Uigs3w2dRuqDm0z55XulagDjt2gQaldO0aZQeKXWE3t/BDYqlvvGB
MzYbp+MHWw6DyLssHYvs2rmFje5a8MVitHDaWblFIC6bTWgFS3QuFBQgPq8MqRsrtFtQIQQYCZid
LrKTF2u/8pOaSQNOZSBKJ1xfOyU7E7VkR/gLVL/sqRm3nruwEHqOSgTHXbuTQ4LpryzWm59YmINQ
mNIhPvIGFEDSiTWXUya4XfAcOCITSBfbDHNmvAzd1KCSo56RpMXd/PBsRTvLa7i2/3l79VGFiZA3
Dxz5IoXzOUWiRmFTjxlRW8gvPOYanNFPCIOzHKgWDkkfI/l5o+l57PhmeBBa0Zu/iqYD8M/GOxIg
+s8I59636zQtSTRo+s0VXdw/qpUhjGFmPu9hBJ3Bp8+KWemVcQLFsF+9udaJfPQibaZa+lFitVwd
a4YtwmUEuBagHIibSDxuQbd/zSHmR5JCYeYyXoVZ5Bl+J9H7/BbaJpg2f4AIw9md0KiEKZBeTt76
zD1H7I/5OtsOGFxnsi6Lvrgq+3FTzUcDpA29PpgI9FTbVWKQdU7aZiYTnRL1AlKLXDXGwBd2yphI
nSy1z2Zz3h2j5xoPLmDy6XA2gn9PFwSaVxtuU5GTR0V3CQ+8kzPg3abaZo+lhpysqN1FobQljaDv
pqlGEzC6P6oGwQ5P0ekbx8epK9GVv97Mt+277rbrkozPsS+BjQRTyqiO5Dg15YcvxgoSleobPIpD
O5AqlvVBxRguNOwvvO734pChC1Sz4ATfRUsvCjGurgvkY1FQXr3lBeeRgACSPWv7Qgj0viG0oUeO
w2tmXgTntObqsMYMo7y3PyPZQychLSlFqcTWfxlfm2daz8yqJDImAYCf9gaeSAqAbdKSXppd4nzj
ExbSMvb8BWb5NYwlgF3gr3FLR7ZfL7iQojK636mQ078QxQrC0qngR/ibwUHSOgPzwolhYwKfwQnn
/WPxlGV4FbfJFujzYWU4IQCQ3MyCvAcSuygPtZB7j2iEGwna2sxFFMYJGVMn4VCdJ491RmhoUEiA
qheCxuC5q3sW34mkgyKLBdRFYXlJWPXKRx36IfKswfALlsRuMah9v5UhcQqFmONLM55orPZb7w8o
5O8ncOm+rGJOIhYhH1lqJjcKuZlBeZ7KHv9GPd6efP4La5hBIr97wQWlCNL+tkE5bYNZuyxw0rWm
qCbVC59dAjnzXMkCM3K351nqogd18o4b9AVZug+Xx4816fDnUitfk+kFNYiqg4fs/sKM1Hk0befQ
6pXvVjSAh53uMexVJ0n3LD2nbvU7sKca0GUXxLl3iI2yQ400W04v1gLZiA9dQ671nIz4Q24404Wo
LiI4NqhzsqRSyYcmqiaYlJh3hwM327njrfBZ9CV6SNoko7KIXDdL5EAFQC/P7V8KLHpnVfJcy3oK
K2ezMpohL8tm54o1X2FGIsfphh5APOVCyVwN1YZWtOlA46qMrcxGre85c3Q/4Ua+qbXiCcqhzWaN
2PBSXq09wN89OB5TTY3Vi6JPKB5TVd0LTd3FdBaqEmdGUjFWb9ANOd9+GMUk0GyZwDxDlteCEkSZ
HEJP8ReDSXdSZ2MSCbk2RnMusQJFyRw3nZ05ngvwmLtuu0Obq5hCboGo9d6xnDK4o+86D6nMhMM+
jEZEPECujVqG0U4dLWJJggWPHrjksFref6VdDr0nMWwpBJlpZKllD1TFOb1c1RsS91sgXT013QQP
YuLzEnjCTKCSTRmIEFdiU1vf063+DTqrPFgOub3o4MGVv3CZ3qZAHIciSg/8IE0AzKL8ZjBjMFjO
90f1YVu8UsLk4x3BvWH4Kfov+WRLyJdzlyiShlTCQ0vzQG1BdxmNQu8xCWRSg+LvKZFp5W6U/1V4
5biywRZRXxJ1YhhkX+rf5DvdzpI9Kj3QV7SCFnd59aVsJFNpT9qu4iTQQtSYEC9F3Go58py/vZfC
EbFeE+4PASfeq7OiXznkLWGiay82GL4a6mYKKiyJ9pcHQt+2BUXURrq7qcJS56VelmWHXC+JRx3A
BB+AcAG6rZ+JGgZT9UQHvebJyKjL7YGrwJbidmO3FTJC33mThXQKZrfAFZigqXhMu89kGCu95eMO
5GwpyZs37DRdZoK2Fd1nhpYv9y1XLhjFvoQGwTsxlbkTz5MlAucWEjAWVHbJO4K0zQ/6O+nAZmsz
gTTxv3Qs5U5z2neIPpokLrehkHYG64IzRw+sx/XC04PJzg18uYIsSMqdqGLzp7XrVPMIQQNl21hL
mEpHrXRk6QLf+X+lvFeHSFkAZVzL2Oaj/AeZOPTDGN3ku9Y93vgkQaV8cim5LORjQWsszMavhwCi
3v7S39230QX2cc77rdwWp2LuC5ZwM7LTtskV7sxHOuvIJCE8sMl38fLjFOkGZkfFb/g7W3GPrZLC
ve2aBaCKTilhcrPPqzmDhjKf4OX+/OiEzPERdB8w3YFWvAZ/WAI7W3UvtlEJYFKfnhynbwPActCO
VI2DFx4B8+KfRAdUt12QMEOM0j9+4cZgfwvjfpI0zi8aac4TebaQhgHU3SG1X881GbbkjJrj9MDA
dc359zZTCeEWK4WDRz3tJzpMwEzdyj5LwCgQhtJU2m2OqEd076f/9hXStqwR5lmAYxTpwxKO0TG+
H/CAyxTvyWTUikcgpPlZMVIdIlgqNVxvVwGm2PTE72rqrm/5M5CX+kUMQQk6gXReLFvhzoTK3kn1
6MkX3SbZI2kRbvmde+Ns6vrXhJxike/TzoTUOcvT5DB8rm4tQRCwnXAAW991wDaplTduddw+O03i
9+K2JnDI82BwA2Q5CPxPcq/CEQgLgRAjEI7wGLMXlVG7iQlhDg3OG/AMbCKHElxGr5pB+1GLPF5n
xw50yc7hrEs4C0wzRYz0ZNu7DcEHddglIlJ2C84RQRPef+nlp/PPxLODlB/MAe+2DR0p5T5Of/M9
MBZLOCRp5QyZPnP1trHfuh8cRhHw31BgUJ32u0npuCu+XvaUFpAmnk0PDNtJSLnLEUN0LWsXjtP4
fNZgVDmthZ4CnqCjRwjECRoZNZy4+ytkM/crZrUJeWoY4nqgh9YAnrcKTF91pOq0bT1/6XOoE7HN
HIypikFxZZXHoZGTQb2NepRnrUs4qxWhTCxv0O188jcDrlogmo9br07Mv966BCuKs1JTjIVEEOBq
kuX3W7eEq+dRkiEooZRJLf6sQCXXjUvYOXElT2zBI1UAGNTSU7vtLyZCOziw7TnGtv+tNSIKt8KQ
apv4ydM4lcTbCML6ww+6NDCvyt4ksczHx9XJXBzTd4UicmOLSbahVmk2y46GSkyb/g1MlMax2hCM
AhfJK3U/4L8sm6Drd93joamwPxTZ49XAxUAXlfCqdCik7sceAATDYohN3BscW3adChQmrJcoCvvr
6llxxoQmSp/sXSsQzvPOsCpq/rudBYaGlAB+wAydj99R3F4UZwfqTU17onizio5x8rkKiFkHu9k9
WyO+VjVUe9pJdYj4nMzqFWtRID/IUxeH9WNTi1SJW8WQ+s61wfHl9tLPNpIlI2bRSBCFqPdJONrG
QrkM08drbQF6I7UmbNRhq3AhQculYCgiFWStJFrCTs7K5hRqi9XivcZvuJpNOREURsWiUIYoIBph
2zTqvSH1lDxYrN1JxQKXnX6B0AkC7QOr0aE6dq1WxwO8lLpH+F1ujVVUbYDf3aD4Cddbo3A5tPVj
Eu/bt+dAlAgsHk49DAeKIS5Q82a6J+gsoDPosFZYRMljPmEeWFknfz0SKJYS6Wk1SDtx/KRVj1tx
u3AOlHzdZ3TuVwvyW5hZVAfmm0uNmiV33QT5RwUMLfg1idomfTX4kGk2WjYRkB7NPmJT4ya8EDXy
xh/oZt71L7IstBtdjFpuoiJW1E8cRjnyO9WIdTXf30Ra2PtwDGQrPLDUoJ6L6UQJjwYmsHDGGHp+
f9DbN3FLMUFdXU7kJp4ofI12M+PNoff+6MNXMe6dpBu0yDZzGa+iZnFXMLara8cxUffSFfRdoTgJ
p/+1+NuLcWmn6sI61CKp1SOKH+Ip+4+fz4kEKFx+ZjkenB+MDd6AsHTLW3OaozSLfIsGJA1mitz3
Dhn7uHjsB9OuYL1KKLQto9Hc2gZxm9sjR6H8RE4YXLoSJaHRwoTSyZpRCaT4FZsoU2EJDA8RNDJO
9WHPpjsnZBSmZBqM479LjhmrxYoYIdEshjiT/qSFTTFYDsiiOcuWc0dckKZmJIBUpOp2jGc5ab53
lwSoN8Zl2K1pUEFy9SWWF5ZgvD7ScFHWLn4+i/+POlRR/KkwXtvtHQP4FU3kulWWfbDKFQrZ+kBR
3041Fp7l+UbjwU+fYkpVPhqeuVFQiMMawY42pspYsVlCVIEDXNWQq/yt1moFNzenAGtzi5zc+sT3
EbA0BxeGG8Wv/B6dxXNgGyLOxBofF7yt6fk+DAzgipO9PtVPzBBgATb5RavUg8CSKAikiVIytVR1
IylmrFpiLAjIyvGyB+IAGnEnOisoRF4DiuGNM9SVIVckLLM5zC5c2XTjJC6UmnmaaRF57a4AYEJf
vTy8fIMzc9/QKYLM45yYkYKSCF10bvIEVYInGKPzqMWoswEPO46EFwzlhkdl+KtmJwpJoy86fg0s
GM4Fy0hKyG/QK+NtvEXxsvHEQSyIbmedeYMF11odAjcnZrTLYO/A6L+vEykBKHj2VGTaJPrAuTz7
i0E0HFPvtsLfC7/3FHMoPIes07LoDDkpc4HZZ5j6h02jMX0lIB96t/a/LWJxxpOa2mtHcxG0gdPt
OvlZHnIKK1DjHNW8nwa5XpeWMpM6Gb1I/crpK901mCi6qOSyNdn4RjjlcjUm1mGfvyCaOw7D8+X2
uVLaJB00Mw7DOlFioRpBjiPo+2hNawEwotMQihqMttWn62lzMcc5cTXRhFPauffhCTbG7B4p162W
2YpVlMLlLB0nhFBmped5L8GIPlrUmdV0B3ShC/aVQNuB2uNHH//QORAE1zbJrNEBTL/0Dw3jZVh+
w7X51r2xrgVWsKlxGbcOGqPYBCwpB4ulMyjgss1akbjDy7Du4k6Ga4zatZtQjSCorj8g5WsyuWLP
mf4lIzq6qku+xuO+lwpIXMDYwPbNI9Dgkkzp1Ff+W4c9X894i57yFHslQHyzmqVzNj6KFEG5VnNO
IOkdoQgBjOP9VKNK4Jsm/h6j8xK83paRFYMLJspWxmhoi9josLpvOxQOdyOtplfiHzGLi+PK7IWS
J8apR+CvyRiLy8iAAQmsLpm7N4/v/5cE5/qN8ocxDjzsj8pwJ/ufN/wxdCaBTQ61XlY4sAiv9jYO
0+b8boDlIJBGUTRSLmTte3kXMrrOhR6NEvaOFzpSKYC5JCjm1alSL2BjZcQfn57mm3P4k3ZYvSyF
YgTf+pkhw3s1XTtWSkeJOlHhljq+EgKWJ4M0IQmtbrj3zd5pt0/zQrNI16USc8AZ4+3QfDP/riIf
0KG/2tvom9tNjg3EJP9hHoa0qX8X2TtLsFEwFfEvhtjIjLPmrfnOpl5JYbN1W/tXCDI5IL8kI/U1
vgw+a27v7/I8EZdzNOGsTFZfjzSpWeAwrLjEUUv6h6Np6kJ/DlymJu+QS/9dsaIUJfpsyGL8xIPh
he1cexfXljvKny6cOLZYfRbguw85U5xjiKXDOuX8cTbdgOTsBkDnn+NZkPank4SBzGkaNyDLydWY
AvwGTLgRjLswg4EuqE6V9FyZtRLmgQVUQ26kuRUKAAxXtN/k28B75mLyNMm3vJAN1ieIQqT+CG+l
REg3ZzDXcf986sCInR1LA9+QpwV8FKiaRp8L2A7MJt8LFvkPfc1ZRLbExSQNdjP5f+gLQg01UO6C
bXRlVAKswwuPwZSWZfSAG3A2/MkGDoSHQ4BP5J9eyEsqqeYK3/Il3/OI7gQ3nZz+3ziVj4RYrvyM
MiVO/I7SwLkkRlOwFCgWt/uyPxbN5r+RXbwHUW78I/uMnOPuaDjgS+pxa5UCyUEp/6S9poGfADwe
PCAtYl/C0dLjFbGNuL0N9OjzO41GCRAmcTjqwujqITNwpOszrq1Z6HUJTXhDX+krkWHaSZS7WQ3U
6WGaoLWPqW0aJzDuJIDNpopEDniLViKqDmiPdBP15ZTnV7WtlN1Wkq9p5yAQfnFQpHV21TZ3Fz9y
5poauoido/Gp5NPRyfgZ4Q1QIefH+Qm0kIlaN9+5RBaaf9e7+17dEMdMUHnCtYk4lGFdBTJJQQHE
yCfQmXgMMqPOm1p3rgdPqyQaNTjMi0kLa/e6ubU6Yqn7ay828jispq2Q9xQ8amtJzTXdSEGZWPUg
Da17YvecbnV09zvAOVoKTLbDN+kuEZ6R6skc57L3Lp9PFHOov1tzgZuz2N6DXZ1t1gr7QnKxS1pJ
Pzids93bcuDcLDZLgDqfvMIxHldLzXZiqcKZnZY94rYaVOI9d1pQGPde+De8j8AEOKa/hsw0ePZk
PgtGdERrL3cOMZhSJgYiMVk1MnY1L75ZJgXTWoME7iluxvITs0NaUkppNi2spPJGfUFZMKgfXggd
szfp7htUGHSg+dfqLheGqpf9n1uP6sYsBkuMVHJ5pgwzU5OitViESfIrRbydVhGHHmzx7NXwnUgx
kG6C5UTnEgQQOUvcGORXkd5KHsbny3nAKS/g7yk8jxKCqK7gndTLWn/Jdeb6uqhnhwH9Kc9oY4+M
JsP2SVAgIfTjlycSgZwa18dFnJVIZYk6mKKAwrBJ3AiipDX3ix0ixf31ud91GKZ28N7guCGkGux9
s01OdEksUTRVeewIXlGUDKNOcTGqiUip3QL7XkZ6b6lj01XkzBEXDnxNFGdTqJVHl9QCT0aJaMkS
G+d2SmlWEDPYdeU+MmsRY36NSLHlPt21vFdZ6WNZDz0fJ1NCRHGp36wk42i+vTEeq6UgKXLpXBLo
qKlpVMpGDYC2zWyuMcIpHos/6m7Gs9IuZFetp7GF3azcs9bMTQv11mRyPT5F5LqvGEO35Lkarxk6
76FM79LW47M1GKlj7JX9VXGs6YUGWmZ7C9acLaL5EJ17qQ/4V4o03/uPCCU77OMNW8hwGAlYkKy/
zSDz/gVIW06VuQtB5HHXH6FoPLqY5/tyUhFbOgEisJ9ajcS6a3DKvmBzh/qUVZ1nFGe2iAhPsq3x
NjZP2BNkkdFiL0u5n8dWsH3CZS8ljCzpVxjAIAGCAWqOosKIPapA+UOWmbv+cov2z2JqY3bw/SgD
CpPdOS4DeHBJXENjH0tp5bD3f5q74Gz20nC8YDEIBDhiqnhQs1W6LnfW0r047FQXayk9mdZufOpd
kv7ZH2Z3YTGMMueVuSbcBku6ar1kC91U7n7HLFEbUsGa+qcdFvS5QGMn70wFNItRwDLv9m4jKbD6
jQTHQVfj6fNfguDa7S+XIsCXyiNe1/T3ksYp6mAeWNgyYWDsqbrh8FDwxl04slnzkj9Ja3pFW38J
wmAN9j9mcntS14QHuLKvbJnDrk9pipCUIf/8bGSp7VRLyLTSAk/VkrXIiSkf9g9u7VMqIRND6ZFH
HK/yGxNJmpl+se/3mmhu4UIEgettmhxt9RUAnFdnOxwYaK0ZdNQC3h0Krw1Zp/1duIzFnyszpINz
sr4NQ65UY1ZVJhxmAWTlaRbsCxBQyShXaqZJ8FicIWCfymU6xMSdJp6aYyxO6neCdNPjcZ8cpzLm
B3irBJKqv4z20wM3obWikn48Rw+AWghvzt1nUMrG7AtRQPVI736xhINB0rAsf9u+DjqAb2SV24vR
MULiMF5WENZCFJmYvnD/aUKxwB6u8v11ZNatjgVPNtFGfAuEWcvh/hCTiuKorkKg8GCZp4ky41MP
sE8UOJzmgA9CFjTD9sWIJtwg9H0d1Bio7D9UsvqG2eUFXk6eOE5QbSPFubseoztAohZIgdo7q8i5
ZyFun/11rShozAPzTsSN5bUAQlyMdyGd35JIzzP2Wpdt6pOHEUqUI3kwyL6cLwWpAAHDpJ64VGLD
48RpIMNRK6q6scywMiOV1AVKxaZWthYQU/ybExhrF5CMBi7RkMtRphy3Fo2i4mVDbVec5bd9OXvU
T4OIZmedzCB3DcGT4kKC6LOtSwFOtyY9abaKUu1gqwXx4GC2eLKNNoMWm5coZEQUs4JcEuWnBTGJ
OKV6A8lgvMmtQIP/MJlDHZv1YGFw6zJiD7b3S22RwkwjWTWN5TY92foZIwZeAgaK/6JCazaG8dyK
tH4NcEq7Nj4ao8ueY2L8YSxQHsa2a9H7tp/zecvMjpXrA/n8628MPKlhYKQYnJbKhxQDGoe5BJ3F
GYaYU8K1HkUtEXyqYGh6UTt80uSonrMz8/IzFSczV7BF6VJ/ZFHc8suNvFrQxrVtr6s1F1yaWTW/
cyCzjs7MJFvLF9CQO8Wq36lkqF+FrAo8FFRGmALB1qySJcwt5+4IogPfEGdpP+Q/y58rjVEaJnla
oGotkFYpV7Ti6nLW5rtx8NE+qX2lXj+FsCAjJCWCnsTUh3DqavZLAZdLIhTpoe6aC+mgDZzCxE2M
DLHeK90GmG/PcbH9xXKOaB6g/up+oNNlP7W9yuAHt4xkaXkPo31IOjgOA037vrSQojCjYsS0Od36
zNwmp0jiyEv393eo2lusG7jZIXd8aqA9u+p772fZ9kfVoBw4yFnor6rF/0w2tjYRgBS1aSCIa7TP
4b+P0AcXlIDRf8jXkMAqjSAQBi0+91Ad4YfG+9zgD/MJ+knaQz+d9yl2P3xSQ+HFJHn62sAZYbv+
/3VY98z2XmjwB3U00IpvwwZ5lphNg9epEbxIA54ThryiKOyfi4XcBjQodZ1SHvfdxGP07NpuI6K9
MtZJsR4FqoqPd8yXiqJ4KnQrsdovr1xwxA2iFJ7tBLqwKfODAY0ohU5nPuGDwUxKNLb0Gl59b/T2
CF0XpU0ioqtr0JOZlHXaLWNJ0TZQQVNCG4Fka/5szjWKGMFlf+Nsazhs3PS4trQ9hPkLoMUMMlGt
foYUPULRBl/AyFWNB42GajkMGJPYNLMhZoG6UyYIfeW7TDgS4LSfP59TBUubrawsMFlu6Sz/F2GG
alkonuF4oU5mxIIQ+Pi2r79p7cTDXczW/cKiMElnWjD2LCxWlvdISYfrsl+8oYpxqqjprr241KNm
T/4uYj4qCtXiPX3oQ1p9qyhMnJP4n2dpK17HcV6hdti99FGuhjF1AEYBz0mi0dxSeMk5WvW+Fb/s
WHqTOUEvSXoldZhgttVK21EBqNuk4uuDRLgV+/JveZEnW59iEkmr9Yqbd5/TDXZWjO3lnIXugd5Y
ZGtRg4skO7EqN6968jRm3f+nICHdaNBtbxc511vhgnLl5aW1ANmrSYHDYj+yZ07oY2KMb6wcBiJj
ycr9K/OMRCk9S+cJtH4qjgg4zl9kNWQtpfw5TjZnTc8gVvitGUnltRH7Z6RgH4mrWCsJrn5NBOoL
v1maFbzt0mce9zKqKjDAMmRo1KqWNnNkEF9Ni62wvZD1YYhbX8+36pGTy5S6HhLzNE60IRxK/wZZ
NYWdNdYfAelmQ7nTYhhb41FzJJzAQnnECZJgVPisNzI/G6S2mgLKJjLhNtsed2r9jQtX0+GvyLb2
dNPPYqSM4l81JEH41ugQ+euYyNQBM752X3j7qFae7cgXgIY6l9cDS/l6c3ebLlaOIUWI4r3ZZNEM
P+2/DbTkIeyEgWkK4DX/ayZ2cu/EN8UlJbJ/JUV3dsbfozfoWIImZuaOBDhqr/Adec/xep9JOf8F
LVns3O+CpD8sqJPvLf1pAxG0QB8sWrCL7wTj2Q9vQ6sCn/L1lRPQ06g5mIF2TAh8l4ASSJWN63gN
Y89s98Ta3uKMs36QvNF9Dgtqh1JS8Z9vSQYDCflIo7HvKiZAN93e1lzGZXIcHtMzLL9YuG5jzWHG
KmnZYOfbJLghBRkGcUuJoH25zDnaWuwSUQ0lgWmRs9rQk403jFIpLmKmVtRk2QGNdWR/TS2Y/k7c
LdlKXNho/L//iVugg43Ycc5qTWbzwcz9vHypJhgF/c0uK3yLVxvJuE3+EX6hKVjmdkOJ09zgAh2E
GVrucwXd/4scCgFu1I305bA3AqCTecVOa21QoZ950KN8vnVvYV40UgMIi8x0J3IkBF9GRBHvIw9x
jj7DhT2sfIupc/HXm/mLdImAiLuNC4ASqIeKX1YwlU1SqLhveSclCbVAqQiUSQYD7cl0yPvgbM5Q
i4t4tcSUm5FEiH7ysTh7DwrG0iNF/zTIig0B/3miThwnwgde9+abO18+1LO1Y2Vsx4DloE0Y4cUJ
MIx+X4D028AMFL3sMwMjlLXZheDaYlvqjkf9CiW5ONXnl5TUzXscKb6dS5RVayHljdapb47IkUhz
0zn+t/zTbKEbh2J6rcyEpMWxPAVAhGW2tBNuv/ukAuebWiZuV265XhaKPDil0qAm28yHWmTf205S
5KGSwSIrPqpjCoCbndl8vv51gyJODPbQeRGoYfwFE7uYZGjd6sgAX6N5rDMsy/OIwicuFI/uE+EN
5Bv143Fz/Z7b/ZIGAPf53HfRX0CmNTJLRji2CCmiIXZLER1dnW7tQT931+WA4i72YzR7mirwKomz
Sz28uOiQkl44CtjNNyLg/OzgZOS+Ti+cNSlhUOhi1F7mqF261ZBl8Ym86yauMhmSxqmYw0bE4q49
wMvmWljP14HBrD05JH52VhJjqHCUhi+B58EoDMuNxW7aDqfT+ZllkqeQg32mlqsyigZn26Z1yCUO
THSQgyxBntdHmujv0PSFSw2bjL6jh/sWC/b8Un4jusvJYqyk2wNMOCzTsWlZ745bHaS7k+BCHMPA
Xz92aE0skgoeKMv66XoD3PBhz8+lPUCJnBN779UzWAcwOyPUm26rEzBI6HhrKWcQWVv3i1MxNSL1
/Naz6Smunv/a/P4MVPpo3AV3fnA81HgXFHDK8U1hv7U3SWukUNDNC6F2baWodG/j5WmXeBpNX4AL
8C9lGU4leksdOjMj/3Tv3faLk4lPHuJlob/f0/GA7OLv0wWPsySeQyIEnRcBOVXPB12WIxnwc4aX
xtOUGy/0qk+eRGLVasUoalfAMwoMaz9sQFlSehNlkY2DpSYprIE6nFD1r/5L9lWy2osLhzXlg54o
43I+OCTAjPnjVqjo+N1X+wiRal5uluM3AA2UzZBSmoXohyDfTyRi21ipT4iDWZLhdaJ9+ZRaH2aT
yFmH/W8jznkusawKYV42NvqfzrqyvsycyTupx1uRDkaRZDp+g6kz3/GLm1KYmBFQEZqDRvIZNwLc
lin1kZGNbabhND/BDS3XiMhCJ/WNOonaeAMP8rG6G1VBTY4Z7G1ehs9ZFHF7Gf1VP6zhDa0wSGgz
Ps3fHlIiOlaoXxIR9vACZYQ69zNUU3sZcUqEbrVlNnYhzF7eM+vWmWEsB/bcIFrT6b3BLEAAB+hl
zTYbmaTM2NPHQ1qLw6PX9RIg/XB9O5Eu5Ck84inTrmdJWpV+vvVM/A1bdYKwhqjO1QYSNBgVI85s
RHClcB/gCaQkENYB5+gWJAYOmMGvo7DJyrRf+s9RGSzzgIityKQMJAwJ/jOIdvuOWALCVD5nTjuJ
ZIucF0aVLsyUAUUOaE20f5coitdhe+lkOAbhZLmyCTXNwGxIePnXWSPMsl4/VVJHV52Um38/UiQ0
0kgi3jZEMMBAJGx6Xa6khUHdfoq7BP0LpD2KiRCurYQLIDKZGwAv4i45cPjxXSGYkWQPbbWvlh33
rTCqxc+v0ZBEY6U1/CIK9ySjT56g584NMTMoGnlnnWdtaBVze6MX7EKFgDppBE197/+EWcLBxKFK
w9uV5PkIrVHuZy+MXCIBLvIi3mN3XiKjr75GonQ6Huz9NJbEOz2tOr7ebkQGRAtMmBPbEQguFows
GNZ6ByyxMsQ6OneklxHud5uCbnSLAollQZgQ6klZBQrv/DLpHR/xFLHwFmpzZd2jEncKV9agIKi+
lJrS1p+UYpXzCV4B3YD/357jXdxTuKcPigmtFKgG0OMpAZ8R92zI45yVEiQZgjiNgDxo1RcmOEQV
rqmzxiB9HjhUbHGvlUq9xHyCqlMnm9expaVyqIPjczj8Hhv4AarjHy0nZgG1pWP0uvQL1UKTAS0C
u1rt4V1aCvFExN7tZPUbQx/pv4vCfOcXqrYBLk6DBdB1MN5awesNmPIL4zh09BO6J7KRElq7KqNn
t0ReeWTXDhjK3U6HZcH5velrWgNg2mN8Hs1E1Iigy2zOXyt9uYETDempFq8+7S1DytV8L6kF2fwS
6qTN+DmXgBuqNxOpD36c3HWD8RMGMVAcV4dOIROb/7R9ZszqhUcjJgdj49TbAFaZ+0G8Nuc+3IpT
hxdrcArw1Ci86t1y7EeTukrAQ1+pLhZ2Q3RqkmeqDnzU8bbKAY/1rG/n6ymMILYMPY50Pg3i3FGO
hlnOzK+XkT/cBJsaW0eHGWUcwqQJALry1cpzeEBbbEGJs1XmzjLSksnCcKWGk6QjCXBt5x0ZEdlR
6tMO07TamQNw8XA2321JVCy+IOAkdutTaBK9ZdkdynxXZ3wSAwZ9BEU/7lO5+fgHPZ4Rssv5VdZ5
Tey7waGXfuMB+XfHO1QCaeLLwekTHqYoKXyouz+gmtJV/Q2nGSXkfvuoLDaRdZc6D0TzfLak39Iw
ogWxzHYpgIxbAXcRjJbSERi3ya+KZBl4og2GPCIULAOCjZf13WtWmOxSNpzfF7GzLT3h9x2kW94t
TbZhG018Dt1UuQkN8idxopg6pN0/hWq6YmitLwkNRFg1RiM/yTWV0N0tS61+bDMmQunvZOsO2lzJ
ghpBJq+aAcIKoj6v37BPO1L2XZB1yR2ccBhAfjqMhDQh1MJPfoZ+u6DYoCPMS6P5pXYT+hJiJMaf
EjBVLtQ0Dl8jlpgh9EFRpmtPsoQ2seC666aTXNV6o7tliDjDHSG2lJJfBVZ+Pvu/0sr9+PaodJyU
q38iAHx+u9v3dJG8xKz5GvGLY/JNeoJfY0vtZ7unZNv51snTAglwbA0CjRu7VtdqMiokNSaJS7bu
oKYxhWf59vWpoqVDh/oAZMp2XycwYCx7iOx6NJGE06GInxt6K6aOCEvA4aGaxE0EfU18C3CM944X
i5cxf3vhXOXxeXkAQqT/Hz6k3QXIH2/LX2/Sq3oQvTJGWdx9wUoeMh4nrz5QJ7+k6ErnOyzG5wg3
T2kY8cgnFPVSHtqssWORhABa+6VaJNF8Z5S4vdnv3mjqYe+traB5DfxbHXp+tH1xVspYniE5P6wk
cf36LDo8oWNGb5e5pzanBvW8NUccMc0tpBz2xxMsd7cx5n66G4OkexUmypLV5CKDWSOt/WJda5yB
j9BHjNCldWzS8NgXU8YKhL/VPEIQ1/PifG6k5uDFE34TKYkLgdF7iFMXC01NgIkmKf4L2LrHBM0P
kmhE7Yqfs1jBfct/JVF7jKLXuknClgQVDEFiJR7Lev3tgzJC3KSitoOggSbCKHYTkFYu9xlMVexp
sKlLwxm34KrzGL2FWWRqJ1H6mIVaWUjORYSgNdfE2aPCxXU06/Lco29viU5UCrHpWBtFIR8jFbEi
3EGYX8JJZSqqm8Jxjp4CKQuBhmQZPyEBwVudLbmXigIKM9DJDpNKDJ8bmZe93lmAfR2h8Gt74hvL
Xy8jFJsBVhQTkcTq4QWG0RsWFItX7tVZwf2vFqPvMw1Y28blhklHxgsD4vs7e4YN+nUDNrSdylOt
73B8Irghp38CxWEofRY46uZc5Bl+AoWscb0On7IOpgJWzmyTNDqGC1ihWDOo0v1Rs3riZ5aeiWg0
b8WmbfL9UUx+xrvpuBBTSAP7ASNIcrmmS1xJvlZ23n7CzHx+bprVW0Ue8GKWlqcCI4zSm95bxUoK
+hA7zm66LyfYCFAf4MFOK/HwPaLXilJGLeD51dOAHA5Vf3/xX+Gw72gjiDeeBnpQ/NtFXTFcMj3Y
jFVW/c8Lw5pwiDVDPfUaP/EVZlIhkdig5nUPOM1p29R7mRaMpcYRVNFoUj5aRR7+uBgLKU7q/gxC
ASAW7XcccYp1TL9l4/dZ9bNCBHfkCzOzCDsPSkqqR0Htwu4FuX/TtD8Sp82I8IIX0BGfcFSgNXjj
PuwnJjhOghHUQH81hOjAEXn8UjVmd6toMhH3LBgViByu4rBC7OUoa/QTHCSd240NWNfmQvlC1nNA
gnRMC4Tuu8Tr7HSZyGc9mZrsYp1X23SCVpB6E4Q2gSseZTEKjCAhiiJBiSEplvdiZ/fP2MzjkZ4D
uUI+0r34sA98QHPu3rIYE3ugQYSBSvGVE9piLPnEr0Nt9HFm7IruzkLMXHZWt4iuuDcs/j6Dhh1/
MCGC/ljqXpqweDLTvAFN0v0I+h+rx4Gbw4yCuGJ2LqPP29DAg0u/rfH9UjHN2qdN8XA4RDsEFwvg
Zf1rDBZw8A9RDnk9dl0NdhPQH2/oXDuHm+/NOwKWBxhAA7lEirhJ5KOTfjtGKU9L5ApDzyPNxCm3
5Ydv6Lf8rsZTg+jEKcSlrVmSOuewIDiw+Qcj9H0LCPKmD3R8f/s8aOMF24rP/bhkeFm0KSMpyZOn
qHQIRfbGeSgjB5LO2gCUlN6bhxipzUAgeIcHnrnw/kYLKOXbUhwYS6bms/o0hCAfwCvn49p6dH76
I0JfGQRs3M95ZGMySV+wScn5Kn1MMmyMYyOUXwqDdISMlbLYLhjLuqjMzgaUyCCFQV8XQqf0lTZ1
K3AkRHC259mx5G3CRdpcwJOhkjopfURn3a+KLEyKnmD5jHARP0Ctzye5TbxRHx9jwhuZ7L6fo+GW
+N3GS0YlgKC1Flxy4BWyWSCK9MHJahmXisixlF6FMFvJ9CFIKNEd7dCMkpzqCQTs72BVRTO4HZPr
PQVdNn7Wz6xzeZ80EdSMzVhaSH9LwdPk7BgDX6fhPvgxfIim66/TBL0mmvyS05HsIyMtTi2pV0Fm
TtfdMBjE2gdwyIJ1JFZt0NxRtEZFgcvNq0+fOQ4h/aR595p7CqMKcjrTF8Y1s7Py49yTBNtCSALB
7KfCj25e5LavWpl9ysCaW2/2jCiSDjfUE9Ihme1uiyf7SXwL+idaN7TWlWwUGcsAonDwH/ct5ljm
sUwJkGM6b/hSkIrkEQEMv+aWMszHuHxvN58KGm51s/pdb0sc93Mng3bU7UfEaBSwRio5/qXMEA8c
KlRYmtqm9pjDw5QKdfqLlWdIojQ6RpAgbbj2OhQnLDb5fTOko1TOpH4VjQrnyB4n3k0r++CQP64R
HLV7oGsfFLdhHE43uzLilAV2pu9Mmmk2XNT6ptlEOuJN7pjudYD2F+f9YKeCfg9ChUuBUWVHAKLf
s1cvdYM57upi/yGAXzpBxIzNCKtqjswvUi1pEewCWB6y1MGrAghTdRdLYrnUYNBl+tYcujaHWx0C
f9L/qAn65NWHrGvTn7Pej2aEkezahBz8NubTcd24yPCELC3cNo4jgXOFLqxmXTdEsL6twGosCj3N
IPSTE5DivdNkK0qMof4Cp/1b4dFfF7SEDC8NXh1OoSdUmb3fEeT8+8TGiviF7iNbBUieA645QaXc
4BSn4RGfdYiHHkMtIe2j4/eHJ9wJocIdOuCmIjD2dVMjapSb7hJBXDu30+HPiQ9f3IxIJWvbLyKt
+roO8aBhIlcBT2RK6+AsLAXFnG4c4ikDZ9c9T+RioyWFrY8LDw+uptABOrbQ5Ri+nLWeMOVbjtHN
lRvBzRzXEPNnqlI/WonW/5U0imjR+1AuwzqDNTkOrkDWFZo7wh/aBt2yOILbeGzGtf6In1AJ2m9b
bRynmM9BIgu9KR7AaZ9k5XsMw/JjO7sJF8mmj3fqWnvsmhfOp8VLXYpdMrTx9Ye65n4+XRkHUpJ4
FlTqQX/iLue2mcBBxcozpi8JmFpGxVvoKrlUSk3Ey0/m6PxJ9KUb3cOYUbuikd5j5MtsIZ2hMSqT
8Dfr34Zb7zRGCZw2O0uo15LLCg20/SOwpJ40JP4OypBQx0OtZhO7RwcoSgwFWw87z6vkxFDUcF4V
6DeumBxT1K/YCxG11YpQyiSJMDQ9aafmSvUFv88aH12ZQ2XZZz/Pp//spEttBVnc4VHMSbsg3g/O
cM0Qf+qXGaJc7UP4/gwhcqxTV2ck4KHZrCaFYo+aE1ytB3kV7z4lgSKiGZN4yG8novsabsRuLuN/
ApaMu6a62EFZrZfbd7tBvIrhR5AgXuzSFiaESYdApjYPRwIpiVUoHQXRLY1JJ2ISj6kpXvdpE61l
WJwYjA2cgkCOPDq3/gt8Y0RRXU99w7xsAmi+QBVDaZF5yuHlP5wqE8/rhHwvtpQihPPMQmR+hc3x
9WHtEh85YcjQymlJqYhgWO+fVpLF9X1u4btWsTl0tp/mCVFUNEEb5SH8ORVFoTDRpZ3SkQxIhOT4
Ps0cLtzT+AIJrxRXkcU8uxlLw9izksRWUHMFQi9Z7q6tSOGyo6S8xg6m3G61SMi0XQZUOF1j/x7B
PRIVwfikCTj4h2d8nDjsbCEgCQ+68phqecC/inSRMp3F5wMgNboyybySvdYl7rKzMmScvVoHDlhT
sqdK93/2qe7JiaAL51n05e8h9jqyCrY/lvyyDi0XwnzhMxP6g7DuZHDGw3KMkOf6xW3Q+CHzKA/s
4L0a5lYzd8fGliLha+ReAs53DgSMOu8XMUNpJR6xaMv2TzmVpsPBpIQwLQ+2d9gbjtusrUPVPMp4
lu+zGMqKts3EnC+j9y0lIjLjQJMEq9028dSQ/QdoKCm2hY/36/kT4IR3qdy3B4j+Ou2LHf9LyZZM
cToC7/n5An9bw/cfLSCDZdgn0Her4KK3aTOJo4S9pDEpkbmIT+0Yh8ed3pGMsjtxr788YvcZUemQ
sPsdm5E5iXsxeVpM5giNve+N5qvfQwwbP8a4yYSwVwwcj4tipEQJ+i99re82kMTrVGfxRwJr9ejN
AdCf2xvgAhK9VabJwDRAD+OR1YMHdWuq2GTCNNzL9PQHqtaM1oRDlgP3AIg+lDIvyQEX1R44Fzz0
AKWp+NehEuB3CoYe0H8mD0vvrdsk5559JkQX5NoAzRa3oHZPObaPWhOf90b1ujzO4QE6sVsaiyeR
zLfA/eAY+ANIXMD3Li7P0YYsSMNh/YjgJ8xazmX2IIoq9OZSgc2g/dXW+l6fC8javiADI8jt1mUv
qaXvrOTpxJ0tTdEoOW3VR0PLXb77/AEQjccQlCvFnIhz8M8EETZKR7GTX5kPacuZHeeQBG1e50d3
rRfVaF1y1DwtBY0RT/aMW28pR+W2y1E6II63l300gMZcxLfi7ZGb28DwRZYMqGC46M2XQc0Q5wrS
/EK8ZInmGbzdkJo4Do7kbT2xJiUMQ4ZrYycwyBYTvB5QEQoqyul9iwmrFyTyS1RZzJ8iw7dV9aqN
QQNvZey5pHTE5yMRMhjFzVXE5T1FuFu/G5N6vCqF6O7YzZ9FPmQAPYpVKBjmiqQwNnpq5d2ZtETd
bVSyOrH2TZFQNn025XK7zz5Dw+Xd+t8tFwwKTbmvoQ+ng17R6g7wVlj9MDjWRzz5wcFR9MS9jyFo
3z4Q/Ucft/o9vT8nNRzaqRC73AP3N6nVST0yi9WX7kJfs3SI5mNx4UelGZQKN7wKDzcEZZbZGWTz
gpBTEp2T9hCDH+hlscV+poM8yDshp5UcgMLb0jJh9JZqAqih6OUb7EbRRuMLXckl8QnpvJpcnQbH
bNb75DKJKCTPczMP5I3exyHPKyqKUQTMBj3Kemw6ZVJ9Q2jANjUPVphHT2ht2IN/ypayyXR/C2pm
wGHBITywaF0bdWrN7XS66vzLonY1gWpyUv38Sy7gH0wQlvWgZW7jN/2wyNjoGRCOnxzsHq/Lvefm
njS4CMEc57lizWddctqHRgWlOLR6A1S/3sYt5CBQKMex6tJaBMnk9sFJ4+nCHkzF8Dsq/ch/W447
EE0TcCTX+aGjTJm303Es//Umw8Zaj3YaUO4+ogeHW44zFBbl7CaatC4Y7b1NuXC0kaxHrEHt5ya1
n86DLgq9sY7BGqkJAlC3pRNQXCQj0cEPzWgMFTCU2zqH1IuPTZ4P109YaEHacb4TqKyKJ6Xtq9/f
BqjslRzsF00vnA8nDvWbdHcLVhiBQB/fiwmmJT+vn+T0I0KQUgxvlwdBk6Pru/SUnqJh9nctIX86
AISglQYuLao3t5vafC0DV/wlJL+0n+vFtrNbh7O9Y1nzA3O7+wRuxEjNYqs+biKwjO/JClqVw9FD
gicF5K0XD+XoRj7EQbyPgkA0ssvvo15G09wUkiHHsaBgMAQJi1+j4TQFw+tFBoM62/kTD6SGFaQU
qRnmF5spgkWyrA8lJRTfDykUB9dyrkWUF1ecRfBoM86PEiF0HXd1LplligWrU7vExE48SVBN9+9W
Fj3UD1iJQDGijHBak0fWEjlDcC7Bmpp3xNe+HVZxdQJIOuWJLsJhtxJ/Sf8cQc1qdGNY8IN9CN0s
vn+LX1pLnimAEfruoQ/yrPdK4WdxlFdHoYboRlczpWLH50giMtFlbXYthLsxIweBgGSi0oF5k8Ey
gVRPKRJAC/FjCuKW+gwc9hPIW5tcO44Mz7X78ZweOYb9aeCxLx+3OADJYZ3v4fh9OL+Qv1mcaGsj
Kfwatj2gW5TUmOVWM60eScfREB1SX0SwQLuf19KP8zCIxqt+40GurLWoCU2XRsJSYqqSf16HFqo8
7SOoXna/EDUAI9XfqMlXDBEY3aq60FMVjuIct/atrDtikqEzm48rjqcYy3dOPD8A5FXplOlHsL06
0SjSVhr74XKKVKM6aZgHeenv4RKCROo210JQr26AFsWUdgdQOWItKAqICbwrNXUqd5iKbafcw/15
qxXLwGmeMctISp6PI+uhGQ5sT2RnU/Qdze7fVf3hmlzrHiwRHWGZFBS7i7JwlWbHJ+qnP7Kgf/wj
FJlSmr118FuyzS+N+5thnvkjEeJrxdp/5qFjZFXzImmy0FcVAF0dTpl428R8FCFS5qPRmasDGHCs
3X27jDuGUZ0YW11yzqdHzZjS5is6asAZGF2MCh20gPDenCFWMeAjNoGDQRgxuSqT/MQ+J2jaXtX7
GH7HRrC3aurQJpy5TPYI9zRdH+4qis23akaKPN727y+bD3o+rRElCasK+paxwVKXTowvsL/QtFGj
nXxK/wNYtzSyCNCM5N1i6EdHSfRdSeavk7vt43UwAx9b2vxuOZZFb//ekUZa5/WNkaAXJ0urtb8h
tLsErt6X8ukwWoMJdodC7BjV7CWjoUpM64CPyGBtSPa1JDLpldXvO+Y8iWqBlN5OkBjvuvn1faMu
K+8igwG7/3oSJjPwrvZaJ5CYecIPOcVUm6OUlRPzkYVikp/byivgPbDRnppgc/F3EnMWzY859XzD
TUuNMKjQAne1ifTmZ7Bh7unuDajL/5BlCa1kIrMzh7yWu2nmQGfY5G1BmL5KiX4SD5p3FDjmeI03
881kjhIl8SV+dvUZlqwt6ifgS6YHLPz5SB6zxyGxRT4z0HEkd7KPBkDGxpo/yZ/YZV5GDVthaqn/
pC+dzO9wfZ8j2scdlL5Q1ADcNhElfKok7V2BScxqoVS5SV5VOD3SAormy2Sa5pVkHQubPuhKEZ1t
gwmEsPvScWhAEIMb7H2iL5zXrOv6mZV90gmitY/wRebDzeJiI+q0Fd3P552PqvjVIXPwoZjEfIOH
GQMFy7cDwN1koXzKL8mmne0WY2FtyWcTvDhgHrDJB7fv/9QUiYa4J9BsJDsXisYxtsoMBHgwkJWf
8fm/n11uj1IkbFstDO8jRHsC3NtN1GJl5VtrIJWsF5IhDnRMY8TlLz9EnEGWpuRJPqfxHk6MYvfI
9hjOSsTr77Ry09MEbH6gEeJqM54qopxgRa40QPKuEMWXQv7dc8WCnWzVnBJSC3fWo4n2lUkJwSmj
eBUevZiQ5CTX+1KBPCZ+wBRQ+7PiyVGo4I7hT4bFKxdnTy0vC48C83dXUC7DwUlHtCaRRIGa57Nx
mrCprh/CPiSfOJPf7qHajgXNutVyksLzL59nvi26cy0KJF7wVvwp/cTpefMvfiRuIMaprQ01Ewd7
24oushhsZkBBIO2W0nW2SUCbICqt3dja/N4U7JlyDdzecGkpd/elPsc/0jqdIgfrG6HLy+4SlVxQ
zKlhZS7Cs/7hZt3+AWNjvgy9xpFiHFLJ30hoF1L2BTf52TcJ6BvTt8bMZi/iArkHhq216SjAUT7a
JXtodm8y1w42UMpuOqfFW8115qGob092bVQ9DWYs2IqOCOsGMZqnzZrvI/sSB4HqUAXzpOUswdSa
evey6Mipt8HTIPXOMy45QlEOju7UETUtnD5iua6XDU8BVvt9yhpL70//syERU5709fVjVT6eJKfU
c2sBfQkqmBOWDuWZVLancQvrfKXJPAOeaKEe8m873hYBAv9lz8qvbhA2MD+Uq6rPLj29HUdTbwTU
GYtwFs5wGJYwlQn6Bd2xfa7fU03sn5vyjQ+Y3DpntERnDrm4u5thpP9jZcT3TTIXfO4vnygFHXTU
DO2IeDxCLydRcsmD9uKCEv7Z5Ww10QKgZMzaj15IYGFDkAr+5+MO43CCnwi8W/aP9zRUt8v7mKS9
JwCujj5kR6UYf42kc/hdKmVtSXOpaJ7JddrM/ljv7+oABl7hWKGT99Bo3Tae/ngfJhWyFWBwCdUV
oLIlTUQmdXt/A7Z4x4Hw4vZLFtEjM+KMw1KkWwRGwLaTYcJ7mIxLL+ZJ52lJz3p1OGVjmeHsgL8f
Wk5GP9emauEdfXnWkJDAUhObmM6fjp0PS2k1nFyyGTPdhjGE4eRfwSmHXz/rM4Hchp2YPih8N+Go
KRWBnLQwMnoz/mOZLWWFTiF5JtkliIp4pAjLAdYYwtwtSK48fPn27OUX5YWKSKOY5nnN79Jii/lv
17UnKY9KFGXYugiKIRIKsSQnVoD88idFu5hRMrdGNYrh1SfRs/xc79gV7B3ullR5ubNokT7xAFD3
/Z/o1InePI/3/0YR8fQ0fU0rnlOrWy2mmE1Q+b/TyDGlmlSIUkEfpoaKkoWP0mW6NSFIsw2PCDK3
GMaNQlfE8gEUcMrfBJVdcLjAo66kBWqa2K7u5f9qed+VE9C1HmQ9kKNF7PjyR25Z3m/xi0hS3GBp
YBf7PXOvJqZBODSzqQ0i1zRXiEGc+3FT/1AnwQ/odYxbR5kfaOtQ8+WAC524BaNHsLTJkMuADQHD
PSdUjACgi83/kh+PpUbdB1Vn9K51ffUyHS1u8oNNn/IG8lyWpH327Q5H0KsqLfofvj2XwLGSNtDn
kRNvoiQktrNkkuytN7Q78ZSY0e6k0aizgx9MlNw6cTJs1SANxSUErF5tp0i9I2K2WhIg3B2ztTVZ
G9FNjIeNFs/VRTuJ6FZVCo7dvBkMOUmbezU9u9O9yMC4m9c2J5XALMfRlJ6BqAwRETzhkA6s6+S4
CL8szS/x9EjczryFdoMP1cMvtizFePlVv+yTvF5HBkWhUGPAjsLZGPp8pOweLvM817z3cuXejtcr
RCUOTbba/pWYJ2MJUKg5/D7SK0Uu5Sc99WxBLDOFEQmnfjsE2mx17083KDK41oHzGw0Q2AWZ5Mm/
90DxVJaWbzA9xVANUU1ZVkTleZhypg/JX+Ef6FhTMncro3LcCCw2cIZN9UO8ZsgSgwQxNkyNfAIQ
djuO8aShBmJIH8g3+QDMVQRyICkTjAgPM0glr1uBp+uRYo9M9naU4ZD0tU5dY4ryzGkQn3XXsiAu
YzoUVOVMEGfCbzTD6c5A0pJ+LHLQnVVsM1KQu+QcBBIot/XSI6OEF4+6BWNfRD5jv6JOHG3nz5Ji
pHZoiViBM3KQvxCRSq0qqIvQs8qI38l0kG6iMMQQLSlkmiTiPsxAFGNsLRqfT1q8x/fxsG3BkKmQ
cmBe5MFFtpgq6feN1HFsthZ78d/d2WkHlyauEUx4hKVvFw/RQb3S4TzXe6GPPNWrS+pnuXn2bcmr
jmNWCnnZMJlDq/1UxF7itcV/OjdU54PXx4unCFFt9UiOWkUX4x0TEkYElw+HyjraVupEZV3pb0dO
lZdiLA4R6VSrzLRUradedwAi/FmDa2Dw2cuTmni6uisNk450sYqkBxGbj93Z0bR3sQpDbsNX2UPT
6RYsZX8tphlrSI9WZGXazYkjm46MMVIJJ0HuXdfYMd4pXFRNABTqwhWDBekO6mnZ0bCw1ZtgqYqA
lrMjj1VVhk62R/8ghWNUUbD+g1ufYUoRPMLnavXoRdtQhMoUuV4WYvUTNXSNmE4jSfdbC5UAoHWl
6oOYNzXqpKNLaaIntzdji8ebrnDWDydYfO+YzXp3NNMmPKulZB6+Y4pjp+BfGp382eVnXrsKRaG0
k+bIdTJnlD2z1phfrMmlV2In80RAtTevorHs5Q8jX8YB9ksdcL7loEpPgCrOIUqz0oIZW19l5nbL
b7y5zyZ2GzdnQC+26ikQU3vG2MvAF+TGc7nBMK3/0ECFt8ajNi7Le5FI37vVtRpziTxETO+cRGZI
mlmP+KteYl0zt4DHaKTg1m3B9F+oU7G1gG6JItYSJ7w0y8R+3SANYWwCLDl8hf2osUuR88SQ/6rP
k0D9sQsjYjuyfdutlVGTDgDZrk33E99saQd6LrPdikC8oAwBOuXZsLgWUL3SBjF0er9bqiuqrKY0
fbqDxkabRgZOLkCOAVOs557AK5vCmnDHKzTOv9iL+LP427BMGOJK6RBDknXkz47m+uN9QVw0RLj9
2t6MGgCGGvsnaSK/Fo0/h9j8ES/TYC6W2IIPi2qMHpkPGwJpYxE6jxmI/Hjt7xSbt9MSWJaA+wAp
wF2EtAY9MZHnSQCmx/ZXO+s1C3pjgKe+y6r1xG99NXFrSocYsQryHJ5izO5OMEyf1P5yReL06cpP
KtkYkORHxsEkKxQUA+P+5Ds5KgWX+qiZDwcMXoyxY5A3NT2I9dgrQCc98lMJxnqFrp2Z1bLa9uQ4
oHQFJxFyXMkPUizvZ+4T8Bmj/W3JZeV3E7c6gdYHZnqEANEzOkGljMr/mccUN9xFQhEprKl7LuE8
JB+Q4okmLUAR9wswzcevn7Bz0H7wl9GmAVG7dZb5MBnXO5id6ftSd2BLTBNCd9KtKP2NeQwF1ubV
JJ9ilmYVe/mH9X7iVOOCujjN4Og6lhbFExQ50hNzNr3O5EFl4/gYoOjTERJJ1pMwOPJekPpnCD5W
zXN1hjEUEsd0/B9wmVpM/CxvfkTe+7B3DM3tZgCLB7Iempmy/ZfjlDQtCVBp605yC1zRpO+S/kbA
D9PlGvhPzndfQ4ykM8toiMZFjK7mB3RZlLqajNrQqhCUv2MugLOkmYFZ+YQ/taprFYROQuUjUnI8
Cp73QLbKMBWwrVlmpPlKk8In73cPXaFOLw3lg3BSGvnV63UE3Qv38qhIyHYxWspJl3Mr3Nad0Xdy
QMcb5bKNB0c1oAua+dPCWDpCXEjVShgEawhxccHhz6XUSkOhPcam/6IsBxCxNOXZciQTW3Np41RJ
DAlQxcyuFL5R5LMY6mDHECBbhQkJIwpJqAgF5SkMj4m73UaBwEPX0KXoyMOf6yRlSaBem7ck40PD
drsvDbdpnabpteU5pfVB1QnIpf9FpvsbWP629cajOo4drHNcULJ6opdmlmdfdolzzDYnqwq//JQH
g8AyMwWTnFQ9fs4dfnb3mSRT2nSxB1TEPrYzSzVPruykNVZP4yarJhLK5H+RWGZ5PEOu18B7Ab1W
O1De9TIODE3Bkp0zBUjGMUSdEvJAqkgzWedhan0VFWpxs/LKjmmi0HHksJSWuzsr9dBPsH7AYpWD
vYr05YIFg2HVu6hg4mm5/O5oQCkHH481eZFuW0cMdrnZDE9Y8AsboY+rCrYD4oSZS49lWxWjzAuE
76JWpLU9dAp1ypxwc0oaOfvV8Ae8wKkSfnfllvxym5yTsdYfiC79TbJZUFTU668o4WeAA7Hhh48L
cDBH23LjCEPliQaibou008ljiCF7QA1xc+SR6ILmzbOetow+TKAS54Fhv3tXva02GB5xSHyjf1nB
hbLTwJ4WiVsqxf6SHQCWUrDmXLXrDOLQ1sCs+0CZbfQvYXpCD+ngMLoDLkq2QXE/S9SP7ltft1ev
gl5urWbB42Q0GGx20E+x5GBCPDCT4CHRa8/FTY+/XUTpH5hLp9MtR9rQ0qVNu37Q/O+9CugRes7/
Swp9rNd+71KUNRNZN3K0HKp8g13uRCf1drG7JzJWZIizokKUlYCdwz6+xYUn3Obq9v+SiwMcJ6B1
rdqmqb4GSgVaZTzlUc2y4RORDlhWW12/fAjBkiYsCBQwO0eO66jdTdnkSu7pGCZaxvkJYVl6uHku
ws/taz2BW5IMDVa4/IMht6GUzhskwZX350pNV14NQlDG7YXjWwhPBgTurflAYTY96CcLnaqCk4hO
/a/hXLrteEHFs6Qfg9TR4saj4HklEULtku7zLTyR5Ufppjqg+IBIpquCPPUnEZc+v9GpUqGMiHBm
NSX0cOxWxxptfM7/kQbiCkm5X15AEmM5KbecjAyZekh27PfC/jFi6jmRjWMac571OGW4nIbkRthg
tyOa5+FaRAyB/9xlGW9yCNmn3JOoQqjFmBdfjVQcZIK6CzltO1rE5CC4TV/9iSnxvCqVHfvNiJxC
BD/lbv1jocxopgefJF0GivXnrM+p8m1xFrNcFBS7skuCKj5rf/8PuJ9GPBm407SqDEz5kcZ/ykVh
AHM/zmlCWoatB5AUXDRSeow92PNDGO9a+eiW2HUlTo9fVTM/0J/EpzdOwuUlHodGC4VGYsnlVs/2
1OgPGy7LLC/GV2RQl2nQ1Z+ARKi155xozxtc6h7ZxPcl2JA9NaPHy673egFLrK3sAgp/45RQs65i
UWmn7MUlLZbNJpBJWy54DH63P+YcLQNuBjnVSuu83swb/pYMOyr2rIrEEjnN/BHEeKC2tauLNKMk
FgS0qLMlERFwaJb/MA5SiyaNnFrkNX8bfR9MMRKcXKB3jAyXNcfIgkhEgsJLmSWewSXjUx20azWd
uynzqk4fMbRcFksnGpmD66dDLyXEnvQUs2BlIfL4auJ33N5IQRT3ogDL+zsXFfrl7RzBpmmQx5tk
fi+2fSd2L05K80G3bnf8yi8g1ezBEsi05yahuTIznOi3dmVTjdqoDzF2VmjvzeqwRzMzsVMyHxYq
DFalxiZDuEVzFXF+fyeaoDRTCD7wa7zyw0AHnU60JAeymkOaXXg+l0vRcDzEiKyJnEGsjLV0d42L
Dyje2wTB0YXO3pKfSRVY6hhzbLlCDnECansKCnTZNqR3+4h5sR9/Vd/lJpcyb/VhkERIyNftKZsd
q0m5vqKGzXmKu7e+POcfHSTARnVt53uLnWpb/umGr3pGTHwC0SHXdGzM0lc0s47FoETh3o73G90e
uF3+KhrATkmMBnRJ8kGGIb7xq83TmcSwGR2XQxmYgIn6aGXZUYEq30ULVjtCybkIzDwCg3i3VQti
BYcW4z58JLHe3Avs0qcjLgy5vpSzmYbIMLuFfzDif8dEwJiJp3h2+OAvhYawDzGbZXpITE+w8drh
mmqTiAg9mkUxMnnfKP/sPPIUfWuhHNEO8+6eNBghhf2OCETtnyA878UtgidEnGnIB5jicnHs8fH7
u87VfW/ZMc7LsMEe0PU9jBWETb91bgqGVBbptnjEZHOG//JJTRpjeXEsgHkv7xaAPXdMwLgYCu8I
pI/6Ab7n4xU9RIRoYMdURkpaAeTG55afUBCXG7WV/F48CuD3iPhqqoqU24uRfLXZoHXSIpMtRoPG
S4hXhh0WvlGNzLOtnIhZAIlJLU0FYeJVZoMajay+Q2SjLlNFxJUEMX40Po58Vt+q1WNrg1F7zyqH
4heySYcEP7zNeZfa3jtc7dsA5aGBCK0nYDVO48lhmuiNE6vu2Tcw6W1mGniixVGb+4xoS3x64QEE
smCbeN+Fd48TFs2RI/EVb16Q1Z0rpUguJcsetWgxQsUOj96a4BwaxgNmcHr/g5sAQ8Y77E0ckOk6
NJJG5my5ptcTYu8k9u6I4SdNTUU86F6HhLdwhGaHqXLKtmkdVGbsKgiZCZxLac2RbddsKG90aTgJ
6evXwRbTI8ZiQugR+zUqUFjekQD/Sy4zknJHE8hkAmFFAyycw8ft8s2zFkeqgfJHsMiYKnjuJ1bl
EzIcdS+eLbGF0EvsC3aJfoIUqCoztbQNxRIotTyLbnN1AK7rzwmlxPi84IoNqqeVRnSlMJNH9EcG
tDUw/hEgkawsc+1Gja1kNfmROWxHEliIv2QoNN8+PPrI6Je/emmIBn1DUroj/ZzGfNTXfKFrerxA
4YyqHs45WA7ihUiJ0Ez5EIrxM1GwNlONqqJF9GZmOFF8NwqevxS157Lng62CIjBsxqIYrdN19YQ9
NZPUKBbKRJ2KkEY5aL5vp7gtEiSbup6JGEJYIs/yKlpFQjczIf/3Z7nfCSWggLOXr+eJnVlOOkx/
CNgqdm8zi00CHVCVEGl+LKObB1P7o1iV+bmgF+G9P6YKDLY5FNbqIMakU75lM2s/2LC7E/zDSzEV
xPFoo3jlUaP/FGWfzRA6gnmDkTRgeH/gnTWz55WqBkuBSWNtqOxaSr9cmT6XxjDa9fVI4fSBSid/
XEIQIyosWaaQrPH5qwMQWrAnqC/fhMQsX7mwAg4RPCMPJdPWXycZqB6+VOFakdJDzp05XiFdaW4h
TvZ2vQ+Wn25frBh2DcOhmBJlxRd0KuYd0cWvgBy2scFbgaS1HrzLRd5vd4gXS+GVPpXWQYe5ZJUX
+WILWAo1R9LoyghTRTJiSj7gfdwXi0v4zcgG1j+lbBz7BT12xrBUfkox0jKZaIbmN1W61TafrVZj
v9J8xNGcQFzeM5oO+WwNjEAok1IWYsdA0dfnloZh/QhJpnGnOh+ewx3uVekOWFUCeFfeyQx+o2fM
89/A9h1wyIYyg5eZKwFXSX1KF58lv9MquWs1dvM6LoOuVa83wb1HSDJ1ufdCYyxArWuXlIoB8uOi
Vg9xw/dDtY13Z0czhMXxPOQxsJtx11vrMsfMB3C/RhAgJFRMazhDm4TDGQA43eXKSREldxxeZAWp
SMiOchZwJ4yxZ9sPQgrEsnXGnVsx/B87vpRPRKEjPny8t6QipetaM496d5nfYqoU1Nxju35Gw7xw
vDLO9UPMZR5DGGEHcSunkC5Xu5dCCpLs8oC9hV8Fzrm59hMgy3BXBOEEs3gofW/jt4PGVhF5mVM/
gjAstPaw65+2Yps9C/obkXBkuslI7632eaabUHmbkA3Kq1nExltZgtIvd8piacAh12eLuxKNH0VB
Z3KLm19pCtBXPwrNlkMMEXQm2b4/5dO/xvEDMUHRfr12Lnhhocaesa1a3jZiZoRKMax3mpdKFbfB
1ucvmXVyp2BPhDdfpEUgQVbQt8gS36+Qv+95K4uZkbUVVxGF15xZBN4pM7vVo6rd27/WraHnjmWP
66wAUrG/vAxV5GLaFDJx8r9oaMTwmbEQFdfAOq8ayEYXS4evzsTYhEor0DQSOfNHWWbCQ0vTGR99
4C1lNySbjeOM4Yp+4hetaIGYgs53dRRpvMjOytnCqTzec0jW4ilTT8fr7rsB50+QrxbQGfYM044Y
R+NvnbEaOzPwHn9r5wuktT+hvDCH4rMeICTfcsK27s571v3rBxxbBXWyTMgxxG8LFALQUInNl0tr
Oli7KRb+WbsER/yg0SwFATnAix5iqyhnud+aumoW5pdbVs5SNVJAUg+mCJiNr1wReIGdbv7ypVJ3
j8XWtCnJBf7gZ7UU8MrojEQ8I+sd81Ap71Hv3Eq0JFN1zr9Ewlc2tLjLphaORLWQEz9VhAbEGUfa
7wfSY1nljK6/xNeRgun9CDcle/JpI2+VnH8l1Qi/eulk7zr4P6CcZ5p1ze+fuxhyA+K0gxg1j2Q5
2wcAMS1lIUlpvwWprgHmaoLhWiAATxZq5QhpSed4vKk0azn1d0w4FwvaHKX3kcUGmMTHFW7GKPjx
VWlO3trLgIOzHFmFxaO529iMu/HWk50R746wd3DvvDWPPRWKnO0U3rC5Y5RikIS/8cCPGz3IhzXv
rCQLgd+zg7r3KOOs+pReaLR+sHRjxSUsUHQNL/lEAHHGpyKAEPoszmE4v5QMNYzu07G5cOpCoTH/
DWT9Sh6748xjxMsulQE2KHiVXxxBYivP92cI9ex9vhacwtU1u2RAr3OAqWahuX4mzEfUAhNDsDAG
6fmxAw9Xm9lUDs8xwXCp365fYE6EE314hMIYR44xpg2+pvUdDJ85ggX3gB8u2oYJr22VqJpBMZ9f
racnuu+PtHhErDj4plSGovSQBst6eZHBC0CoLvOkA6jRyfOEKjh4RaQA0xf5XbANGxlPMQMCqLtL
rRCKqsB/Z0husW617YtC5oTed3QUhIB+1Mz8690zCco8oYGEMtHEq3IHOd8xtAf2K1tC2YE68Fqz
1BL2nX/IM8xQAvEO9zGE2mv2Im4EzZNC6ozp5MqSRN+q28UdXaQDeWIg1cbviA9BovRT1yWWdBcv
fk1O1SjhKEjkB+xdxMGVQqnthsssvEGCINXclTHif7yiPKc5BoQh883aycsS7z0GjDP41HB/yOnW
nCeha3U87t3FFbrbvkOk4nJwoRnqXqXO7VzoSoq1B8/GFgRbQynJgYO92+VsDz3yJW4CwUGi2Gmr
GYnJYSphnZZ5CCh/9Wvj7Z8Gy7/6fJLrR9g8T3YmbvSmYzJl2lGVsUiPW3QbrwBCFZchT7cRuWKl
9CVzmvPbHZUAt+SOXOVupGru5x6Tx5UJ1+oD3xxF92aUxTuyX68m0Okl6FJG9ysUsbKJXo+xGTmM
54y8UJ0pgo/22UeYwKslhdr+ppeAxse1UCncflLu9X61d/P3eP2wbTMFrkla4u07RsqBDWcpdT9V
RIzF4tzE9wOF0dcNT3U7fQnKI3PDUait9Glps30yvQrWCoPMsonHySfj5OpemXU/mhZhWDmqeIGH
p7sgTLkBsWooXQVvjwRdFynY99VI1+5/thvjoPsyVe9YCgd0skSpDoKJNIihFk51WdpyVn66EbGo
Xg9h0b6DOO8yyneclFXfhSsdCyuFZVB/UJd26PQimkpJGSxzsZVCLkcQgS37vIdBP1WoSQMvlydz
/wJ8vqZBAwgBwic+ZapRzQqw+gsJ7xAntk87Ce2jsugJl3mtH/C9R/gPrDQOSJHzcDw2fi/wf7dl
pZH/MxBXwGc/qZ31jh7LBBJnwfG/c+D3+FCW7iuoB1uUf7s/tmyVQNJC5Wn96CcWwL3DXK+SrwZg
eDuvIlgMWnM/Ci6FOVQ3W/TENoFGEM4EGrmw4rQyNucivn88rQNQjUNk2nlIW+H+ILdd89Wvpo1O
+OD7B28Vutwenwi9PM8h2wagarPJ6kQTcKPUsMCg1v5t+CrA14WJU0DmB5YH+N32/2MsuP30q7K9
lIpsZ8Tllez5xjhJ8e3PS3D5Lzw7dOo1p5HY+9DNHon7hMRO0lnedBWAPkjFDEMtZCLNMMMK2Zl9
AgOdKR3NdJqH3nda94fR3Ba2MC+zTEDGeNjGMXWjsLJcod8snHI/1Jk4NARYnGkI4SiI+D31et9x
1l+Mi9smYIAqdxH3QMwSApCLunPiZfrqXpJjnRQs5gBE2zFDyza32Cr+J+NKDxSnmPoVmqry4rdK
zpsR+B6A5dPiis9yE799wmQImKg6tRrnt5ATVMrNa3d+fZXBjUccR62RXOajnMgkgnu7rNLjp1xL
J/fNyTi/CnoU97qj2oALclBfcGEfRV5cKtRwKgWlxjGQsulnTWOrhKclBIu9Gex+CQJMRc0SABIn
tMBC6Aq/PGGE4OtbPb01gL11r5dd2WpLPHeEl3BG6L36HMy3Vd54KfImVLIihR3Emr+a8IDMcQTo
wxkuBL2V3U20ApBbHjLeN4e8abXC+QHN4Evx/t1GovnDVbuQShYbBXIRRWF/Sh5+E+YjSeefpPAj
nEXwGrZFDxeW6kEoT0OjeaF4XuLI6odQB8UncRoZXcJ0uo9ekRN3aHB/S7xSQ4Ufv4/tbzwbO6br
D2c/vM2rFjZDJl1dxexi3EtaVrgYP6GBjXbFcHMds6N+67RSftqd+jhh8/Z0SO7/0+yOVEmSoAgT
8hSG+kRDim2EnorFPLv4x7FHPpnpaSGeC43xlK7l0uX+VREziALPHUy8RbHEKPMZ/xJXacS9Lxbe
7Xs5N7J7/+2cPzzIJjPcQm0L88qZ4/aeH0/dH80GJymCAQsCfpTRj1nk9MTM1wX/2WRo4QSDBffL
DQxDmTPAHb6WmxeOmjDDiuGSbYFpHJFbcZXw/bwFVTjv8IqqL5ypeE1jbUV7KZMfbfJOThigLguL
xT2GVNghrIbaSsRsEltf6lHojsCPG3zyKYjRVC8o6usceJ2p/2zeGv1qVNt9xfpRQRFM/mGQndYg
Ew5PsLQkYeE2jSJrjED2C6Gi2iXGaDWB5GZR6xRdh3949J3jtjpRm9ET9fi2VuBLrj0CHmGfAgZn
T9BfWRbbrARrGxLZ9jCQ8F5SO2sICAB+P6U0u2HUVJk01XAYwnaonyqmYwiv+X7GF6nJZa0UHaEU
rDHnm8r+7Xo3rC9INiZh/+vWF+18+a4lhjHjidjv5ucI++bpZI4VbXILw3m2JQ30kMa3i0i6vvua
7GZFgUj6MIByQa99n8K6YHbHxpaze9uv8Xd3LTQSunpg/3B3kOodQLVOcCBM9JOpC7lfwrK8bq30
5JZXedNMCN6QYNHAF6NYlQ8lhvEWlItASt6SnH5QWhsRIeJvRwMz1ns1H62p7bOxafqYdyW5mTd9
KWSjqe+TjGzpNv7mkwUixAohRJ/8XbXQ8ea3uEoRE0kGyVyTm4EH4eGXBRA5Cp6liTs9tc6VBN5k
ik2wR+E8OtLKTpSJpytu1IMw24vEVuO9sEGhkJhC5lrKu29rwh3OWaYzkyUg7e7F/dxwa5FAuU9W
IcogQUqaaq0QnLq6v7DDjwKAHCSRQwHPgjjU5rzNRAO2iy5OMqS3e1lL01nNCaOXMSUICZuYVAGb
YqAcOjsq64+SLi2/cEjjd7ZyoHgRcYd6ipuU68yG/l01GufOkUhwD/NO7zun9Iiwb246n2AEcGhh
Q7C9vLgggBey9pWf0NJXIXNYp54+AnZ4Zpxr0DdbqSWazhTQr0P4ZJjqfGYFkPyawwoaIelg23E3
+Ucm2WaVa98MYrA6ECGn+KZQG6KWF1zw7nitaXbeKxin3p3X4qhOQvcrBs47NMlN8Ldc19cEdXiY
SO5eW2gC/rcqeHv7s3R/YjID+RS9suXK0hByNNpcZubUyJokelsJw3u9r6QelG8cWbTMzxQSENBg
1B8UM/qwvObCFYZdrVHFV5VutR1Pq1EW972hv9Mr5uNr9ga8rz1UgbgtyaOR+x7xHJeDZc9KEnN2
UXdn4yIcJ3noOKm1pmz2LPqV1lyDW7+V1s160eZQ54l8bdQF34oZbRtIaMiYu1ylD5U1XmAhJIUN
SJSIFB+INdL7jyH2bHBBYG8tzkiB3ij1ntRFymuJjHEUihup7X7/t4mDYFnYt7cnzAyDH3ZlkxgQ
wFqwgvH5sXhR3p/VyISIlm59llluzU7Wd4tvNjuEZifiZcSgNDOsPle833L5FFSNhbowkzYCHZ+R
zuVudkk3z5h9KvougZA0Nj7UXeveZV2nj34VvVeqVaCLT7gCrFumQL19WtOGplyb00HB+t7B6V+J
SF51NJvuaIevto/PhzKT/nGZZ8H57cdeZ5njXDs2n8y67/sGjkCs6cRgEhWmQgWVgs8dKH815I2k
Vq3BGnwzsFMnPVPLSqUx/Ol3nWkNaeOZxjydE+jqmOfSfj5EsI09MNJBdyzgVO9uB9chMUSrJwUo
c5qYFQUC+7he94b8sL2Aysu3wkf4ja7wi13C6xJOCq0zyi7gyEKYcuQ2nSJU6vcRJEy49nlJBMvO
nC2HcEjMD4Y99f0qinzCUWtFsm3epJJKHG60ExUFUk1X486NDRTwlV647/sZPrrNjUU75ydxCWaJ
QIcAjt7juDeKCIIUM0AdHLzoZ83pSeP6famvGY+bWtS2FXvhHvt1QCbTRA9/jq9uP5+Hy8YIOP2T
3vXd3QNm6WMIdGeKSh5S2349ULQk40ldJh7fttwRv1VOvg7IgzjS2QbPYc64fcYlsvfvXfMrZT3E
yICuHi3+YVeeQ96LfYVbQ3x345R49EZRgl2jXq1T7PD+AQE01Eg02BV17ddlvNK//8Ig5kduutf5
JJcK6kZY+M4FY/Vi+v3oxflosABe5MYv0JoyLAuKx+Y/dUM9Vc8IpfE1FKT1A0ICTyDaw95ExRP/
npy7IyKAC4kK7J3YTsp3Mfkxar9iZ8e4t/bCYTa73AlC+6UYOm4sVvXzEQzIlbIyUGBt/2AAjCRC
KE7gBk5Sof5uQmx1m8hVcDa6gzPHDq1h55UpSAQHIya/E/QZzCa8Xgm+uMk2lelMwtqWyUevDc6C
AyDEq2mnKZ7wq8FzDuJOr/7UPxnBt9+IMkyTLYzY1O8s+LAnNhSjs0AOiZR9ayPuAEZ1qPkpKkRT
t5txNyRuCSyxXjc2Ai2H3s6/3nbwU8UFjPZfGGBJd5ge9g9BG3Ht/HTTB5pza1iQOrCZI8TAG7gb
YM/ZTHaDAcmiQa/8f4PGwmRgS1f3KkBx+VgCxSaqT6sF5uHeeXb6P+ZAGOiNSU5D8hytSq2g9pmh
4QZdE0Y0JC2ADQcxpraPGmgy1Qs4T6IZ36M4+93adLUppGfj6yTHI422rKoNtn2UZktiKFeqeGph
wPQ8wA6rbxRk6MJjtBD+I687oBNI/EAmoM84Sx9y4FDz50ntBSWLJXHJEvulf2NzXcnQ4UM9MkWg
9EfrDNd3sv2bTTkkekRSzvajkL/krnukt1dfO7bQHjQhjFECE+FfDtCuhK/yvb10t59wEPe8hMXs
0ZQFI6C2aEeI/qgKpBcS3s7YlzmXsWvjLu4HixNqdHolW5hEhRagJV2TPDkTt2iuSRjNIdw4yc0g
W7Xa0SG5bZlgPEGnP8u8ADRyJXONYuyj5Yo/XZ30d7X1cIHkABktkdINhQ9F82uRsCNOwf6kkcIF
jI7evJehxGdH0XJzRBLbftnnNyzG4rVYZWYKRCsj7ITAX2EB9XEAwiauN6aIoAYfV+tfwbKdiB6x
jVkHuiL6lvDt1C2F3Lb+LszNDZB8cs2jdcT7CqXzmwqP3P3qJrbyBgU1ahtsbgtwfVcXc1bxbxY5
R3n332K5o8Xh7Fu17fihH/E+WhMgyQshe1KXOMZ+1Fsj6uXP+5vQe6vRThkEFEkhbkvgGKDI64xk
hZjL5OJjU+fJ+AHBIPUW0PjqShs9Xbw22z7TTsurOOu37lHtSbMOTA3nyLcWTeUYeJ4ehxTia6Zc
L/7K3zOzo1ml6mhiZJPEVmvU2ZQRdAObmHbN6ZrtgoqXFhMMJc6QpVqPA8sCkVsieN6484z+o/JM
IZp1Ze+XvkLuADYpH1LZwOdma9zoHrUO0lbgvKFi3L90pVgxHsNG8S10YUxdB+wHItbAfiIjwovI
K1ipKG56GsKSL/+hL2TXm1Wb6o53T+yMhl+EO56RgdUklES2eT5nNRhCCkBuP2lhlCLnbYbHigdm
biAXLLRVdbhisJYLf5CEBQMav1N9shDNBfmhfg3+bX6TtePU9syzQqQXFBN6kEWZloIzQuSHZBxu
tGNAXLdLs67lLoQKgT0XAElBK34Ygfp0shmh1LO8D1rgjRtkGY0KLUtPgaNTHP9cOI1rY7UY16G8
NWGlpv66QUVHELQ9jTgvXrE05TiFSqiBu6nqEcT+82MWCPqDvoCo4ja+MBm9y3Iy2zkO8u0G49Ve
bgckp/BaeKctaudhFCqjFEuZfKtYes7JTaR4rE727WCbMU4qsUJRwvpJaKaJOIMKrQM8qw1Qr6iN
XAKCJhVibBzCxqR+OGzJaOIpqA+vJOzRMb5vOPKto3qQ9NA55cOE6pL2UaSqCPjQV3N+2wMRibAN
+SfXAWGY7BVBhJgoez8EYI5kL/U4McX0HoIey62sLONn3c4oPeukgWmt0x5snuRWQxB+baCylbb+
HjHqDBXm8WjPcY4GfONiUODUWFyaszF/Ca52wbYoHc/3XDrm3bb0x2N1NaQkpZglgZaYN/8risDH
ZD6ZfkAu1nI36Hm5nUAHnG6/Yot0i3Mw54fUnUfbrPbV8i3CN5uH9EaxmITysFWsgTFRtsIDFgZ3
xT7/QUka550CHVHR+T/CB3OVIe0ZG/vXk8JfZmPNsKNrCx607BDdd2j+TV91a5w+8wXag2boUGwL
J0uG8sGFrftjNVLno25dyXKb1/0/5tqccJR7PaG8zJb5L0kunigUxw1pV1avUMSSEgy8pGazm8aK
uyRaDdLBlnFySnJOn7Ft0drKXCExkKMuzrhdfHGoTT2pLtnFLcbPU5LRv8N607LEkwoFCGr47d8E
DMaawhUezWasTujzFONUFZW4MB4g/ZjNMprZ5Kgd/HtXrkD8Dp3PoyD2honR6iCgRljT8KoI+g2x
0gd5Iw5LJdeUZocBacyH5sXU11M6bJ+5wCPRz5CsQ0puD/xcG4C6nzoWxmT2ERBfna7ewfdr8ZNx
39i30392RWj6yIVu8fPKzP+v+JGiwW9NbyVnc3LUH2arTbseMWZWmYoyeBjpujMbeXOK3CJ3DTwg
4m+kM1iiQRbaEXuzfS4ZsvSpX3D+NlFPaXHtiDDW8ZwsAvXRAkQ2kIxN7rcPeVkXDO8DEtka/akQ
T22DflhxQYz9vOQIps0G9RZ6SlEjbu0LgTPw1afI7i69oXZHQjVtxgMVthgbImpHXUNSvoaQyOMf
3qXRmr2YXov7gfA9e2o4mQZV0GhtoyIbAdi0rGMrL//XPwdZEtHu1MQqt6oFgJVwV694EbR5+tiD
77Tq9C8XiYzSf8rCwsO2/fRY+PNSjoDzaZ76iW5w/pZAY63XulB25TnibTM9YXxjFRkDl0gW5Ep+
M8+MiHSdfV50lWWQKuS8h7btLdVZvMKrvwbPl1Tbes/o85SXOSXoTRjTNBINxshoP4+7DnOCnHny
BjmXBFq5goPCKqBWjih8Omfi2LlRjJ0B81JaklyCmN6bBxHdsu7jikWRpp2n+/4wXgyfCezwza5a
KQhpzdgEF5zWrLa0hfg2BQM9TcrJsMJdB2UdwYKBve3BJEqsKOsNXmM8BgqamgwQjP8Mti+oz2WQ
INXZx1wrrv04S4RaJzYP0DCozrHsiWBw/AizRoglyUYbOx2scpTS4qc8iIuGVPZ9xDU/T7NZRO1T
6SXBATlC5LVK2PM3zyGkTDrM4KMr05UTjfRWySQC7v3/VK8gli274CXEkheCHWTfzDzQzq2W2Klq
G3sl0fsRxzY0e5ZiyyVE5FUW3qHMWTQ/6y+bafZmqk7VaV3VGOZe/rmH6xMFl5xM2e4voEcaJLP7
pHjNkPq4p9vdxWkAVH7ABzcEBVGPdO3R82lVMOj4y2yNyewwGiPvEtBt6eWLSE0Vc3Aw1tvHgSr5
6Gb/YJ5Jkogf5UOf3luVeWOIhuztln6iZzgur+JMXXvfU3FtVzm3m3zemwrQ+Ium5TT/Dbs83J5o
I5TQoKPu2bDT0EOEyC1+UXguHuuUaPvZIouaEg/Ud4X6t810xYsbo22+w121Vn3ELyEXTfJ//lYZ
9kExy3P3X8bGD4acCFdXRNogWA0kLXXKzBfmfGgANla9PbAUbhqhwmswB8npL/mzoCIr4ByVPhyB
MJwx6pHzhs0wxLmwlP4d4PoMk+nFUz821jjPoenKRs8UGBH7blAjmwtaES3MOZr3wlP0aHlVxigf
JVclNyEmJRPKgCxcWhk/1WE1ZC203awy/Nx//5bKqNI4+Cp3uVQpXv+85Vae6SxD9oWQ3Ii1kUt0
O9rsXRTJl6zStX58x5T75Z5xL++jMi6vTEU/EJROdBRDPzOp3Btor/wT3FmHXVMUecPxC6nPtEcT
8WowFQtIQEMfxW6hXwO7EoN4xIF0eHL/l5qYY8fbAVs4Nv+mt2/Won/amTAnZQo3jpQzzMoTFqlX
Spqys/A3SLokPDJoRVzWwK1OgBAbVch66LyxG4J7ud5V6bTi1Aac64ETTmW18EusZSfIm/Jv9bye
7T1R/zsB8/ji2rchUJaSvi0FG2DLt7txYy9CSQVhJpg1CJ2Qv4Jepcxbgo6wxXnhJdeMAaAMvacs
NSo08AFvb2OzFI0KxSuOWr5iXfFKGYlURNpm3AXmz9stJgW1jrW8kRBVsvh5EqVHAJ2r8OUJC27k
2UfOPFHvJuzjzxF2npdRF8xww4+StX3xm9o2gyyEhIsERvw5fAk5CheZKfRFYqaq/4UQumooGH9E
mgxzb3F4uL/lWPTKw4wUIZXAscET3mS/llk9c5TwMdh0r7Jtb0Yse3aHrmpXiS7m3RX3TFbZLTWJ
4RUZCx31h9rcP5+3hV8oFFYD64V45a6V6tnStY5X9ytOrDkomkBkPlZh/Ng1a91kMvD91D/nBVHW
dKfUyb/ij03+Swpxw2o56YxcUatVLJnW5SA3d9SeamnnFx7knG/YK3/2Kqs8+8jAeyAK0Xx+Q34/
rjV3AcGY+iyqEMKGsg2+n7+HguUWxMeb5/XLXxSwscGEJiaE/uG+U1qriXCMLx+XGqCne8aM7iVI
iCabqyzhWtuBO7kddK+I/RUoF6KhIpeIrevjCSSKXEjNMRZ043VtMgqaJqbOdhaNFrE43Vb9YTM3
3pQRO3yfAd3NwmjCBsDerGXT6tg5EJ7q8B+amapEHvmzhN7JD9ZYbrOBSYZf1lHryznHjcDqq3aa
7cBk3W7uqJD+BN6WO21pZV+XivTS+j/te4GVJJF42BbrMFR3XlfSLpdkOwTeBdzdar0w8J0TeShm
7x8YkogEd3BuPlc2LHXRSPEK0yeDhjhed+MxDKxbohkzUZXZhVns1Say6K2anbniKGhBb8GWyrpN
L346iacU76wjANOC3ZYAo7qwt7MAV5yN6UktgA8UXVMENxwduoiqAWVVDPCQzCcdg3C2pSnsKVDV
TXWAR7tkuGQXYDct6KaXEep6y2PdgQeGPfdvOwj6kOZ3xAqfn2UmyZ735UTWqTCYlKhahghh3qMZ
wLieorP3rvFwyClKPN1VF1HQGvL03c5LHN6XrRfRA227AXZr0/PaBoPtQmn/D+bYxzhb8i8HV9qd
OUvlnFPc0aCPwDpwKYcBY2DsZ2f82UZ4yZHWJLxXtXUBLXl+TVItJtfzk3v1PD9icW+Rq8Tk4f4p
wQuO878lUPy6fBIHJLU1cDIRm3P6wmcnQY9oCkyYBzukATt9jwWktfCvv4L05AAeu+0FUAJ72neX
MPrncCwoVkeEw4emu+uM2GoIUPvMVpulpaG7qHEU/1R5dqxbzjv7JuoAaOiF9iRw3vEyIwrjssUf
/eRkQbTMkPz6ACDNhV/+bYksRvjY3bHfZfBH4JWbB+dH0AUkdif3MSv+MIGYWHAKGoxBZsMacUZK
ku+U6rybNN5ip6prRnBxfqzZ5Au4pmk/gPMgxwFsCjgldie5wZ6EuFL0HDYof2m4p17NMUNTnObG
9fCxP4T8fgDCrsxp6sSQHjgg9YTXgwtQvo+F58BpVqeth56xsvbopJqADfsrKJ3qrcmLlcg2axks
YZfXb4RmgaCaSqmKTsQ5aRRUmVsBCkHxK9WgJqWf8+pLV22WnUGpZXMYaT8j3LgLd5YUWvkk8vCm
HR4+r3PKJ1oTkR2ghOTjEdyQjkBbGexNcemb76Of7mDSgau8TlqURhUv97WQUcI/uGzHas5p7ujr
5Fw407hvw1frDASIbXj2zTdFoeETLI1TiFqjs3ZEzCa2o/2r/NslJ1agvlT7Uk00yPcD1n14Kgt4
EZa0GMSpTuTZBIgQ6BvBGrOtlK1uVL86ahscfghkq/U/H88IspvFswBKj3G2r2eYNo62QkVJiE0l
g+f7buIJN0TmyG0y1WYHANDWSqXfJq1F/VAzfoh/nYEmwOGDqOvB2vCqxgUwO2pnlU+WFwh/xP0T
iYLSCDz61QnUgkT7qXOqjqkqYzO4kPWLfV8L5GatTAAFFuTapV3x2u9OHAJADYq7LYu0kZFoLTgz
oSgrTNDUmxlRgnxgItFVXpapd5wvRZfNvnlxBWUJ+BQIR7mUeBylvYsph9K3LLwKRD2zudmIESMh
nnoudY5AyICCSijRGG0x0o1zNxkKTpu5zYM62PrwnSkINg4Li0WxjFA2htoy2olh6EIYFdviYwwT
pA7EVHiCcqH+cmSj0T95YhgPlQNboWjzQio/TrQupVIp0Ovkm559Nj0mnnsy3WPgxQQZFUxfRHjw
cfHO1w8GzUa8P5oAI+G1AiNK1OlfJIR/1BkIAzjNKrwnJWuLx5U2atF4nGJzWsm22x30eGWFAjH7
jJ/lPXw+HDuczrXLwiujxHHnHHWCOYZ7lQdZ2+opDukMlTEhEatgnFhylLc7wKsZAJp0wRfhS0xO
CFFwxIXg0mj7PKKwXrel+YvBgilxcjkzXJztbL02f1ve5tT+HQOvwtiV4LdkntyyAUvH9tQTfEYh
xpLJO7s712lvCnYpj2TIwQ5kE3nPfppgcy8cD39+LXk3pXDf4Zzb2cOhAr1rtOV+cHrxJizFLILG
D1ThAw/5Gr34U+rCYAHUicu+3sfsjzbqmNgk/V7KXv8Cnhm04p+CMw0jxKQzyS1YIpQHdiHLgIuP
DQk024vSAFTo+WDKjIiCcA2oOu0Njx72NQ6ZJ4tkY0r+veRNaSlAS0oSL+9GiccadM8Int7lYhGL
3nZ9uNTWvZYJozKdX6LGrFnZH/uwX9JMeSVtboIUYh0Namb2AJVZYcsdZbTyDo0RWr7k0mk+zLKy
V0kosyM5eFmq8n1jb/vFBubg3rLlnMqeqkCRyNDORoz7lQ062JkG5fuNLoXBsXuIlOtNtKAkh/hm
4MKERuRW4jHVVITpX2khyjWH2bs+V/bG9JPFo13PBR2rAizASjs+5rS5jv4WSYaETWKuep9x3mqK
A9L9uFcLea9Za2G4lQ2yQWIM6mwKHItm/FAivBzh9lt2Bbtf9ixy3wki/oYMTowCtPeImRaHWR8q
gjUL3k6xDSe1jiR26wt/G4bOTZcTsfvV44EQ3Oy06BFcsECIrhx4hviGm6kodoHSKHjINz/4pARb
91q22QqcjxcXYAVQfN3vAtBmwWaVjh3wsYiG79qa0Id1lcQbXQU7uqZTBQl+OosnKbKQTBh428Be
gqNzWzgUNLyt0kr0QRAZ1LE7SlgbhscCZnB/s9tznUEkOxdoTDAA427BWpGcnRh5WjjYWVnmbXHn
4eYMNWDetxVQyz5FHAR/nIThokFGjZcPFhkLwJ3Rp6eZEybeod4NetUymoKdK8B2n0fn6dZX8P5N
NEih7CiNebv4F0NDuBBMcBwa9JHDP2Hi2vNfCt/NE2LTfZIhIRBHM3bZ4ZmvWcGZOBus0mgSvEpd
aVTzQFLFuI8yKi0/XUWPjMPme528OuE/SlIFIPBZZ858oZx63cdqexGW0WUwprXzTX0J4wtvMa+/
ZwQVp2lWFGqmJYRSdRkY1RpJxiy5OWKJ7GL9/B18Qz9kG5C3Lvbwtxj/cM0fTjcjCObTlR6EHyFM
vI2Vt4HWKYi3Z0Q/RHqXkoLAqY+yCY40GNIHxKSkGCxWCORgnYXatMsABZfzMaa5SsVtCf9OBK6M
+0CuMeMBIGSRUUWFZ3chxPd+auvmMIOszryu8MM710rzFfjJb96k2xOiChHxReL6SJw5IkTPcH0r
TuhvUb3B+hQ2A5bY2wAasCQE5OEMKWAk2ZWYpqCyBrDfj0KVG4LtB9+NWPKjajoP+Cul9HUCHWVJ
2pUI9HRAERASajbtMsfKxnhrwm4niYBamf48DWezg1JLvrcBexWWlaFNwymkcJbu2HaiiDe/XWRR
yTPw4BsC7nSPv2D2H+/lhPPhdtDDDV/OmxAxKJWJ2mwfIoTJ+TufWW6LjHS8r4OgZOdjMpZv9lSP
mrtWUrhjm7FqSE1l21UmtqYBsq7+kX+rUkRLGUVeG5EBJB0xgprRSorFJpBfhCf19qIymzITUtDe
k0Bzq9gw4EWW0zwtjwnGZBomVNVH0c/uRxJiEeiqFbitlvwUZkbWkHt4Fn7d4LBlnZdmD/g8Dxze
qbyoVfez0L9lw0uBWNoSaqJMfcBHybV9lbDlbwPdfJwrjHJ50PgUOloAuEO/hmwRyzYIr6w7cMSD
cKXwxz6nJJ0O6fS1JaQ/UZ7Ka5twUlEAgN0QVhRdU7SIwge4jBkezrI4zejrBUTDWwridRydbM07
ELHx5DigYrWUIchbQtmX0A6ampy3wXc1Q5J5GJLQG/NsLP+GpFffep5tmQCYuaq/oQdH9kqvF1pP
VCrGezV9RXvhGgWgzhR857ID2gT35EtgK0sQziU7QE4+1ZeW/Nfglx3TQfpU2I8WLhQFha2bZFvo
JKwAdjZBLwsRz92WresUUfAkdWXcKgwY5Npws5+6bEtCd60uEXj6BxGffQNX37uNKwCwLNAvy9nd
9HU1jmCOV8jKb2sRdFlYxBZfkweYIcM51wcg3XrvhHJ+7viyCAu/7CEP66kSL4r9jrsxpOaDKe48
e9ljlFJBxB9/spqwlOdzhtQkaRtoB14mIERcPgqeTgR9MK/UQsP63m/1Z4qISqPdxg5aY6lcNQN6
3TmIsJNfkYAGWwVxBck+lyUpIYnZiJ4jVtoDbczuRjKQnsfvEBCB2+tfRWnFgBDuodQGoEiPyk7X
e1orh8IK7/CbJWV44X4JpDaRAirDg1guVGd/04uoSDpF5jK4FmKSSx/rVsojo2bL4985RBQjUL6D
OJDObU/AFP/27Dfoyia0Ts1I4hbg3RIG6p3Ygz2/glVpFW5ED9PZzl6gx+ZgRZS7rUB6k3NF9y6r
956RCrCEXN+z4CQLFOb6lVRk4REY67+vwIZfprNsGJCnAvRCjMXObtlbmTwO45kJ/+wbG7RTcI0D
JuXXDgssllHIWQ2gQKn/1LYhyA9JuENeJ/Ch5VOzfSQP8ALOQHu7QW+oxEW8arQy7aiaeTCmyW5R
By8hWoRfVIBqT8imSHuCMeqELi0H5WZK6UeyZeRYeZ3ZSbcdGYeiFhuvBsRHIioawuNhm+0H4/Hn
ZX7o24zFBR91Om1O8LurDQLS4COipiU3miNoE8cOdWMZfXMdh/a6/mqQckDBKkLcb6RtErMPUPc/
aRd5qdIyKCWflT5Ye7Jyq71hGemQjM4g8WUa742HJfyhE1esrFMHNd+zoFnomVfbVPRy8a7fzA0j
4Q8fPgnFGMk81wZJ99ieYVKrvJyOppIaHUw0tf0m2jNNsk11SVKmneGh0+uCUaNhzV3K2xl1p4WL
QhCXBBzVEVkVsLwE+nG8XeV6ttX+d/VOiKsuzrS7Xc4f06wdxde5pO/el5J5+hfU/+IdFyUq0k5j
wkNBvz6UMxoc7xmkp+he0u8q+ULPAqTG2fOjIFRvheVW7XssGUWQgdx3hsg2rbWrkRjQL0kQVcMR
xqCf1wKgum+93GNCG5lJxYlv9eYCOdIpzav90F7sazjXmBwznp8iBx//Crq1qpnpioy9ZUG55sR/
CTHFZdMNLOZcqp57/K9alr4ik2VgWlP/58DclAswWm1vkXwlgOw8R65SPak/xL3EyAyHkvcyBui3
WEbMoEu/L4PG6IohWMIll9IVq3nIG+3h/9VGOG3oLwa14qUSXDo2fmPUr5KjTxqJbC8z8qbIE+Eo
FSy236Ajf8mSPKkGb3uqMVDV1iouFXTxBd9IVTtcNP5p7Pw/oRJHGFJ5nOanq25OY2XOmbXaDY/i
jncReYmRV80MpPKCVJVlIPEnRWk0hr2LTj0uO8Y/XKtUOO1LUhCTz2OCYtx0pIiOcfGkzbk8/9Ze
SthBOQew/E/7ZNzgEhWwnuTay4aE7ldoHjsWItWGqU5NZBaxSrUvV4qQO+a7ufG9oM4AYWZQUvjX
i5zuGSN9z7tAkm6CTWDKu10Ook4nC6soT3ORZZE/m68TxHPAPSwfmvCphY9jRkJGlALtdozigdNs
lOspS1GtSuqft4OxezF6QWSZxNfkt58enCvt1yrLBVS1djao3GZo0WOzdVCLWU+46FNlzQp/ahPv
dV13wGrEm++LCzMBQCJx+K5Egx9EGCFWfOXR79RCIrxmsROYd3F57fEqrCsSBBT5zSYTTu2opi2+
H1hUt+ip2/7PppJh1SmZWxrXRLOpYInJvlB0C8M/Xr+qoAtjKFy6q3b/l9IV+hNrQp+14c8qdD1s
vjhR36AVhBq8vuO7bbD0vz9eYmzHLbA5Fafoh+OvgEppp6bjuMd6NSudSXzEiu2l3vGjzx11Ih8V
lcLjkWOttUzlQDZQfh7EHnXDbL+M6b4J5PohjaIcj4F0/Ww2zKZE8EriJ0qL4IhMpUBNzTJlGz3b
TLzWtrOWBgcligQbgZpP2z64546tKgQUiYSL4OTsdUebJPOLD6yWglm53YckX73zccHKBeAFsf83
0EiERSX2OlxM8aNZD05SIwL6I/R+nsudseqooaoMUcSar1yAPlnLydiYM2MO8q5fep7MMgG2vXcX
/xyQQS6D+MFgxcDfRHNdlLU1865yElloIM1QM4Kxrd0yfFrbzzP9qCvenhjp1R2lvwZD9HHZGtre
6qAqN97FKIok7W0qKXy/1/V74IJ4EMg7FdC2igy2YVJ5iHjjv5VLlz5gQpvLhpNEd4XlamPfYY7d
JX7JWxOdYlVo0gZvHXyfz0btQstRqx5GoPbDUNT/ST2G3or/db9Nyt4J5KCytjSCeh0UU3PW+7HZ
MwIsk5vtcMDZXPCHT0r1+NX4RUYDDyNy45v3QAHeySGx/VQBZN8AFDKGkrBR+pD4d4TcZ+w456qA
k6c8k1GH8fxZknluqTXJk/8hj8Fj56J+gqRgYftz0RMs9YfHal0DIg0fdnVkS841aod6uCr8ynkE
DGJpCA5C5xB2jVOobvqxFjsFpt02ZXQsx+Dh3mA0zZxH4YCPk6gO0HhB0BMNCF9yBLP65tsV8PmI
Vd9R3qvbe9qngbIzUG9WS2EWnzYtqCPoKl5i+NmG9J74wZxs8zzZaUIGkEGrAFNbV04IzyvNb08D
9dJGq09JYgT7CPy5IwypCj/e80LPCNsg5WBm/dkDgMihiEDXMTtJaSH5nw1T8uEZJX705AjUYL3e
YCxTTqsjpNlBXMJ8p0XHwMHH5p1wfC/7Il5+H9oPYGndp4zeVYkcXAQAu/0h6AebEio8WaiPKxQ1
SnqDYXo/rShzdaKcQCRo9BzMhZc1MxzwZkYXJwvaQ/e91HPG+D0gYUfsOl/+eUhkOZeLmW8pA594
W9p9yOFXU0R6hHpcuW0uiUb6aYnPxKjVUvIjL0M1nkjbQKMHryG32tkJCL7o22axTVNVpuMw6TL1
Zp2gSn80e3XqosRMXKB+oCSpo2sE9/pdfWD/V9zL6nlFTdmGiwvpAhwtKWd8ENdkXuXanl69GPWJ
0ieHqYP/5Vxy6qcLKgRZeh2e0lOBlcXf+bbQAkRHHMW7dyFqmp2MZY9zAji4WZyHCTze8JF5bHy2
T5p8fQwXmz5wDkZ1cd5OJnG7jQ/39FZUmb3gKUzmaiLBm+Npy0fKWuZCdnphJWhbaht1b1mttvRH
cuS24vrTB3W1sgFwtxvXkB2XED7ddIxAHmCvRXz6+hJhNPdwuvzNEGDUYGCnLy/Ly4eQJm15oJ/U
idDDHxOHgWGeDkTA3dcMb/X5wPmNQ9dTX7mEtZpAryCFy+FcgbISnY9QB1qHiBWC5Og+PHFnqjz2
JGDxDQSGl0SfD29cNYJNCGnbiL6egR7SJpVbjaWbk8/KeSgytljn73q7X8sHRDAVVp9sNnICrZvy
eJ2fD3vA6UX+XW85Fw42fTtogmVaRv6/7JMT3y62mCN+RSkhkA8eUDOYapGyaOzkntuOdtGIY8wY
HFmHBt846K/Wuj3KvLyFD4UPA8eEzXfPZXeqEPKeK9e86BDJHE5dJyjh5dnMTjj88i6W6Xq8J7lL
5P/EF3ounC6CMOVl+hQ+qZreR5wI74LMVwRgdrqbDWsiIw+43M4n1cPdPHvooHZwbpE+TRIf9SRi
mgkR7yzwnLU4+KUwe8lpMYDN5ZTRjHAEWxOhNtQ4360kdCQmrcDQiTOfgi4g2waGuSD5hXCtNBd1
H6eoFsjkiB8Pf6OzviUlVOM4ZkyrW+wNIs9Ed9bUoIFnk1tSry9wz3HmYYjsoRKMAnb/gj9+vFYn
5TnznZM1IB7lrUYMkgBn41Z/rvUQl/2Havz4N7O53BRtxJUIwePCVbkYQ8GVo5Y5yVRo7HMu3CeW
E/QZcDX8tklK/Eo1d6n2g2Z9r40llyDA76sjWIfToQ5rKhhvnoO1JoMDtCYq5MjAEn5iWWArOZFU
TEsxEHIjvpe6PouQ9jd2UjtUDJ8toQHXGr4HZ3Sz0hY0bMziU6ReDkWdwabvRx4+qqCpLKjK4AS7
yhMYo9cqzQa2Me/k+GZ2VQ89VXRLv/d3FbDnrhvah1LOO4mrapDnaecy4Bh4awC0uBlPjBHoHl4V
EeeKidsF+WobDlciPxDpJRxMdFH9BnmT9wbCaC91ozJ0EpeYU5U/TzK5jqE8ykPnaLYMu77VSDWG
3moV+BowAc8TDrQHsqmpO1fHTSrCM2gua2zUUHcQ/cgCiHhJCUYxMUPDhk4Arpnst06WFSDxQg/4
4KQ5gCUyASHqiu/KlFr48oVxEUu9DeL9ll+N6CTcYPuAPoEM5wz2oDIk81GvOsU/BZ7lrQ8/Tr6+
2QyL1tvfqzlwK1eOVz/74cd4iedWymt5LSleIxkBch9+tSKgsuqLPARqAYwqLIDrV2zHY1sOktVO
EMcz9GlbJmJGudD1MnS2rQfBL3+8fFSVwsR1OReGDo8mx5TJVPzHL7JMgANUdTvfQbopBsbKi1aa
cRX2HJRwd8k1gRpWIk1x6liw1NC7nMxe4XnPtM/eHI6tgb/7+rAfN7OzBLA7ryuwglHnFyQwEEcQ
/1j8yfM+pSPjAvvb2tKXNdBnTT5trDlBNt7aF0Gyzj5T6hlnocq6UYmelVW5kXEdXC151OCiqcVY
yPwlED00a5oizFeEWVFNfKtkd7Lt81P996UmDKwBnVRkGpOJGltMKZqGnj7v4eC9aWR1+2fT25f8
D/N66ULXSyok4BpsIdyQOB78e2v4J3TM1eqMS5hwOs9ot53LOGrESMj2D+mkNqnDzs1Jga83Hnaq
z8ie1i9tA0dQ+0cl3V8gxnj6APkrhagrnb+GjJhE9azuzI/xP8RMzPymrGEXMWzeclpnugMaQ38N
yRJVbPCnOufKh1v/L/D1/feITHxM00NR2NUjClRQ126RXyj79D+5kAjAGK6otYbtXcF0TfTF75QU
GW3ZNNNLeGGlDT3h4iv4YbjpKTX856TwZ/zLSE+QW4tRzzflCmYNcA2i5InYDTLmV21icdr0kntl
klt4jDKj3ysHqaGW6lhyoEF07yeuDx2hcnCPzj/RXyM34RicVKCjkSyCVHHd0HRN/TGkcIFeWy6K
fTsIF44tyG8oycbvHfFtARaThkkMlQHlp4WnP8fNhA+RsmY5Rucsn47zLQeJ3qxmFkGDsxtMkAqu
+4Zg9AVl22k4JkqRR2H1Z8Pj0n5KYTgotaycldmYrpKkRr/QvFQ1k6q6boM9trp1IpK9qfwl/ymp
ad5K5XVusFP+wEEREiC/8w6X3czC/P7SRSFf4hBfPHONG84XgMsRJGUeRhqhC7sPTmp5eohml134
Bz0fpuv1ocGX70ZjyNLMG3u+XVkU0G7kZQGpMZqUWnWVLlLSt20fwBTTWdHlebtffBC/PUzjThvn
LdoILhCHeplUGjbF2gqxxU9ETwbeOy8E5ug1BC7Qqg+zT2h/uHi1cAHGfszH+fEpW1Kk0EWYWiYO
pKXHCV9M37dJ8iPy9ipfaVp0g5+burTLMgWstDqX/VDK+biJMaKuoPTfj39kLOZEph1AfYVjpFpG
d8+yL+/xsZQN0/GokEg4MZSsATA+9InQ4ZuOrrWPyB4h3WLpc7go1F5MW25IrpSsgSlE1W7gySu+
8hn70tVFMDMuO0AmSyJhxBsjviLLuxa7mTw2k0zFQ2VP9WCt5ipnwiIwtj8ZZPSqvz1QLO9FVu+p
XqoqaEJs13Ywuj6ExzYr5/SiymIi19ODTi6AzXyDIhLGynyDd0h9yHSHHwxeyp7HVQeW9XwVfItq
BxzPl+dVBxucpsvPQTk/1TjQDZ6kQeqx/yhj1kSfBQoFGRyPm5rtYX+VO826QhnhnD5NuvkDj0lJ
ZGGUkxsM5OUA6g7f3501KV/ClXjWaehZyPZ4bW3eE0a3tiks+tnNSmRGA3T+CeVyzKx6Netcag8g
wm3KrnRIeQXModkR/k5Zj3uI1f+JvDkf8MyJszKenyBYtcIc1I8oX9w8dCEKudHEtcgiB7+LR6pJ
l0JBaVxL4IBc6ESW/2aN0Y2s3pBrzdkDqMitHHNilejaZoxZj5kqiALrJI3dkDTcgDfmD+8RO2AU
i2Kluswh+5+kwCF22zdNdsEv322mDSlFs7S7nXumoI7lS6dP+ee1Z9b4s3rHOnbYYxAt7EGq8qSY
uaHiRYNHTbApyXzFCJE41h01OLmb5PDrxGoRneSGhaReEyJRDIqZfbaxRglXSrrsTQQb27VienYW
GYhI5Gpfb5UmYp8tM1z32DSJl6tYmW5Ue6I74GI2FhnguNRoUuo5Oo2+7InQV+bmauu+r+x3lHgi
XdlwpCb3ExczyjzAL1brP0ZEw53CBxgOVyUYBoMUtDZbuzqIbEmOSfjtfvYO/LlfkP+QTiJ85QfX
0T2TRFBotFW05lXVX6twahT9eEeIdWuoiHwQ7tOzWvGS0BR8AupT3g3YYWVeXVTBMxZd+MGrWq4N
DKSaBTHOteHb33pNU7FfF2ufisKlY0ELbZ1FsSvxuHmw9T4xzkf7B7VPr3CMZGbHWEvdQlRytpdG
VwG8btrZCDiLJEcPbx2XxRI5/QmESVfYoNSqPB8wGOBGiHO2HbLKn6kMxKI4rI6DvBrIjSB2UyyY
KUtzFPP5L51nphETs8yD09M/SLHxNHjnB8H620VFN5HSJOF3X3dIAwNmZsFHGa+b1j5shA22jl7w
j08svca5LHLKwPXbCgkLbEbi9GEsx4Lp72ti1r8//ne04VnPkMYS+6cPVKRJdcsYtPZDPstO3k4n
Fu5nojkFQYmdigZr+qmrd5NDljDm6NegunIoM0tHUKu6mZzeqTzqngjzF4gJxFaUThiVJGi/K1H1
mVbF6gNF2E8hSWj2Nk4p0cc6/7l/9JPcrdvqBBwTMbKOo4GiCXm3qlNYhjGzkxzFayIGzvbnYuRA
Y/MFSufEu1DaP7q8GB8M6EmQnnlxSM5uoGzV9nho8BWydfFvjYk/TeP7QzG26V48Mul03WI7Nzu8
0kG27xlSCJBbKVz/h8rIJH8bWg39LvlP0R6/HjxyyRnOeGZ0pOWxoKlld6FEGDvyh7zQNK8XTJmH
15p4JSe8rsjuxjURAM7kkjk/VoGMev7g2ltuTKFlGEWmTnvSDaAs6YVHc/iVtfLXcz9fRp/h8asB
fQcxnCDqp2GuvcZJ0T32XOaRoZxj4nr/6hihQCHiIXafE9akBduSYrRNpCCZQ/u+USBQ//OG0eA8
rrUaGiCIuafArESbNdnl1C9XuiLRUGGpZxB8QnxAbVYKGtAwYx4P8GTWLq2K8kat6SY98AZmq8zB
y5svdUb6tue5cwNWVH3x2bRIftVMNKAyw+fGLNy9AZ4P9o0atnYjFXQi0ht3m6WAJGkIyhBsvBt9
+tXygO4bR/WJwTUfu9u5rZeZWhwGunaf3IW6ueg6/NUL5keLYPaGqFPA0EcaxQ1iPI3v2l3k2p1k
gK1mrHe4lBfmDOWzu1EfVsfCalSyGjKs6WA70isfkGVxq2vATz5op33ovs004edPrdtiUkNwDRw1
f2yKTgqFXgLAhB4Xn9s/p5yBLKx/fSJJXokHtLtp5rHGbXIdVAS9xxQGOH+puZ0AZ8tpr3hlaYX4
31a0nZLYYm1fVPG8Cm9yZTp7zCjp3ICswlDaF+p1APGYEJp+jX/E7+30qneKd4XEFN+YOYShiMXL
+l3nSkHw4p0wySpi0csBOUMUlCv6rGL4heilRRqlw7DPW0cbHZ1hXqnN6at0tLDGyAm9vEg37GG9
WimcCdACSpstFQiWkG9rTUki6Cv7cxXnCts3Igdp6olcYdYcLlQYD/XwCW4BnSoxfiC6vJXtFllC
PXW2wrMT49d1Qwt30jxZAme/XD8v3Zs117BXUIk8bHrYHh7kG6WLP5CkudTxt82U/T58pYd0VlZc
jT+qQPqn7GbeWobyI84fBd0bmUz/02Sma8J8beorXl12NUaj+7X23P+zBm5oFFBztIR6iyZTb8P1
wZUBi/rVP05EfN0EiVCmCwR01cR/Wr8IuipfEljkUfLuxL/r+GXrU+CbnMeEDeqyqe1geOL91BN3
NoTcoXi+pn6KTeIR2h8C3lWkjb1cKnfTuvRxFEgYJtCy5+WubvpsZ9MSFBjjReWXWs281TnPSKIu
U+uCvdKMe0/n63ZQ8UNdyEmfhwy0+Lg0/9MbGkE1Pf+q+WVBhQONyfd7rhQPLTBSh9c5gAtm0+N8
LYjVfJQeH1mRk5UYVaYwW83JWy8wOpqY5ViLRJUUzxB+RRkdzU2X+ouGRWtLAvUJ5P/Ca8+Y8d8Z
oEenCaev+Y9HnT5NNefC3jEgYGLt5eZZOI6cog32Fu4CNqpwvbEj3VT4P2xJvaOKr0aIBadAF30K
UIPFyScfkOq+A0sF0F6qff29tYnuU1x58EFSIVa5QaqbA/NxgTK1j54PRb03GFYU3v/E/Jo9WyKk
jl5HAUBBMAm1rCDXjHN1VMj8j2CBZXzmPWh2TZQ2Qh2w7RZzu/8Bgow4eaB4o+ADcjTC4Sivuhfz
dTOrpdwNsajU/GB1YLfjSqGU38GP4rjSzKP6s1i5OcPq+J1bMJ9Voq+yZ0QWrT20xGVpiVAOBFah
4dtdHKBvm7EzU6KHfVfZ8aiK1LO/FOsyTXKGKIWB/WA9+iXeq7aFp3dbGXQzPuutGmIsypY9yMa/
zcD73KgXYvkt10Vu633P26vtGUhfJngSynUJ2AkeHDXyn1D5v248ojgOLM9E0uox1y9+/FQJ1uud
+EEZf4CIxCLY4YYmKgI7eL21OzqtxRK7AV3acvXvuDfWWt3qJSBNRaj8GMZXTOCBYXUY825c5iMt
2k6qxKMQqZpSIbG2qSdukN8GnLGFHitt3QksbA3M2sPFV1y8GpXBnr5qlkVbxQHrF0DlC/HoLjPG
tZ6CaLR/W9OaKK5qqv8KrsSqRwIRY2ehLSw/iZld7MpfvtSd6hmQWaa7uwLXbjjBgvdBnB8lpuQ+
HzuANKjyQq/CntcOsP+SrGcsIn2I+SDtunDuSq2GNBvfcN0IXmdSeMcxa7PQzCWTJ1QTHeaAh49c
Tl9BN1CfjNpZhKtW+36wHzgEJmMxNbY4tvRLCiYlBWU6eeyjQ2Bwr6+4VwhtON1dq7ndLImF7E0A
WwFJs7ypBz6gi01RaQzk5GYTnF/GctDoTVUHT2sR/pe7YOlYw9wbt8pypQNO+QTKk3gV3BnmRHah
OfrfDrwhrgdE5PAPhd+LnutxGND+u1+se5q+PG1W0cbJ6YW0iFYgBEEBkkD4rLM6oucXUmewT444
ZZhrKWU6JsVDI8+qqqYcfk/HyvxeMqelVmJxRJ1goFnCK/71Lpgm32VIHRlvVrEVUL4ncz2gNL1i
73lx6ekBaqvsbZNixidI+yrRY1XSjfAOaxW9xA/tnVGiSGrwLM3BwMx2YkuC7JExHRQo8LlJrXOg
0uVlD7dW0B0T+grIRKdVpOUE02nPWl5cKJrHH1+fxwkgQC713h6WTjUWSUzMsaTL9aNRi76Yj9yW
Gh4DL6uj9NdGJLRrxMXIRPTKBjA4WQiK6lK2LRBL3QTRgWX6UhcCBS2yyJjceYpcPhtK3XC/IXXu
QBnt3jrb6Wmb6I2Sn8bofd8KFy+uF94hb8iS0aUGyCkBIeNYV0lr/TA4RaYBSXNkL5bGIPAjtiGp
OZAU/I+0OlTmFFxhB8ZWKg65No1y0VnSL3dPfU2Z7lhBPEW/Qf/w2fScp76r3PXgV4E/rqZHHHBg
Y1hpov6JppTAWy48ory/jq+e0QpiOErQ0C9AJkZtlKzcRjQuWMra3XIT2FaxwYbVGYV4IrYyPjQk
qr0giZEPe/40LYNDcDgaTJRFwsyfyfwvnndFJJnHCe9iSYto4/CSrmX0LECm4N9PJIS2Op3Z+QnI
S+XnPz3qmlPmoywwkeF/MsPCJq4op4GdH8n8eZWK6e07H8NxO74LBjYzkUHL1/lgt2CdC8y6sbuH
klaFzua101/RtBdaIOgUXplwk9JciQAWSrU0Dt7gwuMEKA0wEq5zDj33vSwM1z/xNALXQp+01+gv
Ci4M/Dm/ZyszmoGPzU2uV2z8IkaYt7PDoQM1HrZmGErffT4GSMJy9DrDqOVfvJ/6j/plg/yTu4P8
DcX+tmP9ReNwTBv1sB4N4Tm/n3zBifLXxad0zRzaD20Smkc0InxnkNVGq/m+UTQnvPKOwUrJjPuK
WAQaU5lZxvpHMkrWQy6yaRoVDfR3p7GJMmUBXlgdkN04Ucwh3ZBHffjtWabSZrVVgf4s2vwuiRIu
aKiTGeW+mSD7AB619quKtdbWB82i9GQewiBrqTwRVZOS+HjjgaJvxt55KQKi4u9YcX2ZhR7K5ERT
3FoSfYHwg/FZyOx8UhTXk07o17ZvQcZeddj1Rh9ghi6HzDtXH7+EmaVR1cdjATi0wJskOoUisrNl
DVQ9CzYepaw2NkHI3YwxDGH+6wVKUVqoqWbXVjfVJ3/1Yj2iFAdu28rImiujGQHR1vv/ZR7pqv63
8TtXtNTC5B9lIfkOWtFX2+eTWFyTynDBRF/7XehStSI1f7jxZDo2vAnIMD7LOHSCV4tKbRTJ1Com
zF1DpTgK7/7VFz6C1aNQKDoCH3c659O1hKFUnKF5LEqwYRY+LCmwLK43fw3HIWLKB5LHGryPt1Bx
054GP2cYTKLaefe7Ba5YoC3s5rGr1nAby7ksQ/CkIfD8FOX5MFGF0N1OHVbRd7/rFBKvwIEOq9ho
j7e84YUnYgornDZ0Qj9Heq4M8Rhoh7+/X2gxIULRFkYkAdfgmouW4Iuq8m21DhPQAUzGdiCFYjeF
SocwrXiVPR4MDyhPpVBBWX1kIJAESNXVoX51okpimYLL+iIioRKerNTdqz+QXhmy1QfgUxjmcKR9
oRwcExYu8eppQ2a3aMZKqJo+xgFOftdbWkRcck5VZZQihbQVvSFPspbk7ergXaLxFQlgP9dfpwCE
ToQW2gl/ktpZtO/wN1jQboCUKjnRmsdk6exXdBUlfDQrmIzQ112z1f4Df0AkCn6WNxSCBy5K5f71
U4iKEqZEovNhOUwLOAWtUIDmLZ2cmGuhF56RZvQQwDhSPNXZqX9N1ETvdr1v9RFC9AvBAiu0id/K
2+BdEAKApuhOPtJxr/Sw7WGwfYxS5CGSJZpFQMpvH3V7wwO8m2yIlV+eM3CxivKrGsPIM8CAQwji
xDgwP22s52zTU1uC3SKyDn9rzE1agAfHHL11oyoG/EhwytxLVA/hzRzWsMK4PnYuQxKWFLbwPeSg
GIfmm9pGDP55ey7YuApqMiPnIrkkLpOH5zZkoJLIViepCfIAyTw7VnFycpbDLf8lWRdkobkJSIPu
BkMFcyf/pSbdOECW8JFdfcujdYSmQXjX+E2j3mWQcDGEVh7hBYGbutTbcyqvydFBjH/5QBkQ42sz
Cin++eS6xmJg3WsEEBUCM3HWdiX6JHtR/rBGY47Vu4WLA9X3Hh/5eY2q5wfCHaC+lpD6QY/RM+nm
CqAl+sbNKPuAZfNui59EBFizkAN9QDhy52yX0OCMTZgEeykGlDPomURV00wbTHue4gWf3a6AAlEF
Vo3lSqFaP1KGs1FVdwHdWvH/VFmzQoaovnIu/6VFEejNOE4qJwAwLYL/BmxotCfpfo7F8XxVAgsM
dOMKAIe/0VGcUS8C25yrv8a0GgvU0mzKPUQUxpyM7L4TKuKOtWrEdPjFhusxmuluODMGo+TMbR/C
HM1qIFoWjUSVxFb4w35c3Gl2I/kGODovq5VbwxIhqOTWufA8ni7J5vZx7BDA97my2YOvZxLa7X6y
mNZkbTEdjlAfssjYIVq3qAKGA8iw2x0Idfn0gpLkapAuImswLQmmD83SbQHuSM02QqxEkmXmcyfR
dIOOayi4kvaEMRHUU6rijFPCzc032GCcXmFEg9mCkjsOjswlYJ4xGhKTmXgidSknRg2alzd2cnvn
RGAVF/svSXJABXcsj0DCJdC5aC1mpGocxtnGqpl80gVhXnp/Nmcc/kUZpWOiqOKVSQZgBMB1BVWp
0CceggPICqwxrkerDzhRWokOYb4WHqxZw4BVM79rO1ZuPJeoQoIl6S68EA615Ks6xccR33UaCJy0
JksAyVXi9aBbUCbTcBTlOdXEUlfaJZONtM232Ft7MH3+0TWPl8grJn0Q1+YZrt8IuvuzTb+mXHGG
kyckRNhHS4A0sL5OijjBf5M7H8kter5Jzu4HGdk0RiwbaRkLChpe2kD6hiJ/ht7gqJmQt3Ggx7RL
B/NUlfpaN4zoAly7zrk/CyK3aLA0e17i+/NVnXNmqqno1Xtuw22tpGAecskgYSGu7xv8e1CN8y2N
cLRKK5yFq1YY6PgdsxcHOxWK2KtRHIYDc3RP2rRWpCsnmTimStwuiOz8CLJcmXfWf1vK8DEpn3bi
+vR5/fHgDMz6CHDGcWJ5heTOFQ0BxvkXwFd8b9IpSCmT385XzQd7csO3r/9tPCGjOTqrTCKZXUTx
lcbkPbmpvR35ZIDNOZLjlZq6PFbzs4OJyNigkrvwX5ZbE2qb+lILD3bUNIaoY0AESFXJn1qr0DPY
XiiROxgykHZjXvEtLG2ogdA/KIGu3i048kbSO7FjoDyacJL0Qv1eDY8jBz+LE4m0FOnZyRbah3oI
Nq5aacUixr5gZeURNYPUxtp8v/YlpCh9iJyWsOto+QodgidUobxTlCHOW0uco61NlbhbNw39yXpl
ock6+vFcM3Nwz7bebeea4xypvCHSbFUEpOMjVYLoTF789JPK7FzjScQCEfMQXoOF1t8dOTb1cxX+
jv7/2RMWV6LVZGSitZIyyeh1/CZIj/xj5dZg73O1j5t9BNtUhFtAUylYhcyJSkX1LGyikLyodeda
I92VPH6aUqFlNcynk7fkxJ/RuLnT5EXg9jjoQg2X8PfZ92HTVlifqi1drwWA5fUsvB7B3MjpkOnd
aUELVuXqmxw1FciyVuG5qmaPnxqHp7zFIfr088Do1JEGfp0gljefUol40PSwAZucbsA7dFoSWCpw
KV4yCFpt3ZT/SbEkrEoWVAprL16AtAz7NLw8DU786uR35GzT6E+8Th5H4Yx5TqsoWSgkU+2jx9sA
sjzUbQcJl9qRYABxpokaKm6WvNks7w8jI74fUHQrD7sANn7bNqH6RaRfp9egzPhGKyX+qWb3+254
lhPnUXwBVHi6x8rcKokQou2QXNM7G3Z7iB62cTHlAwhy6mZuuYgZjOXAKzNSIhHpI8q30mrVB5Id
7glhOOp5uxUFJwouXk6WHYeGOWHPHNz34Y7qlzlsAgqgVwOzVfISTpw+XOcX2VskPEcP1t2tCqbp
8ndzvjLeW4FqNgiNXjQ+aWEISiVp6n9PO7Vm1Y/BgeojSakbwbOnbfOYmAAjPIvNSGAQWNxNTAY4
DufSzdDFPN7ZbYMLRr6fopLYjgmPxiNCAccmCf8kSKvKrKLLmQBS56yjejN5BWlrRpQlqbB7axHE
4LP0up/gVapVnpraJ/ncBBtDVNMSbs35pFu3rYUYnWhlMg1HEYCn3o8jSJD7+Sg3ZG1S9zK635ir
PZOx9V+Idd7iyQu4dE8XhDV2+PaZg7Y68ddiTFWghdeTn4E7EBfUnhmhmeDg5IgPSSuDkdoSWPC5
1ID158LiiHCJumfilLbzr/T53q+k7EMI5swaLvafEKPwkJhUok6Zbo4KJia43XtlCXp5qkrcrdC1
/elzvfZke1TrlD+hezNea+A7ZgOstFjhWWHj7k15+EVKD8hu6V85J/4JPdu+Dy0I8cI6mO3SauBL
WpecsXJwoeFZUCSDWz6TuGu4kOyzBrID9S0MznBiPsO+8sHhFlO3bjpXN+sytMlYwqIRj9WrmIzK
EpJn49gMxA4GJwq9sbSsHubVNI+pK/WYqWKJ6v6ShSwhwyg5ZSfTD9BzdE4LU5p0M2K8SuYgd71m
yiX3NJ7esuDaUm41ZyQTlrQOSPAbQkkTVlv8tEh8wisP7m5h9/ABdL/ROG3YbOfgfeosn4TeYctE
u3jrUTwTU+ujzNOnXl+gpJL14CniH9N9jMuwevgX4dZ8YiTXdS6gMgG1qDRvEi+egaZP3dSLNj6H
dLU9t5mml27QrFqYubRoqVpyr+Jc8e29aYl/Wx323B9G+5TmijQyn+4e28vGDYTlmcjzwsd1z8Vh
8oycHAZFzp9Oh/hq/iuWBvR7SAhfnwGMg8thWZ6I9KUBBVwfyL6pLb2HQbILF8B74aKjG6Df7heG
vJc1WWhG2oCVK/sJh3hZuirmBMjS01TAVuleHCCZt2C5T4GUhNOgSK9a5vG1dL+oESCGVlNJJrsu
Vbg85dMBKkoy7r9V/NQ1JdyZAtRWVuZtiCd8kV/vCjkIfwZh5rbzvOmEX7pULSWt2BNNJOBWEFlB
IIk8lScf52zCfg62hGlgSx1DjQE0XKsX7fl2uim4VBZPLDuS5ZGttxKsg4nnk/yT7kSIopzQJsfw
iaXGNBM/TLmGjCdW8io3fHXsIUjHOSo+PF/91r2kuek9jiaFVz3CkxCmtINL/RI0uFArg6DeOp9X
avWa8lwlywAJ/X5xO0WADLiP34GEGkvYwQHULECHPA07CDTSn+2BhBDmMF0ezpbw5DgJ5GL6BGNZ
oPHJc2NYL5Rx6jlw0bFbhc69cAhx9kNv7HiF270tt0dpcWhQWoneqlVEAEJNL7WS/meXf3qr3lw1
8y2KkcQDUjIVFEO069m1mnE6qIbl3AeoSr8bO5LQKAdwt2dUX208cvUcn0P3sEAZBVW4fn4AP0aF
WCD7qTX2FKVteAdhXkJEa3LSOkaPtHYwN9ZVuXkeG1NwxevJyogZiXA1fvyGq1o0ZbPsFEtOybcA
VzJz+cwYfr3+ijbQ47Ms85Xc6QqGb66r1GLbGn+k9kWUt13frblbyi5UmEtn0UJNL4uoh1YxlPME
IOUKiEcU6llXWDtmbTVQFMfqOtnlNI6zboxvGNe0ebsjG5pUJmkSzWgfWIUbKNzAfUZFLgEt0ZM3
+tbIVQ41S7cTbpaIy3IRPUZbfaZX6BdLdhJwpkPpLVv4ZwSYSiQy+PTh5ouqi5wytDZ6ICpnyu2v
8Dc8d/vcqqUWEvpYt/gWeVGuL6KlugaPCiNqD0jEkNfPUon7RxgSb6w+eNsU9pH2aRqmnDmeAsQC
X3lrR0b+DEALr5YK8kLHhXbUVNYLwr+9wAMQtZAb3M24yR5z1dXySikkMi3DkUZjY0v5aesBK6k3
OY6v3MzqLHBq5uo8CdAyfENZV4oaedubRaIRHoLqNWpiBFQ3a09EkU1JC1QGS2gMiOz95+dYedgX
am9q+uvbiFSJ8gBqSWWUzRPnehieJqH8nBvPiHa/6ge4FYi+FfL4t0K1Tsp2VKTduo4dOvPVdYeS
UQL6r8TOWuzisL5xMJCZ9cCQClVcSugA8MpOHM8dUd755EQfUXgvCIDsm+kd149+G/WtREsDBIzp
U26ZDoS7f12nUlgngGouo6JRqZrSy/Do5NwJfiXeKQZzDVLMe3VCvgu5ip5KL2PsOBjyla8I/ohh
zIbg5KmS3EJVr6cBnQyx2iPwKYdMn3k6AyMeVNutXiNkDeTL3L21Q5L4qfTr3prW5dcOPVcRkz/D
VJBYhGNrjsY/AycdGC3eWocPsUZ1b1fWz13R9l/lV4Rq7X06VcNOqGcYs4D/a4gOj1vKSteaZhqT
5bsMHP87Wi3Uvbrm/eSoYdT+J5SIz4CJ0TB4+0e7bjdLs4BJgTDT3MS7urlkG5hi9aop+QBCJPQQ
3atAsFvhX9ugsD+22l1jYiEdnc6HS+FNuQU1ssxkKUm1uNXLCvRO2j67YRwuTy9DRfqc5nPA2Fgl
P7pUsECsFK4jSh0JimbBVvH2Roh3dWjVaJBbHgp3kqiH4j2F91HhgwjfR0ZF3iCaH6SAXvlgCDX2
z2HRHrkascgc6iFbVwLB4gTEycsWQKOJ/6uAs6q55/4QRqhcfMWAKdCTvosy4z66LU7IkS96NK1d
pdOWNOz9TK/bHnQwAsxP57A+5sCdAjIYiJyol/bh5JS998nPwBP6CuItP0mi40iiyTC6oIh4Ohsj
Gg46XUt+pPsCEn+kjlFopBc3zQePZRShvA/gMvlWhsPbIBrRAOlFYg2+8bFVJdEt3wovjPB2TUrS
kkDp2OHNAYWg/QNmwDovr1Eyf4dddr50nr56rcnUCgZixFIoluwOfQ+nQdiXk7Cedq/NIMx8VkP6
R+BneEsvIGnShTHWFjd1AfAlTz6tkPToNLoJnw/ViKm05+nugbqv4KvC/ETNsIxXqP7/l/mAzR55
/2G/f0J7zeLrLvGCIHEspsy6UhR862udeNz/yMn7/1CnCwy6OUBqqyoKFt/VZEF85BtJEuzqT/3i
qwSuIqbPn7+Fecy4PrTB+/HJbdTzBgirCUEVhUmN6c6SfaDtTwc0og1XYthC4ybjHYypNk+YyX7h
c7GBXU100SrFTqFRdyQZcuulmoRdthcRpM2t1bHgYRL8I4Wfg3AoCXvq0iafa3JRoKW69ise1abZ
jhkhok774SLHw29/23EaOYNs2IkWIKGuxQvrPY+Y/fQCKIvWAxeQu4/dCp5W05vAT28xz0J3Hoa0
H6e5vivy5ielShvOSGB0TBYyD58znuL0oKsqWBfTaIymBTTQMQJMMBF7mBYv7JmVMvWLpUR/KSkH
JUexiV+6YGaslO9nFidzTqcFGJGbQMjm7aBgaqjcDOwWeC2jyDH6Ssa+758ROB25nN2L4lZJrWOm
6dAgTMiv35iEahqrcTCmKZDh7KPq/DkNBEgEMy0zKHCp0Zc10ANpsoj7Aso/hYxp0t44kQPZKJFc
EYkHincXiqscX7NIaDAl9U8kLbBqcA/fTjSq5OdlrfIbJpT7RgIs5RjZkVfSnWpHV5RxxfMN2U0q
reClte3e94PMiu+CJmhqqYAnAv1KgmCoqQfLNuufjiLbgrMjRyblZcQ9p/G/q+UevpyC07GpOy2Q
cAgPOjNjGwUtIltu/LYhTOTHjEwuVV4ZxvC9ZehwL0/khUQha9DJp0sl/n5sPrExuyWT1ZeNaLV4
NvNgHsvulxThEYFs2bmSRm62g5ZnVLVvuFnOAgq2zRsmUEJZYnRyr8J3QpOo0/LcblvavaqF9CQ7
89xH9mAxAoyTb2ZawZ0+Ym9n4wctPQFjsPA7tYb9sbuG9TvMuaKxAJT7QHl4Y5JRVw6x7fLAZAX2
FnEd4rzwRuwh9XIWqKi1hl6C1fkK97t+14rF/L5qWXL45FDwY1sDDbJb83t6OumYb8hTNJdHhdsW
sPpOwFjGEK/I3MkTS2TF46Zd8TRs3D7ywYsxfhxQQBDr8iXbE/wOO2MlHyy9eq4f5cerhq04O4qC
V0GwoWWJgEC3kFQPvKIYlJOL0APJ9Tyzm2zyP6Q7aCSkge0wy7sCmMWAYHabxhdd1SS4y23dO3ZP
NdepdN9RHqqxyYhc7EFJCnD0Bz8rNVzI2yND3DZPL4QBAxpWS17s40/0r90oUMdAMu/o+DSMGchA
LAdVO8JKCTUY+L7oKPfwxdYdcBs/rP5MEWAasTSdN7pgvtKypW9Rt+5hhgTRyuu9HwwF7YBD9lNG
mwDiyXJH13L8odagADh8FQyvnlMJ6aN0DZMfWQm/HN3E71xz5D11QGhg3yT1fXnBYE6VwvaZGf1o
WcR+CK2E3EzqsZCtv3Oe8WOZ5mBiEU+/C6xuVra5LJYyxZ1p31I1R9spWRRuufvIzF4Q2N4SooSY
HSafX5VPzAVokGrWeeYt4iHQPMK4CCa/hOVr+V9dXdZjETQGiTdz/AfUzBo0/X8gkWIgNhpjoKAs
pm7gQY97cknbaYvY1RY58f13wG0gR5VyvF4cccpQpYISZqRd2ckGm9tRhHr0Y/j5mUlngu2LF35L
vIxAQ1niJUDClnYUCWjIzVXu/kFk7NPSRHTg+dxnQtGMSt435GwmwMcRxoSI4B/TiRIh84ItXcdA
DDMi6DN3eswVsjbaj4sylka8Rg5BnFw1rSEA7q1GNzfE4GVgG/Ck6uc+dAlzv1qr1AUhl0XVAn+i
2b4B5QLO+5hipqDhkfWRsN+xi+hBhKKiHtbiovizQKbPCNSarwgvhed1IN8Qnbv4YhKm4CKtSc7j
QPRNc2w+WKv/ErT1xXP+lxMXUNM0qhi2Si4o62CIxjVNkPCzvshNLisa3ahXfXHuaQn5Gdbxp8rJ
ANsLsIHlEHY17qI6HXeA5ARHjm3G6LEInCKz7TnQWFfu+0okuu7Azb89v4Ycm/ZHqPrTMPkoG24o
mLRVT1lvIPlaoy9FMSNBPcJGxQomYbOZ8ndW8a/kl/OvzHVxVRjeL4eduOj4j0bxnPbSJ530SKIT
7nw9+5TR821ph4oSw7VfghZxD1hcTFWm+pTDx9tKfC5ZBJevAQc8G8S8uUcGfa6Iv3NKC0YgvKkz
S0Q8ZquHfB5pB+9ico73j31TLNMEgn70d8l9/j66/uz3SLJ/aA5kDUH8s0aHpARjBsfC7JKhvcBc
JhZUNdtIpOTn4/+pPx8SDlj3bSL0KCpG/sS4uxqk2ukbaCoTANdZ5WZIv7FC+7uEwSSt9qp+N795
v5VseAoVsuCzSI8sMJGq2BreJA3ctEqGECZfV5w7YkShfBr5Xvm9oYUUsbXjRcS90wxmj3aUuebE
P0tJEOTzPG1+dVC7Lxt60QtGjkzGaO+veQQ272h87WDPrnKOfJMFmqRS6i9Omp+axUe6VXsrlBMc
8FWC+aTVN44P9mZR2UMDEuWmvQVw18bkwYea7LE1p/nKRcj52QUI+WXTkgok1KxbsjM9IEVTEvR9
6Yofj7+H/fTAuKhEPP8V1DGrxPbFrqzPPngvfu+LxDzh3QXI3QQEVqo0o3GQRRNpfZCpCjb65KA9
qjMlAYDBLHppYg/ZtGWJjaRFHF/AiWBppKzh/0ifTyMVOVgfMV669InvZqb/AFa6oRdgiVeXJcdM
orHpi19Aqh1dddb+6Mlmv7cIXaWlVtWoApcNe4NclkJ5cmwUFpUzLHqDLStl75bOyPq5gd00kj16
Utxe3zlHS/ZZ6407W1O2L0cDdf+F0dHrf1tMvmz9eEErl/KyiSIM6ienQId6XSIL9mgquHErXbK2
/GkCN4GNgo1XtV8qegl0xmV5Sh3YIfI3q/GhDdh8ihwFyI0oveCVzYWNBNaNBcq8mBVrPK0x8Z8M
ihD+cPQBPMiP1/5gcQEFIxK0/zkHoQm1/4AnKiBHcL4ogbpKFlhJB4EGwEOJrRMyZiTHn0iPDQaY
UV/DNySycxZIk3DO9VjT7rnk2mEg2KGopz4ihZ0gQzNW1a0lkXaTwz1aNz0fqpzG8QnuFsOj1nN8
skjdcG6Ko/9aIPfJueGx8PYArQ+D5on481iWYiKFCqUPNj8vglnAKuo0//QV7dkd2E2P9p+PhE5v
CeH5TqZaORcagjaXD/P/ob49q7Mz5TEK0QCH5CSZ11cBK98am0CjDYRtRpf3unkIU2U8my6oICrR
ggEBwEzBbOwlLcr4h4WKe+IiA03gTJLq1n958bxafF7hUAJ/XzU0Pnp+R+U3Xl48BKcu8l2ldOQg
LgfA+cuN7KRvmIQ0RwXiJWP9Tw5crIiJN1fpMx99vaRV7tDJQvKWJJ5MExtCyQTgjT5b1l1jS3Bd
fegHssphtSpJzZl3bzlyIW7WXzZtcwIRtWP3hE65sd0u8plzwYIlpjX/+vjVqmPV5qq0g5jONF+1
113Gl7sE4vkJBmKfbfDm9QM/fZDM7lYsniU+5WKIMtUXEbp0N2Cr7jgDgDZXqsdezhBVV6yD0WzE
QFN1cS2Yete0aEtuENKoHhJFYRkCqtPMyP5ePXgovdSiW8K8eFcakR5/bqKeA7QXETUkV7A9sHTY
8QA87E0tWCnq4wKyx4TYY7D94CINUJtFEzxKOQGmUAoz8iUd5lLm8874tVaQ4xc4Qu3Lip3IYywn
ZIEPgXiCPOvR37t1C2hhhoQDeB8GGV548OV6uPrS/8DksxOWNOAhnr5YD+uvMgDnIN1kQmuxzdOb
9iUkT73vf0d9Yv05lIG3HTz7+FQ0K0XP/WUQJkLj1stdjWFC4ReAF0iU0FTNH93L//nRAgTK1aCo
VscvExe2bu6iThxM8zdW9iwj9fgEWm7knFmrMr4Gv/w90Pf075WJkR6fj77w6uIS2TfOyc2cpnAC
/W/3k4i3MB5/s3HX3Wrmdbku6P3jO0lOy/D1KSfEd4mUCxyHJDsAtnQqbblDyx40nsUSvfAixxzX
GMOw8eUZJlipJhy1TnfkibFU49nPUq6EDjGBYRCBAEDqhyDTYx7p/+gI3SEZalVmENj/P0f0poxg
OMpx+pPKny8krxcQbaA5p+1cXnyfQXLzLfTwhB9qJRLuFZfZeh3af0/YKqPFlIfH+LUfQsX69Lht
LRB0O7zlW6NtduNZ+6angDtfbjDFHOhPkwaaMKokKyR+tqpreXoYl15AMtkauAh3fIr/3gHW50Al
ScsQWYybp/tC7RXFQylsZqDuYtvkMQbBFASd3DoFTtIFkyO/+leMfZDiSWodvRvY7Zg0iuhko2al
ksohBjBSRvUJJeDCn3DZC5enGc71IK4C8L720fFipYaJrwVRNZoZK8kV+D76EjThTtrYRRQ3wdmc
/cQjHNmwacnodehMEQ+3GrIw4HpNXkgqgkvMdDDxUMthofvH6aYZzvz2wQ1c8jwSbeRQJ2aF+UqB
6n8KzwThOLIUIrl9hB3BHuvMoJnoZZU4M4S5jKbh14vpNZXfqL0eZpqw3JkT8/EPJF5GxT7qOlP3
Y/jepRmPwef5FHdX7jiGQ3ggXJgodGLp8aNQkN32kcuXh1QfKUbIbjMm3HPSXnSDiEz2miTL0B3u
SwC67Vboiu9BQecxRGzVG/dPY75h222fMWek4t/uwAiMO0cOSusMJp0B1r6A9yy9Z6fBN1d1rXT3
8IzQy3vgDzxAkNkUU39xW8BHNYFqMG8QpLYdSGXjFs+DL+TxW7Lz7DQXmGQlamzXHrzx00QcXG+a
/iR3gO8Fzu0ubfcURRsrG5laPF6netTQ2jtwGkGYVK+uSz+v5Z+/riigmx0QAeMZ1vBi179w3RhO
XJcEUL38xoSikFcR4cnXQbWzUzML3qLFdjqd5+DW/vpNI01U3fbOi+OG5hH4sUMVinQyNC1AMc3X
nQw3Pk0EFva69INP/TBfuWe7/ZzhOx1803CzUq300eayD0ehEnpdXL9xNON8/P+VulKCQ+XSG7zO
7oahnzYj46XcvTxWDYE5CaSm8shKVScQki3xguxcEHtuFPzdwtonA/nEPutuM2cowGtY0E7QNXmQ
EiSYFCGNvEON/rI0TjkIQuBK76DsFCnryRfsfm9Ww/JjBHtxSkuw4yFdExBoeEYAaIfbJJaa4JtD
OXq/0YSf99yYdyjlTOB0gZKtDAIaNNCU4xwGtGFCUl4irK83bBgxVew+3vI47LmW1TQc+hsdiT+p
Tblpm3b9wzg01caP3j68aO9rQTpq+wPaTw6VeYkemEj1rhvxsc4ZsolWglrfjpU1BszsOHVXGtAO
ErFhGpJT3cgPrwx6Q1B4sNiPJjmdQF5to/yzeDCb4mz4HlnZNrYhg/DApYkti99RbnLmb+tI71iq
tskEsX5/dp4+Vj2FwHtUOMtmB8Q2lOZMZNb8CluHSlas5Cm5GN5XA3OQNRnijKcmBBpIyia2DENZ
i9hTUgGNVawT64Y6nAyhYAytmUMthJbdXwAkBozgXESnTUBQG6FbeIvpRffTFhhFaMlRecrCGjYe
0dekJZiAICmkRRk3jLYFtifMuw4jzPRzCnG9l3YDalfTiaUj5y5Ct7H81B6AcskmjPD2sIjcXBbS
0UcnMkBIlDyXKd7zl6lWNOyeYP//RhH/aNY+CM3UlSCigjYHrsu6swbllwAocQ/kzEzU9oUs9kOf
diiUGimduqVvdu1llVFwvhNp+X9zJFGNCkj2lUJVMl9kIKLbMoST7K0AutRa7m2DkDzPrlDukgNE
GItj1iDkorsxssmmCSfu4KsuWxxqPcfZZGpbTONl+IQJxDZIiTDUDnx+3c6u05lbF3fcMmAUIsuP
MhOIJlFEkzQ3UcBqlnckBcPXYT6LnWoSsN8J5/rzzIwxG3yuti1m9W2V0ePF4kYzV+NDiBXHUNdb
e5E7siRqCOci3Kj+s6vZUnoTW7X8iQ2pFlRpLy51Etu/f9YAUX0DH0hJTsIfYEmzkB6U3ZrEdUQP
jMLMLN0jE2DdIJuR8RQ06fYF3S27KFBkH/lrKvLohbGN5CE2gxUUB1rj1MXtGlX02YOrYh8EMb3N
qz28704AXUQr2HxuOIHPbxBRTC0OZ10T2kIs/DSGqQKZH2cM6zQrrtvyHcapeNttCeIlY451PrxH
wEYwZuKNGY6ahzjCPy1bnFxfXAtULVVvzhklsUwfhH53QrlYSd89dX5FUtIpLErEtH90jWkV8Dwg
bMRoKl18NVyameEIPkvzWXhXRFOyWYOFVHqAxOxpYFsR/7wN7906S7tub59jr0IhYf4Fs2LwvUa6
oU2z8Z1Mux/itDoszf+4mHyqCZL0SfZHiFbGNY/sQ8I4c8Qxcna8xUpQK0kq7YM3+4UZuyvOrjm/
UDVqEpGw6JGz+bbDXxrG/qqEDuqfvb9FE6YVfvJ7QdSvaX2FRR7W9NK6mOYdw0hItiZWNIFD7DC5
9M/cD/Abiko2JIMFqxVImjkyJ35qTGpRStO67RFkngHLy9ioJrOVU/8l6y9/FHrvaGCp+a8WJ/vR
HBC0zUQ9m5/o7SLIR1FaTj8a6YXSaXGZ0l6Dj8RdaSmsHe+NxG9/SG2I7SvrKDJxTiAlswZzybrx
VRKdw5m+t95Iv1h36jUlQooNed8YZxoRRzIlN4H1Ex5LykdpzBQUODLrPxS9aIwt5RQkvXXort1g
Jce5MDP8+N479nUA/RjFVpuLN0VbsQmg38jNFBbgkLFstu+Fo0eE9NdpAJr14vWwjbeBVb3hfeMs
l/oKaEHhE4TFYCqSU8kj/dcL7L4dfs2inzTgxZEJSU52pAHTWzqcJmOTi5RsXFNg3oyNREIGl6Ju
bRcgbNiRki+of11UyVxL0jeAZ7anCNBub4/oWvANP7W5Tl9SQOaj47rqcvSWPaxCeNCVT/DvO/82
zQuXka871oP4HeEeGtftZ0PdAmIxwY37gwsb2B8FsWb2Ip2efEYbMm7gZiqMYA4yOgnXjp7ALILf
ht1B/1szf/iXbdQWp6/eWygfVHPd6MvlP514iRPfxBDDsmigNGhdwZSTsdAcyy4Gzg5dBCP2zR6w
KS7RYw8zOMAKMElkZkRpQEFKq+pxN1ZCpJi1FMEbacCvyr5YYG47cSDzTLCedGvS+n+//bbHNOe4
DXkgv2iaQuOkT2VMk8GAj2eHPoRTHypOptIBs3ah75ZYc1nKl+fN9uRV9mIsNijF+0W+v0YQXgWs
q6oNiEMMSU9pNuIV57rCOx9TK1lFQ/y50aO72nSL0rmjfwYKQfjVhRmM2WDy/5SSTyE94TCTBjzd
0kPH6F5jGUDLhvDEwzvNXPr8oEJvLudZjMBgPb5F/FtfB7DvzxX72/ARQq+maujh1i6ZSh6oHkbi
kLb/rpj1XIeSu8PAy4tvt1NiL8XpCJ4D/JZt2soSa71I+vwgfdsMAvWB3Ax9A2Xm/GRvqKcqwgXw
CC+qpsPFVxwrGiZ8KF17NXIl2uBCeolexXLjsRfscYQP5Cu9yMgKTOFFDaWgnD1+fZbcZeXTxSnt
A6liKR3Ckhq4nt7ia6oNUVT7Hm6pQQ6DW/t2i+LMs7Q5oScrjwUHOws/+3xvln8X67FzD+CYBut8
BKIIhJzIp16pc1JCfgJWH1f0KUadJOyHr2xwTmhf1aLf01mgY6aYfCzMD3EFiBARVmpi/KGO03+4
LhrQwCe6QICC6uPPHxWD5YLcN9TIEOVlVHQYXQBb4/JWTxsrKtylvkU7/WzFiLebatJLHm81ZOyU
ds0AuUdPtTNburOaBZ3YWPThhPskyB8STR5E0Bk6zSeYUMn0whwNEY02mAX/6V2PLQvWGBQq5lja
WvGVL8d8yp261GwBHEQ5fmqi/PJQK4Pv2WyltRriDDbi+oIqGBw5aYDHYO0UsYu+ykRdEDS3IG/n
Qi0Z+lrITVzCR3+SfBejK88wtSKRm1Hh9LtQviiMuY4AgxruXACL3nytfU4Nq1/4JyfJST5YyvKr
PmNxygiclUUUq3idxS61fGAZnnzEF11N1eevdNFUMIuTiJZHi3YRbOG7uYH9q+wvDqCvNb2Agg94
ljXPVYhTR1F1LIiwlV+BHEFr/l3Jxp6dASzxIAK6yenO5hsePBJJN9N78EFkXNANawKB4FBI3UPV
plnaIGddAoTHkpcpZICGK1sLhNcL71MiYQk7+t3WLPjC76fnuY89iheN7bT8QPZAVhg+E6Bpm19H
1iZJKxYQ3syVLBom1O94+riFvqzlUFWjzzSpWuK/T29QCB25mY8hDtjyMVr/XNVeRcrUQcCyKM9p
RjerJmJgxjEXPoSUOmLfIjbxHoVXt2t5vVGXMaNOWLdECDd4YT5FS7yIiC2Gmr0KpcA+NoiSP1aE
HVV+s5I+Ld7gX+zanv1Cc9EEseLhPbA5BD4qc2WdVZwj805xKsYCgc3IP9nFQd9rDgDUm2GjlxBY
Fj0EjE0TM9H5PiIbAlX9tpYjTzbNP0N0yrCBJjLtV4WtKwgpaoIAi4dGdCXSRPqBT962zz9QDa0d
a65rXaxEzWJhSHGKiu07+wYtm9FJr80J81JgajZEWBHh8wSSQaiuWu7VbXKdq8XpvIKm9T16PQzd
Ojowr+Lwvc4ad6gseahAL8vIyjJoG2UVCadO/KeELTAMdnAqx880cV6oXjhXO7trIA2Y5SH4d0/Z
sHgj0pvJsBSFmCRpwywMqc+p8zsDb6bX4539rfVriJ5UA2bZHLJMMuh38p1LyA1e+byxI2utHC43
BlBwkQXLFFt6gq5HlBOoJc1ALPu6FhBKJFqQSLwsyNELetn4XifSb+nfyYKRAgWgJ2VaqbtHgHo8
GkgY4po/BAqxzbE88sWfeApvVtaBwpzz8KEBM00sQDzEdOba2nGnacyAwuCv3tuhZZuLtI/nh50U
oknNuvy4WV5WKgPtyXg32lML2rcr5fon0BkxxV8tZoLXEhFHP0WLH2b8zl3t6Taheo9rJNo2iRC9
IGJyw76WWKh6e9mbCC8MvD5prl/0K91CjSlHhP7JkTNyF0ObbgpugK0huq0I57vPsKL4T8rDG2zN
Ie3V5i/v/HeIIUlP2Fj/EOVJpUIJgki2ZLGsvM4ZvEcFnv8fNIuAFICDSpuMPveGdlRqKWkQYluK
cCg7vKenQWy2SIqFdLEz/9KfREyQ7ka053AmzLdUkGUfNcUFU7BEMNcNGn4aYWqqyZP9AsFSLxJi
8nwRGi/0YWUPzGyOy1IotUm6fgHqzlymQLve6AwHwuQF4NiVNbS7NKAsFEbBjuREvLOj9A7+agfA
7/ShqeNi5Azc5u+r9kmAULNHHFUi43+JmcF5g8T4G7NtxJFPhojqUcgqIzDM7V1a7KYNVXM48kPa
bd9sjEqxaKgzhWve06qXEExi+/uh9IpQWjNwZUvR7mcYPUwRLRL/wTjOl0acauyL8AFZbLmtCFhN
H4SL/UkkI+OrcvPOT3es4GK4i6YE4wn7r35X5h6ef3u2r0CngGkz5XVYkA/tXMlGT86lYIcnxnBH
oc7ObquUc6ep2rUPG2wDibogxHPG//GjCBhmjgEo6BhNYNXbMbpAl8gqpgdgQf2IP+9w5bYeDTyB
uQ/9dCtM98/WZum03kh6Avmz9K2YjHJdSeRKphEISaAt5v6GWjYX/3smGF89R0YbM8jq5lEgkx30
LOZblsUZPV01StXOV01QaSZDTn4UpnPa6Vj9hNHX7QODoxLcewdkZpSSKSE8gztP4vHn0n8atXSp
16TobMPoiESA0D0+MYq+jqnhCuHxAYpSAbSHB1ZdqJXyyBJ8NIqtfBrrg0RXHigTQlYgC/R5QcKE
itoqrxlgJpCY/NECohCUqqgrY6+WsyIkQzHOPyalCJYio7q2/F8v+cq5Fa3cIs18mYPBNEkw58iF
3FDCxpbIxKm2ObV8PCHD48tWpiU9lL18xJJCOLGP+RxvAZQyYkg2amMxEe3MMVjfBrJAHG6YlhHD
3Cx1DTAUVFHna9E4GDe7x4kTZEc7J9GixGgbuOiu7MvGA0vt0SsL0r3WZpveLVct3l4hQkMTwprI
GvOZxfJ7Q4zZp6UwPKKdgcPPQoopuT8FJH8Ek8FCx24ox8fP2WBsyYeXYR+uNLfjGr34LVK6J2oZ
9NKfN8ynSI4Cs9a02PPHyYg/bQsxhTepexKo60Bk2jz+aTnMmSS1VtPD20ld97JusBbXLL5cda+l
+Y7GbO/zE5R5lfFbKns+8Oil2T60VNR29kR8BJDgYipigbKxTtzqmZXOisf8caq03ZmAo7JxBMRM
7VGR2rLNwmZEtojqwevF0S8qxtGxdLm9W3QK+e4fcvUpErnV1OPnbmpz3UovQuQd48XP4wAhhhYz
UMCgcoOaWqpgJQ0BiKg6ZlJ0d356g2LRAeAkYbP36dyYTLfQ4SKvjannMNzIvy4VicrMM7+akt+o
Z5d0eqHNnqIos5G/pjOSDdlVnPtLUH0ZQ2mx/atdO6lkacH/24BZgHNB9/deQSDAlmiGiGNPtE3v
Eh2gxVPbXYvPVnRRxkg2kYGhKow20PfGq+ZLQQ0YAEgGYLLS9nG2O7gGdHc9B5RlKfwvDyPyAGYZ
YGy13f0HHS1uCML94QYhtrhmoMu6vemcSTXqL6w5Dsq+b015BY3a2z9lH/vvzEHx/q4cnJwPiaaJ
CE81VE2bLinHPMo4/I63mxRBCm8eeTGU0jqq55Wo6MFaRUqQ17NN+zZRliY1K0W8MNXFoymX8VOL
S4jt7DlHTAYTAfgKgglRu734D8lj0HWMa48pkAxB26GiYQyfIhHmQU9zR6v2RXT98FdRVU9s/UbU
gpnEad0w4yxPl2kVl9k1saYEDnYml7LxE0d8fbQco3MY9sB/K0lK5K9qd8Z0U8PY/I+dqdyaKT0B
ILjolWXPt5TFNLMK3iOTGFSHyo/TdzLRX1iC+EyO4Q8Ul/JT7LWGCRuEhzOEbJBwVgjIhn24Rcyq
PJ6TFkg1P2KZOSjrrjesYEj+KZmzHBnT5ngP8Lxy0Z8tNCeCO1vQ0c6jpP2DEhXDOiZWPCaWAaxX
iOmZqTX1zicJmig2iuroOhXGnsBAXOexGs22+GPmRV3sBoSBLTs9MBkqwhVmwIIfOH/x8jzwezXM
P6y5yWi3TwuE8qisFzqKI+S6ZUSuieAVENgyFDFQjI6VuUyv9tSjmkUlo3I6MQuTFjTBakvsDIlD
cEQsSkKSjG467wrNbZdcfhGue6QD6k9Rl1F4uP8ITf2jhpJsaZKJZkvCXVOBRVj1gHBK3GbjnChF
NcQ/zr/IhtZCNTDf2duVTIqmZlkjobk62gpI/H28wcjIiUm4TBLdVlyl25Q5qn+G+MPLq/dNos4x
QUgALe5RnQFPubwFszG8xOWG/l0LiuoZufQJgd1VD6EfkQhrbWg6FcdWE1U4th/MG7/UROtu+UUD
twvZk/I4jFWTbpZU28hrwF+SutE1LmTohnBNfh0grH+d4StkMGX+iRdacHSnslcaEf7vRAp6aZLN
hlxHmRS+b25vvhO+iZpe5tCAqETxkX3Xr/4J0ZX1DvBbVtC5t91TVtx74V+2wZqfsTEzXNIBEBdR
SDiRS6FoqY5UbhNK9sdB8R+9Me7+be8cqtwKvaMOOJz3p1iRN4S0+Zg2DVCEjL93gsp1FinYnWX9
7sQSj7S99HBZ+xqC+g/EUvcGbM5uBdOXosK6+e8VNmrluM4A9w65LnbNLkWd36pLNNNEttSL0L13
vnOk52n/ZDzT+0JSgu5ssmLbfsvP79timI8Gm1/dGn8/toccka8tnSEZLZJ+nJCDV9fZYrHsfZO6
nJJZIMzOp2uE3ViPKCpxOMxyDbwEx7GBe/X33CSewH5yrojMTgutKuYp3avkLbM3BJ4GpFVsiADS
TI85Yul9SU9EN7Ys+0tKFGgJnkqgKuIXTyHKxT/XuCKZww61hcqPkc1AGCjbitZFAMK60CkxgZKO
aH74Lak0+Sl1AIiPRPsEWnAGJjeVf2ynRx/3tvmb0TvnJZC5ZEPO9++FTyTc5woRpfQLLIwCjP8t
SO2Ho4sixy+n2JspqyrVJsgHLONonnnK7rZdv2WzLtO9vzi4MvWWH2N7yWY8r1vDt8OGRvEt1F4R
07WiVN3vyj1aLYDcsMye1QTx6G9IZBA+JDbk3MN8Cbe/fDB4md8Lnk3N64IpHmhpsJo4xADGRVWp
2Shw9AfC222147PL3d4DISGgcDbvpN01TSuNuwAuB/CLt8JCX7y7WbhxLwY3Mf15HsCuSPkvL19O
XBbJV7Lm6WnluwV+1nT0FmQUCPKMH3fmt0f40I9C+KvAJQw1SfTJH6B1BxsA56XzDGNQ06h/RaiQ
KPRaUE1W27di1jUVVoWrtvUHtCEKNGGx3vmF481QTNso89M2qQDx+7rGCYHSWiOwu1fuOGwR5en2
Z8amt/zcUQn/udNheofaBTU/skSugPgno/72SnsbbTZBwvkzwJLrVSSI5awyWYnlmZqnHA6jOlnJ
gvRgkAu5z36OCRYPiuqjMyXPBgD8ptwpk9hDgauRpS1RWqwkfs9iH3sn4ipJshyVc/xkagSR/K6z
yVNCx7siwrwDlhzRHGl6AbQJjMP4D73aIXH+uJzLnwkdGEHUAcylL1/vOAXOT6qaokECgWsnrZsh
UPPXORsU4XuJkN3TKscrXTDo83a/39FlzknIs+5AD9Gkwt/JrWeXMfHW3uqDsBUKsSCGb1+a2eBo
I6xx+hYwp6R/p88hJXKFtT8HwwglsUzgfpDC3nhf9ZyWq8hUsgFUSBRqPOS2wAt5UhoVfYGlrl7u
vzWdIY3V5uHbmQte2Hk7Re2IFVehv3mnRkc0YvTe1GabWF+pf8i0+Qu9RR3PD9Zog2rQSFwLSThg
ltUK/u8kQGAZf0451gIUzOfZ03SaehGBrz2ymNApHkcz9B6YmyI7SZ/IU3oS1f6st+1fdJ8bDocX
CeuJTrlJ/eJrXvyaI972aWSj9926k2j8bKAgHh/fSnFsWcJ1Y28W9PueCXd/yPGIT3S134oeShL7
2IF5NJD9Top453fouhWxkv4JVVF0sDkKF20C293zpwH6hKhSRNtkCpLkCsQEChqZDQ5taDXhSvyE
ZY+0MhfJeaor0fn7MWv0XzvoKHPtU0zBD5UxCnlq+rNAasHyN+BEEk7/dzl0lppWmoD/hwo+EhWw
MrRl30Hf7l3oZPrAVa6NLGqEcQHznx2X5nMKScAikkp0ofClI1qVGVsFOAPsyNkuMaAcMvW90hOp
Ll7hvpMa3uICa8BuwJvt9K3WwkySwvtvHQjZthMzCU7zGqdBh3BI1uaBV8st5glcJtqnZYG12sCG
LH8kgbG6IdtQcI7YfKWXUD0xW7cQzjQGP3ITccaVEL8/+JC0SA1+XNnDSmvo6xf0DB7E3XI3prwW
CauhU7gCDdSmKSyNqoDBgFWuIdYT/8b8rCYOzcqIsCIIu+MGFTYIYfiXmmtLzE2CEVHWGAwdyiBq
REvJHicDwctrE67cA/zKhgEYqbGBNzGXIcjdRdw667PXewGzKYLJv6C5HOEPLyBvfOWvulFTp3M0
sEz6pPfRDNdEAyUtxVNaZK8BHbyI1WPEiEbgV4nrZBTDeTG1wWUeVzbsK+H5AXWJYTJIsSArEDw6
SBABTXqHbzGbYcJ4b2Tq8gBzTHLgSdeYOb5l9bozAHqMNoT/yFIq5HSgdNbXN3JhvpFhtiSjixHl
rirh8aB+nBmWSUi6oKBQ8Gyzlp8pRbDSmcPYIxhUSoOQL9jB2qKU8VJVyFZ+vlV2rXUlvYBfsGA9
n/qNeqS5mX/ecJj/Xhd+Max2DBPdKrLnoxVtEYiq+8OdOXpMJ6siShj9uj6DqjsfCsvn9EArOCd5
qjA2sBlMyXQfjtJgxPY4C2/DRnPu1f1Opv6EU7M4I3x3zcsn6Q/KPZsRFtug89lKsogMvYhKVetF
CIHkNJd/vk+wPUYotehZ310T2Y/T2mel6NtKvCYYTeTcutSWXfuUN5J5/aBdKwTFyiYzWujq9QwD
Q4S44OJkW07iLgGUa4kysWgEAxPY/u0DiiBaqvYuieMcR2HHkmFmoJ6P3NPhbHvLhPk6LKX/nhZx
uQ0vwbATgeeKkv1WB3OsAZdJpRROBwOPebGIqYZAhi7NIjX1XCfQilg44QUcnAbwfEZVlo9m399v
p1eymK8GLCNtU5Uwx94+QpFWShBnCAtC77mh1jk7XEHMw89fm4DZQ6xCyqvI/k6gSCZnm42TQjwK
B1gpE/N7HphDf26GlgtWCO3HZpz5p4joTCF3cIaisEu0IhTmGfvF3MJiYcwt7Eotb0O+T9Oti2Mq
kQcnA4eQ9cdJTVBAejv0OHdF+tEzFzMHxGP3FaxN/74hRompF8lgjbZp5+9VCTUeswiLQibfp/VD
Pe7UdX8pzjhKbubfmOkWWpDvJDHefU/kDB+4OJ5Gsawehh98Bjo30IQPSF6XlIXt5SED6C9PlPDx
vyE8W/1GYCQtkYEA0oCOXHct7iimDm1BIfHrMjCDJ1XhkQu7rIoRwZnK2k/yKdzWdIdSeZKLxfl1
BnmgFolhzH+cxB3eAcEpie0v/uh3tFBfsx1xyOf1nQW1CP3llHqtxAezTjzhsZJJ4M6fbWFMqoK5
mNA0Ppi00DF58kqD6owLTDEJxyYKzOtU5nF2XcY0O5gpVuecH0l1A+wNhQxg6BnfxmVegA8ESk7y
2w7kw0NIamdqL4cGb9Ha14EwuyctiY5iRPvDNKulHLi/tunrpgVRtlzq11ipQxKSm7Gi7wVd9Xbp
oiVYbffUSYTgrKoj4QJj4D3uVL/sbcvIzWIxMz7vDssCKi1fnUEXnj81rnLVNBuIWT8IWVG3/nKV
OLABZNSyene1Sxpp81fSv7h5Xqm/h439LtHpSiAKhS1F/BiCyNbNOSycVZgd+M7ek6zi+BeePumD
PywLtBkeNvl5H0nKXC+eiotcJVRork3cP3USLDbsPzdKGM/9rVaoVVqmxDnhsaewFPUqtNH/4Lod
+kE0Slr+FwlSzM7TG5/9BhIRZ7g95SwXJwvfe15EheaA4ItpHScpMR0nIdo05OS+/95ZG+s4tP7u
4081ap9qXMLRWLttueplhUGOLKjH88mPoR48pCev/W2vJvIIWBl5TMOlKKQQ0//aB+abDkPar98/
L1qZsg27n1qZ305WZwfA9EZ1g8eEwnmYkcv5VEoKIweI4E1Tp9BNf8d8zjW3XDihTMA0Ns9uTeyh
XaDlqbpGPMS0cuoHS+WQW/gC8uT6CdFx5dy1ptRWT2lX0mmvzbWXD1jeGWbSrw2jIxVUUFx1HCYD
9ioDk1HSmj1tnKw65PC7dom4ce7Q88WsdZ32Yf/sTu/RTG1ZAfFk74N3GG32HRN8r0CGwQI2MA0q
g73fSglmEkQ+bNpCXMUUVsQfko48sBHA7f/f8yK3rqEbNn9zK7YOQ/lW4/zm+SIiJkQ+sYRevF0I
Dy7RQk4Z7gOIDPxaq/EvbSGs2Tpd4wPxEYugd+3uUyUkfzuoD1zmQ81BQ/C48iRONlVzy8zdnlW8
xKmUzlMrRi9i3Yrs+BHtLiGTtUk28OM2t8QX6ky4PG5vuKfBzFvFhON6t4Ka60Q7L5C/JyPy45+8
w99YOT5PDRPaRXPCYmDlEBhlR/gPzFt8Kty6iCi4L52bZOs4qXwJnBF/t8B9Klq5+Ixz6tn+/6IX
Oj2f+kEOzUjKSfdGwm4hF+HzS60cvGIgZ7fSsFSOuTa+DDhIQLoN0QRuXabfuGCvOnBolWdIybPR
YhtIGF0lb6NyY0XVao9bD3SV/vnEC/hzHEH3fT7+Ly8RFw5KE6Hr8K5z2D+/1XQ3xqNW0O6XdNmr
772s3RV1NJhMBsudJt+b7Bg2blU/PJBPmwj/tWN6c0Q2XUKr6sQd/Lse1hCVdDKAkA/pXkeOTxsV
dTzYX/hagfZGtUP5NyytgHKJjtl4HWMzWkwyTHHMMExHYACzI5Jkdax2Y5WbCBudGUcBVCpYBL2K
9SkNHwii9xiBkhIGVji4X6kRFrjTRu3nPUxMP7qaOEt8P3dLA4Ud1J1McB4fBxEdSDUjE2xJ3ia9
b4JRhZ6tUOJeq2CJixn89Y1sMR3S7T2Y3eGqx3lnITFH0FrNqP9/QFr//32BTgGFTJ8yvcm/tbtG
9x3889YchZeHNrUOWGqJgsj/UqQ8+X/BeC4MAAYgOQkRMJFASifwWqgrm0mF+UdjWDPdxwkRLXyu
8PmlumMEcZDHmTA6XXQnAIYC7xGQE7y5dtuPuy/jvpYeyFBg8BN82Vif7AtgvhjAlFFMYO99dEZb
FFkuKFOKk9yUqNRGT3ZIGDZPp2ieuElqsr0CLCxTyWKvKpTTnkdGU78ZpWIChbL3rQfjqS/FC0f0
XptSYGih6YzbZbVLC8WUwjjKpj1MdXOM86XJZ2rH906kULhOGntD+mv6/hVr+pbatrKzAJzTe/ld
6bGHNAIYm0INKj14CGsl79jdcj6zjwfjScUv0UXc/JcFDfzYYS2NVotrfJfrKdN78/4ZiIBdL1Hn
s5/IefsWEQcaV0Aq3A8V5ZSK8OHFA0pIt1l3Wal60gM4An44cS4Th7uT5l/+/zTJ6D1EvMIjmGaO
uIgTA+qfdixxKTTnNmE6cX1SgdEYTdT+es6DJIHZEiYcuv/A912O5ThEQYC4b0EBmZAjCbAkPLss
Y3yMW/A0hxde4LrHvVFwJlaqPKnY+Ppa3WoimuE75mvmF3/NfbXu0XyesYJpyMQtk7DGXwmTtiJX
tal7gBFRAGfxqblEypmVddy/RB/S511RR8VxoaQtb1/h4ffKXRmSwxquuInBn8cLPSw2Hls24FPR
8p0edHcX6nwGMQ7Tgeir2Krdo9LexRAY12ZvScupoC2WmbxSBlZjY53ZLPTnqBTUgwde22cNyqGT
NUxk4XLFxNgBU9sgh2ZG8dm5eNnfrS4Cqt+RsThBz/0ANH8wytH/qai2HfnMdhP3dM01zur8HYzH
1d6E/e7yN0TIhNcpvC7uA02n1ne9GDh4Y+TMnwzOaTPjQhzZ6PCManzh0dptPei2+lm4YlBCUA1w
JDFRaMaibnDMoQcB8X51ei9hPa6f8t4VXAXBPK1Ew53bQGYuG0UxMw8lH5WThbs+az+hunfW+Cv5
KrUvzd98iygSs4mmbrA/P9o55LCnRWJb1ZdqM/L5YAP6dT9DDHnqAAvnWnHeeWHoqTZ/tD995CTb
+LYVdqBtrUKRvzCUmjA79ZK+S8zslmuLqvcFV1ZFjh5ssMFUSMYok9/K5/bYscCQHp8DO8CotvYC
NT3W4JIYDJTQcOm3gOURC74mEdJQeb5NzLKY4yL9GnR7Qx4HlilgQ5Jxjmp4ZC2EA9CQmMeaqx2O
VCxdP3xY+TTDDhudeApVyT/WP99i1ogzFuAjqP8v43HaG1X+QcsM8wejIaubb3dz6MxfQ5cCW6yV
CorTYUioIAnJnl9fqSeQByYo/lVMYTWTJKelMgNstJuYXHUoqOQeDxjw1ZE3BhC3qO7dHCuKiNJ/
kaO2EWyHWnQK3AS6y3tztea9uiXDQn3ZR+/yErWtd3P8yv03OkKaDkRJ4OD7w8nfMM3dDR3VGqWG
N6KMH7pNWOfeUqqW9NN0I6S65iBZeQkOr8Ebno/MjHEE2lDuZJLMpXMIRPBxJcMJ3XAciIYVClba
FaMksBc8mEJTIolSrFvX18zwLpPsRx1jftJLh0bW4hh3E2SSgcPylXWJWqnPS6LLUsu4ZmuxwyQh
6+LAFluiHH7ygIbcVjTyKBlsj60XEUzO9Xz4TnwuIdpJyFM+g444BvYyExcmeITNOppQWQ7IgGPw
Q/q7Tr8Wy892pOiTJStgIRDpeWZ1rDCOZhIouUFoZ6zbZ9uk2l5icb61V7RHEN1LLrSbAmFNfV8I
nrFwE7oXENFThaJr7H3QEWPltA0EGlu5xVG0Ln60ewAPyAlCaihGCiAdygRTv05rbfLPsU7GHR2t
pOQHUzlrar8Bb4+trmWokcD8/qLICNoRoaTMMFXMzsqcEgjXHOH/7jPDI7foOQslA4eSW9V3IFPr
z8t+Pzi6o9i3OIhQ3drgOKMjRiB5ibuSn4UnXWv0TJlvdovYZazd93RnMGQtBHpfXo4wxt5UmkLI
MWv+k1cF13h1/H45r1Nc6LLp1kGDoSGZ15/CFISwROeC+QOh69xff4rRyRZz4WvjpCbqep4HiFo5
m8uf002r1mFHlTkus/ZWoDmZX7hMATa/yA2WIiAus44Oh0+NC0wr5jBR0ST8dhA/7k/B3dOVWpVt
upawnUb+w9xR2zYWk3HZBKSCKmH/X1MgLrQM1jrB+nHjYy+vyyqqFZm3N2zoD5k83GPzyIwPBC7m
7qVrp4VHmlmCKpRDIWARJzSKzbfhw50R+dspm3NiftqYJ+G7MDs5S+JuT6NJml7RKbMF1Dt4Okvi
oFTWK8ePSaK1HZkgTW6walb90tOJsfBz7RECNrd2xHTHKZBenIqRCCe//F54fIglBMh5ZpV9cX4v
tY+GExFrSxiCBMYOsV0mJM89KQSegZujQgCcoVNsEa68TITeze29CY4UzKvo84P6ZeoZvq/OtX3o
CxBoQYQmFsXrUOd87szGA8DgaHZXHfwXx3MHPcPaTUVL2CVFp4oFMTnmli74OSucboD/PAZlQqSg
LxeXowk2kQlDXyZUW9o8VsLWMESx0LjSuz//AydqcpW9uN/UMFQeaa6qWdCxOWsSbuDfbIAyJkcE
Vbnx0CWdxar3NaVQJnLO0yB3K2192S5xK6rqTqzigmtaH898sDdYDspblQ1mQDLa4TgbKW8BGoY1
1LmWnNU3KQ/43OYDZBUOSn61PTZ5QBJje7RY7ocBO4vP0aW5xgfaZU9mwTUSBoWnpwLbGvWxTQzv
ykQVpYM7xxJp2Ry5lYIYeZniE/U5eXSCkBIzpZ/QArXfsPmJDkRTk0F7+Pr5zJrV7rSRWeJwYM+t
eo1gfJwEodiRg8Jkx149cK1LSTUcxzXjvrvepq9s9AvoQFsd9zVaF2GeBTNqC62spLHmWneeQMoJ
a3Kk+WO8n3USVwtP0tuGTCOVGjS/BC+VneeSKY+XZGPd9RAgPIH5jqLYbrQJljUWJOtDlNk9Wtog
AevavJ/XDDwJGOrIrKo8LyCnma3092lTWSpmM5wgFWrOv0PedidPE+zssS3O2duKGDlwb+mfu4pQ
iICl20JQBu9KmQ1ftuynjfWNCnmpDooMFUxkmQGO/TLIYy1QpNCaGVb3Y95v1YyzpsKg6r2ggNxJ
NYGh1Rv+tFxaQgyxsyudoQX7Y6pTA6TpRTemr8EAK0ULxfnmEitVz2JEaWNqG2AWm5CNj4J2h8T8
ueqw8Xh6WsnBk8mg3qs/f5EN9WHH9y2kL9OtqO/fH83OLyKpv8qWgMUsGh5gB4CvlwqzxXqjdSni
S/RTyMubHe6JDPOe2sTQUD/4r93RFHmBnfIsFuJiJX3ZXXZyRfu446YUkwHUQvDL3j9YbMRoGmCp
tx89nxUgECblFlgvKT0X9tpSAqtQXRu3m+1/r8U0yo2P8Fw5nv2on1+HuED9fxYYKaUcjrhrrRFn
lLDt29w7P6TK07JhngebBJgMLIx/7/g5kdrdcvD6lY1T2H43aLZdv68UiREUlKW3HwCRP4z7f4uX
xQHiCah2tJL+y3Dp1tDMtHO5aTI1o4I39lymQjXvpIf7uvuEGg0Onu9WJd+fSTFiStKZKxT0aUOw
9rHt1h4I789XO3ZLIXrMKsXBFrwKSYNQW8dvZ+NalXt4hLCWwIgutFrVi1nPqxeiU49TpTuKpkiQ
+Nr7cP/zm2os290yODeFe8eJAMCKddUyk2HchL8dFiewQHygXE6ujXfBrKCRSRJy/ZezeLX/ZB6U
HARuYwM897KCPjZ3SVT+Qvb9pP1fBCaGLhqu66Q8DcfI7rg6GfKi++BcY9aflB7cCRqmdMZiX3u2
k8AkVn8IFb02xhEjM4/VVJpGunp+0fBCoE0FV3RgowehWg6FuZfEhlwi4I0axcqXvt44a8eYuvw5
GQTRTqRltwYezUv5q79Z8MW9qwpPqD96xCfHRtTX2C7biTSREH76+6ZD6g02YLbWZE5wmgFQ5Tnp
Svjca8XavtbFdm+advLQfzmifCSoRTOBN2xwbycN16fn7B6c/P/YW67bypsMOh2jV5yPHqHCnZKi
5NQqrjqylUczh31frM8K6IJir4XqlJiIhReSOzMecWwOLhXqnUmGFLkj7UxMgmlu3wKDh+da9r1N
CTUlLlT29aXSfeKdX9ADYdEykIDNFzEFm98bv6uaKPj/e67cKZ5XjvD372RwlBqOk0fRRkcWt4Yu
z9+iYoDSra5WTdK6+j1yDbPymd6w1YAF0fF2Mrw5aDJBWWnk1eHVAhxdgMtxmFiq0IN6CtGz7znB
0iaBuRbXho57IXINPymxqISTskJZFDo+EqoB8L4/hRtk7XHumLDgR6cWGf4nH8QBPRVWzaoESqvY
49tAAE3Bc83sVTjTar9zYv01Y1WamYO2A1NXsVtgFDZm/nMJSfjmvqr5gBBJIF6Y+pCAzsz1XIGF
7GqWCQoiKfiyxNXtcRIVJVilr3iXX20wmR5KQR3Z7o7LO2mbeVtmLTgRs5CggOEmnhpFeh+ft/LW
mlXOUwBKz07sbfvD3bgb021ynb/GXHJQVRoncySWSy85/CW7A6Vzz7llO/wYuwVniEjIdoZ8+dzd
59hh+M6+JU+sVVaz+YWE8owH8Wf5skUd125OieMK3VRq1Lc+x3FwgXnpNvlCZtmqxG9iO9Dz+bv8
CKPgVY1wUKolsnbRPcdXRmYBX5HOazXyA+HsFY/F/0zQKEY45ZU65WNJoyR0Gq/1hOhRZE5yw/jk
C0lg6aupki5iuI6hTBmfY1YM70XAjvVjv2qhVfa1kgIBgWgH2GUA2pYcGRFnEl6NOgewYEsf+UuA
nVrbLGp+mFPEGpNUkyKF2VVnawMSORpYKnauYSBtJF7OXv4bH/eL8w+5WQT7Lw1v6uvFOcCtaXyl
1cBBZA+N2GyQgSIexioTo+rosXP8bZJG1XYtbMwa2nnpwLXT88uX/XQ0yGHf2XCskCwSw2uiOpys
JYP97oJwtU5V79yz9Q+E59ynzCOf7TVebcnR2fyDQqIurw/iz+b5YYFgrCriA7gwh1TxJ7COAWbR
q6hoyzgVzIRjvWJqS69UiMHWHpLKmaEUPGd0XFfWkYQYSM2FUEyzfTWlA5j186doOinxgimWw93t
6+WTsDr3ugxmxodQpkcEWXgM+d6B12WGSsXwn76EaFbEk1Zkj62+8y57yUEnSR1JQtcUtQjDQjeQ
hWkS7IghjvViD8amRXIR2uBbVKtygD4JmFiWmNRG7ZrMJHFN/AvMOpDYICDOjEZcexo2UNTAqB5s
uN69Zf/yedvuhkV34BFUR8OTUeZNQU04PV0l8q5y7e8Xd7Am2YnjvwP2NI0/3hGah/yaSzDhqFUO
LX2ZX12HnEdhCiB/R8HLwrR+2gHGhEnTYbu7rXLB22Bi6q1OyDlFuiIMnXSqchSuGxdtuaDSecVT
torNUN79ZnKojncRpKL86Ylth/9vxMhfIOVVJp0Fx/s94yptzTIXHpac8RVT0F9yVQlyUh5iWaTc
HHs8bk6nh37a433yYjLtBVat6c7Z7cN3BOtApSLQLrk7E/wc/c9Ws90lwAovENbwmDk1MCG4jzQT
IExayNJtlX0geKMu7qziiUnv8hlkClmXbac+XGfDkVUrmphn3WwGfJQ0gnhXUQAz882idB/h23fs
FL/horlL9xjQJ1zJi5+/8LFb0dJz6/AoX9gmjIWaVRN1VIpP70vMuhoL9KYu+K92xS9bFJAMxP5a
RdyOxARLHXr+VWjpUJv1Ri3uBRrIRLXJRwKp/mbLA/kgKA86PFysgXjYMZCUtE9YZSCgo4k3NY2H
Eq9jm6b7PNa99x3Ei5ataqM6x0Xhigdxo2McKEeDGK8uLw/r22xr8EE+fSf8sNE6B9L6zhuME7ZD
xFmT1Bz6gYcWt3C2KAxWBoelhUEa76WBex4mCsKPeo9T7gaANfd2e2yJjR3bJZ6chbduMYn60Br8
+1DKeU/EriyzEg6GhrHPpeKi5JggnJUlNhtnCwAVDBcxNw5IcZYhZdZUHf1KKIQ+f4/5zFqmm40v
FyNSv5GNL1x5uuBiHvzDRROyEJUfd5VPZCi0k5H4OAK4jz9HYDVmkvOE6EkZufwOG2DlcR03jjlm
CXCQ05rq2eRoLb9CoIfZDTgxIQAIcO5H43pxB5JqD4Z7PMxhZ7imtPvzu3qEbjH8DRhwQxkWB+sF
e2dQwOjSrA0396yM5FZlkzUayxHHc20dgU3VqiCNUfkZ18rbHdX6MPOeXJZmYwn8SP6sZFUGjnyB
N2Ieesl2Nv0mo/8TmWuhyYHwRrsUlH2fRGomdJYUIciJWoaV6nk+9MMTyXHwG+knWcSVEiNDjVRc
VN32ITNFLnPUXnBYD2Kr22lw4nTAnRgjM/ME+daKZSqDzm20bfMyVi/kOuBvw8C7NKfZqdsvNEnD
SX3efjwWn93oIqAO5nU9sBRtRJL9cQcYSMZOTzLGE+cIGS/lhEDUqmW/H5gya+01p8XJjDsk3zuU
JPlcy2nudlaVvASvSx/jT8Cv0CpVMXiZkzNPMJRuZFQdFRV4+E/bY9s0XmzY5Z7IktypIwKcePCA
tY0+r9QOvax/xU+Y6mD76nqqeeQOTq5os8cQ0Mj3rwSJRbVeyOkpIJlgN1KlXNhjlLWGwuvkWnyr
zOPree2zUkipsj2IB/wEQ3KTEz0yBk852Wcrt+wnvFIc9LLlToa2FlIV0ZJ//GHvi+746XRSfrJW
M7Df5J0JgUOGnOTG+N21+Z/GROD88j5A35rAv4L0Me/f67XqGz6y9KQgwOX2y5wVNi3WQEMncx5H
ap8ywWZV4fLmo1LoIX5KYSYssuRpPVpJ56RxFSux8J1I4C9QYELF715id82eU2juTwboXlNfdU7K
iWx+VBfpUfOs3MUTL9ASoNbnR9tGlaEBXQ6UdJztf4dS+qAm5guSYOQ8jY5NOu7Jo7eiY7gNHqeY
vHb8YUWOoAsi5INJlpZr6fKFHqUitfzJOR8d9jGJ/lEqw1y5k6AppBbJinNfenipdeSmZuL0My8x
o1tppgW8FXZBdqE+NmpeOOqdiBpZTA2R1GdnIHH5PYNT7n9nYxpFO+jiAnHanvqYhfmMtoL6wKc3
FXCiphSy1nn1f+Fw+ggrTG9teHIK6wzIpAHgtctPKkpPWf7apj1/eBw6l7vZH4oegh80dzk5BE6P
nfQGbgG4zfqOnFT1Q2ZkmDBrvSaTPACm1oIZNTS2qI+iKODW/Txd+8Vqnj4c4r7lnRVRNAUBzlMJ
WQVQ3dM0mkZMOn0xcpqdCOswomjoKrwn7TsKYgH8sS5BEIsoGnLHL6w+4ri9LTrYFZ2nqt6rbFGv
7blogMzC4LFoOzzon5oSSHQZ8UQ9rndzQu724e/9o33x4fu5y130UDOliU01CBZQ9iJbftJpGKnw
7SYvQ9sWyCsi59rVRttuQ6hTWhSSnvHgA4/HSYeXo1+xSuasqcV1jsRhgbpB0G5aVfBghZZlpvUS
Hj7/JjGb/Si7PGtGImuF7j8+LgN6Z60hMmGmnFgMjPC5QDYLtLvfy+5xLhtMkMZ7Bpe43pCvLPnr
vva48FF1uLQl+afCPq18rXstC1KyIwU+2+652hecSSkjNwSI9ZQxkHIMl6XJSOxp8HSn0Irjp9HJ
MDKIflP12ZppBEtpaaKhqWy72xyYMOlQiSUeo1P0z6+LlWnTTjEpxEz5ibIlV2Mr/PRbf9/DKY1P
AyO5p3PYTIJaQj72m/aZJmfQbb9Xq39wBRsJjgQTu+gwwjZgC7VLzjJWxhyDeatMz9XnnNghCxHe
XPzzE3NMl/vrkEOfM9nwNhxpPaj9rCkegtrB8PWC6rLhZDKYucATzHAYodUqnZZrunwojii6JO04
Qx2yGeva6aYxqstsXPRdkmkJBGISvElAabfkvvlU57yzcHnBFYGhJIu+xBzuT+C2YL2ZSj8HkCzy
OYJz82r819+PExUKVc8C9eSUYRIO8zpXueaRTKIXfLQ2X+Z3rd+7Vn36aeLVNBeKvzp8v8Lz5eB1
/FEg5yhShJOwpOAZ5d5iE/nMkh7rQzUuW+zG4rVua6snLAXrtK0AD1fmpac7YUUFQmlSFgkyFMRv
z+zpZqnb4dhwxnAOECUb4QDPpdvWANS9hRp5G/KyXcQoZsiATD+k+U5ShBmH1srr6uG44NKrpN24
bWJ/yvEsUUWYI3bM65NhVJ4sfSgesIFRrol+R3oXxS28EaE6HFHoqfaOfoFPvYaxKitalVZsUHpX
iUjEwE485T1HgJRqErq/M+o7VG4c9MrvpTZrjwZF4nIMXv2sPrkzEeDiD0/G1/K56E7ofLn5WpoT
i8ZG/HNeVcbyzlyJY7BWpOnA10+PnvbxNUay7JmlaBGGrbPuEyhm9mvhYXjpfPbc1AxDv+nirZpE
ik3KsXQb+cezylGslqasViVyqbyHlsBZyi6ucUrp8oJ7hLqNpvsOcVLZwKecuIK5npOIGOaCMlcC
fFYWb7wDQZpazH4OF+75btLu/PAJuOWR/NrXYByJJ6X1iIc2NX6PFRmEGmVMCUTDMFgIy5Rysq3O
i3X+rPZd+1ihzJeCXSRTtl6lDnybRku0qA83Y8z2qN3b4ii3nD0MNtUKIRYNvFgTzKa3jLTYHTpK
pY6EQUTSAESXz8pbLB3tbDPwbSuvBcJ9TLp7czR2zgpfcO1IrDyFGaIGAYocl/X4SbvrJgRGNR0A
Klsi26hK23jF4MGPSgvCIYqJP8+HhwLUINhsaS6p4ifSERIjNOGZq8gymjaSbOdbI1bOzjzlaDMD
J5LgabVJEBUvxqtWZmqSCB3n5sUeYvX6WozpVLym/JjTk8aWkz1O+lo8R6JTTlV+OMXKcQLU4Zik
0juh3UkwOgxIly6yCMyzePSsZ/SFij6iZMDajBe6zxkmKm9TgBx6BpJ2cFH8KDBD0DEJ0g54mY3y
Iyk4v2DpANikO6OOWY0WAi5hTJK9kdAruIJdEGw3t3T60rx+B3NR7d19NkYQe5Ko3vAWzmsaN0M9
M8WTIEok4fnzNs4OzXNA6O9jZFW7yxOd1GpmLnYYE+cUVUi/A59LYcLxbU5YyokOTeH6m+1E5Tc8
qE//xLgSN5ziMZel2/N3ChPr8L2E8OGwICSAZRnd3Y8mGwVObMRAH9v5r8hKYYp/utkQc7tiJACw
O9OZmw6/NBxZb+C9sPtvjxukZc5x57A7MGwfEX93LDiZnoJGkUgWCRTvBOlDHjieh+fDlVtKZvYh
I5y3tVrHTncbxFniwFA1vskDVn3nnWnf9Oyen1FKaCeI2+EP2O3+a9rkYW82vu/FzK9aBeCzaFS9
ZYb+iX0fItjzA8wEXGL2n/rNGC3IimLf4goPe9tJ5Ml3+pX/iNSivnBfd2I69/yDSCzSiLj6mPp/
DoCDiNRZ6gmIN8xirEVSLvNJYPAUS7MsLKIj+7q+FuWaSnZHbe2nVec5qlw6gkEJd2JgyhQk9CKm
GNiZK7nOwDpyLCGabtLl5+8bNCYaAlFVFMLU0tuHTrKPVfYKBOTpFdf7lgxOhpwjj2hkbccSLxUj
pInBU9I7owyfLT+35iURDUXhFXaA6pJDfxZwcsAQAxBUVIdyj8kNBW7pqyavEpHbccB8ym0DAggg
YAjc5D6lQELIAvVu0X3+heMyYkZ6TyEErvS8PBR/JSQ6/usobZ2ygwTUT5/fRbwRBTGgrNd7oPD2
vE0q1QMlF++bVW14izVIYBs+TeHaJ3Ll5HftzDFYIE07etk/LbhjpLLPoBMp2CYtv0HGiURWluMD
ggKKmVuqnVwH/tHGQXRFKlrTUprqNkYSaTbAvNO8/zeBCvhl1vPmzvR8WwKp2u0YkTWtezAMBz/x
a/ZC75VdJFaTA2aDOk0qZkkRG6H6rSdwcAxY/Zy6lPUni/9RQxnekBn6gDT1lc9u2hZMF7c4/z3V
kxRpORVFKvYEP/VWZF1Ippws+L7pBMun++nt7dICGpIgpd1SgVq8QGo+CRxjYF4q/NogLCX/Yap5
u+5UE2UJnqc64gpAYJA4Uo3alao2Juso+td+pfrgd2TU046UmOwN6/vR6WAtvYh6cqLQXNJDFeGn
oCpV5NYpwBK44eeFfQlcUmnaeQjMpkRbUSNNINsdFHUSkti3ZZob3hZjn4yuwpqMSZcY0yAfAMoZ
4twYNdEsrtfR8C4V6+FnT5MNbbbmXcPX6Zjn4QzqacA2lr4Et3TAlruXr90aFVTjXNjqCovGshSs
un4qL8TRKrfd36sTFCvXV0b5lTH7UF2h7yJP+AnmJidqu4OxlAsI4C9QuYXyBi/kPHe57ZgfQ5QN
pM61ru3TLbUZhWjKLc/JBQiP6k1RYSrKteGKymlRcnfxwYkpl0v3D2udguxZFLkIrjlQ3K32Xc2O
q3tFm1gE89z3kx1rAza+lkMgxcpQe6/z60JuclXuDFql/5pvV/OpYApTPu+5lPX7b9YceORXavE0
9fHvftNzFW5CvpNpuAnSVRnad3H90g5KI5cHQF1mlwVf1inPBifcRCXu9s/emwhZy/34p70NQ9N/
hkhAypUUSmt+6b4JMwyr0muPsGBoEIMm95virSx+/lkZU+n6Y7ZM27cPsoF/XrvrHZ46VJEOdRNv
Gx8Yza0Y7p+Va+RFxf/DASrJ2HQTPKe49+Z9mainzzk7CS20vWCoN+VSpnh38THBPW4d0jtQ+GJg
L/KNqkqnswbKxZEvCJQvLpSh6SEtz1Lq/gkayxmAmhyulVc6k8ehz5D8/+rMmieGAcLVOm7ysb5U
Y5WkAGQmvrBOPQQ7bDb7zpn+Nrn3l/dJh4kwj63Oj18J3akQE9ae1iHY7mQN2UclXIUmUuqWEOY3
U/FTalrESDVaOvgyoNOIOHFnHbC1dR2EpyTzCrmwWRnPaTqrlA4tUKPonqhgBC6D2tyr5eVifVY4
Eq5aofnknOx0g3dQ8bccGnV25N1U7StzsaPrgQtEKDiJqSoZbZJnf720XqX5SBYoxXSRynmOWwlv
Q0UUeNSx77Exfs3TMxg0nfV+V8vDe/3YalPyNURVU4abCOVaeGhPFaeRzGm7+dKbQHTRTZwyMYFX
6CxNrUlExhH7YS4AtI7i03G+wBkXRTij4At+ufkKQuhm75OqygeKo95OplYURPpVK/T2jXt2srcu
Ub9+9mLrZMJeBUfnSpBRk6RCnaN4X7nUY7ggJ25gK5Dtupk0Srqka+xYQb0OzyEfwiPggA8z2xk/
G9rUK5hyBOYr72aei3XMmaatB69XrD8cLQz7aa7Q0uAuOBw5FzJQliy8mPCXNk7PpFqPZ1e1YAkq
fITQX+Z6EHPZF2HAZKwXP4/OimE4Ba2IVQEVLglhLvA5Rn0WGMCQy8E5VaLD2y7Dk5lP37qcf03E
e1evVVw/3YRrJbDYc1vGSb35KfmaA/drStl9cVJWx5vCBhRhqukKCkJELfnHOqY0WXKX6ABcovl0
AwamxSXRy3g6FM96o9fczfEPL5EmkP78iWNqNxkP62z3PLGZx/DRWsz5y35Jjzomes+OSoIBIb6N
PjkfSvVudfeHmvb2XDcXqYrMA7uh0R6Q6vHbH1WsVlCFBi+uIJNpCTqziNRI79yGvCSkWSypJXD5
ya6dEpjZqwNo2G/jaibjzxA1N2r1WkzBE8o+IMGuRfCAKEginDyyvg7r/0yusvpvjw9fT65NMF8P
C6NR7vMMehtcB525chNPk/Frv+A7CQLgBUaOjSqRQLRYDeFpquvmgM8Tn0Z31QjWCI2MnIREUff+
dmiRWXrYPRfbnD8UmHJT0I8K54SFO9lJJQXzcfFKJm5TM/kz4XQyJvMXqXIDRQ4HYZP63sOvD9rk
GR88X2xV2CgTupP4IS7doEWWjv3qGumE2NkfmvhL0nkU/bkZ6j780OxUtVXEdnBgjLl/f4ON8Noi
z3PDtkpw1Mwrqux3sydg/u3vh6MeGREGM/HZ6vWYSMAgoGWz64mZl7Qtdpe26saHUoOr25NZHFR1
XE90N3Jfq36L2sJ4KbjtHotdEMAfRodbEJSr55aYeSBfA0eLLGfXLrDbz7jPx1SGAyy7XNPjFUag
buBLax53mOKUdvBXn6MjCQbKst1AE7Vs/CFD6ap4Ejx9p9CXdtN/yDBBj5J4fdJwUuTxU+sf7n73
QwTpJdkW7u59eFK1ZD2ptWTWy2KDHGvWnSfNc0dGLQE9/jr2f98TVJOYTxuDf/4DyMysgFooDfgK
p+yC2mvUMFkdtNPBmiWTdU4axnbNYon3XB+MND/yOz+MXmQemhtUfuhrUnofMpwN0Fw2J7FjbB9a
ANtrZZ7QISV3ADmBHRwGiQ05JLjWf5fELJ+v5tLr5VoPdFLc7opXLTMHfBpcjvgc7sgDpYgTApyN
Ej0Dv28wplxuLgtWdpKSa9yOeHX4v5AZO6qr1sWVXCB7qcFm4TmL/Jtmls9E8Z6gTyjq6LW4OfZP
jTueSzket6CRwlf3MMVQWNO0q51LRhayYGBw4+inQMa6U5EKD3CKfikyjtNwJOMKtENWN/WBmERo
Q5wrlDZVsFvNFDTyQw7+2zEQ1lQiuF6ZHMFGg3C1PTMcD49E0L1yemfHzAI81+XoUSN2lbSViznP
S5srxnt66pLhbsVwiS1Hi414zNSTEvcDD+z4Ef0PBMbNsQwCjQTbCf2jY693ChUDJiEuW2bGQQJW
Y/5gsgRCZv9Fq5nZ55RPt/+A8aN4dWBoLHdOVVqxjAyjnEeyexc8yHZtP0BddEdPKBfdlTcWBvFF
5mvwrzPBsxtOglpa229xv7CDCInNgzP6TrjhyGmGpb3bgteeHymcQh69K8InBHD7nHudkblA9huX
r6RA2uJ0WFum9kCgQAPFyC/tDgd/BiR6oKWUNVLZ5zsEdu7qOVZEpjS38rLSdXFUp1Vsn15NBeTj
2Xeittnxxf5fDu1X52L+EgMi0WrX1CYBazPY9fJALaegYK6UP+okoEGxrnfcB2JFE4zeL55MO5lE
fT4BmdoemjXFcAI7RQxMuqv9aAMmx7V8E7Uxyf5CH2PoYz+7zuRNPCMK/x0OS5TfGE6iae1hxCtg
WCIMS49ZlFSnVTW2EAQc4uchkmGUVmTeaHp4iT42WKQgP5yO22CeG7ETfAXZdwXcqWCWF9DJMIVb
AlA0LP4EZtGT+9IjZ1L2xZXW+iBMxaxQJjxfGwxa4PHJouS/Uf3P4HfUmS/LsWMO4ZiU6wgufHKG
Es+1np8esvElHcEkBiQf8PHzczEfMi/f6VTJQHlLqNb9TeiHMUiPx1vQ4hy5tjkiws0S9zBDH6xG
20OWH9EOtgzJGEpN9V/3LT+UA8TuzH977/p9G2VM8rb2tNt6b2/yycirfaJIQJSV4ZZjb7eSKy64
OFxyhYo7HmgFHM+blIqSdVJRnNNEOCFTfagTWzA6HpeXT9woegPsVGVsIUOnGbqv2NGJZdIqDrRZ
fMD/vEVXjme3umU7ws3QGbSLKqK/dci+xwXbyyDdP7sxbPEhgmtS3JMG+SvH7CiAezW8WBQ1oUT0
cvKK4iwOaYKOQcXFARLz/OXd1nCXeoPf7MhsmOD/hK+TkIzY5wyDrOA/VvLyBiM7fUFIUgEN43si
V4EQnGZsGCJTLtv2aNruyEj/Yw++T/M5kGYr6ehKBnTt5wIQmoGmhgfi3e+QxgWukfFuMMJM9pQY
IPxh4GS6dHgi4mngrtNmN5rUwG20pSBbQZkowjtsxwqKqpqu1NH3vO2T3uZiZBjfhcUZiP+VidFT
/AmmMwCdxTr0m/y+o7rLUcDbbH7Y9XRVXYVA9hT02pbQKQaKWSD2puv0YUywWrzgXo8cSIcLgzpa
bFGPpwEAvC+zTW7QGkAhoB37Qnnj3RRPKZSH91RdtL6D3fhR3cNhs+/DWwbw8Zz+EbydcDjvr7L/
aSnflBmDU+dtMu7yxfHUF5iZ760eTlyllPHiQmdhIg4Xdnp60Y+yDwE/iKgkNoiycjGzLkX7VWuy
D+dGlhtqLtuE/oBgsVBUetQUWZsq63Lq0rVGvrcqt2xiCsda7kFtS76h7HCcJwJywsfuQzVgVxy1
AZxqEun125p1b6ed3UIb6Bu82LAdZBkTQ5nTqmphCWoB+KxBqbnbJ7ihnCu42HD6ZS0jJL7IVuYV
tDjB9LtSS2hVD9+4+EYD1g8zo+EmWh4oZgRIT8MQyleDJLvEtQ2QbRM1CZx53Bzkf/W5BswbntTL
1rC9WIrkqevZCE6y+oMdyO5IfLU5YZVzDT56JOlK0PhUqTw1oDas/68ga2B2PoJVCCzLDFTso/o7
505C2MOCmODQLJY5dh7gL3ESknKl5PcL5TQ+kFtStApxXZtGlbHVTPrpf/JpPQ83Za6Fbh/FliKK
bie6Sa+roM9vBRfgjWG8mH9IWJSd6eOgBocHMzF7B3DjtdTyf0pFuNKItUN4obm6Zwa3+eOhL7oc
T++BLjHkF61ingW5xC55lZ+fEILwhJdYx0tfR2cHgpznZqvJO2EZTmTvLdBmnFrbLt70OOutj3TA
3bpdoBnORkjN+4WTxLOaOn1UYdx2wT44o6RO6qLfUJf3eqmLj8DXDjU3Kj0XlV1VUdhZ5U1zf07B
MbACh74yH3N89oj7exl1aGAqH+7QNr+Upj8ymM5DceYMpP9U6i5GoBGmrOzjYxfYJQuSbadduM67
xCWHDgqkOMHntlgOlnOjP4lomYmEtAXdBBrndaNZhAbPiFoTsPx1orrrum4Ifp1oKmS1U04dIGvD
UcL5b86/dIrxL2sObQyymrVjlDrQXoFRtC3Y5tduludXWvEGZku0ykhW8vdorfyBA1W9i0S2wqPC
tQu/6jtfX5334merj2QkyyZISvO/a1+othpExhqcmNfrDN3CP2kF+XCA4PGoc65X+N94f/XZF1jE
/mEdw7BKwkVxLUpuxUb2y8WMT/RbN0CcNlfLGUu/fQDGiApAM0pDmWVWChHY6NVbxDadUHMMR8Lm
//wN0IJyS7KdgV9SHXA4vQ2A/VrQcztDDXhJwNTADaYGf+2YJJ6/J3UckHJe8+c7kZtQO8IfMsaf
Gy2KVql8xFlvq4CGkUW8hYKJtic0uYCcMyJVYyZxH0nm5ewdoNW8Z7gIwvHTDEAPJQRmGTrgOW3u
87TrRNa+OlD1gVN315ivObcI49q2VOwp2nQJfcuhrrmNpd0nUvHFpBlJeqzajiGuN3sVfe95Zz/8
HkOpcm/uiuGAzncQAgeXwfZW5YZxo7ecn8U87HwatRR/1403Zkpa8X3kmGVYNiJgr+dAWFOEzjkx
2G13OOdwSvoi9i0INYH1Ec/KFtSBFvqOZyx2uiobui915iz3jsOIAVXkvu3FFmsLAelo2xCUJ2j7
wKAO1oEaie9LQUG5AcbEWnsY/NxHOyklyXyeDMyUEqO7dAvfhUDEoHnAYn7P7StjDph06GyqKd1O
RGhzjCqepMEJfeKnExQweTi9woA05tblbb+KRnUx3HYnfIYxIC0uQ1w25PezJvsvYRDrlW9M1HOU
mTILZaJIVP0/uvyEZM1Y7DxeiYYK02OIZLgGNW+7MRbx2xRAsWQ4hnV9THjIIoU9o+nezkY4t9RS
h1ny4Arq1Nj6HlHYrDahwS31vyuowE6U3DqNknRL3KHsxpe0zxqcEbAwIyXR/nhCyWk2t9TAtcpe
wE0Dk2XddLZUEqCNS9V/w6aJFgsWxvrYwaaVfhln+y5ZOxS/mAVOsv42pYQY+6snWJLiWc1zjVDB
nYM25eoK3tlsLI2gb8t1htGHgxm7fd+G5DWNP7cBKGdLMaNFXdELLG86ln3DEnmhlHa1rtp1t78l
Xkc7jmsnJiiUDCrSTOrYicWfnQzTB5nPn3tW3XAwnHVU0rM2N38XGeYmDDxUynKsKEXf1NPjczr0
kVkNfpO4apXIhvVAUwki97VSxcf7YSvsuHmX20nKdlG2Pwm4Hh2u/vXNycR3pSvCl/KsBS2YPmep
E3pF/1qpJ29Jdb2EPw/dCRA4k8qbQ/ZuqRwDqcOPjjm3mzZhH4YxMcDVw3KJ6+maz1U2yNDpXzhY
dplawUF4Xi5zF7LmK9Q9jajxvqu92Eta9tnz3zzc1ZrCu3PmuLpwitmODGjjSwEcv7Xq7YJlcTk1
zMVaYbrOsKs+gtnIigQ6wjbpie16DE4TDsvgpsz6VkU3GFYIAurzvjzSFT5syGIAVkCMMsdncqUy
y7rVvJ1Z90XnMapMbdPTCZvIAZIS3Ii7UZ4q90JycBsRUlI8I5Asw2PbtvjmpjlPbm711S8hnun1
XXvPMcOMRMG67hpaxbcKoCl1DrEu+zVR0+YIDT7FaxZnYWYIDXR34t7PxgFmeq/dBxuQvJKS8cwX
YWVl/AowrSiIhIRx203ZFokmsxt+mriAcJxMqny+HT3VHwUx9GZOC6lEkBI1jhVupyz4Xj5OMYjK
nuTAGSL1nmyaZ4VMUtFra154VNn8O42deUL90rGnSRe2Iccr79e6n70pxkNkbJId7x4uH4HQYmHE
Id+19klvNM7ZS63aGWvxj+rh+sFdRLxkdvRlp4TfC3/vqjDnp97lBQL5rufDoK8CV1L8vWDXyT5E
u0aQ5yLOERoUck+zzZdrZCcKUUXGmvqQCoqQs6um6wydMXT/GBkbJxafHcsydikJshNSVAIsHHnK
BkXhMO5ccXFMbE1OhNb5XVgeLGAHwwy1aTJkWXJnYW56yjz8zQGAtVCVzK2Y3wm7iNJ0LeYFv1qg
X4G3uyWoS4PWHO/GdbOCh232+toe0ZhbqEgv3/CZRoA0mpCH4a9Wxh++afmGuxfj40AkPE/zpEVJ
Lla6Mgpcyps4yaQlAX5JbwghiGziq61llyg1AwS1zrXzMi/iMBu2rKjaUc4giobECVwwwMKzdrVP
WkPpwBcpLInNwrFP+KIijcCO5KhBFXh14oO1X0B99yi3nZ8a573PaQdz3S1SoiDX2F38OvRdVlbG
7NUL6uN/rPkbmj8aLaeEkOz8iUap3lfAYyAMnRoh5hkAmPVnbmWkfrwdLzEdF2yaBV163nMrbOdr
T0PSVRmFAdPRbqnDVYmUFk4QuXW3j68hBMbLMDTb67FjSl/ksqmv9+UEa4RTXOQIBIS3QJnKggtA
vagtETRDtFbhwrfqlArSgGMZkNdsMhjeXi4Ek0gEGOPC8gxSft5z8hVb0S0+OfmmAR92q+T7XSa5
I17bJWhFas950K57BF7daYVxx40REoVl9WB9ktlstDY5BIK+YBxl3xWqvwZdO54WUbBWg4gndOd2
yKcszIryfl6KxoYX+CjxtWMOv6t5dRX9f4Cum9uTGTGumk7P9VBuLyHZWsTZV1hK/REPttjDA+P5
LCX8QTtaMiLr2/lu9yWkP0XgAKK8DR/lB6SjdCs3SpOi+/Vxcg8LkvAqkxLZ2On6hFBdsGNVFkKH
ApuR4bUHKZnGSxKBOX2ym0I4jByuDuR6YSLBSKmCp9OFyHfDoO7bSLPe5ZKA31tPUbG1emgla79v
R+SCfINjdHwgGuMhJ+MNNiEKo2p906B5buCb/zIthlktNuoz2RXb+1IpVNevYDZo/9boTX8C876M
RfzjnRXwYajJIOKfb1Pd1PBXyCcP9RyLBBAqn5/9VT4QC056OWdkjxwpc6rGW9vvirUF0JOzc5p0
YkNqgyd2uObtKxDuka/dHl+WOehBPFXWwnSW+ER+gq3JPklj9SoDHy3yKhCMZI4j2oJ4NMaK9zT9
nFxKljdf8AN9rsjPN1IYIh84lNnLRjBk8qDxAl6LqjBryy3THJo1TtYLUzuTMpx+C3KmjdXMgzJs
aW3fPzzqtJ1UvzcrQzUIKnrGGJJe/Jmq8hwl2lgPD21Cj07Ul+YEAP15nW3GBmc0owFdH6jVmhqo
z4cdezJPA76fetw5x6hz0vTXftN+CG8XgTuubyq/ShW6R9SkqgDZL1yokCp5TmxrXWXp0Yi3oRRx
XEGgXIHf7XJ1PFlFhDeAJOQVNFPkvgjdIjWRbFUCSp67SqTN2Xg9uUswcjbY0X/uzaQDUZpRf6xC
2nM+pkg115+7/7DDCRv7OGHxumiTq6hZ7UGC3wumJ0oQnGVZVVCp7NBgV4ktpwiSjc4bRzf03tm9
ETa+CuVVXVSYNnvyMRdK6wgNBjJLF2KVcP1sBinO81wsbMeWMVgMvv0tfbvw1j3C1C6FzuKYrI2U
FqxuaHz+QqFpJ9mqbasPafmHrGYL/7v1IoMZtgk4UpLa+TVTyvtPJeX75TMMUyc8jHTLvcTswutJ
eunOkIXKPvW0xnygWSj3d5w9kSWaNlptYkmRf/FnO1b/x9KPMQdshh0rbwyNZ5NMm6w2WbRICKD7
U5h/2CrS9sAZcaeDOgfnMo4vhS2sBhXKLRnWGV+HXZUEIR3hn5q5VSSmfxJCR2AQ3O9vZu+krcOO
l8nd/qE9l+QxSFnDS6rVykmPsQG98AiiZS9ZtMWSG44GlxYPPm2c+JnokMv2eHVEu31MiiAhPm3M
0fzN1RwbhsP1l8EQvKxlV5q611pLczHx1GxFssDsjpc0iLdARenPxsbTdqNp1rsvP+GulrgzG291
Nma4Gbe08Ynzd6AvDXX+6CPSlLZly987z+inGB0NhuYbOrvumb3X3dMotLB4J5+oe5UMRPQ/M3zT
rJVMIZcazZ04i1fgWk6es0eaLXXcnidgCxHeO2Qj77sc3Ha0RQvEgNzE/+6IKmJwvunrhLxS7Xne
gMNoLpyMNZQpHzlXp3TokwlLyrOojCqmn6RxG6IvrMsQ+Lmrb7kbpDgB8PliuMQovgjeX1ovpNbw
ivk8unFmbfhbv02ejIvzdiuTiiCwcSH2BYQHayY4RsNCdPhdPbj2JgrALcdTU6Mr49ctDa3H/wfV
HoNUYJVrJLQa1oJ2FTpno6UkxRJS2oWdM+Kvv03H9AS3fLdjSLdUsLtVi0p8mJvnJ8IwzSngXB4W
9pNG4bugwYRHkuaMUk84YPfSEvXxmfRXgQFphoQOYz60wZ9cvQWrV69CyAXtZ4vZHwtDa475Yzj4
z6kX10M1YGNtnFTKPN1R7uBnXbr3dTkRBtnmogmbrpv9HQpyAf0BPUY5BqXc9hdO7GGiFAyqbLGj
SDLAbNUdFYshFXIsHBIWZvjrP8iEptDEVIbiSj3egd+s+oZ9CDDZKTyDLCptno4NmzomzCnIn2Y6
sjPHQse5RphzM/9V/GRsZGs7y1KN9Bkf9LNqoB2n6Y7+PQAPWtvWWg+y0MgKeF9RzegHWGci8DvN
bs3xIm41uNlQuGJINTZa9MOq9aZ2BFis/eTxsbdtWovY7keC/DtUjnUHEEQYE3D1UsdAe8az7caE
61PeIgnGPeaMrS0469r11Oj47vMMWLbpD48SOoa8buCZdbTw2UU1sEa+Wss+g3XV1UcTZT29ZETN
F7uG+yHTEir+86yKz4AbpWVTzus++9E1Mad/CenQFIelGjVq5Z18CcqLRj+zy0a6zoMVbTd+OvkS
sev/09uWHAbJ50oUr4OIYs/1QZ6EfMv0xS82o43Ad0ZRXprB/2KF/iEj7/TuZNDI+uDteLJPd/QM
v6rQS2mJ8II4Okv1YFslNAGmjVr7xkkZhO4w7aN4bMcPeImaAMnqON865qmJepyOhtCkHsll9+/G
+k8KaWxbyTlTBVd8X+Wp1FXWuCXVrk3NEg900SQpomG4MHzwNjixYlyz3YdiuxOd8KyLnuP7a7BZ
5VxF10jZL0Nqi67qv8dGPHRxvfrKdPVcm6al7uaw6tCXCz3cyC/jIor6RYBapLDIbYHE16/ni80w
SrqUZMHoHr/xR1C1TN12QEBMjMICAGKEzmULulDAM1LVToTPAKQPoEHYGruwbT9kLy11g1F0mp9Q
OIoEP/292mq+js0IZLchP8IRjW60afjvyBylWz9XewXbr0xQ5jxpi+V593Y6pwZNQozUvJVyrYMP
v9IWOR34/d6I1CSCBRgd8iHTFLqRdJQRSMYbFPQnx4ytfK9oyKYigzg4N2/XIuH14lbw0k25MXke
hS+uKDBVtgSf6GGtM/tlK+nQj3dqqi0WVyKlp19mG82PGsQ4pH/yLeSlqecpEF6fi8hTXSkGKNER
UbKvzXI7Oo82EF7n7hUnF87+T78YzvSh6cDhWv+zM9j2td2l0mCa7CRWlsY69peCMt6/HANsbdDv
hG8slyMMwz4pvimhvbe4iXL4gkxeJgJOrXwYdseCL3L/qqlbHpbuQPo4sz/su+8pLQDJgFh97x8Z
9NnGZbeRzL1eFSC8c4eqWIhPWXqksfxQWpIT/wMzhlmztqPn2GLayi2J1I2hKs7bd6UQEqRyPKFl
GdoldQOu6DFrc3dTU/7UZ7hLkRC3Ol2k8/WarhdM+/GUZEEagp2Dn4gMzdPw3TOum/Rp0Oylf8v4
pErZkDvDq4VSZshuZ7ys89IOcInn8KdMaiK6ovHk+oMqBXvaZjeetIXxKwtJJIWzPrI29afYHewn
wLWechVL7RUaAQrpBasLLmjHK2mNToXu4PRQh/jJqgIg1nW/dSo2al8KwxvOfWYcG8a2OqeXHlOS
e5pkxVhut/JrGmjp+RapNTskoYUz1qL3nCon0PDznUi0szTMz6cgTD/KWonhnS7zDtpym7f0U8/K
z1g+kLJVOP5oLUWqN0/ycWR8+icc4vx4wgXefO3aRSKVD+kBaMRgAZ7SWy0tAbaJs1gJSiWVfKsn
px4T18qOJtr+jZFbqVf8iwGwSUYU1sLoq195RWWNBntjXQfhrq+2bEeWuhFt7l2sfv/RSDy+8694
bHae/OL/3LMj8OMIfYhm6Ls0iqyQNOwwlRAvkbOTeUlpjHHIdTztBSUKpEBk265H8dSGECkujEsf
hA4jMD8+1I3K8W1mQK7DFhbrFcQU02QpewwBaq+t6yRvMvlz49np8NaYrSsRhgoCoLFPuCv2SfNu
aULqHFUlGy4UnvdOwgE+RDS82lgNorB5uuHlGJzF2iJxKfUzumq/llaqL7tmwkbfccmpL0NVYHhR
E8sFTNZx6NliLwnvA3dMKSWJ5evIJ9TWU3nVsL9p0PyaBzKFlN2uDqsAGvXeDTUxdEGNvIs160Ph
eYtJymdkEhQ2vGq6dy4AaODqN41tjTM/c/VU/5DMtE5fS1NNM+MJJIodS+q2+zEraD3m9l4z6IQA
OhbuI80USdfpC4RyzeNBWfDo7EQlNSMsy+K0Azh3s8VW1TwTN4l4FcfRsQl5SAiiRfb5AbkHSCvk
Xmh92a2CJtaEnB3jEvsf48jBiGB8DV6NqPl7o6N2MMSf/1wtGxlUfuy5OOnb1loOzI0WdlyNLwxO
YKlwzfC0VBL+f1a7n37ablbSd8Fq9wZzFluiX7jzlNjB2SiYwhpR+Lr5EJYBmqUkS2XvbtfHCMmh
A2lu0Y09fdJWzZ5XQCYFsOYezQUvoZoyzlH2wxSYAsnbiLHmWQKw2nnFlTadzwEqfynutfqJ+BGI
apoV4IihDD93TUISRUeaF6ill8txRG2xL/SXIrmlg78hMzE52yXnukJsOc0GaKKUUEC9XHjMlrpH
yWw9EPHFce6Q2Nr1UDieIMClqh+jsRYrD8jvcsgrWXne7oaodyl8kwyGJtKjZo+q/pLbxX0hAgvp
uQPT6AkM54HNN3lDjbK877DkUekW2AoY/u131ZOLB+Q315Y+RI269SoDBVF90lfEn+wh0yYypJNz
xaU4S09XvrjbXc9/t6eTE1HO6wQ/QByuRkO9xM8CSGI4I92HkGU/OTcV3HS2m9QEzIVHEU5z//3p
jDpggbtc9l0+zM90C2Cu94knwic3VSaZU7zm1aobxJz0O3v7Y8ML957aspjSCxXSK8wn3juYxJ8G
P5IGDYEzlREW0711cgA0GwDCTDRS7WVEHAMVmMn5mbswJ736YUq6u/2GH4hS745YGz8zREsy72Wf
ig2LdfS5XGweK7eMsGgzObPVX5vI7RaBYyLoR3sqNI2rKnhDjf7zYwSeWEY2uiMk9kJkTo1pV5He
dV8xR0arlutJpaEQP6MNtwOZIJ01cYzmuv+D0M0w77pTvpNeezmt5hvL/4LVj+M0tMW9qGTXNilV
Diy/FjY3WK1KNj4XNOdIRGAYFRUk4M4Z3KueZWsNEphltVCUW/OgN7yzgM1Efi3/Aq8ynZN/S1y0
wy0VnDNHlpGXO4sEAIvF+qWdIAco6vapcm8Mrcm3To61t3/qrLJsaYTWDFyO26XPJ6yR72/0gPSu
5dDd2oqWEZuXipEONXAN3ScRGFN+GjAwsEm7zabLKz1h4ALusz5opDVsK6b/g7xUBIFhjOsYDoom
RBSSCvwp9Q6zlpc2b5oUPqIC+YW3VaTZ0cmvVRJKRSLkaJqiB8LjjaqQlP1DWJW/pE8PoI2/biqN
ZkHDJhuyPlsVFS/l5Y0RivBAXYpSkJTrYD4F2oTE9O1scT6WSX3V6YrzCBRxqzAuOTCwaRmT3Akr
G+vM0Gu7qzUQdGwhqLtRE1pYVQIy0SZY8y1j1aD/ZbxW6qNZB+/XA7kmstFoy2meAw0LtKfWhwB5
higBciwihAtdI5SPmk4t1ilKGP2xKyZbqFaLyll0ONczp6zwXQQQo6mdN4u7Qtw6Kgd2elwt+m0A
O/7YkYaZU7eQcQpE+nS6BUOQbjlejE1YP9CLeKmTmvlmpbZWAqSeuV5AmeV5oX1tBSjuRgB1N0YD
Vcm7e3GsuEGYDmKWGiIlLcLWEwU9xdhk6KM+9iixH1Qcp+oDGDCcPKjoHRXbTe4qA5ysOIHwIPXX
9UPek7AvaPGRnz61IwPvPQPXZ3JGMepQv7CJtGmq1hzm5HbiD4AeH+kfaAaMrYdrs7lWwjvnSd/Z
VcYVirt+y0kKxCa3R2pEiotYKRbUPmceJr9m/ZbyYQwBsRFyhyj4Zy6RBmLRB2q26xu6qQE76vSD
XhhsPLknW0l3Wmo0GZ/E4u/b2rLMkHqDOSdmmaA+MLuuBpSdtzjLZn6I6BNHLfGjkHmfdog9i9ml
I+YpBUyz+JhLsqE2iJRnD1Qo3YtXek+r2MnsNXDL2fzUt+5rnWl/PDlhCOFSwE+9h7VVn7vAgc0S
rh8+LZweyroHQ9KrMO2pGhbXZfbab3m9r7KhJniHIOox+ypXdO/Cn6HOWZ0oe7ino2XC/R1lMkcP
0JLlGSb8uS819TABJSIdUOJckqHvvneVgRge7i1q7N8+MkVd0Fu8bef6KtX1EuSFfGoTguPaNInE
/LWCN9EBCc09k5at8lk/3syjpqL/qoQFvX3Xwpokxp4WRjyHNgGHJVw07KHrgND9fLZyTQ27Fkqd
nqPiELpJEicCbnpLWWqK7U3pv4uB2JRKt7dV2bBGrApsHeO/+1E/n0He1vbaIeZgjn0jF/FJTM5q
3/4zO42SR2/T/nr8QrRJ+Z8HZx7C5oL/YXsQmkD/Dp4eBZO22yPxdnR8n7YRzTpxGZVgci2DHt7O
rmsR494Z5eIHcky4m6ecCXCvmjliaMwPQTG3K189uVGbHSRcERQaWw6nLTDZgPIQ+tTBdyxHrEVd
K5Polw53bJGbYD/gFvJxh/WZREzjQwHleEJev9OwhFO5pOnX9wq7xcTOMf2dxwQpdA/aA4hs+za9
uld+slqGRalpszorsqtokI8UnBiTQwgpV5jKAJS+E08i3sTuzNOxYzCKBqddW401ZZYcVxcn1SST
B6NdCbiZSOtBNVGxlokDZdSZdjzy0N5vliif5SH2lGgXTPqZSjVgeLM2PZKwvn8pSizRkwcgQxST
H7N5QzkSDNSsgKMpTozsIbIUoFh/QktOrGEazyl/Yi94/xFd/EhD9l83SLrM8dBvm4Wyx+zfgJ3r
Y0/kFVqqkn4BYTNTFhB8koRVww8KkfzoPcj3k5qLxOO2ecLMc3n2lNAT8L3UR8qxIS/iCq/mEJZL
VQjXLxs5Q9l5jqs5yO44qIt/x9ebhf1EtDRsaCEfUg88N8eB4uAFCJ3FPv1oW/inWJmx0H8njYG7
tD6fIgemKwlwVXGvjyREC7SkUqrQr5UC3sKBsNHSiyvfSZIC/bs1atyXHYkyNXcSCa26QRifMtD8
IaF1Io84w+1pQpwHYGsjr5pR+RRZpTC7t4EhmIWGLl0AyDs6WRBIjrrth70Rc4ZRewRjZ6uAOj7a
N/WCHBDiYRKvUIMngyH7ZwoyyxLUoSEOtPb/8quA+xqoW8Exdv20IVgdAOcF24Uli4LTVGgBPebY
B66DKwYc5XpvSn6kI0o7bxFtqMJfmcvmwwPQfOHUBv6s6pn/qxE7BFq1L+Ksd1lWhCZ98HM+9zKJ
piQdUaoI6PHIYNVi3qjiWg9TnMMuUv/2Mi7KwRIBuzBKCeeTQMTfCkSkr3KVoTfT2+6cVZiJFb2f
Ze69Botcw20gihJzimOeReueOIEhjG6awnljfMvwmJAlcHOfEwQRKyznYcW1JOmRlFQOmyU/y7+w
jo/KH6Pn5zomuzwa0YQv8ChzrSK77S0S4yVblaYuY7SIZozKxi+jcKl1/R3SPdXBKlxSvuKETfiJ
6yKM9pUcrnhOosmMByUxxHnMlB0X7UEfPJSh61CC8iKF11gK/OJVsQhoAcq69Vw9Bfe6/xJfuyYE
zqHNJfWPdZqAGtrqL5ISAfdbwsPif97KUlQMJ0guO4MWABUfqAHufE0Sd/1x0karRP7b6MLtx7n9
k20z0qoj3fMB/eoTniNPjRkdsaJjY+WaR/4kRtdHAoVl2jCEuHYiof61fGj0UxrWNQua6LkN3BlK
KgbCR45LIoQaN398oHW+xbVEdz++3NqvwyGrEstBsPin3WBtl2waVUO+IOs5DzYKy9+bEwE+m0r4
DcEAMasD7D7DXP7s4D6ozLKiKrNfhOwgyAXpLKdta2dZnfw3YIZ6gYc4pRDyA1OOOt9amCw4Ln4o
lp9DmJldzSiubQ6gSM8XRGfswZPsL+uMGZt7beKKME1SzwgcAMEHiUpiQdYzhBD2fBpU7mt4lLI/
WrN9D9sMCrxG9sKCJv5+1n8YkbG/ejMm6YRcskG5XTd5nmOhNg6n1sk+KYqacJZOhYaSDCJKR+GK
7YWS6TzHpXCnjfbXTO9j/8Nmg5a5JtxJCDUMMYeqG8GEarDnzdwkU3ogR/J+Mtww9ZFCu0FBMeO9
5xfxNtrB0vl1hkObEUSw+7ShzNRLl0SGwVvuX0hDW3TE3JE8XP4IjKlQKmX1tzQSXbvqbnMW8pNa
MgDBp30oKv1opW7I9A2KQjhSAbpQQPR0c1xAy2EKeCaOveypJj3H4G11VnaAOuztcXmIhzaGqn08
ZJ6SdFaBTY4Y9ze6zMQZGn1/5RFtqteMt5o/Yuse4+qaLBSyZr5cV7tF2lTs+HURA2Vn7kZlKyt1
5NwS46YM9C8XJehDPFVa3uZkTG3FuMKFC8XhyC566K82wOiSbDvnlEXUGvU+sMaPS2o7k05pCCUi
cj0uWALUlppVU/3R/VnMTVW2VrUNtgpR/TNpYTj01qpdjvHZJ4RhZOMkSB5u5Q1lA82TjZwLBj3Y
VAXCZPPzvnixGuy8wZf8r/16Ex1u7R6IdMuiwes5eL2w4lYv6rXw9notzDRBfUz1VbWIvLTJ0Ru0
XrjJAasov+0zf/tcJyHFFq4MB5on26NQPc1q797oQP/pQQxpsFn1QAT9mT7yeuozTaNYRhzSXl/X
CgirdzP0XyJTJqyPXWnDfplCN5zSgnTRu8ukO03tjBl5SYf8N5YuWWSx9I7SjigLxeVjGjWbXq58
ss7Xymmkm5qVlIp3n9XjO88+LbdUAxYnIXq1Yospa5/ITaibI1ZsZ4rJ83N6FOq2cxGAdrjpmLMM
DsPt+0Z46o292TZmwUQ1X+h+5VGVuWRanC+r3HkIo9YuHhOxxG7DJ0JOdi+RFuKayyYmBzh9HBD+
JqsWlFZZ023SIn0AXx0rRsRNnkxjckSZwgZZeRBTPAplYwfrebs8bg1bceKdkAZYlrl350/fjWRa
eYXMBHrQYB5uYN4mhpQEdZ0CDMB8eNJZ/ZCvEIH4+83tBMvbUQcDZn6hIDpiPcSbyMMasi7Rw+Rp
4Wxz84g8rFMw4rOo6ljAbXcOtiXCbc7cccBG4ESpCJf1VMqVE8WU7ZOQwwDvXb+ujWKfuuTFpWwr
ha5h0HW5Lr3KmI3WbrqKOXu4BoHXw00iIXHFhTzXqN/+SaUVMHpQWH3cJMsQlSvGKAA5XDg0AZ+0
ULblqHaWgpvj8Had1mXtcXuzf4RIbXTlNtheuRcnYVhf6ejf+51RqYfpjEY2dNCjYL2IrInM2GFO
TYtfBlHgv470x2ulIWSICiL3Hux/+NhcDMKebEkKZ+NTnHSSIU5aceoZo6sl4loCQmzFermEpyo6
kla27dBlRMKRTx83aee0fxOjLuEFHVCN6T5pqOZmqviV6cJuj5325qTbAEEFC3wRG3TH//Me+QLj
niomO3Ixh/YbctumT/r+NN4cil2I6vA+3XKNAtX9pkr2RJUcqSlfqUSAVhkiBwjjYvRWYK1kwIw3
y9MCXJtGQBIlrJ1f/IaOayhZqRBbgDdk1c9/3ChRG06ruH1HPbMFWat4RbfP/ylHt7HEpTQpK26Z
5xFCJT1piVOTzSXQoGvkwR56/4hd0zq6WnlGpC65R7XQXyp0awCaCuOrrwsaDsBkOJaORp//JwAv
bFKpDP/wWs7c8K7S90CBovXCUObnZ6KQAaJ/yCVN6Nshrbp510uXf9ZEyJp8JLiCFwlsflgnwCRU
RU2dNnzSZg+V6MBh75eILE9e7o/sPy6R28+ecYXfg2mIXLFzg8LidE+KIwTAdsj2/oVF0fsPqWXo
DlvyLuCvtWkk6lwwEUGY3AG6+RkqklRLnHCadktJgxXLSDKj0mr9ZCEviBOIQ1IX2m4xJj6CwJkB
92iZlWopSMvFfYmanWmc/wLxQJo7lG4y2k8NRPYd0eHRhadt1uh5Mc3MVN3N2YZPJ+KI5yqUI+ga
2jFACp6TgeJfDQA1YSCCD3EbrzzVzf/vC3C3MhYe8c8d6rzln2ivGoXkgwQiIXoRv8/s/KO0kvA6
UEuUU1XW7WRQXkuA6qwrA6fyFcecLfzqljepogXF4xr3r+oRvoMCHuBj8GKaC3M6bLXug3Q2ScJ0
Ey9nI9WKPTEIcVxt3iXTuL0VYvXR0x3RisFkITIU0HhO592Ww+pQqUy5xj+5n0Oa+FVKjj0gdpxz
MrdsPTIJpJwVI4F13woyfgjHfju2L9R0j17zTvqvNywbDd6aWEG7XaemD6RhnXUEjBSTykV84Ky0
dYLpp8uwyvJAxrquHcY7KEqnYHjuRWHMsIpitlmg+z0YOTFR0GsBy6QcqUcb5paUPoz7W1M9HDYw
f//fqAmx1n954950VKTEdlT0emqFrd3VmsD4oB2qCFNEJZjKcy43QS4KGv81ruYIW44alXsebrdE
GfQKEbieWazBbDG05xahiWWahONokd6QDp9WNtBTcQZphVGl0PND9w/1r4OWGdC+vDeRoDgoDVjw
YZruQrwmmuWSqWK9OajZcX1L9NlTl9xK6HDPGDX8NsBONDAxymaQE7CGKbkMzaeDCS8s9hHm+jW+
Ty5e5s5cB8MyhWPJPwjI0OMhHBtU5cMJeTDxLLq0PNE0A+KOM6AnzqbEEhLWxXurXdSupTvkxhfG
udfKJp01QbOAMgmQkqfW3G6YizkGE3cEdPJJLhEjtIrKS4l5wl/b4w1S0AdRe2MuKEdNmkYtZrn9
RuNuepBJZxMKyJWuDO+NrHFvGUTFzJsmpz7Yp2R7xRAgX8gJqUCtRFKwP1cXHF5T/+gk5qyWjy80
c/gfsOyxes93EPZTFagjzAJW1kJ6CuhoAM9QY1OJOF5vQQXymeAFNb19xjynSKBA1iL5gaEBBR+j
PYJTjKyFUALYLCkGmukJKyLx2ZfBXyyYzFlnsZLE9jVo2/mncHBf0qFKaOW+jQ7l56UK5L60G3YY
Y7TcNzLcyv9I6hkw20F9hUsQ6tpwZD91Mkf/f/DCPCjdTz6tWyCS9BNZoIyqvBNaUZtfUqs3YD+O
EideLXuyKSMRqFZObqjQPGUnKu7VRiwGtIXR7azJt8rfgZTUPwRwr2622363w8LMAyFqMyJFpHN8
dMhGeVlmXD2QuwRcSVV7UaSrBsGcBn/WnpweI+WX+yBACB3C/uEEZ5D7yNmdjsUCZNSzWgsaCnh0
nNuBdiAS0Q5+ZL8zXCbNTum1lWJki8BX5ozTWtU/1PaGatsfiJv0TMUbj+qYh2MDjeQF/hqUNrj8
3+x52g2GbLjX8U7EFeYyBCONCPJN7DTSQtV00zuHHD4j8I+rUcN/DHlFQsPQhNFdD4T5HZzjkFUg
n7ijHdvJBUsD2coA1YnTZgIF2Ph68NEwLe7zPzuwCp+msbIsKuOZ33PSnVOdGmEyH2oFv+G/Bffj
IxGcmxYTGqlSmDmX+vZFiyzUeP1JnnRJTwvxhuK7ouJLO9MB/TRSt4loiYY7G5Mwx7mcPs0+LZ76
CwOEVXhRGzX8ezypuQ9HKbrcLY4hEYPWzUQ/fbDxe/2k8e06duXcg+IcJKKVEzqlWwk4hoX/4XvW
o6Z11rLp0WQfbJGeSOCJO4srukjapyqVoYkcjYc+N8WDWOtT+2V2f3lUTcUbRymkJEIJoXi6S2+b
imHSUcUt5G38bzsZ6KCXVOSzI91uVGLAX/rIy+iYdgTjNr2V38MLP4qV4TpGZuU+SDalWksELz5q
FVjHMYPicz4/Xf9/N5pgqUJPNHev3wYxKweMBfPtR1QOFA4TNjLdTmYasXYOYkQMbDxnBspA8Js1
z9Rdvff+zP+VTBowe77gFxU++gKFchZTD8fD1cgdGlNUUxv8n9NPXh2gSnyxoeLgqvELi/FU4q8y
OG6HKrtsgx0n2PEPoKQklKcD/Ld64ZUj2pkUl0Kz9xzIDgXzxDTyta2rmtnH7pDEJnhA9Pjw4FLW
hkx8ck/SwvhA1AnqbOaivA+6JSsHenCb18iwyxz7G+4KdeOtxjPBveYK4PCbw8LsSNuefmX+X4h9
su2S4/OF5gVnb03w9C9ccbFzIE4ed/NJCMNlF5ZvwowuHbJW2MjScbhL1nwXjr/gCHbVmsjiPFHq
c927D34WiBib+rnHHPml4SDWeHchJ7fXoS9/jEBMNbXH1olhB5dxIAHyDeQbqqrDuPQtVvPHvvIK
RlXhj8cgGQ79x84e8uyhLfD/UOalUcSOIzSraHdRWdAU3xdQ01+CcSXaG222IYPBJM/qrEeR6MOB
Z3htvH9zn91mu3Wv1B4THSnk20o2dFM1VaXBX2vasmCYU1c1CQiGCrUGMrCl2dHDADSHcluRGyKm
RzCUV2SeitF/blOW2+23IpksJEO6w9ypcF9eo2iseCYE6mnmtv+3j10z03sPek29dcDfCQO05gzK
qRnlfXTn8PMt0rlgY3xBwXW0LLWvmiV54EJLMZi5WkyDybIbI8g+jkdvNX1oa17ETfSWfXjI9N7g
C1G7QwYmMQe/BWF1uREbxxCFA7s5GglkP8QQIY2PVA1NRnNprhALolC05cjH5r5Yw5WdfNbS+sc8
yHoo5hI9XGIQYZM1AWoDTPuN/8Zuj5qhzdL1CV+YrtB1a1FDW8pE3233zLbfFhOlwGczjFmt5wTj
WnPkwuzPoBo/GDqCVU7Wqh+xNdd2ZA5ns5zSXaMQUXgurbehiroEtWzFOS+xTEAWsWoYltAyH7lI
nFjvax0JiwSahaFU1LNOnt0F2If33O10JiAe2tUv/EhmQlLPbeW4SMf1kxylojQFkYsuJ9MubQf4
oALekrm0oMkUwb9ZyXYmQ3bH2vqn5i++j29MuXOdfTg0VvYMHTUwFTkEZMRPbdHwkmXa25rHa+iW
eaw2Jqv5C6LlR9Zbfg2186YuNgZEhLk7T3V+c7u4abPQFp11Zk2ma8ws4ujvLmxF9ljiFlq1+k6Y
IkmEoy11iz4IB6ll7n7cuVDyfIGUn7/lzZ8zEfspWEeR3LqIw83c2zY/H5BtH3UAkVtmXzwlLvoI
pYGVgD+RhaV1zBNnHicFxQflfcK1+VKVdLDCGKQPNI37JLcPoxN1L8i+P9A8v4TY32UPtfFqb8ju
jU+X7+qxlXTlK34Ju3AixChOUBZ2knoEpSgO2s8Q0tg15BFfFMc32FW0iCAo8Oy9LY3/zcfzAeyr
Pf+WtqaBqEFsPjDdLV8lJ8FCHQAiHSq1sE/58T1QDLQyY60cR8jzRzDOYftxhPhRp8g1q2JKp7SD
VbQEbX5mXt5QNmaivnv5jpkIa5k+GsENxsuvWewYzqNRlxCUv8kZa6cR1FP2poRImwJsw4KUIW9H
vdbFwPBRYn5fkq1Y1eSvcR1lV6WpHp9Oz5vPrWjPeW8IRDGJbGzxuw4T1xOzhpk136SpFBeo+517
5vxgqhF6pHcWNe60fYAWVdwyqDOCbUCl8tJu2otn1gT8MdHPJVIefRQppE9RdZEPa5pFKGv+Yzom
+N5I2bbWdhQlLVOHIMPRbfIWHtEz+Ba17+0WBQzgMR9JLn1wLN9iXTJ47KMFkgyZyiG4sKJfW+6H
H8cP9QW46dvazcFhxnG2CBFv0bIhgz3F41wJSt0uV8lJKxPULaIaLXdSPZa8q/3rvmgCv5AV8e2t
RR8sUEo6KcBlTGz+zBP/qn2eBec7WtkILSYCLRXVEvxLLUJfouyFWSY6HZkjHWLFVqhngLsdNOte
qQb8BVU7YTXJZjS7EBinFCMzibk7NkokeqMrgiaEDe5f7YU4oLilG14tY9zunmacFYXaqY1EqXF7
s1rz5HXZy6iOH1fR25PVPyozj3hDrCwITqsxX/SU2QVt5XRkgLXD9tvownJP8c4ti19TQtpKSeBa
SRJ1L5m2yxyYwA6WtWqgZ47UPrw2TNhveIYZvcj/UFgy9/CFtp6AcsGnSx5PWFNHhBLaOTstw3db
AUly+kMn+qB86X6/nxVXPgUm8UReWewfny7uGxZaLnSSof/srvgi5P3ApbbGN5LC6rCndS110EpI
eWgnUUyPSDMDQ+owJYA/SUKZCNYt1gFTciml1d95FNOE61YFejc6QKj3ghLEpmB99RIZCuBkLc3K
Mb6y/NADsb2JK7Spclth5ELaaQNqONYjvGd3B+Uf0wxmGaF5/V0H5hL5pFu0m6c9Pfc4KPUAJtlb
MRSwmVOSz/oo92fSaOkGWMk/82lm0r+8+Cl/5bW4jFDyh5+i6pc3e835L80driMMdPE5wppETAXB
IjvqR7qEFQsIK3Sqo3oWVqr7+LS8yJ/v4wAJ3WHPkH4hSeXIBWU8XAA8nKNInGexWLH/kcGn51tQ
v+iqnHTDwfPvWzVq+7Kk/wzvXYMKazV+5biNakv1SJxyRD0ua+1qhjnUexmM8yVZqVLmO4tJYjBQ
952qKF/dt+GqM5l4vJ2fgxD8T3wypblMaRCCOKFYnaTDPI+gyRmcmaaM4BfSm2fjMTotp3Yo0lEt
XaJOM7iPXE+2ukpiRqTpm5t5mr6JGCXEMBaL+A5r9BZuuO6D1lwcH3YZlPdrkrITV5ZK2WwiN7e9
8iA41K52Iwrlxwwl6o1D/d583dHN7abpfrSOek4QRQLCWfP8H74BmVMXXZQI6GcYmaoysLCr3gsW
SjGM1vLZCP6KLDxKdUcGwYb6NHNtotesKc5COF/qWRcfmvlwtLdvYTOpcqDS3ImZ17C7zyWBVCDN
BTtt4iznbaUkSvLKxeUx7uDsANwlukqrCedgAc9Kb/1J915X2fMDWlMqB4nf/uvRrxGTFJYVDFka
k9QTxyOMEBQzSEyFJ2knpax36gL7Sveeh172L4k2KPfmWbINCHmiApwBadObolXDXv4cOgsrqf9r
7H+1lwXhOHDPcBns+ywwVr0pZnff0U2GFoCqIJ3zYFZMDedlUzvCGMqb9K13kgclCkBEg+pfA1O2
LcQUpdu8Tl/r3Vxb90AlNOGlw4WfqZnx9osN+dW3c2nUaIWOrm/1/sWeFhO1xQQcHCHEGmki+b44
CZSWoPL1h0DkIYhzV/8KLaIZxziknpW8lvK00SNf/GRRRRpyZmTACYAGkRn2S+p/x2l3mGBI0/iz
a8gHXlZWfUPdU+CyS4jA5Jb2qtz5HSwNhCAGf2uecJrALLKM37PS4JuMvR3QG5rpj6lKIP4MO5Hu
VZoVkSR3Fk7BeUSdRhmDw4TBWzHKxvo7SETiv5/jGewul6sc/EH990ZLBCTYyIjB108WqZxEe94x
iK/xReYt/XCz8+UltIb1klby+g9+ViYYVRKPu0SgDho/0QuqAUdNvGsMuE15VNlNb1N3ZSEXifX1
V1ikbPfcYlmSWPsMqbGzYGgHCQYO1EzPg0czdsHianwhe2LPM6A+Yb1Fafhr0pvMW4DmJR0vieY0
r9gI9u0HIHPs5mHnWWambyHMGEKIUjG9b9w7VWnEbjY+1O30TWErYJ+kDfBLDtB8hiyXAPQMSXYd
9sYjnXtOeB36OOYUBO0XUja3uuIKdW1ON4vqfXz0RQYT7A7Noj6Iy+Gbujs/kCyqHYLAGv8Rd+U/
zgE00vWzPE3RnY0/odgPuHNb2nLUqITQ13Z4mPKzNMl1GP/fUJF0K4r9KuKtqKbgp9MeGslQMU94
t/223FcH5vo0TtaE/UV+gRP3oIzj8GlOkMuB5cuV7em6rJI7hVCcI52A9a0VTJI3JRoYMkACpWCw
65T5IcxzeOtu4l9fKu4+QsUT8saK8i5zszLctYwMrOIiT5HDfdUNpHs2uRpNsL+1JrGZjyI/kq6c
6ejav3ZhYY+npQMRhpMkHIXkYowrP2J2rbFDCI/KcztffzIKLgGrMsmkqPC3a9rRwKJK9VD3JGIL
0yB+1rlMJeEioND+sGWCQwOsUwRIpYUFgusrKUit8z4aHFSPSkBRi357NBY9Rs2Ul0bS4BeUEb7C
B+CF6et27TvpyE/K9rBKwYyv6fRVYg215j3T1M4abpjdRX+9+h+qoLDFJwWFM4xHO1T46XGWz2BB
dVdqwG68aiQGWPOee+t1EeppE6NU676Khx5eLF/sIyeMz/pXFKs6wTVX++8wdnd/d5J0bigf/HCr
Wsojp1EJY1ZjIY4rvm/HuwNiohsDQq1yNCKfv+LHlsqgEtarDN3pjAE0/gTbaUOSqY33wiiHYfPn
2X59+SxcoP59TzZ9UJdFdNUWAiNwFaWuUh/WcTMksxENXckTVXhVgBWR7rvFIAa5hrB1AzFiLWas
ierrwv06EzJw/puWGAPwhahV5HkK0SLnQT5Vph3EJvf7PnNgj5DVjnhfIlARLHc3Bch6bGzVoBN4
nCwLxsdGGbLgutu4sTVSu02k0eH3iLx/CZwWk9YcdXCTFzwOaCCbO2lcm+LrP84zOBx88Rtvdab7
j10TqzKzqAix+GWGflGMEvTADPVjEpYnOsg9lrZ5jTHOybbbFM9k9NmdV+5+nEfLS+wtxHylsQ0E
ndCpmN/LPHpED//UAyeskqIsbquKyJR57FoWzi5agoTV+EzzhwMvrtg434R7amZgEWaFU9F4np7G
Hn2gxKVExIuuEpKSslGWYU/UiKe2RMuDDcMAJRwe3eU4sqLUg/WOXQ+yDugZ6RcNk6AW8+LXQN+n
Q7A+cYFfNorTkd4CcW+6tjjr4pdLFsjEwCu8lv/+dSfXcURKfrhxL0ojSVcgKivKytjunD40fcXT
yQBhLyNDCgq/Q442dn6Bb28A7FWlibI4d/6LQt86QhiwFlzUkGigMyDnELXS6LB7XGfwW/xXqCz1
MSP88Cy1VSM1ABJ8D6icDW0zhhuC6JjyMMRin/EEaQW+gXiWgeZarpTRL+m2+5OV55aj+C5GXgFm
MBGLYZF3hcrASlVd1hld5kZnhnf2xehsmw4RMIa+qlg8XsMesWQZezHPMod8anCwveFZjnE22gJn
57/JcvUsVBLaRiztUNgIg/9Apnt8yzQoIsQQ/J9Ois0k9cNJ6FmWJkhYQk0qvIbRMXAPY+lLJg46
RxmiyF2HS9g8QofcdrzaQy8v9EMZcUis6sHgYULr2zHEOnQWTFeSAmC7cpcS6jRUCo0XeEezJVso
BM76gffBPX8PFmP0/HPFg9oh9VlzVnz73qZchSfkZPoJ4cCG8e1+GhqoAUIy6XK4eKmaDfCq9gXn
5RlUFV0PDjn7bJCisVQblTbD2Mk+YF88lsZEo4SnBVNhIGXI6a+3L2XNBlAtHLlcFNvNvl3nBtK3
W3NIN+L0fVtGQcu7ifiTy0OPP/caYlrx7gdGW60xoK2iy+syZO4Ilubs0WRjdmZSIN302jiNcIui
xgm1C+DRHQe9nNJNkSzu+oBo2Z0I81E2DPVjuwLa9WBKBX5L86kPrx+hVkxqfnZf2m2eDiQzrEYU
xOWJY16/EmmNtfS+hNWfr670naAKn8WMK2Zb4cK/Jox9RAnM50IOHVN9fdt+qAMz5oT8iFZGK+ht
tvWc162+wCExEHS1wM4qwiq+dWBMGRFmkJBi3Z2Ymvszu2YuWFDYB/LRbIn0UE2w6gOpw4K0g6cT
/Dpc2gqLg6swh0iPwA3QJMNjLoOuVSoEgSiolCyd8/ivd3VmVbYx7yhzd+uxKQlTaWEb33ZsThgb
SSp2nPCpyzRbGhVuyLF6kBgiuhpaByDbDZNHD4S8L90ZDnpMbcFzSeWFqwQduJJX8FEZ0EL5SEIc
/uC02WaVe/FxmnNNj5MZdg3a9aY5x4maKvMLTjHDIxCx9MCl25PoDP8hOjY1MIfwOXOFfqr7sueD
FenvuPjKDCu7YRSbewLI5Bbqsdr2vn7CeqPYxVoN74euGLPwPWVkWfQb338LW1qIxSHY+wDL+2ps
qhM8WHQleXetQKtqka0jxaF357JqNgSTcABbxxdcjiwwHLSlODyQTrIxykU+ZeVw9dJkUcLmP2vP
cQGFmMrV6r+DJ+HQatBtHxXsb16gC2hRfTV6Qv25azastLkAwgWwWi4spD+VLVdTRi6M1q1e++eR
0ezb/Emu2KMkAre9+n5/i0DhTsKGngogFBsDlTAZYgZo+hN3+LBpTm+j5UIrUMYjZUJ0l1bhnXI6
pJb2bSKnlI7DEQvxRND531RvnVxo74Q5w5Zs/ADO5jxgDKM+79m244KlUVPCxnpD8RMIGryxJgbs
gBh8BPRwIA8QOrVCOv112ln1ws+pymQa8fQ07OxZqxWm0CpkHx/uTTivPPzlTuiAzCA1xx3BCq9F
UkAyYVxv/5w65D9JjWMehw/adY0Zd6FRt/m9zjHuqIE/derGmGKVxHlQj3+/UvCl1Isehpbv7qdT
H7bwEAxcxJQyOyNUpYayAOsjc9uRixPuvxJIBaUsLFguoQMv0AxS4x7/87yinEWKY3NeDNCCtrpb
jTmeEgqhtEnqmRkss/XhZ2ZtJnIUSvsAzJPUTFuA8ytQo8nakgH/6qcL8y2si+hKdpx9iz9bwewt
9AU8JEdwXpFr4dFYVEaQGS47DXgPVYyN7zUdl8RBTT5jXzLIj9fXxSUUM7L50N/4FvOzdoDdBV6L
+5iPKbRBq0M98Fh0KLYyK0ZdrLEuh30VTFAAj/6lRT4LL8ur1LHDiLUrNZIS92I+3+IzSgLnRNdo
xADmKEDmbgazLGTxEDS3nohWQx0QTnQDOyUWC0YGVAOpxqGmZjt8mqhQVRBGphZq6HzRm/ku6NtL
fZll2qITsOLDrhohTXjBFnXgDW9FYDwoEgVG3taB6xxNPpoQUSaTI25XJ/9Ld2mqUJplo4gE5gqs
wjtYrt7rNLeUoCUr9ODO4KHnuIMHoh01bpOMabzDDtKOPKMKbx9icEd5E9LLOknNB8MPtoUD/Gxb
AyxdyjlBVFYqDRspupeubuxUNaJYe2HJyJpekWwBzF3f7YlPGUG6Y5MuEgI6rZ01sGLNeFRqJODv
VVy1fyAGh7KgMo/6gFTtsxLiDVM6eL/vgbBuKQQzhJOC859lcGzwD8jVCx8F1TnOlSzob3jMhGON
rvpme/WgRXKUc2DptoPWANjOQFj28SBZMp5RoA3asjgJIANLXddfY7O7j8UMlr8EVVYTr+KEpngR
20VEFfRbiRk997+tYWrRyDr5j7OpSFPn+IJbF/fosBorcUzpIvF+I5I/uppfrPxcmjzj+bLZ/8kx
V8duTnrndjhKTDQ2ZCJt6WoWbfaA+n7tXs16Z5yeWIYnA53isAazhmmNEAhUIjQdwtH6taXs4WaE
5DGW9d1VadjgnrAsoL9+2h+C9mh6K9D+O9Snd2669u/E3RBTozj/ybHDVZitDJKK3edj/ogf0Aa1
jZ0tHMftnNNRSEHe4yFH+0eXV8As5M84XuiDgMJEQ17R/xeEYgPH+uhLmkJLwReKv65sWzCNVEp6
fe4ASzu4rp9LdfT3mx5Epy7MRVkDOdL5N2zyfLQ6M7uRZaeNRG4/gQGFBNbLsKu2DvHkECRwh99o
z4++0v0/IUARnhAva7FdkD5l0C2KvYl8cEay1e8GZUqMVyYTlHeGeu1CNbq2bSgoOelQqY6gqJn3
8WzpfrOW4pPuUnXop8z/0tsVfNGS4ab13rMDucZEfx6hKHYU18+61quQib/yb1Z+/k0sK6XkFpiq
JrJJCUprP7U4thfENjxniXg7kVKgjaIDUidb8osjSwhguZ1F7FkfqNqfm5fU47EBHVKO2pE6jY7c
/ifY8H5rAmU6oCYNNPtfA/wuXS722zMoNIIgDy7uL3Y3xdGCpJ/Jr4zWXFbUqEtCHvnxGxVxD2q8
mjmoGg9+1Qn72aHPbcHUS68Jm/kCrN0JCM3XqDed1dOJd1jYr7YoZV1mqSq/sUqN7dmGCU1Bq5kg
35rGWUMrDDhA+Luzd06Bo5y1CKC0+gZuMVbTO4Whp6m6D/vw868D2AZhIkK5rvdYCF5SEEJf0Zmr
N+yNILyH8zWQw8ef49y4cXVD2Ak6ETItXwJyqtCLA1ttnW/FHI2/Q+E07mKBJdHt1JgcimQad19N
SSRD2C5cuMg1AMdtnoNIHZOXUascty6nRYFOOFYvltrfo1mjxw26VpLz0tWx81rxSWO3grgyNVA9
nGDVLitOSQvO2SlcleO+43CLz+m1WTA1WoD31K4O3aNQVaDbzxgzooOamoa+qmjODto4PGdhDOnk
uhtn2/MAV9yjhaYIRZ52gfudxIUfBNwt/EXTe2fOQJr/70fxR3tbtYVJO7Kcr/rryuP1a+G8Y1s6
JTO69lfDZRYRiVGPifS2yCvOfKEnmb9ysYxx6nLt8CWrZgnOPAOUB8tsjTQ/Uglwnu6XLPd65IRD
7XDnkyBDgrnYgMw0QQRDxRRr1eu7o/M2atRIJ0rP1rTiBhe8omJ11oaaLjGs391PKhTKR0js2exd
mgFvOAJNetrPvX7r1s0MZ3LROm487BsAHihvGFbZOLkoGN/DL4oLxi+vc8olBHa7pTGAKvr8N6jG
bKGxHsS+MGIID2PX+AcbQUr6sMNV0FmzQ7BsMZgu8I4Pn/GSuBu4KBZVu7lxzHgwYPte6C4ryTaV
yGELDKZ3HBFSS1KrPE44xoE/9DCPnLkEWBT29h7jc2nIemsU51+hDUt0gxFL0g+lvfhkbj0DzkFP
3qfYCRYy1ihp77JVUYjjz7UyX8WHTmyOgYD35L4fq7wosMU0HHGjeaDiT6RAY6aL4vkz7xaqLVBP
76tyZUbuDIJkpW9+B1ZWJyAKiKPXIBMKrVyUVWIdaZ4O5qDDIU8EmYMXwY5Py7ceA3J0E4QBl4rs
dQ8PHmQA6f5LIZi5lucuUPNR+pY4fujqmhgoRQ6G5fkE56m6QESzBJNwuGJl6bHsvXTGvNTIMBn1
W1tgsZQfoBO6BcPiEkHUaJ2+4l+5z2FDgzndf0eMALgAog7DSKsj0kV0KfFFZDHITjUH0Ekw4Mk7
t251lyaiUnGQdpFBWoWQK11HqCTRDXzGvKGI3eqsaZWBLzSWqUJVT26nPuzmbUDYwd/nOkwBBpjW
/s3RPbmEG+jAPeLRysR/qiRkqyxx9E/o3Ld2cUfdVePLXJLQ8XfvxVMkDUmhSZSZRvOWt5CYw/SS
/G707GfHo2DjtsVv8YdhCe7mK94q0BLYUE6hJxckjd1umzcvCINR11KECNN/gNSJewMqRDWTYSFM
JsU/y/Bu8QhbbJ46lT14e4isfOu9R2sor/QHKsPz6sJpxKC1YDMOkDkQPln1OSZmSr3UJ8opbtqq
bihrWZvUVRRb+CGjS2W2BvMBwAqfEu6hRhAgLI2QWYLd/bfEVOqQFNjmdDuh+IAEKY0ELd60E9hX
ajn3ejJu21RVAcR/qUmDTN4SsOwcIuO/BZRn0hetspm1QQzP0yRhTAJv7JEpdfgKQNPXa+2W8Z4x
kHwXqeQEKo/kWBQbWm2zHzUJOSNJ6/+OJmOlojcNQD+8yvvMDxirNn205GDMklNmeSoeyoowEEwo
u/Qf8jMAbKens81cW85P0hFMR62exhAlcTj5ibz5df1lukznRgdARrxtNpb9KUIimF+Sw8zOs6FU
p98trGRLEa74uKsct1PXvz3FvbrXfnuroB3BWam9nD3YTfF14xGHI/Ll42GXCUjqWkZlH5Sa76Tw
2WyyYj8Ft7Y/vnzv4gpBNqzBRPdr1DHqEQW0TjvqFsY+7PJjpKhMVfNE+cFuXtIjFVjRv7nmBnAs
YMN6jqa9hdOLpFO2jf3uJ/kp9/Q4cF0YGIIaHfVRjGD4vMBpvUERC5566vz5OoNnIv8cC36RVRjQ
6UAFvcyne+XJc4p+2mm2/1P4AUh38yc+4FORYs6QnACGlNj88CQqSVqiioseYqSHQQdIQNswKyJz
VPhcvkbRpSohXD0mjKQMs3Z0AYKLlfra09BBJwyyloiQg6+4EmF6yoyD029at8JBb/I6Pva0gT8v
+YmW+GiV6ymQq377gtwO8/qLhzaJI2VnAr/8yjuM/K7im7N5BcYmBNgNVM2ZHrBevOGviDYAlMLO
NIO3FEHny7BDrYf6+UdhdnargDimHvC5pC3L9eKWX2lDN05CDps9JfV4NmHbdJCxKDBCJN3vf4/Z
HmOpLSNcQpQuEzfhjxl8+pXSxS/t6cpXAWGGLfk+zj8R7lPy1W2IVa8zNeaYh10orzzuRtdhv/ij
ORzrhgrljewd8d63BFg8dfGwg7V6ffx/Sv8hqycnuETJd5CGJgYiT0u7c7vjNoRf2ysQ6Q6XAI8V
o5kaUt9l/E4kVKqObJmSO2WC+RA5Q/kBtEmDozZSawvuzATJYzXyYBjWIdaLFNXkUtEtFsPbFjRJ
a4MhTZcdSLOnX3lI3BePt+Oz7mMVt++Ei+PSOVOLnQEYNzaWtWAcCX1xCi1tLfU4hq3A58Fh/Md2
yt6A7mA7H6fmYjYGTXbL2LLZds/h449/dfnNvsBQWh2Ep3tvBt5/5YnPh+Ab1GK1z9wl1PlY+cV8
OYeJ1lLbOYGJEzeDGbCWs/8ZcYY+h/2w9eTxO/MQhf9y7jFSiu3Peyx5szdKmiq1dq9fwdv5g1os
yBQJo7RTG58CYgZDW0Lme6EleOOSpAPwY+hTvoUqcH1QlPMAWaXEq9N/D6JKhvxbRacPsEfZiDGz
Pme+S+YmqjHFQrGHBjdLSF+0i9gSmI9NiqZmLWprH76BwyyONiMqBCdyXfW2okR+xJ+8GueusZWQ
0uf4YH4lEcOH1x1NkwGRmXwT4VSOZioo/gcbsfpspXLmPv1yBvUQXGj5n/mB9P+XpabjDSSto3Ba
eZ2G0j8+/rn9mNVGQ7j6jVhXGu2ggaf8yzMrV4uIDUsDSJtqGuv8B8CtCufCX0Uw9lOsraacI9oQ
Mzwqj/fpsXMaiEhFyXReT/cjV3kNmYRKq9OacH4Bxu38QT86B4nC0ySsr0nrbPKRLBbicAHb+pCD
yLmMgw16NAenmDJD3KklKfBBsGxC1eSSBWiVA68jqYc3Lyo2K23tI8RS/ai08qbH7mGtfmrS3lvp
6dsYjFCV/4U0hc5+1NoQyzd8Aqgyi4biTxDUcAyKmMz8b8oFe75jIkKp6StPU0f2iQcpzfXbGBow
SRn25DixKoW8iDxlUx5RgpDqGy/kQ8kqBBoHJXsS+pDx95ipRQeXw/e+9VZjpDhWzTBua9Qnh4Qi
1A/qdWY4W8eIF6nT7jjKPdlkznsVeU76aa+wLgldUjRYO48r745hO2uOtxHQ2p/PfIIqOXKPLbpx
rNT4E1pPHjVl37RhIT9XHwKN5ibRVl5DRug1WHB2Kb5uSxEBXPzQowjTRffIfxtDE6wmsSIRBtaP
V4z9+t7TWBNcfd6bEmtlks6RsJOQCvebeO5QSaK3niT+IC17b59ZLU8LVp05ash4v9aw4rcOl2k+
N/kJhvc3qgA6PS7cE4WsHkCKoqGgmn1q17ZaxinJZj5zhWP//OAs2ZMSaRzIuK7cWMrSOQA4mGeK
RubZWCIQCzPSZRNucqTxCxAR5O319D+Jok6BilcDFUzH5CNckQo3HZiiEd6edeDfK2u/1umOpbGP
TrZhz+adJpfMPQrU8tMwSozmb8/PmrnSF1/ShXhJDxb8+K0IxiCbqVug3HNPaNrLBv7WNNv5ij2r
ITEVbzIbIXEfaLkCuLFtCHDOHdbccOhHp/6s6USUX7Vh9lOD9u5UJi3NTTIsjWC6+tUszYDwTRZf
mBx0uJ3DiaLbg9P906Z3KdLohy1Si4B6bkGc1An3rrxdd212AThvp5Z36JzLzD2V68WMmbX8mZ2M
+eMfxzlI9avRjDFqW3wXJT+qg7IhiUhKHvEp+a3wEsu9my6ZNngAx2YCTD4hDGV8v8Fxw1XaFAGe
S7tk6F2OepMf+auoVgn/0UCmEQIyl5tQCMjX8y3I/zxCSyk8FAd1rqmdVWbyGV/M6Og+2tdFZpd8
BU+nXiATAWTG6hMxFIiky1CGmoD34ypLKsEE0zA6gA2H5CCGNNA3W4VsT7hSndzKJ535Vvn+N0CK
JLeLCt6zyU5mExS5qR41hXak3eU54QN1Wzhbu3aDuV8cM/C7ckeBmtbBXTHy4P2eMjDv6K/LM5ce
4NFTVil/wUKZo7jUzWnWHYHnHCFm87P2qVVl7HxQ2568xEwa3mqoH7rrYGki0PjgW4BwtfmCQWnZ
Rj5kRV9REEB/QQVz5aWK7MLsG3LrgFEE/TwiWHQfrbnjBAYNBdaTZe5cW56hiiLRFgwaQY8Ftqwx
VepZ8FZEQsjJNCWUstELmJ/9l75687k66zdyib/jwaYKex3wytqCdJJU06mA5CTb1hClD+0qMkHd
JopdqwUB8FEFd6BeMCoQkMlkQVfQNWSeFF5cC5CaMt0NrrjaSqn0Zy5PkOaPSSqdhZzvDO0s0O2L
mLE2+SlaMcNVebKkUrFHRKb4nGx2JDsADlMtZVctoMqazdOecqMzKdKf1e+mSfrST8XSOZL/qKSP
53Jw9xMnSxVEn7MxpJ9qe2M2+KsQ1OrKEBMrsiEIrmM1fFQ8zQvmRk+qWa/7JGqc++SiHw0EwohY
1tBDsLE2yVphafMLuMUAU7vEozGt9UaLFc8kh/PN7/3751yoKetvpHDNg4R554cKJ9BRoesokGhF
El/z0vRm9H7WJBt7Tff3cswpMbXqlzej0Q4QZpRdxgJnt1ZRItaYoe9Wfk/BAAcQ4v5yjE5dktNp
RBTFlh+h9EYIOpzf7/fDxB4VpAnBLf4Py01BNxaQGEMjiNC0yqFCQTFjdLR10a6d6Z7irvIHm5Af
ID71gx6gix4EkNu5sr8IHeMoJwKYq5Q7Yt3sq5dp1qnc9zEPtyu7Dt5zEJ4mDzgSbatbi+iT3kQx
vgqM0YARKtDKbzWik9w05RKTTLC91Nz487m81OQjGoJId99yP60s5Hun+Brck+Nep64lEDcHIl1J
Wq5bBX+pDaHoXbar7Q5g0gbQqp6Y6Ir+YuX3eCdM4DThCDTj3z6YVht9TypxJmj//NxnW1sl5rLi
GmneM60/wr+BOtT5oKBUaywaXqKhpCxX65VbIs8XMtyFljk3Q1pvdaHLW9FKrvTR54zyZUiZ46CY
Hy4ygKvvUVjQAqSHfBR2C6lOg2kANzuSOCDn9v63seByEEW818W9YNdHdY/QG4VO79SA78c3YJJl
loUZ6KmDKf+jsab/SirQ/PwSW3Ti3rXOIKSjz8IGJ8fuKEM977PCYW04oVZvoSjDgGLTU+21IK82
05mFTvXiqRmO8fW4ktzo6iz4MM8gGxBdc2q4cy0sjyB6GLvzo7pekU5mJywdJFrFSihp1QphgRJM
PXLCZ7U7AW8TrMSzgSJLPJ4XTRFhH4afl2vBrVFFFlyqL+Z/gptch4Odr/X9wO1/9wSSVZ5acfqQ
DQ3E2dmu70N2/tu2hsBcR284vuagfRsARHO5pp2fDfCVDgGjJM7mjzSuZeqtMiFHcVx8IwBIbMVQ
OVS5HGoe5f5+nH2Tfl+AEGXJsjXd/ujwJgju+niMiOib4pVJDDe0f6FbtpudK5yFEnilRiYgOCJt
Bfe/D2nBDwHKEvY3h4zcT/looX3nGuwjUf7kkvmktPbjCEHTOFGQsrY64aDbuJoeiHYte7pi9VxI
d8PFNiqHksPFaZcXMk/nxaTKnpAdhVkO4xgkM+sHOaOIxE4gPvANk4uXhgdlkHNYT5Nr1CNbQ+uv
4JZlBmhZkmeM+h0cdoNVKe2CFRUtgSuz+PmW/uYTO35rxJvWrBOELY6Ynmv71wr40aVOoKlFfUax
4QcO3778NqpCKL2I/0V9CvWWCDD8V50XTRgAwHzx/sJUHn/cm13OjQ1bzMxir9/B375cJS8iI7l0
Y6phBUYf1vULd0DUvlKwiKLcMU13cgcNmjR/ZpA8pWqIa6iGVW2n08ycOad9IJPGLtKXj7rmg1Fn
tGeycN6Kf4h9zb5yaqoZLodl/5IWkZ5iPgb21rxrwcSR2DHrSIPtPOAj2g1iMncTbuZCQq+Cc1q3
/HX/UpbLbTUV/Ug52i5JB8EXF3SWn/9jHW+KlrVnpizS+7m96eDLntg/coCf4R6Yuw1fbg/B7Uod
ruas0rdycCJ4G33V8kGJB6J7mqnm/259FJHPPVVJrt1pIgV9RvHaAEaaqTfJULkZzGQQu9VUiYM9
wHQ1XMY11S2fASkuFTGROLOTHOmxmCvozAPtGV9WLIJnaTVuqcl6sSGrTZn67WC/0dF2enJP/S71
712T7R+aUZHuPu2NXNf7VvMSS/VSJ+SHMsN+2NJySv8MtjhkYFjjmEavtgGXZ76oFXDfUb9qV4Ec
DTUxkXDKdOQmvYQowMCSnwqXN/1JQ0TXxIu80ZG3410pLSlJcVbTV/9b6Mhaz1khp5TI1BA32nxo
djJkN6clzVDS/36+oTQYPiXzKcGtNXMtKAwo0rfSy9F9OrBhT2b+/T//M9gp9p3p1ioEB90LImql
7CDoYSj7Yugnm+ZVMUVynUSMCrvHhK2NXWokHWQ4RVpKA5be6vUxKj+VYoiGhmdwAGWb/YLSq6St
wcIBMvx5BscjJr2QixqeJ5gc9MPcqHE79y4vx3UjTw6oxS1v3hHs74fCM/S4kbV9isk9/QYvLjyX
2JQbpVZadkmc1lOUsSV90QmxbIKqWNiz0xm8STETmNJUWmEGXJ9nfMh6WU/WKxoNHFBvVBrh9b+S
O44RufhIdFK+CM6zrjGq+M5YzVliJsibq/jlXPsbuYOHkP0lAprzA8u86gBZahvFtOQl77sTXLAM
IZKDY0yvzxA8b/tXkxXf4XoIB6iwFwa9KxtvUIUX034Bx/aaM+P+tLfbWHpwh0BfnddmAVOczgod
HEZXhrnSESAvq8xCPcqJ7SiYvURvhc8bj/lhrh9psmRsF0geTliVg43qOkUM9OVW9NqV+5604NKl
Gd3DtTVPx7y0Lddh4Z1sBkSY/UCav7T0M434ph307rinqJWkCjq1LKyrujU7o3TTTRubQntw3CqD
Oj1sZ8IpRpPh0swhRKGNI8Q+sJfftUURCoXcmRK9hwWUIG4W+m+MdWiFVdOoBpqkNVZXU8j6wTFK
iLKBOQFYzfW49Az+scp7nAmuCqOA9bLzboJ/o4/sbz5nUoGGzQxm+Qr4mwmsA7pNlYdVQ+/34FUP
UldkKAyNDyLNpoWde4of8bAI0AfSCD1pLIQ6z+/YU+P78g2iwbZynqepcdHEzybtozmeE/yczoVU
8HQS794YuwIZr20mx4mI1oj28r9ttyrMIaciFsm9Z8kGvgbcfV5eAns/F1fK+jjsoOoGdBXooqaD
Mej5C/nrRGxwTg49zasMJwjdN26tX7dfS4I0zrnqW8p7ilM9VkgwWpo6HuBbOmuMn6xvIw0VNkV2
7b+vlXAhjeioF36zwT/7DKuDnK+OrWu5mu9Mf1e7YVc9fARu2EetmxcIROE8UyFkBsYYHEaznrrv
M2zzM7tvhAnTlFpc5D3xC4K55QaptDXvI6gCAkFuyzKWv92oIjvEbyKVdszSuxjbXbcbMU0gb23c
JceK+ishv0JIiNuSJjYP/ErBHYj04ugzz53zvnWXwwkAPqDs+nf2K7OFPJ2QEsXOEw/Lw/LlpKLF
p3/pYgD0yBxnTZao3wmrBwR3HiB/zl4DUqSdjQae+F+MiJmL16YjsplLtU20o9JuriwrLV41bZVM
fM5bkaNdYQp47+u54H4Ez3bi0IrPIh71ey/qDGeKbwUZJp3Devbyb2ELgNJthZfao5aJS4+BefnW
J+tjusehuIlqRsj2r6ohS2HCs7+2NhKgslvspmLx2cXnSHhHVPi5yg2LNiiP9f9bcgcTWyAt2FMK
iER5ntWY/1457lImCS3vxPy5NozPV/3ecoA3ur536nZaJNte7x//nVhV8VsAgiuNlP8CO1VKAvrd
p/lQ3awBPk4FECpCsK46Bne/kQeqwTwb63LkAewzL2/9Q1eq5V89Cp/G5iib/ru2h3lWxViZsFiV
rgkT9kS+ThfYkn0SkKnWsRDtJ0y5ErFDdiPteH3XG410LDTRhjgJOBP0F+izz0DPRWTPLoKKKQuU
PLNg5nzx+LBj0BLzMXRtxP/Tpfri3w/lnzyjeT0Aeo+awfieHthuLsDeX36WopLPgze8VLJhBWfr
rzK5FFMAJQWhDcsuHfJ8VIi+a68rbML+NLPGsRQzcYx9AEBUgFKg48VuA/Rbsmv7EpZHPSB4FF/X
Sg8GsaA1lBVTW/AyKv80fd+SAivxPFHT0aXq7NfIkU8+vvNTxFSOgWv3i8kIyLTS5ykXA0IY+7V/
TSmWXrY6zR7uXMQFJGumOp2f7oK1PKczzYmrFioc70gLbP28E+aGZE14CLuErLGspp4xGrjfho8D
kIX3xS0huLBLnvQHEajT2Y7QAqcQL7hlYGTS1C1Py2kp0lQfTKcBJWSJsgSkpXQiF0PCgEM+rReI
qFkPxbChVBbR9/tZ03rFKJtRP4GSgsD7ulD6e8O+51+qCwQB/YjPs2xLEJd9VauFMk9/SY7r1gBf
whB3w2MKtyBEq5s0PJb2CJBTu8SOI5jFTZ0IbAy8kErRoA8V1MS8RUGCrh3+dq1nlEslqkSA1PmS
Oay+5uOJ4tE+IH0KEy4aAcRkhg07ia9RxMEpXEiIeMfUTY1ef/MDuNBZry4LLNzOnUd4h+YykSrd
l7oh7OGWIhTKvOa9DB98y7YdiP+ddB89di6DeNLjFZvOYG2p0q42xLDyM3LLKiUOE/j7tzfPdrIq
pd2rmRpI0+epnQ1CA0eOsU2EnO+/9NPEwuQzUZoHVUhHuR3NvYeG4EspD6C5VbH2StliRUflW8kn
ldKvCaa866qRZDcETN0q3rMiQ+TT4ZsDw9ByXzxFVH+BnWkBP2gFIn4qlkG+zr1dHHe1LD2I5Pbd
dtjEGrU923ufpjuPmvcQ773QbafLdIROedXanQgVt8llw2EKN0gN6zjJT3sNG3VvzW29lVywxayz
aa/yIeQ+VheWzAFUXD/GtsG0BLPj6UyQZAgoV5+Yg45UB1GQGMWSQpM2ZHoIVAZk9ynGipjMPJsX
ZkoXmnwz4iwiUxGPDiwOkaeoRU2a9wc3JkZ5Az+NRHC1wf3wHD6czMpaxofxOcNkBgQLlojBorLR
/UOdDCp8mxBNoyCm4HaQYW1elbyeECWlwnVaqR6txTMbUz7qvVDl1cK+mkuAeS2hY1Y5TqQe1Ms+
QVa6cyrB6Nd+DkubFN4T08uSG4CoPrbGgvUyZp5ecY54Ws149QtatYFfS65JUv95u81vA59RqFsF
Lc+HxpTsIITEXbEfm8mf4e2nH6xX2THYKTevsJGFdb5zF7IHxuRzH6WqRDHslTN2ENORYWXy9P5Q
NaJfgXdB5qvoZl/lOpHAlY4wb6HefGvL4kg1sIe7DTWWZxnXIi5bFWJ1sQkFmuxh7p7R1sldsOUR
XjNONeGt59L2sq68XHGIdwSpDSUc7quhUAr/UAZsDQrrjEJGFmm65fgTibjoVdt82RsDl05i3Oto
h/PJS1mUDeMmjagJHHdDl1kRyefP3SECeQ+gxRKT3z39IzY8LLMcrRMeAj6wj63ZjHGRAu56QC8x
13Unjo8gHmBGOHYO5zSARXE9NMOXqpT0wfQadAn1lCPK9OK2+gBup3d/kADjzh3dzYS0ZFaeigSB
YCjdl9W6SNsg50NoHkhWVyqsmuLsm4Uk1+EOZJwo+RzvUlza/FTGM6O23HKTuDpO2MkrgGxx2nqT
Js1zZP4ikbGtAgIjMPAUpmY2EjpE1muIyXCJzYD66WEm8WgKfO6CUHowsnD9A0GECUenqaF4z4ZQ
neInR9GQUsTpLHEbKxX+pRK5G9AerrXLj76jUaos0LprPTPtpSSnJFOWJWHDIWdWx5H83ptFKRRm
8aoaCQ7L7yQYJIVfSv0jNnVJsHRzNw8O3oPbgH4yy+rJRESxU4eMylAL2hPayaywV1bkxhNFB5OP
3WuPVHA7LnzzMV5Ov7YZnlAn+uXO4bXFaRLJJx37blisp+Yqm5UzOY+IFQr2wwiTIOk0RoqC6u75
fQ72YUiuqVJHsMYMYPsgSBYhO57NCjHT2JOpM79zEg1p7i/HgTZkqwDEvoRNUPNWpt6sZ0CaJa4X
XqcRrjNtBBymr7kNLPbmXd07xp+j4W/wU8ueJ2DhvQekgqrLrh/cQkE6aYmkDbCHBEYFlHechx3Q
/cUR26Q3bjewPmxz8zNjXXKFg6zsQROrpP2gElgz70DE9z2vbr9P/6bi8OtI70nvIVXl6qM5iWCS
ySMj1ynBsBqZN2T59QcJevcZtEPOvPOfpLV5K6bmdK31Hj1eN591btynQNRm04yqttjgVevNS0pU
F+3CQBgynJuq/LDiYpZGY3Jly2HtvOvTqmf4srZVAjyj1qDSiF5rc9JklLyHL96EzhYPnYNaUKir
4RUZEvIHYbJ2wA1eJo74PD6XHmaeUfSWt8tF92LSsr0ZH5NuT6Oa9RczU5cJxATzmMcfbRihYG20
z/TQ/YDYse8g4j6wb8jjK26i7eUnI/4hnTMgNfTspQZcPOnh9hTKQHoSjhAwN+PWPVRpXEQ6vC9D
8gQ0OLpgUU9/arRBX8yz62sU6yj7FtNm7QD16fKqTLGwrowk7gHg6YxLdUiipPyq2Uh7N6/K5pt8
3wtDHHlXC2PIwArMgMJvNrGflHx9c0gCMOT3S4b92ncaQ1kS2DGUNjmfV6Dq2OXf1Q72cAG1qJgT
n0OuRTCmatUftO6SYJ0vJbeSc4GqrLAFdJdibuBV9V/wC7nQABbloJVJIsa3Oixp5+3Pc5ULI8f/
3UCCBLGW34EXa0XS2cgxZ4te2rSlN+TSLpiii7R/PBXJa9WJVim8rCM7DT00dhb/yQkd44+fuXKe
/mrUg96zs0GA+d7iInMgSVsllLC3OJyIPLErQ7HnhPZg4GdfOTqJOkyUMW5/tDe5p8GmWcEbfDxG
ALmfUX5inBySFdbxmqcMlivaVjZagDNoShkflF+m1Jn1zchGEiu1rU2g9SlWNB8+wDBBP7r8N04H
dHsoos+1XbOdvzY2bKr47Ec3asULKlZhJc73WsqpnrxeDgXuhDzKHwymLrDu4S3z/tmbZyw7dURH
QF4WfWUfAwC4kDXSSN8s5qkQpN0WbWebluETiL7qdpavNf2E9K5K2e3pSrOTKFuOKW4EZcggBteE
L9MsRhxJFKdPePWI/xtKsPYV12eUEAqGkcvNDuxpmkRGY0s1PR9ZVllKqpKQvTpj03583ePlTmtD
QE3camvzldmkWGykTmEVr4yH6A4g1YQ6sUcpyxpsuv1CkngyLLWqleDUl+RLsRirRJTie0ff5jVp
NnBrKxGzKsTq7OSADzYdA/EWjBgVAQxt7MFOrmbCYk7ePnWHraUXtStMLGonGENPbT0L0KBgO5zM
hLuMRhSj/T5HlxqQvltdn2hDMr8G2Sks0lasVsKe1XJ9DcYJI3KdOAvvX3x9l66Te3ACvZrf8SPo
vhPN50rHcayOH3KkgNz6aHy0HoHPr9FFDF2tZlIyIVooya5zyawqzFF/aldFkZexU+wmBIeFOJKr
MkYs2qjELhnggCndeYUMJ2O0RlmldJ8UEOAdPIPX7zlDCvhhUi3ISWu4O5JfReGf4NVMrix+oV4Q
bRgNMFVF07w47751XzmuFf+KEUl4WlUI8VN2cLwVikT1pcy72Hm03Wj/vUu6FaFTKTWUvN+HOwCZ
E38wfanI9eIsBHIZYDUCj85CYOQG48R5naWhuymvKMmgmLe6O1lFT7HGNDsG/xb3hO2rGTGXe2Bo
16j8rpxbXXa9uc3YyIvTF6bMa5slViuYixnnrTrcFyEK4/oB31XJuCJB6gBS2xeMjEwU9po2fajm
Y1Q/syNA3JgvYNXLjr6ahNF5coLigzPSR9b6rL3/XH+7TDm3Wgaf9WzBJllB8jk3yNTMkjAjWvsP
jNeJMJ9aEVN3CuHZJ8TNU1kRGAyHyEIjL8C316cGEl9DkGv3SEConVJNDW4I2RRuHVHz4t7mPuwG
Ts1M7Lt+1MdIQAmdUUwiISDgbzT/U+YbpVC7DblSP1J/BdCCcl8JDQ+wGGCIpMYtVtMp6emb8e2u
lQpJ4xzDT3dhAKOXbRVPwCA6ZOpn+hFo00oScSbL/xs8nmrdrjsFLYLcE3vuvMyQXxpgnpMa7pK1
P762zUCia3kSgBLrpbJ5uoIxjeczmh32axp3h+esSYpJ2hIgarh4V1vbd+XgohSllrYRdTi5up3g
msYYDy2isxuIPE6/lJez/miXq+3ikprkXESQ8Wq61NHkgoZhpzjZMC/BHYPEEj4MZ7ofRYu+U3cL
GNQcz8CDwNzspGgn37SehhgfE48XVXzxKvlnBtaaymWaH9pofajo+YeF8l5/Yjot2k+bILekfvAC
OcpVMn/mPuBYe/x5XFpxHe1I9ei41i7DJ2J14K0q7S/teZPS677BygbreQqeIRlbxos4XCODl2kc
sq2akk3+pNwWI6HZxcevjsbZQgwbkeNRaa6GgNlcyGsKYKbQzkVNH19MikhIVkX9alwkPsXRlqEU
WqLWKbV++9fMYFotuCspwTWuuqMMFLozRV+eyIGjFpCJxbtJ5tA8aHJHs4X3mkPGeWO9Fjsvgtiv
+f4Tyv/XOwyglkZOkiMMiKUmidsvWK0RjLHKU0RgCMeo7az+ujmNwdEaEQbVTs0hBiaPWas76L4K
Ur7xQorzcxDfoFeXqtngKuBjsACtSHNHAwszOt0LedLHro6BhTrLqpEsAICknJZh6/QKtxU8XMBo
oAgG2SEcVIPtwJz/ZqqC74xoIiCdhr9KmYIN5SJvoIgRJn2df7Ze91TgFOI0v5oaTHYATU8z2Lmv
plrD7RRRBod94y3qzFJO03D6r2tDZmGFANylr8bYfxYtf8kN3ikSdLO68IzzA2TTDiy07e2S0MUq
a/mox4aWtv4D0HV7YJGpsGWUf4Ya+sVlNv9PAXx6adZcsNA9Du3Ig5IswEgfjXArbDdkcKFRWnhg
7cZVaNfquWRYeoMO6uQptl1RTaP3AvDB18HJaLeJHYmcoZZDZno038Y2lVpRutGFatsiQrymEiT0
TuJ5kLrtQLpNCz19ct44c/D0bRF4lMg5NP38XHi5BX0nZz9jn36LTYWaYGvqtXNmHzlx+98gwc93
0safQns3B+2xpnQp5JCzypdjYLzqVdijSzUdmBvMrq0Fdaalq8NHadCU2ndInC8d8rzGgSFRDWtY
ZoHID8WASgxFpI+wWkeKR2xw/1ZRQDKcHgpIQqV3otOyUeoe5YxyGnnSrnUHmh04XJ8oAGCjrOtJ
WsP0TuPTkcBmz8DHMsGC0o41EdR+9Qu7bZW2RLXqGZcvoiM2o86UDe9zmlTOgCiKFXW5Lv8BypJ4
TcMddzLLJ0G7djo48lSAF04riVZSyd1YyyKgJ6NusZdyidXbO3CMXOO2bjfc/1iHTBR+TivcBJK2
FeqyVvWQx2A9Z99LuoHfqGVmijFhX0y4TaN2lXIAv3Xqzfiklh+TROOsJAw5IukBxVoZ0315z07/
L8AIFDjDJ9pvyWaKsk6DFRZSKJ5TJJRzE1ImjC5daV1kf0xqwEd7S5f1E17eP3iBis/2DniCVUmR
v3me3860TIXox7nVbycqSbvtwXCNNJXP0acWCO2mjThhElPn3OFXj67+EOH5M1YR4hL7srsdUgjq
s1SUL1IRzDAyG4kHwD4Mg06g+mZIvEqYBMFYjnqjY8J4Dx8ZA/zDZR0+RY8gPMfXN6zN+NWn8ow+
jNe0FWPSGawZYvMzcnZUt/h20UttPNuXjwiFR+xMV+Ai0W3uvjMDVaafYQnvnJcgfNNHOqkpzjGC
SMEdXGj2o9LbDx/JoOeFgYJI/XW6M9lcw4uJxlTHTqcGxzzY97ulExK14aO6Cil6AeaSov0Zc+s5
U6GtSGo8QZZmFB/p4ldBj6wtF+iIcgGKHRLLs33Ilo56WGBxYan5aLiQ1iAWYOiNFHUDNOkxPiGi
3YX4xtf71dlN+z9gPk/XOe5a1QISS9n9KQ6Ary6vu//QoHZsDdHyVtn7rdA6IRw09q0HygC/Crvl
lqasJvlMVyLAIisTbSLhIjKEQV3HHfV3XovCuWMPazGj+DOPRYEFGg/9bSVlcQP1TJ4jiNogjSHj
Pb3Sl3iXEetSaymrrZHZWFipqSZabEFh2+lcIrC4nd0xtbM/6ftNpUHyearZmKJNpow2ffm72Wdq
v4aEencaXrvIcskqqRfNwqZxuAT/T3f4TJ5NwoNNikgjQwka3P+fbs7KIZb3PQKguoYX+wK8DAo6
WfHIbaJJwt9t1juwtELaUVAnGM7pLCaxZbjJGQ+VSRSn4B0Qg4+1i2gNnYcnM83dneXE/fdLt2mb
tF+8p+rLFc0eqGmdf08eO/H7jsEjwJ5HLb55eGGfO2tz5CjjehQ9JtUnzppETxkykIlOhsmVaphy
RG318rbEDFdHb2VYnWt8ZUIyywicV19688qKSoHl9yc6E903AANg5Ptv44FIm3TGhdgqGRvizg9y
4L6XiKsOmi2uNHqmndFL2D/N2L8pZ3ThVb4H09/UayMQVgeY33AnPi5Zi0Jxwmvww12pYBkwL54e
Z96OsboFTbst9+Z+th389S+zt4Sdy+Q6EwCyca8HiZOmShNY3AHzd0zN51aMtqJ0CjCaZ+os1Mk8
gkVBDgpy8qBmWzoVPONb+KvC5UQb+YoQxahOfBHEA4vvKQkVKy0+skHOVKuHKtyQP5SOziD76nMj
RzSAvOwTFu9m4+xIZbLqYOG9awNGUQeeWIdEr/DE49MAdwUyY76KVgRu1izJz8DutgYnAR8L0BUE
vUUDFbZqNjue8+tVyYqMWxF+NdAVW/bg/xRkGdoqw3lqfTSz9CQ29FTO0nKKrFMeoOTzv0kpB3NE
q9odKedF0sJp1mSrHxuTzJwIJ5MjWbaQu4Ttf99BcJjPolvIoDwF1sA+JDTD+eChCGYtyUkGZF5Q
cSe5o0xvBbY+HfcqswN+cz5DzMkhf73d+9c+mpbLXRuVOPF3bp8G+p971u+SkwVguCcTX3wrWE4j
F6jYxT7vGRiBYdU/+Aa8R4n/mfkKdMUhpRGM4ihsbOJioWUK7c1xaON4TaKmjmhnMDWr2eYn2xo7
6qAQNEKog4UqJgv9nBsaEnBF7mWVB3aM0ZQoSs2Vn6PJYK7i1DGk018fv+WII9UQa+6WW/5MDwsU
usFgelAAoxP8s6PWTzhsiKrbwFiUOs0jxIARwcG0/IIL6X38NY8LlQ8x7RdkQprFBlqDzZi5nUBk
0IEDdfriw2gOP6aTj+c8vCSJrg37MSBFlKt2j4Wt76SR3877ctOh35ctqfbGYUs0A6BE92ndb5h7
rouTZh8z7KAleI/uoGAONGS04dGofRfvhznLCcQ/zvNGbLyo3K3DGJEEzmmtTfEYU/Se5TZiCCvW
VHxRxAA8sZ7Of739welU5quXLqvSeOZ56BnMDW8plR4I5+7z3psQ6In4sqX9XXi6+/WuBNogDY+o
RGNKVXe+jtLGRgHgwm9IrxUN0/KwWnZuMm3zFB7iJAjijPbHxKqPCP5ivLqv/88iLYfYUelBPFBr
T1qwKsMlE3m/+MiK9BTXSW7T5LMWfnV+Cg9yltBZefrhNtpRL367npKtGb9CM4YISDQ7iOWh/aZy
6nTzPibMRthQ/umctqNklxUOPpo34IVyfOFj52isXWj8ZzwjHLg40mWGpqH+7VzSosVLPRRpMpXv
vP9FbISdqJeEENOPJm41Oa4mRfQez7WaVj3EYq2axM72nE6vBXsoCpabiQmzDT0zHlMPzFrINJIL
wQVN9Ddsu7MEIdq1DLsWoQV/SKu7+Z1An+oR6g8al7fZ906GbnuKejp6Pt2l3CiwnA9D9YLtjtPV
AjapTmY56BntEUTk+bv+OZu96T4+v9Y2EBhPWf8n+M9wvNU/vRsfziTLxqDE/LlV2t+BhSblKLCU
HgjQ6bfZ2CazZTaTLeIan65CYzl4ViXYMjqJ+yBdjNQbf3FSk5jOKhgDx4c81SGb9kjUxik5rkAB
0kTp3o4nDbx73V+VVT/00lYhoVbsci++PfTy8Af55nxx1T7B+svblq5ZrY1c77Kv/qBtMxkiz/MI
G6NQ7XFc61oPjyQt39FKSQQhnWSW6rrKPy8IJ8hT6Ue70BKaJ4vB2xY63nOF5G19mmWaCqgga9qi
TOSGHFLjcXKzhlL8hy6sD94knwx+QU0m6VARA8iiLwJAdPs/32a7M017Hulevro0ROVG86HWuyZE
g6ZhRxIomBOkW2/Isdfb6D3bb1QJWB5SXfLzEF9DFfwi5QSaPDERp95c3ETCVMlstRWiAqEhplTV
HH/vg7ykrG7Ho0FaABgB8LyBTeAI3OHvgx/vJbIMtbk4jOpzCWHAWh/wHpczG+BdDFS2/G8nCQP1
CdlX5bJSXcipSWF20uRljFrvvcfrVpoRpuQvpo7uvoOExVVY2qjlBVBuYplz6g52jbzWEclDvSiN
uFSbwl11yM9DoBE8ACaJrTYu48aypZYGZmcMNwin534pJ58+wSZKuRO+e7KfWidWM2b7SYLm4xwZ
0XMoFoZACjlRt+DtPVtZw/CIkCs79Mgk7qTAHoc5upoee3zzkZvXkYgHhg6d2EPmztDJvW9qTWK9
ELDz5ffMVj1NwHm5wV4CFMmESXA4LY4FAnHr+hjPt8hnkx3V8/ir7CczcO2UESqY7ZfWEc5QbE4O
+0X0US8G3DkyA/FTRbM/PteyzAqgrJWfhA+t2Scb0Yb7QTDzfevQo7rZsJG8F/jo2+LOT8DRf48K
y+0PA+AfJYQVmvEY7YVf1I4LFOBx4ISp0Wm9d1BsiSgYrC6/0rRQxuxozEdTyAQZ6F+ID11OYtJT
yDnBTYFyC1N5DuQuPEktFvQz7pEAgCYHU6nSxpDA6M+ddcwNsZXhpy9ghrQtW5P0IQyA25Klo5B/
fWw0EExRDjO3FFI4Fh5T4rqmqgtzQcl55ej0Um5JgCcJO9oxuvRYPVm+MZy+Ts4uBde4nythdsFe
JproWJhssXagffvE+yLd6aYi6VjZp0IPsXz/JcHbAyIKzEw9pY3DVN2OVQEQpsmbNNJLErSYtv3c
NuriskK1b3dXqYW/EnzYEn4jBz9QeQb8EKJ/075F/9X27/KT6mw9wvyu4XkpoWrKSQ4396Vs2gWE
X72p18kV3yXqljMfRdFgnR8aWNC+Bcybk81IBFiK+HiqRWsSKddjVH2XNlQmj0jkQdtCpiJrZTg7
AAQCdBJbTpDglLcD65+UPB0dF03sEdUXzHzFvW1VJhDJJLQLjAAN6tEgVdpAYvLm7LfwN8Z3jXUl
ds4GBzDrcMFAwGCEn84R1s7SWXHhLRvSIWRq35RLk2HOEjCp3w3yougO1Df5GCJOu633DgRp0Syg
j0E7ys6AeRovAOpdMEJMw07tu/AJjQoBJPM9tRuowsubnHKM9UpCjxUfci+9NG0M5FAbHOUn5cXN
ewubdqyA5cefeZ/+8KaFTCXTDD1On567Vx/djyjbzMeBhdg6HSatZkyS2f2m0s0eRo/ZKwALEYhW
/Sxi/E8xSuTvVjYqL6S6RfhD6swQ3nuZeouJsY1Y3rqFzkR9FpWbm/014irK6s8SmdigVvrmanRL
I4a7mqi1fSmxa5E1lgJHE7fqyzxHZZ5Cpz2UYfVK0j3hE44VkmzEil+SPcQNyWhGJnrQTJN26U1q
2xx348bo0TruRYyakpiUIfw2jqEoxCUBw5yt1wLpSovgkpU5ah2V6E62tZgcHoSreptpueTNLPWU
fosLRmqE4HnHRN157bjHByQUqh3kB2UVYL63GRDTnVaR8ciVaANDe1mGEWnu5d8xZffqitfRYWaY
QfMPMRRYuxDE2vV/eNu1e++7LiuNYhRLaw3l5diM/V/s8he3S6XhrPYfx29QR+Xe4j4zeayv0ajU
poniB0+o1aoJfcW83aQefVdnl5Hi7cq+qBopfHudK71XMwpuu+rGReiGOFbc1U4Ou1NGwLQMMFzV
8HEvL68Pa3BM+l99d72AJnWU0bUX0WokGKu4wtXFm7plBzlaKz7pIQ1ldJsfS5KjXAjQz3Ar6Lc3
84ghAqAxgRsECTZSSNV42mlZ6ISvYudt9vsfdDp572mpsXMTfT0igYG21c+hnyZgaGish8irf3tu
L8LwBCJFtPs3aVljDzTlsuwSztRNu0/lnlWSaSHhcj1qw4YAsNWcFAHSnD8aP+k9Sej5EZKJwYBI
1ul4n++4k0lewyEj0Ig56+pkLaCyL4+AdHsfBGLwFWihqPL2Ngj8sWP4L/wbgmWiwjwCNXD8CQLg
/L6aLcMmaTrkGJ1ncieh92fg0txFMUa/U8kkHR1A51JC3ubGhSb30mgF/Ldlb9YWxVCvSc2jq0MW
HPPFSFUBFcWHGA4R3Pxd3TbMDOSIvgTwSXjx+EcF7pIsV4ogOCsGHFVf9qK9eqSOxFJmp69RELkR
85BV3d4SK6lksrFgPoD0FSiyxpVdppvMSMODUjWvY6YKZt9s+qRRv4AfshvOBrunh5xHykbgQDQU
ceg3mU1ohps4sPmmFjmmSXx2nbrYK+vjiXmIebtqCPMgslOj1OjmAP1bQ2j3BxslDWi8qmFU6tSM
hxQvjy2tuiKUBqYXU4nFDbEF4OJY7nN5zy0KFu80Z+F3vlmRMfNPClNBSXe8y6HNvRXafi46bPdo
2qaL5tZ50rs4OEipn2hCtR8LuOStGYbYD/o4dGqsgICzlCA26M83NpOnibelF8tclA7uO4/1RRK7
W4vrdcOhFfyTln5M8aiZOA5CGQkY7RerLSg7z+1w3K56lTOlc4YerLxFjRSONfHlrPGCXvmrpBRI
CzpeWtP/2MBSGD7SS2QBd4gqyTMPOYjq7bhtJiEEFKBuiJowOcCb7ZqRlDQTlB9JQaQFeWj3T/mO
Twma8z5XDTGeEBss8RV4nVysrp6irXcJuUlw3wTekhM0WZ1KN6WB+ASEC287y2MPEg1v4J7j2bSH
15TROTK3wnrqcMp8x3ywd/McyHih1fA2iLsuj9jLomwIutHaDWpsFj8L5vSdUpArpJREYv+oK/E6
XLcCGE1nHXSwENPpNd4a3U0ITBRh9CVgxr3HWAwePqVn6pWP3j9tuIaGL0njcGyn0ZSXk0wiWHD1
3fae8z6WAfh9UwbA77rgn6EVDv8E9IUIofiNa9fx3ni6NtXIuU67q9+CpSQcr8n2QO7B9Iopj0go
Wc5yR2f6fZJ3/T4DBFLB6nHWrkMbj+XSDh0DDXIKdoPAtBuMJAMYrr3jqJVXrothV9c/NB9YAL0I
2oWwMP+TiMh0V+UoP5XN06/bNH9V0M6XGyIJlCOwgZ8QqK9SOy502kb91VSx2/PQUDhweOfQiTYZ
YAO4m+H6YiObopxEFcUpDlGoffLISKaTaflsdF97/5iCGFRqK8QTGWaQnRLdxG+SlHOo+0YEtJJ2
+JPYEjVPbWmKRyNQ0EW3lZMGqhLnNWu/aNRjr0ZVFoDLn402QzCGFeMQQhtf0Kyicjm+w5V1xiwn
dqUPs6iuHIyQX4WBlSTkcS3B+KKb91j/+VI6DydBpdkK8mpQ/uFMZUPbn1pUz2/Eph327bd2Cf5O
8Mj3QrYjGmQu+uVSKsQzZB9P/wa80Tuyf89jmss90MZ5qoSawdY7mu0OcF+Mo30tuCBq6FDTs1BH
FlFcyHrmV8JDsT9ETqGzhJGf/EKdG+nPfrElHP8idPoM4p7oQNWLpR0xL8uq0PNdkWv2B19XVb8i
4ChoFbg3onagjhQ7FVndP92m+GpteRL/QFGX46uwuaCzIWknhS4GHe4WABZkSR3rWlGlgfvNq03L
Hxs5jf+aEDufalfNnucptZ6pWcWLh/DoW1WMCSOpgWkP04LO87m8rE1aYztfN/9+nX0ZC1ars4vc
xXlCsaJdzv1Y/HGu76i+HDhZwx4x4PxErwo52kOwGn6W/XI0raZrBjRPJVfuxsvSsR+lOHKOLFIj
x51EihGHN8KA/Bet6wVNXfiJkdeeZ6gjvF5sJtZFhbj2Wy9hKyP3SKoC/aXCoZGx2r3SxQjhVfyT
u11pkR9S5Zik5pJ77KRDz5Ovo6+ALYuS4TwSVl//AaBiNWPIjp1+4GPTb3r2DjG9yetS3qggg2bk
iDju7sjXA+APk3XPonPv3t7ewgHRi11XOxnDqtqcSwfA3KWI5y723xZno5RbKjvIljDwjlf5Mmlk
ZY0J5b5+mvtw2tdiM4XO4OZZ5akOoADMctrL+eGAR6/ILwKh/x5vP0vvYoCLzcjJr4fLWSmGCZn5
HbfjzsmsCbsBTTbU3GEon7QK02ckEI15Yi0sEiR0JY97/W48tP+f3QD/YjiRuOKzi2g5VoJsuQqg
4bSoxBYC2RSWEuuLZcqy/iK3Y7qDJvwc8tfNCcJP+lYxuv99upBe/UfglB6Si1BNH4c5zfyugxDI
rNdUWKoxfc1G21Rl1ZtNnCnP3WLdbdZFwLi2yrRhJ5Z0aS4wnUMQhdQJfhKBgpdgs7ul7x/V4s5e
YRnmOBoLvVEfAO8Sj41ikGoNKTYC7jl1uN4HUQkuLrhNKzYW2VeBzdEszlgRtwSliAh3ExQdLGat
TgOMKJ+5z1MO1W0Hfi7ULhb0TyVw+82wynoGmueQq8bPYh4qWQvKDCYX2IXyyUDHFx5knPCF7FE2
s3YFtgcqYuHzT9HKjmJlc1QT4ZAjEvehUOrbv3Pyo+6Lc+h83bAJhULvWX7/v2nsOTZqmtoq6Nbn
8uPvSuTbtYMBxedoxqrQF7R8Wi/me5uRLOveDHg/dHelDWz4iOOtdCrv1tLFaUc3fXLrPrpt9jtn
besoxNd5LIlZHlrHFK+LXrfFlqQuFr4j2TUx2p+cqiytFl4BP6O3JhFLzArb8qSL53f13asXizZz
OKwZnISH0HGgCPTBZTuk0Bbqu1EiVt+2JBBgX3n6RYgAx9E36gamUFfeUoeIC+L0+MjCbcmF2YVU
QiaRaZ3fQ+8nk4zXF2pVU6yeby0AFE31m26j3QvsyVyiasu7xwp6pQarTXUImHyOHKN1GWaMT/qc
bg3Kg/PEY4RPz90GCuGNH8cKEME62itz2phyXth0qZ6bHjcR7biYNNXogsaDrxNc2SB+vWFPebWG
tIj1CRxJr7Z+/bBxyHopQVHKE+f3+1cxMgGRSJb0VwFpqMQg1j6jX7pc1eWe8/6C275n3HbTYubs
bwmPdrH/vsh0jQAYP/wKooNjj8GRHXP+eNHRNJ7Qph25G/Vh+mTKE6W6Waqr9CKCGCtD7mSp8CVo
hnL1fHV/UxksloYKP+98Z22Ly6JWA6Ueb29860y9jBxfVKcIoOdCIdvdL+wZAiYWXfhZEw3lvaQJ
ywq/fkOzx/sMTiZGOmXbuA93f4UfYi65qD3Y6jlP+xJje8Q06Em7FBYqIrcJBdC5lWiEeolznjWy
cSwhe2Rwf7PWpHYNEiOtjuQVMU0zV6mAy9/jUN23YurgB0G4nC12uOFDKeMRYP7mnhOcWRQqXcSC
nhBI197JQ75EQdGgBhYsBuRDk6n1UgOQjXCen6n3GuZzyaGoBuoxLjAWLeNiNykt3eJWbyUc3jJK
+/WzHEpomXu+It5oOgy+anCM/X+DW8HnEzdqFocRb+GLh+Arx5brn4Em0Me1p6OuC8d2IrSSMqdz
sQSDVwjogcfJ+W+ollvtLo4zpNZwVs7bR93OT3p8QLUiBQX0CxB1rwytcXrlaOEAF7Uf0Vab1xzV
S5hdCVBZDQLLoB3YPfbK24KHiJf7xa+JQa0aUKedV0A+sxVgGnFFSRTLcRE8YHB3riooPzCZzkhZ
x84Isyk6BYgPwFC7+uz1YCU9B76LFd5HcM7X8iq4Ja6w2pMMOWtz94SHfAnkm5ugMeHpwxybGzQv
Myu/SMNa2N+SuZzyUv8vz3Toqm5wBMH5Az9/KbkmzYjlJ4Dj8qb1La1n8wRWaER+RMR8R35b2Jlf
RopAu/PN+T0K7cHoOFnUSE9GB/96PGJWQOgO4oCDBXWl0P5YCHAaOXwPpOjWoyjNShuTd6PffMIw
WJYB9EL10kap3wgWp5N7ObjJwy98C4z1Bo/+LykNn6y5lOiKlj/U9KPGVQu+GGLxMrIGb8G/HYTg
fEkTo5F6NYUnAPIKcXvYR5qdeREUT4Hq3OxB9lNDl6oYvze0nqVTRSMKxRHnM0FNXKPIcMU+o/xa
nMv6cmK36sqWYtwUZeBIb9E5HysGWN8UORPgStmeNoSwbZuxzSCm8ymEvvlZ6m8JTcvV52kjvNZq
TWmpVY9u9HbwPfap3XmW8ufMFzTTrp3b2dv9TZfdf0Kg6A79QdDaAyqEPhSpLIQIkYKfGr2wYzoc
5t7h2TwdpgJW20I2SjCx0sTlxBQ4Sc55q64VNCSk/NDiCd2c3Uxu+Mwgq+IpfgFEo/Zu+0QRpe6T
WJibJyEMiHGsbZpAU/O660/TE1PWOODHyqI8a+GhMajl/bcw/43FsHgKHa6rju+pjA9PUhPsWiA5
FlFyZZLtDsP+O15V5BrljyhwhyV9n75ezgX/1NqwXazMx4kHekQsoGTYvB6Jtk+xI8ovcamZ8oUv
2k72PXGAa6qrXwx85dpGpGcBoJjxvp8oRavu1T0e9ayd5o2vETSu2qrWQCgfv1Vn/wKSGH58/K0s
MdtSf3gGCB2UgtI4XUUZB1D3c02GYcJ5GJWOOVsp/AySt6vfAHEF9iFI6J8ECbZ4e39qtDN7Z/q/
UVKNuGkELlSqlx+EPuABRQYMGrjcAqTFq3TND/bxd2WlJyx+w98XGUaQm7kNCX2eIPRbA9g/gLdE
Jg9GRKrK9azNLlr88Y2JUun9kdt8sR61o6krI1YgYoesN3xK0KUq8U8/G0hxK+GwC+I/+ugSuImM
gFIBfMH6VOuQ0xMwdY5jLgcH0UfleGAdHSC9G/4PMHYc1dVIJMGuPp/IW9NaXUKCB8AAETmnDC9z
X+1XIdU7UOTZhVHSkMJlTqyiJTTWo78QSDKGNNz4uIw6O45f1q80cxO20miBqnJ0gkBYdJYjyawZ
CkYy8sbR6s/qkzGMla78pfHeTaaCcOZni/mzUYQLaX6Xuy5KUQAAcPF26QO6BhFHHr1GDY7QXZ/8
Ouf+CFACuf50NcOGZYl/5fIZpbpBq5An3FFOtpI0BlMHtM2P37Y3ZrrwB+tFkwMmna6AG9iOf23a
0wKrgsTUBXfd0wWTkCNvOxxAtEPaYZcBq7wiNSNgzkuMIdkIMsEaAUCp0guhpXnmQs6drf5tK6Wo
JRryXdVk1iclSZ4Qxkm7QPIko023F1xCjj3qYhPl/AC6dwxqGxsJhK6RD5dJx4c+88BCo6fMwLRJ
aTTRBV/5CzrjXW/TmKACtb1DrwhWmozmWC/Q8Wns6zWXTxwudnp0bIgHWWJcACBso3hwhrnmasWa
x2YBeIme3DQ3iFW8zdtErFzSh0MXyFnFg6R+liTnYatG7J08dUCjcY+84Nk8nMbkBlJMuKhLA93U
aHoemBC4ypgtMnlS5EFktzPvqRh0Ux9SxjgSa3i/HdQDCrmYfIBkHeOa8AhaLAqyLCh3lNEKZtDI
6x6Dp97Kv3MFgUsNQJMOuXfVbZwneAoHq3SZ9Dk4sdXE18yr3fJtYGT4sKUr9eMMvCJYR9P0OGIj
dEq7OlN5MGbYMk55wT+lDdRFAhf0HeFolUWLhFtz7KVCVliwcVisK9/nZxDMR2K2Xa78zWDdrTfH
MMMAS0O/an0qeJuNLYDSYztT8lADrdTNOBp5m5U9ni3Rl7oCSwtrtMHzjWlX33oR3rBzhOPP5TlL
QZGu/A/XigfZVUu8JsU8CdOhDQ8sr7dl35dcJp+i2a9itE0XMXVbwGCrVH2Jp3T5x8B16Ubh94Qy
Z+DGIQ8iABZD1fiF4Cboya2A99dltWDkBHp8MuOdN1xku2Y+WbL/w4aizSNKyJ3luXfjiM2JrW2Z
t1F6Ur7batq9fqKjr0qPYb2hbxpkbZATX52/gJ6zMirpb1A1vaD4zygZltCTBecghcIKEsK33ia8
GKMUuO8D8pOA1ug9PUKo/WAopzzC5hbjIBKBg3q3sh1R9Dtc7At75mA8bTeu/+F95ghnHkS/ES8Q
EhYJzrOuUKladJNaboAPjj7eF0CO/2RIgnU2ZRNnKTRSfPL0GR5mqz+f5/5PEiVmiEVxE44b0xMF
Ej1P+NfAFigPnDwIMX6OAS9yYnujIZX5cnBhha+deSSkc3/D2KJ+Nz7dL5lJT/i6lHrOX/PxADW8
e00dVh3dJX8deuwwm+wd+D9pgU5YNgSBJ6PkvqK/djRHtgArJPydYsc1DxN9NaU8zDymVuxTcYcm
E5AjDwmYE5e8uTZeFrAuUjwMkrPzvlJU+lUbKU++a+kOVHrSdPSdi2DMhTulnJG3cZgwgmAOLC5z
rBg7S5C4XuDZ4gwbp69g9XBRiMPX4ZB5J6qA2QPIrZ+a73SITo94o2c5mQ3hUJ4cc6fZ+6gb6If2
VAAyZwWe/+bePpRUjgR6zpwXFve3A6GRMqv0z7x1IwkPyf65QXmcz5OBLpArRExyTu7BYF6vaHlI
iqo1SfD0M+zo22195LqxNJClht6ZWLEeTyertjxt525u1HisbfhwcMzC2c6t11+oySwGHrCOb1kW
bhZSA/Zuv6W23YCJ8KP3pYSFQyKnIQZQWEiJJLvHWl4YMcVCilk20lsLOwP6PFBBK3JzVSQN/h9Y
jRj6HnI36dj1S2g8f8RuQduvqTNWG9mZWTrpizzN5xF4wC91frAkOZPs4CJ/4YDnBUJJ0zrHOpvX
6PEIS73gF+4fqz899qSHksZIZrfDDd7bNOvx3ZFtlH49ScEPhI3BgdMBxLw1PTbiYEZf+/K9s95l
uixqKzZOMtVFWLM/liT9xsYEx7m3SMCoRy52nDnjPcSwMaSUuFW5SPlbmBzhtzzSqJtMB5livgJh
QTWAAuIqH0Lc0MYKHSKdSUUUyRP8nQGpuOLI5DU1u0GCGrPg9KNhzJ9TD0tESFLql799ZX95IHK0
rX5aNkpcXUNBcBKFZKdAV+DVVOUp9kel1Ib9d7BpJSzfdGwjHu/plDfO6FEmSHBzDyBP9X6wfT/B
GikpKCpKS74mh2E+ZqAlK5APuogL9hMgkixSaKNpAeUo22vdV6hizIl5FuckMxOnhYvlzZUujcGp
WuJY8sd1m7BhYYBLTma3OpkhAb4HxxFWX2hO1u8qzynAGE2BPmP0BASk1ecsWDrEwOeaUqxVXtcs
a3Om9KQsJVeqrcevWkGfxaXPXJxGUPGkFo5HG6mMLfNV8Is8qh7AxoGMlbZ9RE2cNQx2eHThEoNU
AviGdNGLte8RR82B00beEyU4Tlo/+a0RsndnNvOxq7bco75v3uacUviyu5wtoT37B/tBJaDKNH7D
aXi+rBG3MIPh2zpL9YVBd+yiVLCoUZ8BomL+69xotHFfiX+Jc/rapAyvfJ4UPX/RVq+0dgHzGREe
IlJn3U0TUr5fgd9qqaFxYdOZtSiYGQLCmULiBf59yY+weagcwxdRGUWQntEXgLXCIIbe5mlLhVor
7BoJnHxpjnh8PTe6m6dwqnqWvmLPLzYvWFBk89YaODxwCofT9WwFnPUJ6wp/KrviAwY1lsmoQoK7
MZjHaLszoizKhrIcjdgFg6A+xVIvbBPjASghASa/n4+5r3fF+b5nZWb74UVKAkIZ/HPihIH3np6L
ZHMOgdT6ie+Mtf7CoJBVJMkxvpdAhkQZjL6Ispobc1JskBg+MlyehMfBoa8uJ6u3tMQxufpIQoqf
nx2aEutsrqWoVwN7R44T7wHwBZpVRsYTC9U0OOk140TIT6lK0937HVhz9VPDqbr5HAPv5ous+Q4H
+bdWyIlseisoiFgDl+HcSbnMZf1w/viIsxIafJqWX353U1yuNt3Ng/bK0kTfLuBwYaFGDUtnJOvj
QUxo0sSNwDstCFmhxRFJAa6EMoBYgomx3PGBvAsCFznezkVzMMRfGCwdc2P4P6Il2NThUUf8N0Gr
8PG6fSEwrAX3wIQfZSD8VBO5ZzgVi5Bu8U06bP2isxoi5We9wj+b450CqiKNrgEPYS5DwJS0Syuq
KUhvSorb4XPR6FOAeJslVWgxza4IGFT4SfhGhYejyMYQSgNZcnBW6Ne12FtAkLmgStrC4stjlgxU
gI+3KRCzAwZ/sO6kucDY4vAqFvlx47JhQ1PKxQVfOXKv0wJ3dILDpx7Hov+ZOoPql67HPqcLttKl
Why3K8M3raf9SHPHnbKXZC+wkv4fSJIqY9KKmZt10rQiI9pk6G5nldEkDxAc66KKMu6/QvzMZga8
sio8lngBjDAaVpNcHmjCcaOWjgxvRnUaOQJcZ8j9zkTNiVUB4EokBrbbKku1rtqL3qduGB8onjNO
Qc4/Voj+SrHViM2e9kMwHn5FeG4W7gCGSyFaZrXAciDQfUzU/HlMFXEH8LC2pQJ0spOYN5e1sJ9z
4e31INOgmCFL9P49NFTFf+D+tUVyfrTdd1HVNSvCzy0S6PXJAa/cK3HwtOfqbmBMIqmcYmCiT66l
9vO28K9AiElcjB0m/h/EQtIANAjOoXyGjNl0rEUQjS6f/qfLa7v6+6TOmS0bPMazHQtl9obfXKSV
4gjQ/j6LbrHhUyZEwpeQwwGOxEoDD63BkBg3qcEMSGC7UOvC7PNOVHjuEnI6iqen/XfxhtFtTI+u
0BarsBFfmr1XccdwzOMyfGpVloJqkz+KHAl1Bl21OQxDiZXduZ5kb1imvachOnVttvReIUng7xGY
toI3V3wiwlkBlIH4WoqPuOONdd04GXVr6xl0Cm2SkXthIHU77BWjKxgEhIvRqXqGOYQlrP7uxD7m
sPZm09BlwYBNiAF72sPVkd01dovBSm5y6r6TVGAptglIxWwcLqcl835GzW7Y7SCXRlPvlxF8KAR2
iRlm2YVNFAMV/g1TcaBo1Dwss5tnP2U2+RTSG1jkzWGV+KukAobdtAk6EUxOUabhwIXXpVXx9reE
SegW3cdO2gb+dkjZXV5GElKWmDDYVNIocfPiukifkcRaK3O4geVLDn1NenuL3Xje4dl3WdFGyi57
MwLBdZBsmaF4S+Vfz4YfBKO5+yw+hZsyiy9JyJakXkY58vbl8M8+4j1p0XcdFJRu0cjnGyhAwW1q
XkCb+Dxi1X6HkRkjkUFW/UVrmgES11UR5fojhicf4m346KO0ThQXH6Yc/0A5F9OcQO1FiwH2RaCt
pmR107I4tIRIlXAoG5dC4OaIzw0EH4ZYz8HEXYpdD9F4FMPtajbYdzv7YvHF0IwrYvR2dJEHN+rb
GSrUAlOfnC5k7weg/jPQU2iNxv0qNDoJxnhcnnaX3998J6kAwd6eHt/LSuz3rvIusqey7MqpHB4K
gaSA22mw35pH/n0/Q32fDvBdYq3m/sV3ni5hX5BjPLi5I3SAcHBWCmzAIisQlM0mOrMoW/3LPPKb
6uODIWfhYO6MjMdU12V3RE2ZFRhRWAgV80BSFHZgotufRtVdFh1WP2nuLK7oaw20J3ynjieARD0V
kh66ve8LdDV0T/Tx1nfhiIc2RLY3SGxG4E59QtNCCyigOzyhRJ6MF8sis3i/O/8YcqdUCfI4mxYt
JZoFdqgfvSDGEoq4AMR10MVTSt+6Ln9DKDixd60YlHT86L+yDWPwn87FF2K5B5bghiOYNJEnJOtv
dMu+VRV1xgPreaK4DPTgHrlolpI0I2BuDB5jJRpVQ6mi4sZgsxG4kPcpL0XeQQ4YTsGNBDZ4CYfn
ZQKQvQDEg2vusJTUuHtwHMS8i3Jdd//qYTGnflD2ZwHS7AenGQt0ZNdxfjmeJbHIEjhxbdABQjw0
i9G/OoIBNIpIWzkrOaqQGmMrP8TTZoM1v//gsGLkk+j7YlELELK6FELFGlAniZeJL6hBLVnEE1ue
UeYSStBj/m3QEvFoCzoaXhSJg00gzRIhXLtEjLJyMr4r7ZcmQlqDxmQJSaH27X37t10hTert+/tw
nEl2xEwryC7CS1tFniG0as8PQKMsOtoOBgY1b0LhATGTIfsYoU5kUjNNqFQp1527EflaZiUgiO1S
gqUHNzxEGKTPoApY7hPZ5+SyGODI3AJK7dEhDkwEVH4p7NG+WQnKhrhfgY7g4yW98ENcYreuSITK
Dc8Rq8XJBi62wm+bb39clsCx0KZdNYec3NFUQgquHk+a1l2fG6xs5z50K6kyYzaZklnDzt+FrEAS
3N0jCJ3YpFNsSIMFCJRJalBV7DcVTTqUYCYZBHHhpSg2xpQCXZLkbZkE+pXUlVj9pGnV8sjdidE+
QfYYMc4qbsPLg5kpzooa6U91gXIBsbWycQXbAfpz7TT1aSOAj3e274oYLntwvTaaSI2uFAGS71o8
QFyiR6sWFDU5hT8V/BcromP7GnbTQjiF7seI4YIuPIl9FKg2LOBGzOpIa8SrtyBj0YQXZFpwaKUC
qD+DwukDFMEw2alxF4og5UcvHhEjAVAnWnZPQ0OpD+zXw+cpgFbGwvfVrd1DdCbJvsU7kRr3K3w3
uMp7KIx66Z5bNi25byiq3qgySdfIcovmq4ReX+mH5WZ8OkDV8gmCmLhefszdqgYFb/Idtg3w0exL
QdC39xLkrFzwi7dLkfLeCx+IwrzywhCcsbGxd9N8JcLq2pQU04pA3GVvLJTkEoWiTid70VB/mAh/
gH1iUuC2J4OdtB7n6fRbuRLiBepnCaQnH6eTFkN99aH4XjQ9wsjfAVn/h+qFeYRfBbPvrBwN3/dT
oJS08QI0l/RjTUVJLdIi+GB3TYgaGGnBjhWCTBCLQjwzzVudg6TtLD8mjDxReC8f9Z/T/z5hplG9
b+obB59tK9lvkXl+dMVaZtqFgFjHeInTUdvM30ht+qeeUWPIerA2Qo7sBsLegkJe7ZCcDr6OkapF
TvCPOu8NBnk5jbxW8nFiI32vBGYfNfTXlf84Dn/hlvvEvnAmEM9UaxMKER2YtryLd2zWosfonFE5
rPZAaud9nkOUqJeCMrABMUsMcln7/eR5MeEwmjk09qGdPKBvLGrO9OGbE/e4orch5ljbq7suft0A
JCYFgod5H1YWNdqKPiqSP15VgmYAd9FXjAbr0FE9db/vzuQ9ecybMS0P54uRhhZ73Eh5fkU5sMPo
VR3PrOQIMzRVvnBWNi6Ngo3vjkddY/i7yIcfS9k8WW0FFm4ImGbdcY9UXML+zrVRnnkxs1EDV5m8
0q9GsD899AZRflHbVE6ya//VJS4OyXMIU3DY4n+/2RymhFzalaDDvwpJ3PiLQfHiO/sCDySWffU/
g7DS5Opr8Wt1u4LfkAB6wCbpmN8d6A/zchD0/0btiwFvLV4704R8i2vKbECLwLknMjIrh1Hjws2E
l+iyiwdpsfa1jkVmGM3mLTLkJSIMqdQw9zWPt5Sj0i9PfcV59ZYDWW6gxUU7OvIpgg8giZngpScm
AqWyW2KImb14PE8XEhpiSEctK3r33i17MD2gA4sUCtnqWQXcwZ4F+na0X4oSTdCsBuK7jWzPnrja
on2vfEDtNn5RkxdPDWr1NNyOrlXWR2Iy+9kC96B57jhzXXCEN5kKXkOSAszVSs3rrrpvktQa5MX2
i5jbno4nSUFwH+yQacXzZeB4BTncnGSGSA928ryoELh0W6347W84v5a1xc5P4V9kFAiIIGwWlMn1
1LoO34rDU+1i0N+jVjU56/276VKW5Ddb0OHFYgVrgIiiJE+J1pIcjOi7FAYmKvmEBVdQKFOJHPY5
zSgMdlNc060Qm0O4yvKsEjvhpPogByge5StNcXPy0G7oQBm+3Lwgt/WHnujiAUtaz+C60HZXjH6B
qSz3Tf+Z89qVSZ83CSa+3gHO6JzryZa5APqEY13IDo+PXzM7KQBFVAhaWR3vl2vMbuCbE0agXkVB
EOeZ/ICg/+G6oOQu+P+/6S9hkaVvWXw80fhRha1mvGoNtiAvXz1DIsvht4250aJ1tc3yhi1S0Ns6
cA/ddI09dc6EBsPqhT5Bfq8hS81smNeIraysULXqrpy+AFE0fxydVTh2/UrwC7ZZZpcOtgTVaXIO
xYqftVPkjCP/ino7cMm83rZ3Q2JIGgoMe5qV9cfp63/OWjLf844xa0Gp+2zeGTuTdhH0Want4MuC
nWFl5HI+bMEqUz5tVJGBY7gHIOmXeuP9dPrIX74zpmiW7U28epWCuT8eDGRTlOBWaitp08M01Puk
ncY7FYQaD1knGfTx7yKrmq1c2JtAvviqZe3F9/nzWYWuAveBI2qCcncNEFn5A+ie5Bwrp5/V5dka
BkfUpxhpfYrekbEoiOj5sAdDLJrBgEqm0Q+5cHTk7+mHK1q5GYO69qsGLi7Yjk89NdTcAWgxKF/l
bwGSRRgkL/2popKkB/86GP+gEExvDBCndez+BuT7AGdWBCms1iwB0fwUH6LgSE25YZuHTnCXZnD0
5M+L/odDogDQ4xaluN0Jc99UOzxS0JKrT6b8C51mrX/KfFcdeM68fmq0YuEKjklK7qD60WqOuvq4
74yaMDsfjNVv0I5TSb6sjraMlvesuhMlFuzNR5iKpTX67XAgQmPcKTd520Xj9WTIPlbpN+z6g9/Y
rv3FFzJvyJamxHQQlp7h9py/elCznvP8SblkR8d4CSjW9FVuc41zFMAcLUDeggtTfdxjnlF6RVcR
mr6vRdevUoNaO0O40NmMilEFRMKSL7PvzHI8IquAQPv0mYR59lbTp7Y9p6z5U/kWJimBUD79FFDt
mbUYgkj91nr6+gs3WWvSWltdHlRrq2BXG4nHMcLPB0ZvVTGdghgbIp59sFkcmfWyD3Oksc8h9hDC
HZwOeZ3zEsOoBl0FZkSq9nHnWVXYu3/yFnk6D5lFktaLBN68LbSQh+RkgqUeHF3tIEeNnhXvqK19
Ssk0y4DNy4rxy0h5gKkSROF1PI9t8lAUy0mZhJ5Yq/8t4aq2GZ9ZtSaouoQhF6GAaotyVg2OoZna
WVqPHJdqLu85WqYfiLTkBbZjVc72QWHqCaJV3L2aRuVmoIv1Sju9S3LjW9ulEfHBNkHSaLIbKpgQ
QfUmwOjX7Zg/R9Y6r/sVNTiQGFhTAVW83zRZ2tQKhCOGOtr23uDMLRl1WG4GJzbs1I4xD3SiwmN5
exnRcMWANrvXfnsZr1jald02rNTaGD+4VJBWDfLQJfANB0QEPEkBb1Zk+TJVA4YCKqk0JKdrE9sm
9I7y77wjcqal8MofR4ziwGwkzmjLU7vLHK8rEm9cnecS1jS0wUWiZ76aKGupbhLHuTUj8fr3XS4C
lWotygT54t7AlXR5dCsf/iTYJi3ezScQahOOtvme9BiXaa/qIfbH7RdOGfZq+MYR1Zw24+kn/d5s
Soshxd8VV05h8t9zAaK30xZ/kNIaL32sHym9wprxLZzPtJstZMoXwtJ5Salbgp+juiZLgUrSP9gc
rsCFRTOZiimntqT7FBj/oCZUcdR64MF5OgIAaIJx2zeaxGjv3kwyGWHMnQyRIgMyrervPRr+ExAt
/4uKVsUOMv12k+CVWPvrqAK8Lh+Lk5AwnixSxzu9Kp7se/aXhjjWFwndt6Hchdp5l+TWg4JXP9ri
8FjsflbdnbNBS0d2GhLltR6E7ZlDBWeG9r6kWzMxeYYneqULd7MJEK8IWL7q40FAB5vdRerEJHza
s8J16+1FKdFeBLoSABd+sygTTEKzPyEZmyYxDF3S1309bytfegwitVXOc1CYKqlgR0m031zC8dmQ
zLCNEfvqusXyCMD/1meQl/h7FmzI46/Yz6AZvOb4/is9dQhGWpHdw338Pt4vs7L0uDSPQWUfoD4+
jqpJ4z3NCHJ3gu938DGtf7DU3gFZE+KMZzqf5S5OrIGDm6jy2SSwwi48eDCLstUybjUClLGBcT7D
qRRFPaFPJlMXJbHRhYvD/1UiZ7elTDOovXBIUOjJFe34XBLt2+5cPwxAw4hh9cOuN172+RR87HzO
yCTyVo6oSgfC3/HPSblpwM3WI2nmZuPrLSpvzgZzzCIVq9BFWY55myxQ0Wsgl22LdAN25h3kUUvm
ZTmboAOwU0pBykT1dWY3ZT+PV4ZxM9jlS1guJYA5dTbXTcULzfR7HXOQOjso1NRWhsvHTDHHT3yf
x+eHzGEoQXJCJY3hlDZ/EHbx4zr6/FEYQNvHqhgQf4lPrwH+vzyVl0of8lyGD3OC/cE/Ewe3Ngd2
ZlaE/CfC2qNZIDpVcdeQYmLAHELVqeIbmN4xWr38UAi0FeCI+iEFvJ+SAUddmPvy8KOh2y0PTI7D
Gwk9NZRUSJqXvDgrDXJ5BQbJpu8Gf3NFq1/QW4/8b2br+/ez1NWel1RJPYowNcfeG/y02z1JT3hw
7UwFrTDYHpKPSYgxA0al1cSf1msaOuZBOidDTYanSQolsTdT4A9EgHFL3u61yuBJJVrM3CJa6nqF
rlY0vfq7YXbeY0vR89pp8pHQABqzFjsg0jLMv09TAqTpCv/VyXlQr2uMXt+QQk3YNFTRdWc+X3U3
xp4UPUY/nW4cv3DHbQ1cHhGsmxSkyIoVz051owxwPMzgiLpSuQkX2UW0e2tbueIkYIsFGtoNL0Y0
FxPFYoH/BkaXH3Z9Is/sr/dWybDQjktvTg6Qntv3YelivIq/Y7D7EFtXdTWw1oGRJSObMbnt/SIX
w59x8p+VydRWG1DjX+cHxOgitJGzcJo8L+cBXWD4W1wbtLUiERpITwksV2JnKk9jGmK43NyBH2YK
Ee9bxmUnyRNKovAGBLrmXYcK2wF0QVFCec04HW1zAG1Oa63duPoFtpVkJ/PyrqA8w8BgJrQNZhYr
w4qtCbAxq2q83ETbB7QM4lVFCzGeuZjkRZXhLJLAS9RhaR06xOgQnwtJnqlPfJer35q6qqSkKlX9
sCOOSfI5ZBvDHsL4I9ythogswQNzFb4l+Y7Wig/rTqVgEK9N3AYU1drP86SiA0PEjB7ZlEPDuZ9F
4lnPUdBw9y/z3IbG1YP8PgaVwGFzSAP/A04Nr8tZXnC6u1CvKtkTlpu1+y5aRm8Yrx+otuxEzF1j
B45gfa9EO1/qQOzTGeK9nyNWaINA/K+cFWYRDHrSmY59fG04U7BokSSZDAwmx9asUrMNqcaVp5iF
jm9jaHmcRgt2h+r1VMFXfkTyHVcQ1zJOe7c51tNJXpd9JJlQQpfBfurqHsI4eM2zli1mycxLwRo6
cjtL0GQb87YF207S96DpdZSrxkTsYJLlaxr0oFd5Siv8cgSm5LxUS3I/03xzIPOH7kPT5BEgtU0F
juLvGUMrSHfSkwu6SQsbA5J7hnBNxrBXLVm8ue+Pt1p3T80y9TLkAtf1JJq5EZLtCPwhWwLQRRHN
HjDu14pxK/YKTX13mBSCP1AWeSNcBtA2xJHSRssPdqh5+rn3eIeuLk0U69URT5c5WME5LsuJDaSm
EBUhmt1OT6ADuZSFQge6dh20tVfyFxSXAmNwPPhs3GtBxPtVjEd9JIjvefRK/BayQ/KPuNhn8aDN
z1On6JebjgA0ffNy2O0bz0aU+vOsIYb0fbD5i4YrsgyNzrVSCOM4n8VO9cxRcRbdLZPVJrlRxKZO
iT7dn9xfhvLjE2VLpeLNIyNpKc0vcHWJrbogZoQ+0QZC2MUUVA2Jqj2jPgVN4291xxzZlluNWHOY
k8h88KSd6XpfD01TOn16zUePAqdZnihJ9+MqszLKxjzVf5/kRpXko6U4XciafcgcXZj3wcynTmpv
IpVjsMqFTQfnrDiJKchmTA+/EH1ip9auNnhIjLTIAT+3xVTiKoQRAsT2pgDfzb/K4ip547HTgDZy
+mCFM1VPIpgO5roaEV9gV0KZhjz3WJqs07CPwdAFGrZckzBrJ95is66no2eGd+SRkDjlEnZ7LMkC
tEU8yH2APFjcSgNDaRAVv9yoeQ7R+ZtsnNXqPIvnS28SgAZXF28Ho5kQBcGql0YDsyDadb4F3DnA
lk2IUTrUqyTaj5P1eG1xBejE0sReiajI8XRVQ4v71KvicAO20o8ND1JSI2gTBrEb+55GWR0vzfnR
gtqO6Je7k+UnNGB+lTP/KMUBvWsfw6Cs/64BYGvDTbhT+ZWY9lvn7kNReZ1Dri0vWC8kB4we+ZpQ
9wEmPXWIZo6i4WTDPgKAC+1Ro5+fhCOMF/gp8Ku1ZIMnDMaE2yvRq6bnXNP/1budGcmfERuLsFBx
3BKJ5HI6YbkIGrvL2QPoYaADWKv1sla9bfzmL/Ax4ddPolXvntRpYaRnOauAG6SiWMReZIWAdbWW
nUDhUJGTvc4ssTkXEMY1/D6KK2GnDTXtQvE+6eagY+XNAKg0nhmS2Aqm6gu+2NniVGqL0DMZZO2b
fASoxuBNnD5eFxbjx7FtnS4PVJ3+CPCgXJO2BXS3mPt8XJS/6fjjClJmvIo5HpA7Xq6pHI5tcIWT
z757b5s6FHbjbCLZMpI6LRQuK3R5bl5QW7r2sW2C/8xHR53t4DvntkpSfVqstxioaTgg8CgCMXIL
Yqf6ansnPCz5xbeV3aMe37JK2qAwHcflrFBSPuPTV0tul0CVkxB7VFGtNT2lZnucL2hjc82jvPKX
4TATdivHZDpra3xa/0BYp4VatVo1dXLGUZ1QQvo0K7leqeiZgILJFTo0sHZx1JZshmd6KyF9YL9n
Fq+k9FDLUQQFMVBeDAFlqw0wIZOxeU/kJJKalLqYK1JTfdQWlAVeT11BEHuL4BCxq00CeCeeKQCc
GJV0q3xlklwPESCuEuhShdqZvoTzU/Tf0GV0SxBtha5KfVN2ftdbJtsygLkaTks60hui13bYDljO
X6jKzF9jAwS8qufvjRFBGqPsKcs/jc4DMonRSsPoN4JfYp03MrVY/PJGTUl0uueQ4hOKuSp+bcHY
VsC+5kgey7uMmXCsasgTSvk0wJ6ZbvH6uLwiBvKiFQvcfR2JcSGAKTaN3nH2XwbQZoUPeqSGFEt8
19z5cUQkRoAaIBLIJXK1a50lNYhUoh7uzaq+kV4FDL3PmejjBHo3X/90s2CZxx276u6u3RNaOPEi
vNhbS0ZEKBtig0ABnRJpRER1FBwheLiPOaS/OYBGfJRldnb/xwDENwJb5zijLmWTcJB9IUBrhxXv
pP2O+J2BLlBba6JhNELn/YaLooW51+T6jmXIVMBufsiagmQSF5z+o750rrSctSaL6rAn/vuVs/Vn
PwHbNsiBYlhDQ7rZuIXn3QtrMHTcAe+Y+kQ9gVsdRWMGiid89kSnA8hABTQ1/xaNT9ZtgyNzLBwa
VFkRzgK3TWA2J4e2Z21EZ7I93183W8TkWZHsNDtZX1hTGZbSrqLn8qapdAz2yTDl+F0cr8Ew8gru
y4BcTtId2dT2Rf3Ru6N+/sTGAW++q1F4gx4VMBsQqRQ2AXTAgSXa0YFPylq92Il5KLbDzHtJmLJY
Lq9iiOYblQUOY7wyM3kmTRP4yd+yXJh0b7yQGE8EA2++Q0A42B5cUpXo0MPFYbMdeLkDcMDUqy/m
Oqimfpko6KD8xORDsHuO02z2SR0nmjOO5S34mxaeUFN4sj4Yq7fu1vRyNAZmbZvXGjN8UWhce4Xn
4Me1f2wXn1/yNCtq8NfUCTeQwP9+GtXPfpn/s4PX8TSSemRLhCC+cDjvBLksFRjPlBLsot4/MO32
kIjBZ36HTFVJ5d4D2U1Nj5zWKE+lep9tsc8dudlTwn0sWws0vlwD+SJ4+EyoqWeZBiBmdOwM7xqW
8mZLF1/+IhFsh8pVnuOXZQ5vq6lRPXqNS+6AmkMuVY6DC5B/NyV9/Tz2XFeoOWGbt/x96teMUMYY
QsEjaCv/A15RqCxh326plzGF7VjUaURUD4t+P/AzcCL5KRsMZBH4YCaqxFop2NyauDE3sOSHDfmE
Dy2n3U8bECZ4+UxZ4E4wz2hfdos4UdqUtChf92lrOSuHPMQCHEBn7U1Wwj68z9K4XoPk0qTaJZGz
ahr+HOSjALLwYeZw0zrKVN0BE+aTvGmh7wDqkgqgYS6SnB3JsqVGbhp8AedD2qt85uLoywXwPXN7
irFiIiU573v3Re5SImLgB9EsJdMTEhYztLjXbAhS6lJMLbiNAaNuDI2x7OD1GxvDhuz0K5mMczu7
F/kTKSxvNBjc9UQiJfq/J2LMM4MpDlLWlAkH8Jc8nw9v129ROIpCV/jGZDm5yPQt4791Z8YL4V73
lM69wouwq47MUWLFW9cPhSbwkjk7nZBauuZJj9C6Zpsm+pQK0mrvHPg/BpBDPA6c+N0U0q5lIGt7
54hCkUfusUca+155LZBm9JAeuUTvkRstZgfes2ngiExnadHGbjSqgP8I8VV46zNJ0zeZ1z73LKWK
KqgHpti4La2wEuychPKpKQjHu/hnz0m0jM+4K1Kkn7mw/q+kmE30NXBDQTGOwGYljZy9a6WG+SVg
uxqRz1YWytJ6lyvZ9UhrP2S/+KzomiY69aC7jC24EISGYEOahFOAFg0Bx60JqD0iMHn1T9PKLoLH
FqV9AN8G58V4hjy2+11HmnsEKTUum52RmgTTiaPzYeqgVM4j3kOf6cF+1rQf8fj15RPEi/oEejeE
GcAHVjZssq3Q/3QmLzTm3ZOAdAXBtrcVEtkVrziCgp9TnAzIecwPyO0BtJCZHfuiHTY1V6a8fZ6P
mipJUXfUhmVbU2E98I8K7+eJV22NSh2ohWo+tZWa7qpYqNzI7KlFnhCvr+2J5BK0EpQYnkH83fCO
k4rKDjT3UtiGX7NnBKZCEM7hg3urx0HE/EW9yych5AVBGqkdJCJoDI59H6xQwziT+zc2dcEXckA6
pt8fU1EnDpeRblebzRYAQ6TfxptuQuHwlagycewgK7gzcKp73ol7XZDm6f4s+h3IkWoBdk73jYwQ
4zDZuRmKfu+Macp6Yp1LGWwIsF1vMVES4kP8owfJUgh22pNmZBD4EIehGGw4+dJn6ARN7dt6nC2i
Rw8rjBi4I41gwgYBPppgFpb+bG5pEqTwrovr13VMUC6ntktFmsg3Xyf5TNA2uRKMMdt7c8gAMIzE
uKA7dkqzpvWFqReDOfEUy6WVX9K03dtZirRvvPmC+yBvxkk4RXEGy0vg7KdQJsCTddfbGaIoeqBD
5OQyvd+GbaZFH7jk69aQWSK5X7l/IjC8L6p9HrPi4GQ6oNU1c93QG1CPJv44x92vrlXPqn+Oo4gi
u+6GB9N1YeHdgtLVwL/UALwO3ABhP64nIsni01AYvFMfKtMtWgDajYgfIaKQyKsuGJB7cgQG9V7Z
Xyj6HfA00e3UA2FyZ2NrL2K61UpkAixR7lwXjagEMYqBK3N8jMSR+xXgiyphvwYLenwvRXjbYkyu
UUMFvNSseTXgysOii5P5O5SByt474zdrBrbKgAEueKzd/1OITrxKMBxW81ks985/hz7vJpoD0L+H
fp5G0P2pWMSwgFk/Md5l6OO6X45cUMcaajcvFflUVk65cJPvozQt6YBUHTi+hEImUIN9f1s+dKpV
I4pEPsFqg4BklqBke3uovSRivNCj5AQIdfVUmIrIIHH70aQlXNy2wCrcIlAbnkG1lxTkjjRx28m2
xvrAUSCyOCyip4t2pSEDjJKMZcyT/pU1gyrMbIfl0x/9R9eDDo0teLD/Il8leaHrytpjqLs3rCz8
ShhxcXKCxhmJtuPLobSSl6ZuNxS9MHiBRL2Hh5fexhTJucm/OurQ08KxxI2eGoHVuvZa8zQ9shM6
vYkLOL2hIWvi8SUkscRvrf4R9id+jnYu9nGGicrUvgnqv8PmOC4Xn/m8dxXTzB/8ibZej0kCcnCB
hCruZilGXCev3wAm2DK/WsMd7q7uCwpNOLufN5zYxPU/ALGcM9Z7e9CKQ8fIXg/Uipb6Ec568joH
C5ykmLvmVeH+IM7eQMKweqWGBLeipDFxnV+Nu+bZWJ8dvNejUf0CGLLgis/u9pxVP3aLnVMe5uQD
Lrw/VV4bDUlOHsNGuUF3KCUL+jsGuo6Rec3G+czw67u85Ksttu9OVwVXLJ46nyQBAdWDB2+nwsbW
hgIYI3D0WHkiTDvzSzWPX7swyQzptwOYvu7HiqIaw1u4elHePb9Twz0zH1AWJj4lq16E+CX6GTJS
Tmz6Zss6lQKIsvGQnQJ7d8fWf7J2cZY5UDRzOUdrw8Cp2hpoUq1gf/7qOC5Qb3+Nfv5t5/IalELL
kaazwiz8djo9K8i9R9lidz7bYcbJF8c1ckhXu1npJZdgiy8UdIK52BFY65NjFQvhwZEpP1rcq0Fb
DSuNHnj8pm9auQ8Yjdcxv7qdUbf1mV6aZ8zbVEfA0J8Xe+fF8kAq7jge38a8ovF9p8k7k2CoA+/R
ZVLAZrN/cKQaGWbISCIRppY+gcO+c98VCe7uvMPN23xmPxPv+FMBpiM+RroncG/Ib5g5289XUhOg
/zF74Fr3XBrT3Aj7gh1VapjPq8hIzPdj+K67oM1XCFZhXXq7cXiqR2qWIZjNYMxGD/Lu1Uv0i9PX
gvRvYqCy1Sgvd45D1laeG6psYylLFnYP6h9E/APF+SARQTOBVawzeQivoJdb7k2wpxkW/wRD1PjG
WFLaOBYyrNEQjvXUrslvDk2yjJ/mDAgoM2Ig4XwUis2yDCjNlO3xhWrpHmeRAW1WLTfSZHcLAzdT
uLZ60g4D0/ZzdUo2ar8ViuHOO9xrR9MpIsvQ9oUBPVgzJy2qt/ufE/8Q4r7A4kJ/9oCtuP4Szwr0
VFj1BcPDOT6M60oH33IEtU1zOXUK+OMcsoJnGv3Z1WlgmySPFeuP8DtEuTFi8fM+/dRmE2X9qYAc
atr/QhJymnksabSXf3VVofUP98o+GGuylJQKe4uoniAVkbM7QkeO04fG6x0rs+PHfJlpHKSEM8UJ
DrQ3w3aBfEfqE8hMI/FSpjIh9KvtdlFeG2NIdRaMVJP1GrDLLGC1KZ53nhcpTnmaGiYEcs+clp04
LWkU6OhK9kk9ZFwhtqUadWFupSYdNF4+zhgjD18Z6tYECJ0P+pJIL1OTVgC5ja/+2l0s7heAD640
3viJ42JOSrGX3E2ZxEfeK+qkUwDYwqLTVvSFCGReGgD8rkzDLnscVIWVOiAyk5hijnMf11NDnAxw
qcql2F6aSGwLpYnoPxht34w8bCvdPlTKZhmrCog7wBAVIrGX3SgxCYaEFiVChgXqvo1GDRnWEdqM
1Lgw/TPpFYuFx+RcrPG/yuSanb+RNgN5Vga6PyGBSvt1UTi30ouaXVvcOba67HgVmovdahIDVDO7
avzoduWgFmwq8Ry5KQcc2bRqTwiWnmJfmqhPYvWK+0SPWtX6A3rEdLqs8+y/wmh6P01fA/ez1UOm
HTLNpDpyU4Caru5KVe6++WjgAu39tFcSgUcndBkMPvJu/vzA/YGNBmoWhfM75C+7gW2c4qCze46v
ZNQfB3sCiIhJd79q2qc4/cx0caX6ze2uidD94ot2ghHk1zD6VoCn8RnPEwVIo3oIGVezrvzPbeVn
FUmqRZnyyr/3OHnGs0coIbYL63GvOP37I/Fsu8+NkzQd5mc1/5MnXwsxyEqsRj/Nq+eC4bYN4HlU
DfE6bfgJsF4iZdDx3DWGQ4VH99TICs2dMTCRN2Q6YzHV1gXDHxzqqETN3R4e8IFk6ictvkYLmIm1
qMX6/UzJkgpcDCAiWPYQPgmBJvNE8DX5Ltdi2ZKS3g9YpFe8Z/SKLi2ZoWU2R3rGinOSovtYUhki
RqRQepZpvF6DmqIzl2OEt7Ne4GBKo4+ovYOOB4HtcCQlkr+zh8hEJurinTTtRCvdIDhjUlttVUOi
c81SJcQZZJ/tMlq/uYQL/kfFSa4h5euIfhwQGeelFjrmLb3dwwv0xgtclv4iXmzcbNpw/Go1pzB+
76leNbKsiCCW567PnyF04JV+NLk05NT2JCv/ZbRsHxENwATOA8iRi2dOq6ElK6nqhJOgfhxis6lJ
cIzqAJcmjCctvjaQMuOvnHYMdbh/2AXmjpnPM0jXyudvDLJTf689ICkKf8alKmwyhq0dy149ZzLV
bo3Kk51pRChPg6XPPPjl+e18PK1DfZs6GL6NK3ceKTWpWiH44B5f4QYVYiuEWJHjWKyQ++j+htkR
w44oymjMdhdbBM5pgGToBQLVbc3zrKt7cZPyiYPxmQxRArz2f4iktKBGtpyP6SPtLwc9Q8cOiqRu
Yph8b2Rf3qcNSjXLjs7oGAStz6fMSzDnGOyElkM410ZPku95C4GG/Ln0ZjDSeu20+mUKR/IJ9B37
9KO28YbGbd8tvSFbRpWAwOHAdHbo0jOKvSmkEknkLnw0giOmQjbiuKVljiNsOd4YMcFjSQNJL2Rn
DGyPJ/GQBL5nnNJvakIEnCaxEarOosHQAltfS64Xh1AAzuY8pEH3bNCSwTtiGN+sVW5wMmr1CJo+
nEW2SRUYtVjz9351KoPXLtJgONT6wpbDW/f83X5EivH+zJj34tjPogK6oiKXoTU+Qy2GvPtC+zAl
Op/GsqPCUjH+qFpRDwz8abwZ2pHl9bQYYAJvNK2BcaC1ph/n3csajlBy9vwrxjkAjzz1ojxn38c4
C+ebvB4PRe6D5ZPQi12usS1OFZf3x8Fx7EW82naPVMTwW6di4q0JRcAyASyG3P+1sMzgCB2r78VN
M5l/qHh7Mayz1miEB+ApSy6m18LwCq8UvzKww+7otCnBBFe8KpjgEewMNmp083QYlkNtzgXKGQBS
2F5vayLQyJ1sdvQWgSXPFSo5A6M/ry0LIarhO3ZN1h82ZHKE+RhJmyjBHAORGXM4MI8DWdg/7k+t
IUthzD4Lrdpe+QTmZL4d21Skung+uGBBYjld6LaHMmOgb9swQqGIdil3oufg69t14qI8zTa67oTu
lTfgLbTWn9ZghXaHrH59IC8K1UJgJ/6eyF6i/4dEmpKonFYB0eplHofZY7KmK6tcgX65hcBe15xL
KpoIehMIWXQItaHCIcASAoNNGEACyQPurU0YyELM3NDQ4igbpGuyU+fKVuAXC+O5Pyqeo/imTOM2
rnBs3C2fzAbFEd1PcxnFCITXvXAaLpg2ST6EFJmlQ5VpyEf6Q3WGTQ2m65BGW/tOCDP3iUzySF81
ufp/3phlD7ez5qn511Sw0UWDIZZAE1f1S4sVyvXhjCiJvDcnY65IN0v0zPRIsYBXaK/5GEkbb3Mp
mq0rY7bg6LxcV5xTMUQ8QB7DiA/cSoytlz4b4l2Ke4iCcwvpHlW0BasSQsci5ym2ieWjEFWrdiPp
hFi4SaR0eAJHpfjKII6q4TlRnN4f0c9fHN5vpRXcKXp/ExuoBynepUW/8VKM4LkBp9nDrkcvrl7i
Hh/2nd7ph8CmGGQlgQBYrY/W3tCpLbs4HvzHHEFRSDkSc9i2PSUR9unpqsggPeZvo8QhSgPK+V2j
UZaHSbDS8kBMPJulzp4Y83xL03lm+Mb5rV12nXBrVpOCLDVMSuZgudxcIVJ+t/0f4kZtwzBFJCug
fZHm90DKK4OObGpBBEnDS2Oa1anXs4NhyCHnxUiauYI+miI3dGtiXcPfYblRGiEr9M3tBzSv+6O5
w34k24cmwX6AfimQoLAmhIslDeI+TxZrL2Ro8cbdaZGvIz93RCakJatUXuItldBXfG+Biqeq+7Hh
M+KNdG/XJawKSV1Tc2nJ43CjGb/T+iNxasBWRx1XZnNp6uTtThpQIvOw3SWUAHg8c9eaT3fxVCTa
rXUTU/V6C9QlrFNShL5mbDw+82Am60SkhOjI/eRLlfATrLLa76XLjhly5/DGvCzoxQySb+qPam3s
GM6UnjiQrXJRPE6dSqIsx8qgYpt9tuCKzwqdaK8xmV2NnafRAwasshA0O1igu/4ZfSE4ff5gHHvS
VC4SXu6HCBlTH/YSgq6X1WQNbAw59lhYlMkDyYICK6uAaINRyPVn5xvAEBGeTvmx4YeMCoNxtQcr
BwwHhImME1lOc3vHr2qZ2tnPC/7VzwTfsiviHYxcqUV3tJaaXZ+EdTFh8i5pFXyU3blHJ49O8kKs
1jEith2nsFUEBE7Y/hzuNHs/R3L/co5F8pGJNyjHeHwx+4VPp4z3R+QFKQGXLnlErrzo615UBE+2
HaJ+JDq4WHphhjLU/ZHMTXUWsfFC8F8jE9J2sQP5aGt4oH0Li1rOZMwAhK4VlJ3A9BShn0OJgAbG
yZKWXnBrw3lfFTqkXo1lliPCfRNdg9DusUAxtph9OovlKH5l8kX8uQvIOygScsqLCbfCYYHlIX9I
uSGTh3lOHv5UfvKg6g0jAdkVCz74aWn1s79T14UcPagnG0SOIKTLWrfIqDFB34ChBXHa+aXNKTzl
3JBUOXK5Oaj73bUSkXshyS2uAXwVTpP5F57bJ45bQZf3+9MLPYHAJzn0S95KfG9tyeiCECqZjWAS
i8jHoRl21nC0OcL58czWO1jRCQZClUdcH4vVEXzYYM0//ZF4RQn26nyV9iNk8yGlqkBAzEXmTNbS
qBzgoaChgYv3o9hwfoHg3pEV+/UFlOr1RZeGFMeklhzI89GPVW3zBwQ8zNwYKY4eHplXlmzwXUOV
921U7KbvU13oUB9m1QdH+99wozH/+2nuVA7hmoKT/drdnhuC/ev96KI68d+2e8oDxes23unXdiyB
Mx6XtEh3vxZvK0P1nP+CBE7qCvR4M3GlvienuucNHBpSFOVbOgESkGTprmaoC5jT7e/fAVYW4Ncd
aRqHy3HbKsXMvDqTDwmQSr/b9Erkecgn/Vr4VdVmL8dB9udmv78UASjHN6PF1PENa4lkJr6sbscr
aDqodLsctRhPGveuHvSjvxt6WWeXByeOH+xJTMxCzEKfD7yPnzkbznxH7DLO3YWKl9mFMRPU2mLO
A0uUmT639D1JGQt1+jwOWDjf1J+mi3FMMryMku6qEsijHGYUpaW63EMlzzAqWSs7C9Tuuln03imP
Kl45Y7w2aBJ9pAd2z8Eglgy0PPDVpjR4n9kZXmccOxiveitAMQqn93ko/Ror4evVzuouLjUXemrQ
8QNQUJpAoXblxq511upB0VHMqWU9tLazPLIBHC1zps6BWM6XFoe1oYnmp4imQg77P71wmUNPyiJ2
G9EgeT+97d6JmSf4qtvAF4qks+Fl8VyREATlpXuEH1i/oL0SQRi6fsrvH0zLV00uywPQ9Mbg/Ef+
HfXJkS33hJtVcnWQv42qYfNwiyefmstv70ddYd8Out4qn88f4RjFYEnm3xjVEnKBgZpvKlWRi+Yk
vgPWsNADcgqmuQh4yxDd/wxCM9mE2z3x5o1jqZPI/HTAtGDJuprMiNqFAGmzQp1zE51dpVZSW/bd
ZshgXR3rzGDYXO0oxj211urqp6O6y4T2JZ0V30Yz+buhH+GK6AXqTsnriuK0K6TegzFVPod1uW4J
slntbvHE5x8eucX/EdVFZapE0HwOhmTiojDBFzJdWDxoQU9lFdmk8Aul4oA+rnWFtHbWmxbW5YKW
QWeb0xLtpu3q6sWiWgeau+HZ3H3eq9ktkObfZ+7+kcZ2/2joG+U5UD56q3d+e8WIHAJSLr1qqyN1
1onwvfv2jXRhOD3NneVe1yIxYRcY9c/NE00WyBYxz/ttktg9j5pN55UughHW4jEu4VBJ4vviFZZa
drlOCxIe9aq1hoEYRLhlNIXNOXlDXlgeAAXdnCfkS4jgEM72uKfzKjDSADW8vzB28/k8e4UDmAk2
4ZLBnqKkQsTR5oyaoj1SnLRjJqHo0HepvC4jTI2RuH9ZNMF56+ACGXy0qEr3AKD31aGr3L8JA4UR
+Njq1pRv4xo6Tr+RyGTC+Jck1BpzXSv7Z+HcKsXQEtX8NfiOBqzLIH+/0CWRKtZ3/gOycVD1nVyO
8QqQZYSJliukACIZKWO3o/s1Jn5791514uEtC+U2MvwEZbLo2iNVsdE05lscAd+T1S/hjGwJtMuS
UkoM/EmNtckBmfjLJLv1rgE88LiBPi9HMvT2KT9FX4TXq87Q7B/J8+3i3BRmTcM0ADpoND7w+o8l
aEfrd2alzCEn71kUX/vfDtjPcvtD5wPL/4ZLEi1bAz3qCcnR/ge72QOD6gqKaLFw4EVR434WG+30
Zfzx5IcvcmXuRPsAF7UHoMTiFhHNN0S/YcT/6KApJpLXJmC55pxHocsu7MnagplKM3BdA24AdQLb
L/0f77oQrMf6fd5DzHocx0ORKsM5KGS9ne/hLqrOzmlSfz1F1WGnikphX3z5f4e7yyjJUIDZvUXF
wwtz01J9ZyWKKMEO2jFS7Ov2dEKN7vcG+8vl+6miEkEZ8DIpwCJj6QSsMxznLX+R1bsZPuBRbwdj
uC7+v+YEoCFXSlIdin9KsCSUHQRyTa16WBxBGaFNflHmlCPpYz8UbwkbG4FXQrvxeNsFZYfg/RJt
Rl93xbG4C9hIhHM+2On9EUu2ZVlTdYZfoWniPn+rDsgPa02tlnTVpP0TANQ9ioPOoceRYBUydhdJ
ZW8m5HoE7gcfFodTRgCq2aCgFv5G8b1TJWXRNPPR2SpQAZgon0nN3jGqJ7d4Qe7YaWxguqzbIc/y
ZQ+hQPrJyOQE2IhsQhUAi8VT9XjIy7fugCrATvgumGBKG63TrTXNF72DJwFuTVPhFTzvMrrXqbil
W0cpIAP66nUDF9449wj2JFEEgH8NZgT29MptGmSBEMWDXSMYGVPICcF+wpXuTaOMYQw+Pix+fJft
KmKOEhtKZi2+R1rjqxlExirmzlifL0a1vQZmtUTfQYa204vePP8Bd7esZNAU06FHYeZLFTvvnVox
A5F/DmrQXKo6152M3KaSiWcLCLLAOX1HvhAKEe6+unXvXe9XB3XvtEvdgcfn5o9Z03194HnusBLv
mWWQaD0MQRuBgSghdax1fcDj5Hv7IaLRdP40IL2PhY8BTg0aiZ+JmvBjFyod0uvELlaK/c6zC5sk
IowWibHSp/e08kuEDbuQdLYcKceIDCqHMEoYn0I2VUHDcr9TsYbJ9Pv3S/cvgnG9+80HGSJYozmb
y/03jTgfZRFhUalPBdP4ONeJsZLI4CJIJtirlj0Oz51A9bJ1mg3WPZMk8CU3vINiNsLUxOd191Ip
yD9zZOK1eWHGfQe76jcZqyvRgnMmpOJoYgmPbsc/00Bz9HyD0M6k7lrMFzIH2frBMgeEjQYLGIyM
t/CY1fuYeq4aGu/9QtQ/zeGSatPLGWk41El+idzPOmjX4x4M1UabNF7nHv5ct2wX9FZP5hlDHrA/
mpUdEKIWvd7X1BS4WMFGLgp4UvwCn9ah0kevyPi5G8pp9u/qXD+QHF5e/yLWO4LDJxgu2A4moIOV
RfLSYxfe7i50joAu0VmEqUFVSpkg0vo9hcIHxhMQToOg4RQDps4ooYVKJltrQnvWtNcctaHqrzDx
G/ij5cDgvDKxQeFAAwSgmQgyAV4/gRUr2KCwN5zy4XEEx6gkoMP7+KnhwAv62HUlOI+AnGF4h7wL
WaLyTN0FNWzW0eX4scJ9i8Rwa+0M9yY06nsy+1oC765QwTDv0MbWzPDwfkZAm3z+2cBbqhikIuF2
w4nT0PqPg8LO2n+2EkpiEtrTYLCk86DheQUKDaDJ0SZxyvekZxgXRGcT86wCcMbNvu4w03ntFmW1
zmwXR7pDIt7dHdUU3m45NCxO/uiTWMw18MnWH/oubCs3Zo2Ol091BIRUE0GG9iidEAaWPrdwlP68
78lcqdecci+LH5ZIfrr9eaTzE+NArCSlBPS1sL5PMpeCUKxXTwBKi6xmeM3pyjHQNl2O3I5HYzER
/0xLnyFsgWvtLqkVmiuxf3Yvp83UDr6EvFvMTCB08Ya5UUUMocAp60QBZHGHvnNxuHdhNfAf3ilg
wCflmCrwtmgZYEACMbkNZiiKG7YRySQFutwh8qtTpx01foE5/HUV5RRDi+RdK18j53AkDhIDOG4o
reeKeZOFAd2RVqwXt/wf896Wd7gsLu78mNbFbWEkykGKHvzCWDJaPdKXxsgo06x9Umjfs64wXcZ+
hLmyTgTQeh8nVlsAPxDR+/t855D52fXg/xsRUjmFT/C1C+GODiijBC+KBV4NMWN2JREBgWkGRayG
zmh34I2aonColyLQQ1I67lU0wNWy/7bKnTyeh4gvM6WFmNJXiIno+mxkgDrBsoWa68TURverCCHI
EPuSWI+bteNoY3ZlHFSYVyiq7tnGzv/WBFIP19w+/eZuddVdF2BwY8swT5PBIrJdH+7ef14g9pct
gCf34jrVP3e4MwV0mLijqz7YKtlIVhBTfFE0wb+Ud/SNklmoUwJn3Ul8g0H7sWO5s0axIXsWtKCU
s4IBdgO1RDfW9gLXylQoLLJ5o3+FME1GhBlQMcsu4pW+yuCLzfLC1E5zh8xs3h8jjW7H/LjSR3gR
5Ib93pOdiMfl+1WNnhKa3ZcvKCRWT9GDXIdhynDTn8VL5Do7Wj995/7/y2xAfO1KQ61Q6mR8To/h
XMkATN/P8eBLA732ZX6U/5edpj17haIs7fo9HVRUahiNteB5NHAmori2ZUjo4n4JwHCqeA225mFo
OsZyq73DdGB7psRIzR/GkJWXi5YUBLLMuxTGcP1RHcHrgbJeItRJLkYGna+zO5QR2wUDkrUJL0Ad
3w0YVvd8PJhnmOs7sguS9PAnScs+SscOlyL01hUCvsVqKM3UkHYIchlSqvIdNItL77nhGBznbrnh
/DEblcAasz60bnY+hJO/K9+X7Yfl+iCFQl/FdAQWa+BFmJ98zl6x3hbtBkxZ+JCnVDGA/lPS5xJE
P8fcFo19P9l2OpsYxmBFdzFLorebcHsZwVauCKwH1BfbQJy9DcXdY23R7QM37K+4wKeEFLfVcITd
oQFpAM5Jo/rgWIlg3nM3ftADWXr6coJsFrIHuHNtQPVXGQht5DFwcJ/C35Thx23q7zb0/V6wZRCk
HBjJ0/Oc3jeAPESJzjmSM10T3mY3l9fQnY75YWYJQdtDyF7NooTal8Oy6T0Yua4FGj4ZoxddTk4g
EYMNS9byOqGFqhtwLTxZvS3fZfwn4oyE09GwBlwfq2uhO04uUwmyRBzgWeExfJlVEvcAA6N61Zrv
XzyAxxiInjo/KoFN/k8ukmp2RVjiYnRaIbkQQvd8nDTc5M/9XaKMGE0CpYJuS/BgwmImREQW+I+w
8zTcFaS1zyQZEnNflxxLyP3zeTAGiIn5skHi2lkZ3ipJhA9Nnb4Gf2Is3qdRHOW3vmnomzjop0L4
VP9W5C/QRyZchvmrp0MgWGzm6nsVCdR+ftxbpTFNRTa7zSppa2gqtCLiIR8T0KyX7oJ/h7grIyjv
eRwfsglDCXCGJjwYUTBrzdGS0mwilVvAhFZmShkEanE7fSZ6LIa7OjdsE8IavXTtnd4Cj1SaxUfF
yG3GcuhvFC9/Cftw7KqUIf2ZtyUzBJmcWNC0ZqZfSNjt3r0CJ6b10tcX3xjPEwRM+a9iuVcbBu3c
f9TG18XY0eDBI5lGRryf9knjh34V+HKYz9Od8Qi0G7JHuOvvmyHRTZvdt1kYwRKljrGUwVU/ge3n
Tueld6yYSKckx1oMSRFSR8Kau8O3j9JdCUTcSMsyvLUiNGQ6MjxF2PChPqBQSDVQDiKisjecaKN8
cTB4PJ7dq38nF2TLi7L52W6StWOMjPoUGI5W+GxIZrl5dvx/dC5lPCjqzn1wihtgGxpR5KcKB2Ol
m0AaKvSQu6QBOvaaFgzgaI3EoRj2ZrcGIasC8gr/8ZO5yt8N4W9IUiACWJ93D8QkQTY85x2recgx
THo/Fnz/s/fwphhWy8ZlrV4SobZPGspT/DyJS5H2rZE13jzWFSEIdBqy4X4YpZE5SSzb4mWXmxb8
cVYTM6mT0G1BO3xrPpotvqCFQjRWVdakFbEBMLWjro1+ZlBSiTbdGnqx2U39bTiZEnqYWL1kfRCO
GpcWWmYZ4WJAEUDfycNZVPNxamy+uvjayO4dg0ozDctB1zYfj4BW1h3qbjVVf4UnzTtuxSxtGTI9
mW1QoqL4ak9Zry1+G/sZSFoZjfcgvsD2C8YyIKMNXevlnEeUNPaBwtd0U/FVS4LW2ky34ne0pr98
dhjE6DfkY6M0VvRlQHmoz1RhnfVBnWyBslF1NTfwQkNk+vb0xLIAAr3PjKlCn1IJb7U2IPdetLca
PM0Gnqs3+I/dXNCcmbC6827lQtGLuH7XSTjJMEKheYQDDph5dyVQ2zI5UCHYzxP+l7wlM/aJKHX0
7v1Xf9dGdrkM8re2MJk1hw7rINYrp9NfkIs2/bE8TPIW7IQl4MuOcjFr3bd15hxsLDL9fYwmPITC
MgbVo7XJE9RTXBgobxXrGGO0PHFbOng2zspy5TWlRhkImH1xcWdTJ6xVZr1aAIvAiNNjNGAFiLLW
LfaQSK+OOYE84oPtqiNNU5Nwfgx1uieCxahSwCl7SsSuhW7QKimh2jI3CcyPYvflJNqd8Iszpkwu
nqx0HeGG4hofDLcOp3SDFL8SRfpLZxU4+td7d7WdXNDwnXDOXro2E5jqPnE27K19RiDJfDqchMak
Eb/BcE2x8FlnCa1Xk/ZcJ/ddbZ4fjkmTn42LLi+AnQZeImNaUwLu5iaxA9tIktZPOzLA3H2QBBfm
wa4XO6FOYmCsSGUK931ZaDJV6163eMiGdtYh/R4yPOkBX18TLDli/bAFI1sRGGrdT3/9krngSho2
SG3OmIMrqBMdLQCHsDjw7gB2BX/5xCr6t8wcfTmYCuWv+qjkOqTfdJaa/B9Plv+EJgPwV8O636i3
2PhQ1pXzlD8t+wFj5geRpZwZWzFPmXZo4iFtY6LRPkgl0Vm9RkM9C2OY3a8kZCOp461++rPy1zPo
SAETfHCfL8m4gsnqWSrkXAn+NCC8ToyBED2dTbxTj3Nw1yhc8YfZXzdfEHdT3vj3NrxiLKM7t2yD
WB6y+RgFtGpbz8kY8Qdnq6f1kJbnMflHS/xTJ1OVpnwYa1g+qK8ZdkgpTe+WXDGx3/qEUNSRfA/U
hLx9p7AeUZB63Jyq9/9VcEUbUZYVzv1NzdvR2z2xyhQmabIY/Oruc/Lxw2yC6KCXO4cnfkp7C/IJ
Z6pUGEQZwd4XSHKAhPagWwiiHxMqwQDuNqXsqaxynxrchhK6iRgnZx5fx9s+4hQ0v4VIlGDHbmy2
QH94DCA2arPGkGf+qAXYagMDB/sd51ME0wBcGF07+2Nh3yI+MBln14cWMk12BpwmTkyAltCE11pV
Xeo7OqkJLV5m/VyKIqF5pl75fjD9tEyfI8w1dJkE+6hoK2OvYvLDZX/BRk41HRGsjQ4HBHh9mf3C
xjB9PpSNYhU8Y8k/CEbxTWkv/k802HblCcrJuScDpSun37pR5xDJ1zXx/o+tg40XXtKRUkrPhdny
Szr13sG+OHgAa7n3ZjaN85x1X1cXZvbJzVqth8lZc+0AQA9GtIAWzFWB00Wv9/R4DnGDKI/zWpyq
v608VYQCqHah7uM6FHgAsDDE6MumzidBrvtnJ2n92kBnS2vMnP0Sfu0Z1xspIafDgt9wO0ETSiiu
Ncq7JaF25PyiO8uHc4q3HfJ5xDZQhTbhNI1wEuW0cYP6w7fo83nJdgEV9Ld0FxBH6iQNuTusp4UG
rDnSOe9DUFfmfJx+6vHaWu82T2IdPl+Rpp/9EhiGhMw7Uuu4jv7eJCEyj18IBuDgEIeH3d1zdK/U
uvGu3Wb+91nory8zGa1p0Ll3jYACWXDvK9He0O9+67amtZcGawoMuoE34db8z8v6fUbuMD1z8Gml
T/YFFJYvg9B5HOYlZy2TAHGfj5WxOLQ16CwYmh81X7wZtpLw3YgrhD1o6S4YPgB3yNd17t/OhLCf
QK4Ro3xL33UJl/ysMQ/1LmheXGcX8BXngthLPmHeT9dBBBFzsrqeTjJ7ZAkIqIeOucC1aydKThhn
9Dg1W8TWW+52GVkpHduKHggSZlh5IbF2bQtdgQ8zqlaaWcDM1svtKwvXaB+MDTI1Z3FsZ3IVNiaz
szE840U591+UIKqCVkVMD58Gxco6pJMcIttNRBsKyxENSeZeq211K1qpzIEnhVoT1OqGCFLnDMUw
aKdXmI1M7C5naqv3wNNXLwzeMDUpx8vd2/yx4SCnwcQBSSN7M1WgjSiodji1VSuqoxBYMg+nz5A1
4CD+BrdonksKpNCP9KXWNnSiJcUCtG6ERa7cetv7s0wZM4ZTIRbJDyrSzm+i0LkMtl7eS7z+fRaO
sR/scWW145gZ4gJFgEXSPtjc6J8qoVBnCyvwJpEp0aXr2xwFEKH9yzW9pln1fF4fMeKpvHw+C5K+
gJy8ZVpAfynLNRL59NX0qq9Q1PcS03VM9TiRXRR/4PDxczQnrJ1WcXodLO68RUv1d1keYj9T/sz4
7QryvzRcq6iof2Z+SlYGkFZ9utQmv0xrm3PJ/xUkn5vpZxiybx+x4TD4R4NO7MHUQd9U9t3pZKEx
psDrgygpqjgeoGiWq2tzHjzcsxdqZ6EzGtUcH0OuDUjBdKZJPpWNFt5TFPe7cQvsbVCBnqadNlE1
d5jTb6u7Qe5DKfFYWHPoRGOl1h9IyosJU3aqmN735AGPvGzESzuJGzyiPlXj2Gb4WSzI5CinhQMT
smHovpwWL7QdUxpcU6d3Cy7WSnzHMk+FXZP28kCb07/JCnjLv9m8LOzH38jO/yetl7zGZVdgLY+G
PZzeUzBC7TN6asiZLn+sJ/hIrbBUjvb3gTFUUwxA8LpihkVNiHGHWRia8RPMHEnAR7/XEQcKmd8b
LPbRGB98N3DFlH8sem+R/ARpct7HwSswwTTsvBRNk2dQn9DbKTIqX1z+E8NTGgSqe/psRih+PTUQ
J1jQlb9cEI4vWLxiQua6PcpfYVVKPqteFi6n9pWtivZaZAC3Ga7zRp1g0LCYgM/RPah3hf9Jgspn
KdkXG1ur6QjIfUs6VBs4BISHtDGR/y16I6kJyEFvqcR+Z9HtyaNNHrGXm0OsbZG+R2qhFp6n+VGp
YaqFhjg5xfqrqF4HCRIWYWbkmhqcg5VcrRLZF+rmh1ViYsHtljWZxUa/Fs+o0guUBm8KAYkIVwai
oIO5dC8AI3n+gspXBK/UlGzaDxWZxLNOlVZcaR793jOWGphwfePMJAiDwcQb95Sw2CUMmNEoOYL+
Vnn83ZUVfoYWICpVrqfyiB3qYZVZV9bvJ7w8sip79sMBZrHdqtQmoTmZPu3fRTXEM+VTq/IlkjxK
IhhLgPAw+iqKaJ5so6BQXZIEYEfYHr5uUgdqXfCPBPXoE3KRQGQg7RjBsXNSq5Fom/nxyG6twAwQ
6Bx0DHX9MpxRFLt5a2utKYVu4Z9HKJYlfbQpqiBKxplNacSXU/SoJbzSFJ2Eo23GddLZdQLhnb8+
vYddJEaPCEK5/5Hs6DLplWMFFnpJnRcu2hmGSBnN/K587pSRpmUPqXw3k5kljuBLY7FXqJYSx2Gb
x2XFTpmMp9r+u4+v8OkVHX3TQGajZ+UO6dpI81xq7zCENle/IvOjS407oQbRrOhxenNDPi0fx42n
L6Tt7ZgHSshiOOkMv93y67x4s/k4e/fx1ofQLfyhj+BVmpq/guTGx2SLcI1dcf9zgEz76MTo+Q9p
2syJm87GDALaXSv0v9xIsnBN0vZ2OagnQwI88O1lXHNgGBocSmHsMgYQXy6dTj3MU5rnFt4NiAVw
JgC5y+ug5gH35qfRZ3QNRM4oVz6h8f6yOKKqmRZmAJQzSU2GVnJONRBQ67IbCLl46j0gVKBNFGAs
07p/0SmGl62KHEQgfaKJka5y/T+DeQz/QnbpxsKS3O3Mpj9q0Tta8+qwleMay1lXTqIeYBwL7y+7
jHbz1+2g/r78Q8mJcU6czzQNbVy//APl6upjy3kE7lOpCMWvg3/bA6aWJRWi9coyEQ9pgkf2K0Kg
51HlIcsf4vfEc2VGagCseK8QfvyB7eGmMw7D7T7cDrL3fJsjR1ctul9kicDbRp0PXqbCaTZzI6r1
czHBSYsIa7bx9XHBEYmQ6aDMmjRTK9bwoSQzfOKxBl0LiyiUsbqcmPfxlX/eWW07YsyQoqbfZzcF
xQvtNRd3B+gQCmOh3NPblM0s8A6v/i3fZFAc0sQ1KUk5QlxGjhITrI7UMrYmT+tAqHBG9OeCG25d
/wJr4FYWE7JBwGlOMCORAH/V+ja0HYP8Dv2xd25XTpq0oeLutvQ/xUS8ukG2+nku+BUyT6ulwb2B
H+H7Hij94nK+tuXly3eVk5yKnvK5w3hdpUt8HiSQKlU+ku+ZwbXwwRRuUIFcK59B4XVJIkMZWhTB
E1I+NXUUOoMwOCJ7kHOGyEKHAGtZzYhdq70gKOuS7XbVS7JabeDht+8lngIUL1vmAhtPzGEF6BH3
Njtv3b+KsVtH7jj7vHwOxCZILPRwi6EaqS8xgV/MK7lbafipS+nf4wOiWo+UtNWt0VK2GSB003Lz
7gphWKmZaqzmCzD9UzLw8VhZuwrU9q+/5uErYj6I7jzj57VtiZKkYn++P4DiDR5ZtksPLWmRrgUJ
x+hrpIKr2atoGVh5oZhwkMk1iJpCsSY9/2tGV4SDZpy5JkdB5tTegHJu6n6isLBwFuG8oQ8u+P16
jyxpsiJd6hpNmA8+KoRq7Mup5SUkV0+o9iiw19KVcIVWQi2V0QbDgC5b540DLXC7w8i064+y31e4
PTBgHnTHe5BqySxOrShV6wGUCs2Bg5DG4stFbJw8+Pvp1NSFi2kdgQWCTLYv+AO7EIPC+3pu4Khx
QCZO7vPXqL5J+hdJGzaE4Aki25dY741vFXJURarxdBiKpp7aUW5yshMn4mlNWcLIUFuYeZtZ9mvl
/6dmhyG37yp0l8P82taSU3BMsssoOum5CVcp0E59XqeU95bcWoZskOuwdEySUSrhuVkkeHy4x6k3
c1U3fCrEBiv6ICBYU1V6Efh/aDZJRKSvUvWC/VT7wyQvCiU/ywzJU++d5XV6K7inj13vsxa7zHtY
BrxJXyqsFKI1rsIrSF01WWDAI2Jaqq6Y4aKG1ZJxaM9GRtoPixBbrIpBYVn41TZzNhIT82lU/5Jc
T7Im1myNUZjKrto1Ve7rrNrXKCgKGTZtRilWoYFUECLKh5NAzQHK6V7LvVxe/oSgCJtbFb2LdqrY
KAO/NO+LWfW+E4059ESvNMNWKHRn6653wSqfGLJki/zTb0bgqVXQXRHHmMc7yQz9Jjz24Yyj+3lB
S8Yxk03MLxsXdBk3IQYSMcVwWKPTCkPEXqPXkte3ev7aDiGil5ixSgbDboKiU7d/l/4I81WUBvKn
IomLl2GM7jAyQfa0cwJXYNzlZTmceE1z06nEqplWbWUv+P4aW8ybK/qriThJoYYh4AEzKdMPv1iH
augknoA9hAdBcLzRlb/C9Kwo1NLF66YTQ5QONvWTcY34MRZAyXcXjMDSIjrmnYAHOSImsmXtTCX2
TlG0MWEGd76n2vQpCKsnuWVghGSkiECY3nAriQnCaeBpVminuQWRBQYmakzwIS2QaksojnMP0zOj
l7+qq2nRokgslPsxRvZb6SqrYiKfv2lqadsOXBrpNAnlJLYNXINSZKKqnUQwoKnv/Lun1Zhn1r7b
q8Ip+zcuSO9v7CERVPgD/Rek4rXiSueBZ7/KxszyAb2U7d0h2jzEJqTBIhN4nmY8An3deFMMDUb0
yw7knMRrspLBez3+MCaPiiI4IRXDSgM8ZxdpcaS6A0iKfxL7YhsKjnC7c5akVtS8y/+NVfPqP0pM
40Rapkxj+xku2MreE5DN2B/VD443uyZuN3IGrER9/o62DY9HVYZFkvOp19x7QgkcHaSRv9ey2Ghk
pVaXgyXdiAiewCfT/9B8jN7znNomUgIU1FLW4YpJDWyE3537u+6ijxyV3KbJ0RFe+f9XGli3Avc2
RFkBFxns53Jg9HoUR3A8lOuAQQJdI51W2xRXZS+Ez0w1Vi9l9iF2HX0SaD5WSixeklPKgtJhUOuD
VkAkNiNX0QuuySewLr1JtMnFrHCaj/t98PZ8Cx1YaxKaHYYtFbz+RssNcPqCVM72cte7yMuxhIlK
gyUn5ZDq75q9QP5uQhMVfhAMQLZ1k4uc7Zvb1HHkYi/+7XVohE2b4UuWbTSrnt9XVsMTnJPxkj/u
ziAegygQqVC3mu5I7wWeHJiUcsiOr5EwcM+fQZx7IiP5S/Q5aF5+fzMYZKiBbzsANAxLJ4UzsyNQ
ByvisPdgdYNBdrjjVKJVFw0C89UseWG3Ky4wDWx0mb2UZZQ9f/paQziVMV3mA0sFxuur5PQAWUDn
Wqek1NKg05vMcYS0ZzU47eW4Pyz84P3mqHJzgvOSL/g4Da8s5D3CDmRKznbBgjnaIE5jCUyl0JNc
U4l09tZA9AoUemYhtyl/OCrTp7gc3XBts48c6SKUhg7hpaJY50x5ZukvSPC3GD81hOZF5GyK4U1m
fjhYJRqzhW1z+/TedpojVv3W67byD/v8PGr8x7XATvfYpa77hC685Yo3q1bWhv5Yc287buRu4hCZ
QtyP7fjPUJtUabkxbz0QkydWzhsN/Z5ocB+RrKNWRVNC+XEZtJNLC64Rwajqjttfylk20c1t1fzY
iJrQ897UahlW59FadOqNiPfbOEr4CuSB+bH1vKtWeon8A4JcOJQkvJJyfB+sLXi/3iIJ8GYnbCb/
eMmQkmSgDHN70fJlWcsgk7PW7UGyWytWfXnogO5JFOZw5XrGjsz08eFxRePu/yUjp8/wHCYcgXXW
9rzeskbgMMf6qCTSRcJI+pHluId+ZH2WWjwUPJH0diQXoaueX0idD1io71wZVAHfik1D15T8DKAm
OesnB8iWLU5OD20Q/E6w5Y9oIsY5zbxBTgQprytzS1wAoPsULXdlIzsH9BBqIbr180HQ1eeP3cdb
I2q1yOGbo3V65WSlgc697tdCOcedJmTBfVQw2xB9V7rP6KVjU5HtjxuF7wf6Q+XCw2Edb0CXlzXO
YYHVSFKHvx29UpZj9+QJIYzDf3zak4wsqXaodajRfQqrKP5+VJls4N26Lb2BHWIvsCc4i1dmLPlP
oJueyKmWuxl2X3goAJLJGc0Vau9JITTQoXaeGOwB+Lt+m0FxwOW1/mvnM4FNDtQ57/kTgvUemVOz
FjJLuYpVEARuiftD4ihl1ejMQNy7GUOLHwLUhXMZpqIy0iqlC5pHY+WFbReHkNpqyzgEGK23Nj7k
raAV6rhGqmczd1mHtD7bRBau6StDeH0M13Or4rkqJtEqbuhxvFLJq/B7yJUGPxqihWmwZCCJf/hQ
s0S9SmyESLBNMuFSmQ9NN2yWkP0npKFEuhXT/gVWXgsIEYxesoRT0OTtg3gp3gAQ8ootFh8vg2gA
1Z44fUGjdKM08dguZCM7DByMuibpPPNnJ0p0frOph/B/RWbtnZkHiXeXSZfj+x17VbcGICaiDcyd
0VmuhdchuKkR5B7chixQHeu7bHoHOow29fkj1EuzZgTqPI8tcHIeR1TKu4wzQAzFLm+Y7/+YKl2o
7qFW5Vx8sLG9DtFLodliUh/9EJhwzQ2RMeC7Qfgd2sP2NFGGBDCT1y50xjIVxb4GZ0slsssbNu5c
CM2pXUihWYuI9UsSU222vDhH+FUznA3dq+W1u6Qy0IKJWy4a4tIqsZYUsxAYbEJhXwe5PmeKa6DD
4Pkd6AnLxphw3flZQQn9LYfid7F+5hKqk9uRjFuH3EzAbn+bQ6B05GVEfZ1ZIoEP5rtpBd1anLqE
LbH3V/sH9SmXl4TyHQh+UycYBci5e/tcvbCr6F5Er8cqTkGaz8ulYfe6lWY1DnHtgm3OHvhtrTUV
NQ/VnXtlTCDw8ooqmTGHFGo+Bew0YXf3vp5qdyEGZEJ08+6Cifb9lJFEOdIkY+cATqvatKttq32T
C/wK2jDAfEdn2e1uG7yPJgGzGzHdKdL9jn8HmFQxtxjCMSZdG8K37I6wiLXPNdtoNhm03yCy7EE/
hrykmd3n/xK8hLr24MxN5lVcTrZTJG8TjBhxzo6joe+YaB40KzppFNoYex09aWvGeQsqIpHk2yHH
/poTEVeOjkp91Le1GPG5hq+TZF2ip+Ow9Oy5t0AZlIkwe7VHXOnT5e6siUtVh71N+AbeOoiuVp31
bP+N8iL1cmW0P8T+3jKOxdbOiBNU6m8rSDA2grFTdyitEU8jcM4y66YoFABbR8oeqmroNwycgbEO
6eq0LxxH7UNW0Z+v/8dCtEoeZ/VusOSKjzN1iVhfMEpU3UxbediFIy4TOTIGnOnSAf1/MZRBvp6I
nbHcfT/qmsYsSoxjIMC4EshBn0AVuW3GyKuwNttA3Ca0CAhTEGCUkUqOjo012HMes2I4RMwoYgl5
w40TD+cZT7EUW+ed+OA/71w7CFfQFAudMvOJqN1b4Aun8DLaqgurdCOBcnpvMRPDqYICNNONf4YC
WjCJXUMk+4JsZK69uS5gLCuNBo/6ZwsDSd1XfXGwtvSPLKCk3a5FvjzYpVMNOGkAEQTCC+MeCbwh
nFSOE0hLCGoM1PiwrjOZn27stFLi7lt1VOlSzMM60L5Hu9LbUhOxkqJ9s9HoBij97CjmRI1YVh7e
BLGzXMsARzADmw9LNpPIQcGsTMJ79vNkqFV71mmo9wfKjs68sJMWhnTIIt57doXIGwNqGojdx6nM
xk9PfaGOJ4Ej32M049joBWdnmRUoX7ij24gFgrrJX7Iyv7+hvbbyayubcrKioaEZNU7XsAMX/tPi
G2LNWBJL824QVQnJzHwMvhJpvlyW9omz+GVP83shYRgtMKOXbNOFcGsnfgkWpUCwErxYczL63JPW
bil8qxeSECzeuhhmlskkK8SW8kNLYeBPJnonLBM7UEe++ZgY9HAKbqh7lP5ABHufcvv6CNF2I6NT
dX3o0mtqgRF54YKeoQyQ3Vwnngp2l4u8jN8IQ+MMiIxtieG3JdJSmP3mufswLdFnGIO4lDn1b04+
XRbBqieatQwXJWpLjJH5Fv+wqh3bXA7Yjvrxd3iRWBYDIKGEXUVVFqjscPDyvpVKgb7MVCLgAmZs
4rr+HQ2PGMfCpnm37sz60DHf32IIptZUxNPCCBkCAGYsaZLoZY8JyDVMJaSthKhCQ5sR8nmzt7FP
YX552wXOcMJLZmzM5AObG6o2J59zNp2FE7b7lJmMWk7Ccg54hWbJjS9eRu78vCclp70WIGs3t8pz
PnY1NWCWvwFoewoGwImk/GIuxJqpcH+bH81i3dX168w8nDHkqMabxlfAZpvlYSdGx02TO75GfK7n
PsqebGeokGtv5MEN2SthSGQq6p27wdAjCd9lPBgRcjPPzRNcHkM1OB5RYILppVwuCPU06n92sb+s
GoqSBHtOmUuUgLNOQojHbI2thId/cK34gKcYQPX4eqXFfD3o1R/jJrYL7kim/AWZnHznaninwszS
ZnfTM8pgEPw3nPYow8u1RRckQLNkiL5I+fnMChFrt9oaFBgf/wxpc++ttLvB2Q4erYj6OPS5wNHW
Z4Bdhp1gq3IzvNJ8t4ej3P/DBlNUxKPRsPvpCsE3PMN9LQkDnxZsuBsTR8LkmGvX1tXsPvBelyo8
vs/j7IYtUTCmXhjP6PhOJw81+YvgksczqbhQtcl8oQAbNYXju4P8f391XdrJldLPmVFqBxIm1y+g
tDQSswME9wNryTE1IRGz9J+GhDiD6QzP6CXDi6k8jgfB3Sm0wvJb+q/Umk5qDnmitVl6EdPSI7ZR
0N8Q0tPt//6w70dcLOmh0pKTB/52rVpfNxknOlowDBBdqobFrW3tCjNsOabVhz2dn2edsT2dlNrR
74EtCB4UCE7ZuCTgA0BPxVKw8+DUSf0gO+SPCBAXpvxHcE7qSY88W/ltXcfWOjulDu9gB3wZfBkY
6arU71e0KjmUFKhWCGqDgPl6uns0FsEUwg0Kjm8NYjCtOrH5etEDZH1ju84BFEW6aLyKOpKXK7VF
CtkzVw1O+qxOV/rhu6CvrZ4pCPvuyZpg1pdKfvxn3v7XV7btIRGfkGS46zxASvKp/O644MMpI6Zh
brtCTmaIVCLpV0nOKSSBqAA8Xf9iB+FBI7r/NkEXA4jGDgbOM0znuL8akxJisCib4umjvqhdNcGH
RtK83I1TsLfS5g7235/yc2b0eCczz76EEpEwn0/wWr3/D5FB98HjuPZpnpnMalLEENhynSG5ecl/
LRDdkSD4JehIIXcetIe8cLQQSfLZcje5xpyi9rx+QBO7BpNqS+NU7QiyUxLqp+H79kpOz/bqNKXA
t4i0QlJwGmyWF6zKAUJYKAr1nSl0rmkcAVtSUHN9RKl8nbzCJd+eK/uFe3n0ErADJasyG3ZQtryW
p2AEz9puySiKiUKzMK5PMXwsAoWAK1/k20kgdkHSFps/geqcTkMgt+FCWhZs6FJ8wBxlXeZNqMf7
D6jHfI/KPl5UX5ZYpRn5Rlt4tm7B/CUcc9lVTY+T/H73UtLLR4ZRGjOvA+d+ez1+4XFDuiSOTmhg
pWmy6oFB800THV8vyzUWSLqybMrhknogLAO+MrkAKwoWisYJvea7vSR1IDMQhm/1GjHdkVDnjgvQ
oUX36ogBEVYID3/PcpN2l/I4P8UC25yRD6fHbOiSZy35JwR8ZuTHg/Y4uzBJQhRTvMZue/pCxn4Y
SXYBeUNca3VvbXjTMMdzl0+5F12TfOnjS9gyRskzNfOCR/GX/cuk5xsBoBh6j7dv/VN1w1apEuhJ
2y1N7UdURC4XJ5UmKL8MSVL8WmB8FBL+7ac8D/5Aia4AWWR2GimXpyppxm3tUQ7YLbyZTySxkhDn
Yxa2meA3WVWeBeslNt83g6BJFyDOCCon7CVCOol31MR4qP9yNjlQ2kn2OxD20Letu34muCHaKQSP
7BOg0g8/IszbViH6d3iuXjAuuVkB3BBM63VShQo56R3aWJKRJ07k5nclILNKOUWPi/Drblq5C6ag
JRCU+/V6g1SGnzl+L4jD972FBdIT9v86X5vovxzK5kP7I8JTO3+/6+7vXvjvWsP4b39Xi/lzc02R
GplS8A1VEzyHVw0ryOlbjvsoKXQ3u5IpERpKhQz5xDmoYmPm4pWjULed+UFgX/Vs+Fq1GlX3Tq4r
/NMQzulDmqmRmBsUa3ND654PVK0wElUZu1qkUpr4shaMJbMojD2N+sP662lDdf9af1+WAcJbpANi
/Nm1ZZXG91SEMN/3s0nzC/NOdl4XbKid0qxcoXqlMcjr2TfpMSk95TrrFHpPXnFLU4UlaFhbaTWz
25Axh3tgm6WX33jTKJeGq35l1/YHxlyl+abtH9IPJnsO1tjhEZ2unbaRD0riMnoP1mCS7B5b1iP7
89K/S6PiZu+4PVt62nqBOCK+E0bWOZxBAhpQOuof2S7KS1A4x2tMisUGkiTIWZyiRIOv0IWJjI++
A1k/9KQb/8Mzm0uicvMCs2y0qSVRP5FWVtEsaDiBa1GfBaDqTzwSrVcvAshH9Q1cvICz4vJPAwUm
YBNuTU6EjJJLqNkyggeD8Kg/poZs800hlsyua8wWGv7507Lg+zs2uI4bHqNBdOQe2hnc25sY3epH
PD1A2pJeZYMVx2g1u1cQijNxqd0rNRIavcePeYqSzo1mi7UcOsuSN/Ng3jO138ern1xsB6EvjSDY
ZyhK0EYNI44JoSdkDrF259fNaaHQPdE5yXe3oM+sU6wBMqnkWJARL749Dh1+VfP/Olj/4hJXxWL/
dBMHHvJy61CksW8M3UREf3ZUg5ZBJaDcYlcx5XqpW6ScpegESfRdZ6E6mRr+YW86jqI/WE4gPOTP
RNww8GkyZopWA/7lh+Rw+HV6eoHyBVl1MEJkY/gCYnuEycHh76DrS+ZVecNduQFQh90amjs87HJ3
Gq1AkTuy4BtUKlQBkXhY0iuYPEoswuPto09Tw8hq5MvyjcB3xLK2PoJkeqUh8wqVmCgkXzWDfEGK
6Z8/PEtcBp1dAkhRZfxp88SIXUEs2LeWg4aSjgZA4fGtcf6j6VXnu6YxjQAvaANowmVjgk+akq9V
OPpy31H1Y7pKmWvupjvO9bB7hg1gTgD8y2zOOqnv3zQDCI6o7iPMdWd+udR9z08uQduYzEANg2Ar
eGeZ2zbUZB+RaW35hRuvQOl8Yo7Nywacf+Bad6RxGN0Oi9pHPhaf5ozruwQeSn3iMDhXe7JEWViH
ozYcWaIiUD25/nCvBvxQeLN45GgL/sTvI/qaPAJMdL7uGeYXNpnHXcNe9pXNH1DuCSzUw9AT7puf
bZos9OrgoULzRlpp49VeSoGAfn+rYPIlGq00gUzdXELeJcMdGQwhS2GRk0jxSOphKKx1xAgkxQek
LTAITveQx5UTrk2ZnPI7+A2XrmdWvYXa+l2D5S/o4Nep7Mn+8YW9NXmT43lLAQ4/azjC6/Bf8RpJ
dAnrsHw4iLpoOT3FKlU7syHkQx27sYEnLPTqP6Yp/jYRuWXsxsmhyaClRi2RurfZ8bATs+snVoKA
jJ8EYVnwOQS7amkMaynFAkuN5S+aq7XpaBu1eNDQh1+fM54xMYBa77IfTWAGq9OhDl1oyw+t3wSN
H4q65LcKN1IIdXcistKEBPoCk45TuXqEIrchJmcN8sDITHfaaK0fRSO8Co2CMTWlJHkPMP7kSU0+
Dx05AwKUSulsEw87MHYBuChJ11FPNGnTg8oaUz2eI0MP+6kKDUYjy7D5Foo1EMQBIjcp4SGtgeSi
qjEiZhNKSi3mD9Sfylm5jT05HenH+bRmP50C6PU5EpMCxWjS/Xfeur5z3Bpl38MJ9nRq7GDeYkjp
1PFsx8DRZ6oYT4wXSQddYato4lB/jdNXamIorZpk2kEVVnuqawwDGzDNScEf82Anc62oJhWMdup0
PVS2CpW+A2YR+aTcf2XmD2+risLb+xbHoSKSnTGA5Mm2WkU+Q72wkZ7ZXxaWZ+uPBzmxIUYckEW7
uFZuAGjYL9g4+cN4JELccmvy9G4DNfJdF5k7wDjd7ChqW8NYD2sqp2s0GRadrhkIqyEwXV1tbe2g
ZtZGODLNyk0NEzTg2KUsKkU3VE2cO1v+JnIoVUXCYGW6r/KtPCQVNW+j+OiuLWBSu2RKXLss1J8Q
D1pjvE8rhZ9LnsNZxY9/Op9w+Zg3k7KL9kCwNVUGjyHYg25d/O5B8S/qXUQliX24DIIG9jQqxUpN
4XfvhfNblvazloYwuqy3NC2807Gmh50cKFwfAaX1EtlXCu6+s0K+Os5h22KwTyj+g4IN1EHCHQ2z
9edcMRAwUrtUZAmLg1pKdav0nrhMvn8e7T0HChyBszfX5dda7gicHsaTIUv2s1lwuTXRxk5jPTtH
mDJZmgBAuDfr53lbdBde4sX99UV7TwZbjlijwwre9AWn8mZZnBGOGZawPHTwJGrHDYw5zIEHWS3q
wIcyMJ9qBc3a5MGjq6OcQnWrOFSU81+TzO+zAyOrZl35l9HblotpqAG8fRLq6SvgYFSJEC4KQWQi
OHNU+7gLq914ZIRO+dIgLjHcjfuAi5ZpDfBHu6lyOZkIew5IK680YyFiQT/9GdCXi9ndDt0nO/DT
PnaKInID88mXujFnAv05orvHx6LX8WtyebRhBoT/4IJNzVaoWLbf+PntDyftLHeNSwbH/TqE0WiI
3sVzs1Q2AndS/Dyc9j9+0H3ZmfrT3vzQO8IcNjhxWrksNG6nEOVgxabnTtouFOBvj1tNG6gWzWpt
KqpZodgwnkQMOJ1hNBrZCUXAD9MXaWpYRlLlbPgbT4PzMt0AkEb1bOUpEFviqJ/TfJcQGkZQ2sI1
SuDBqx1V5NrWSjHbBBiQXMR6penitCq98VSYDqU8BHEOfNxeu3v8YxV1sJjSyHfS4/vG8TQMzbFu
rp5OF9V12guT+xJTF7teaQiCkYjHaFRYoF87RafiGtc7Nrr3hafIPIXgMUERIIvOxcyTGV7v4Rpx
Sz/tU0QBItj6GW4TGjS7ejc6ropOq707bryDvvf2WkTIS/L8dSNevcBq2joQAzss1h6uTgSrjM+O
FM8DW+z6nvIqNEGzQPP0xszZK2X6vYHXlCD7EtNRhdlYchOz2kf42N+B3ZKQJeuZZ2atTHKMth4P
W3IlqopJR29Volg2knO4rAQJaQse3EOSwvrC6J3YEiW7No2oHKgg0Fs6RmjT30jXF0FR4PGox9cM
B4h+ATqYVPwPwFdWEShMGy65T1gwMTQS+MISx5gSIy3nWoHITtLxw8a2M4p0qgpX27xwbjc5Z/qC
/tFqKcDpazCSeSL7Yz2RXke+yqvVlbX++t0o9xrkLqnQPi0TbxP+InKEsvugzbGw04g9TKQGvbWA
ufgSa1Ieo4e6TjyR5d1p9qxILsk0jYG2+LwJs+orgRkwIuyAVT1Zh3BQu+3m+8pGut9Pr/K6d+hi
uz946Jr56aYoSWwvIHXejGZIAEYOKtYvI6oayVA1Y9OvCePAOnrl2XXrpt3gXzPooqj645/mIaca
y59b4SfQE4bAZ26zDWx0E4IrIYbJICYodjoZ1xyi1VYbJXJuQC7i/IiD1NFB1jAITd9tc6Qg7C1L
ZKfWvCCjzQYOvRXt2ZyO7adTRq6KLSHoDRs5VoALd1HxON8wTiCgthgjHSz8Yk9wHAuoWF1soFF6
6OIcmLh1/CdPmz7/Hq5aFgnqbaOt47OKspUbKjCGyN8lYolXY8WCwLDwRybLDNEIMfz4KwESl+r2
p6ULXU4bhGWlrHH2cJSyEPAS0DcZRvimB8oaS6JpT2dO2iQzMzG8GpqtnApXpkNQwT4tHu41sgUw
/gdR7TRQ5WKkSOkT74drgXvJM4EI8K9dt/LGa9e9mUkSl2I8CDCLH5kceSYV78KT8Bln3tEUw05/
SPG5/d1MO71iBXjIo41yd3O5eDAN4ZVQsiEnn8mMJmL4DvD5pNWAW77sKA7/vpag7tf+FZ7oECqe
Fq9ZEg9GGdiuiwz2UcqRyOenJZQsTm6D0g1yZJT7W1s1x0UviwWmOrxSsBdhA3sxawxO1foWnD47
5JkXXsH+DtNmECu4H1li7BJorjW/G+sxvfPLmG3kq6gpn6t0YOBUw2h2HW70AcA88D36c0uQoZeB
GQyu9/lr9ay1v7hfof/rglv6wAKCdLYFEI+esVp0/vWnbsoa7MBHNZ5XGI3N/2RwVtocjxZ6GJNo
gEvVU3BzJPTnvK24NbKXjIJa6dwYyikOIp9j7dS1Ae+AG45GDk88AuzobTvhAH0X4eW2ZC5GPL52
innLPqN+sKqEhcNKZVMAcaIiZe5mrnoI5L84iBsSLqvJYIHBvczPjVw0BOsKLMlocnZ/VN0yT9Yc
IhefwYrPCHs6UMv4bfUp/YGR4NAKdZyxgtour/Tr2wq5UoggPG4AxYVZ7KR46LvhOyXuUQFu6QKM
lvF1524QLFRUYDuI1osD7l87NCxUNEU6drFrkpT/Mar1IAhrsmlvdxl/BK5kWVi2dvyKQqFzz61o
GzhrBQkvAEQfYl6fkYU71WMeKqebLRvgaHv6Ao6n2/MNRroZZYiXbRQmwDNDT0gG2WF0TJc2ZuF6
ODwNc7pg/YyOeZvYcyOR5zoJNYLeHk9s8bwVYnaXE6j7kgkMxTw/h62xFnVyXv2Jb9u93dJxMl/B
SKn09FglWjUoOPFvJvs9Zo48+/e0AvheS3avekePBOeGAhDVaEtjOe7UcRHPHQt5jbef8UrX4Zz7
MoBF88riWYd17pJ/vRFlWyLqtcz1hf90ov2M5vQ7PuIZvxyntM2mZeHQeHxrJSXfLMgHW+qqCgDA
WPu/2xt0IUi1A+OxMHMqWK8XeFMLtIHu7RVeORy2nMS19JcTbbez194oG2xoGVn+KLCy+Otxh0lX
oE/W4+Zpq3WLzskwvx1Fe335ldsutFTQDsqlfoCVBvmc8qdXnciqRwGWUZWYQb6orIExnjWbER4g
PxtKJ9ounygg+f+vdlY5Du72DIcYYye9HIzZR2gPXW6HgkhbW9JGobibjzeSq+4doOEqRoYceQL7
4l13Zw/jkmLie1lJs6oGARz+QKXqhtMbXy25Hh+098dC1QivlZmsozJTdX+WIshtXvzePIR5NCme
gdaIdAGgUd+z7qxyiWMY4vNco+doPHlwCnjwzT7Y/zs/sLULfLyIXUJGj2QxFdLhYyD7aZ3F/0qq
PbfhbgIJULpdWEe//Ko2MV6kjCItotnhnCqE0+cnF1gCVtHxRAUmuK8Q+6RYB4xecz8QxBJckXtY
dqZdCeCr4zLaU9vJtmhu1tWgkOkg9SVHWcnW74TS0lEe+GrtNQu/H0M/VNqXHvUuRjUiFey7Wm7G
yO4ISKmApqBBgbR45PpoegNZKrHwLGY6ZAHIOb0vkMN9TIE5LbNUSnEJeygHMqfS+tFvniRDJ4kT
U/ZuHsK4FB4V4l7vtsWthNB6pFRiXpCCcVtwOVQikHK31s5K5aa2yAHQXdpR1+jdwzN0NQsXexVT
4VCD5Tx+mdib2yWw5hubF6IlTCpEwbQQJXasPMPYb5ZA50XVVnd24fmMnbBVjkFnYyJ1eQAcwYkt
5uC5hRb3VMrU/mpN7ZkSW7N5K+f+eIrUxiliFhQtwLKL19Wm4soptROUdBvaTb4iXI7od9hw01aQ
YfNh5pihZc4yW1O+JQOhxBADteVoKckXkkbXTUOttD7phKQ44ME7+luJ76s8krNet09OI59QRzrJ
VCRvRrVVBgXVixSLTHPoZlP19mV6NMEm3DJwaKEMi9jB/UvgsNnQeRob3biNhouCeVQLGqYhwx87
ixyYthbN1MGUJvjXReRmwNiTL34UxRtj9Y1IZIIghI3ny4XxleB59tHSBYO52jKHRpnxmDX2TT81
ZVlkmn+lSC8VscgW4JAh2YoR2rXxqCRQeqnt37UIgp6XkWjYJR9npveA5ec4bg50pgBZyQzMZ7zL
NRIHtvxMh3rxAgI71UMSLgtsiG8ykc0NzmtGZNIT9QIY2Om8PrSGUfYTTi5N6mBswZkWpqE5NPUj
kQItqYtGWxgyVVBRmQphCwcVrgxwcCzx3ZgAqPUpHMF+jjIHCRzByPk65zzv0PFULm81XPxMf1K8
uhi39Z7RIdebgpMdPncD6AGEtAB8Z1IOi9+sFSWl+jFnx4bhusLbP0M9mR+ZdFO3byfASrloIJqQ
6fuMlds1FK8hs5Nzi3GmDKWE4NCLl8cgMSxUWr4LxhYiuhFeD5Ef1bEv8SEsbWAtNqt0NaseHM73
k+hZ5QUy5EFOaxZE06Fakcfpyd+Uq5jLb8t0Le7HHX0OfLDWihMWgbLk/FjkLMdZBArptylGRUau
lajoI32lXDHBS7vKAHDzxJuLhjME38GEw8m3kLe9WK2fC5NYMa4+txZzI8Kwd/vfIHfZ9Bx/WYyC
QWcra4GiG0iHzk2O77Q3QXogMB0nhDCS32Uo5mPNn3WeKQZravGmV/c3hFrcYq/H2tEmZuP1hzyo
tik63Ux8mCllk/ruJlkFT1Q9Y0Z1nfekMKAtcLFo2F5RadocrXUg2yuzloAwjAiUwENU5xcIl7vs
YK/WIR0GY35imDvAAa5RnIENoMOHpMyPAoDfDIsVamz7smYFhXMdg58392XVfZ1oV9QQ6mxTbxJ5
SD3WzBzUrqz6TT0NTCvCxWTEssgA9iTTLb++Jowl8RCGa3XdPNsicGf+9FgH8pxSo6OWrQrgNAmA
ltlXfcNCGMZPpaNG5y1D+SSOHqSIogUZuWu//esegV9GCw52BTp2RXem1j46QXm2/b1pExDb//Jl
dsGNphtJxuA8FrBX6O5POieZiFfVsuLe8z2yznZdd8LKVCz/R1eSha1yolEiCSwqu0P99WlACHgJ
pryAivAraQBB04E5KFx2+KFN2MtUuvTdu9hN79mkWQdifdPgztr4jlXCvrltkw0KQROFx9gC1Nps
cuxd14LjejPf6Hl+fhk/Le1AzbSX8y9qLD3PoWNqgg3MY6Y1rOHZ0ZARvVkBeFr0cz+72SKQ4Tbd
qhr4FbaazxPQDMwssSBF9rZRIrO0pBaxgmOPLNbSBKhKizVkfTwuzpupQlnAh3aMdHqXgITmWdSo
QFV9Uen1y24pE2YQIcmCNsvpjuxROzXRE00WZgjo2UzXymKHoI+iGAaaSxvWjzYhszKIC8fTLrfT
vTyzNsRJm35su/eIQkmZG0jlHWCJYRLSi587KCBuiSHP/5I0foESJTys40/vMJUT/T6g0qBrt9PI
NGE0+3ky8EV2sshrKvOEadDj1Hk7QWQ7yl0P0+HjJlEa/1rj82EV6I6KJLPpNtTqpJ3moeZRI/5L
B8FQ976PLlqo2/37i0L36mAZVk0pxpRTxgOufzImCowXsh0K0dlgBIE4vQ+TQYpFXBXa4jvLMrux
SyDUj0XiLlrnfiAyyP/hMCbAx9xlur3XG2LY0IC/nQ3jFb0HqXN9rOUMn7YBacneCW6uaaPLmirX
WScFSxIEwqnSx2iUnKo8BL0p4CrPNsN+krwc/DqgIDbeUy86JjgBWP5hrRFpYRYmKQarHMGbaafP
1nlGxM+BZqICZHM160MkHBBPg3cKli9xLboPwWm0soonFnE3yM0CkVTU6ma96vBLv6uxjj6QAAeW
LkbCW56CqXAj2hXO7duQsY1QGmEHOpKopiIR7/5HzcXcuGW4eQ5eyPys5i4qw6KQtiM1rJ2o0FwN
Eoohi0alrxL7899i1K7d3d1PnWEXeVmrJgM3wOVb7TrKhHUwcSdQHFh5I8kWdihuqWN6v7Jt0Wzn
+UFrHxJX4tFUuYIJwrYA0ES3kaE8Fi++E2Sm1lsNiQHDXBeRJ4ziAGIF0hlBVFedtU8oPYl2j+yU
U0tU+9U3v91p8rAC7GNd+tjilGRqgBTCk2MO2omyOrxXngzMAwOyWzXtqs5vjjZzyTF3daQ/HLEu
MxpCJZj7gpqb2CJqu1xOh3iz7JjtXrKmXkKckhbnmT8ea6tXVq5W7nPAry5jodFRcpihuBxtK0Fm
sEW5Ruq2HAxxajuwUQDR+Rgop0udpMYR+HLSxaqZRBEAwrIVqJKfLYM1OAD3VJykqvnjUbq8vjPl
E1DDryYDE9cTFo+Acn+RSfn4Jbkyru7cRoT85lSIo/iu+TF92IhJtPb7IBIWMwwvA5THgufhxK0i
Vtnpxm8kVTQDH0P35l5HdfG2bptESCatVewSiXZ/vrC6IU2apS3+Vu9gVOKF+Yrf5mAvPvUuFwE9
5jw6ZJMF+F1JGqJBa2oFGFRUy39VKECSV8Pixrg9RpL3tVANnDPxMOkcMs81g588dA5FUJmBSfs8
bgztKjuzk8zCkO8fTqRWakv/BGV3a/YZWETRBsquQv4/Y04Zki+Ae84ahvB0XF4+T1AqFa5UetCw
27VhhUJQ9C8Di/8E3jYB1/nvl6WdxZju863swMnrtib8CGZvwaBudEDlHUWIfZn+gsipDa8d9aCw
kG/drjotl7a2+tFcKcQ3UeCa9dWjoxzwgk+eT6red3YNMxpjW1QOcxBA/JGxo9/VvFQzpmbUYsxX
blx83rKXQoYub5y6O6hQm0UfXTm/w7M319GUnSh5l3WOjav89++6OCZc13mtSSbSV+fr3PnufFM9
6hDbGAdU1oicULXpCrf1dNwCrfPI+mjQG+7A0p4L0K6X46rf0pQXObD9XhZzLKnglMVb8pTx9oGo
laoQommwtkYEtUErNPgg+sdAm3+5olBZ/WNo54J2hTRBO5HZgCLazvanWBXtx7Fa0ByytJSm3aQo
kq17ac5Qk+FxZkSGZgNTdEAljJajOtnwM9yVQ/qb9tsQcJw8uYFMLpFskL3qyxdYFTebT7GmHYEi
nBIxFaYgFbHRn91iOHjEjp1NiS3MbZdtQ7UHwgp0gX7E580HSaOPMAaE8sKD+zmpScUFeYX6tWl5
loZpN+uWmo7/n8iYTE0k3o81L2NwRMJ6wnF2RtSM+hhoodYp0iew8c9WXYy3KuYM+Zz5ftRkS+4n
4C4B0vcSg+LuPFV9EjwtgaiPDjQSme6XUVfTZpmmEd/c4JEnzZelS8mimonO9GFbAGQvv0yLfWUh
LODOaZp6gjp+D2A2aFfeOIIijWu+9FAqawkO2ke5hcjhw6BD0V73vCSOcM8H8+I6CmDaYDzjwZdZ
OdLadGSHXo7dATgKAV6QujxxOMRrB89XLsC8mVPT0wmDPYjJLot7xD6w4fehICvWhjp+/FX2V6CK
wLgJRcM11tqowP87Ohwch2pCBLz0eoZ+322BDQ3fkznf++ha/LC3EFrXnoidHLN+YG/ShL9HhIFF
aIziEMc/2fOIGjILM9dN+SidNl9qUVTE38TvvDTOBw2ThsT+YR/rDPXNQWVdZHQjYGeAmR8yO0+Y
30BKcEeHIk6WU4xk1w/FncaoeyIv/wJONpcST4/UxpMC4SK6GOyuLjm7uKguMpMqhScfILIY7wpf
ri3eUTHVhirDvBu1bUJXJjE8p6x7BkVGx41QuKCK4Kd2Rt8v7k/3xDXA8xXefBegf/3T8ckeD/hC
zproZwPKrUXoIx/d/rnT7LU4JaOFtLZrzbCBuSAGfXjQEnf59FAmRcr9NyHwF25iZugEQxXMKGDN
MBuf47q3PwX+oyegPLPFlqDwXBgAAcEXkxvvUiHk2zBd1hyFqeb/Z8wHXw2Rkw0nVO7VxQnmPjLY
hefSb3obKX5o7GjbZkybAjfd+v4aXPcsYZg3anY1G2aNH8O1rMmxkTMhn6+ZURzx9g20cs7ubg4E
3OdTKLDAbMsJKWDQpEimW2sCftle9VK/ORb0d4KbUVLPKcUCxRTg1ciLTfwgjLKrRXbBRlOIgJuQ
fH3qvPX5EeD/qm9wZFwjnHQG4bT8ty0iRyju7AO7iK1afJLPZcJycatYWY1k6oKze55mttUuAzVG
WDy5UxPvQ0cmPdFzme049MvHRBr5gHCOREQzi3z3zIhvGfd7L39VcRsqtO3rinu82N6OAxOZ0zNe
827SmVtwaUY2nJ2JMDdRkzPzW4JMVXN73wJZBKT7y7cKBAsWk2rc6upKDEJzrkZAFixIm2bhxgt+
HYwidUUfELDRyzkzcu9pXldZYB0Xtmif6U5rCkNJd65VetzqqDS2Ch/ss0Zw8BU2NqNIGeTmrUgu
p+9fCsfrrUIYBAuDSCqukGcaRzn5eNfPnzE1lPKkYeUHyHX+iyAJvX4JybJ9Tyh2b1V++fmXRgyr
y3een+Y20SSnWeJm+aI2n1rwvMIEltBYJ8CiScc1XjJ9nApQYtKz7SNVyp9trS6XGO+PxguoOwhx
bhDdIcPIBu+GwY+pu86J83wly12R7bhkPL9wt1fqSzYcj6AMYFGH5M7Wp1KqGbHUn2ETMp99cmlS
sjg33UylXHby6sUPZuTvfwZrfX/q/WqL2mOlt3XE2qN8Vwo2dGfKYDe390Mx1OrH8XPhYLJ0KZ44
kEvpaAyF3SHbZxG8B61ce2eNYTKCStKy5Az05zWHCzy5PIDS3b+C6AkwyShQeRxw25wqvcJVMpce
gqc8zS7W+/UD4QFF9HD64va+nSdanyaG6uLGinB8+6pUfErb1vS0rGOydilWpd8juy3gQUX7Ozjg
npRcCpKS74RvzCwF4lP9ur/rEWX0SxodJNVMo98mbgvT7ACzal9ZhPQCk3peLlSmQwPxCTTYqZ3T
cHI2FKY3dhssdxS4ANCx+rKn035U16ELhkqJD0LdgU9WXXDtTi5f7nhHQNJ69t/YNULsE9NQ6T+1
YTb6GvHlykj5FIvWDnaUQoYmYFptFjJh8iS/lyarOMGJfJuvAJpAOAr3fDUXRZtNzq8vkyCJISes
eqsWq24bCB9DS3bWzLoy11P7wXlgnOBw5h4dxubkinAOLVRWf5yKtZOQFr1XfhhUDU30dYF1A+jy
z/dwSQ3z0VM3m3pQ3zX604FxwF+4w2Bx3fTrOCxDQo0KOCvgTkycLZZDhX77tQJA4Fu0LqdghXml
AFtADyadBUDUIXR5JxCiO5MbglZfTdUcjGo/6bztLXu7ZLfRlwV5LRPVxGH05Z/0bf005L2zvI/f
xDiMHmZiME8WoC+/hOjABVLyYbj73HbyvzqlyWXuVPi9UnaREfVr4LKQtNh3ej9bqw+H+cwJ1hMG
y1e0YcidcAEmagEee1k96B5SYtZBWz41rNHpdLnPn6f4HAQgtxOtgwRRauym7aUFWW2bIPfkszYp
MY4ELLcc457m7CRgblreYhj1TmE7KqJtjS0nAeYALjTFG1iQXFu9Eih0YzgxjyZvU+02IkdEJg1S
EMUNgsWBrdSmS+wihMBrYbBYdA0iEhYV5+40lkNBZIiGXDfNf4Iwdk0dwyp5c/gdqkONopaTebK3
ZfZwZFUd0LHjoKPGsy439+2KQIZX5Zr1E7JoETT/WtdvVobQUinUbnHRVGELwaZvg7x+zaPlZ2iL
rY3KeELSbnaf0tGsEjoB4LxlBqdgZvuJqYUoz6a93loY42y0/M80sKUFnYGL7XI94TaZA8ZabtjQ
wmbagINVJD3vzDs3iyGbeXxsHK9svCC2m8uYCjIVd1m4Ddt/BBRHZ8H1QNPieAMvk90LUFNMS/ua
DzhMWs7KT3VxbUSPIVM2EVQxyTX9acouLDS4X/HmNfTEw4mDgLlDSTsmFtmDEXJYg7QLnm1+JOGS
a74VvuznlhFp1KWrAQOG/XfT9UeUtUOKfUrzzXo3YDI3y0UznyU41WF42nyrZD/QHF5NbaxRhSls
INZzLjuXGof8CyUArdx595zhUhT6Px3FTAkla01cF89Dt0fDVApu+cuChZrTrEq7dry6IZ0e9Tfc
zX7pizxkZmDlG8DpvAiOgTvpsCpUawgkt/OqU7xfJoh1QTd/a/C891EBi7x/Ku7ly4GtG8t8UTSo
Lfr51IDcy2DK6GKz/tZx+/HId3NTApq4zNnb8nuDYK6gzFgxxrEDbG/d+qpE6gH4HXcuxqzw0TeH
mwUyLL+5qRMTF7Db9vcTOCorfGeyy1ydJeSalpKycDVEQt9gPz6r8Erc2DUWW/yExl7N9azFOunG
KwiiALASE/pay3n7P+/TL5Ne+ChPqG9TArwzKdyKbuQABVCtUJSyPIFC3v1LsTpRmeu0nZnlPLCU
aOYFnj9MPmAEOLenSgMpltb2l9EE7yQkxFtFnIYZmi627KNOks+Uv1FqpfRuGb8+MSTyIRZ/P5gm
nv77jqPhRqvuqX9j+DjGb9zodtntS50/hjHaCTEIpAa0CeweN5SOfx/Vxl9iPYeXP9vklZvbdNme
RUGJ0cfOYT18s/cywRqoKe3tI2WmXR4jdRxIKIAkIDTVSyiJiJtbj0J6cEQMEbMbjJCHHuJNvqWS
u2sw945GFhkY74A9MXS1IiSRoJnQ0pZdG1zQkU8jSgWDUiGUOWmLLv+xgsMfDyKspwIn0/A40rFS
GPPff99SL8QowYoYPUhu8qXzILBprGqJnOIhhNIPaGfHFamXQY1iyY27ZUTtjMxIR4FoI7bAuSE5
o06TV2c7EQ99XNCdaZl2YAGSD4Xd+/9gf81TP0PLULbDsjPu+TC1ODOnzuh8Ge/UTggPbVbrxbDE
HhZYRht9I+1YI/2oenkfcebWBl8xqP3zJ0DrNhC/eJHa2wU3bBgOrnUGfIqBmSKu60xmLrf97f3C
DcVVw0BA/IySVYBGJSyyqiQ8HgIONboKOAqhvSYrdElFaaZ+4ymC/gKGmm5Id2r6vVF0j3fNtx4z
ys0K1cX6WTiw7nvhGiKwRUyCpGieiMKW21JBZxjIcKBeuIVX/A/3JpHY0MJ7dxmNxxDlR6g8qkk+
g0rF7wqxbFfc3/wRemDUOcl1Lx1FYfsAbKAYUckiiqmzsQXTEHutJ9bYNTFNvTB83e5zbYQROQEa
LxbPePF8/qpsQkgVZJTU19wh32cpJnR07LvZnnqIScYhw+1S2FbvrC8F7yD+JBPTQP0Kc7tSuEeC
JAsojLXPauZhi/8vheTTxyaZ/2UCHEIM0qOqRSc+ycr2MR0SW+VW2E/4Y+OKekrMdXps8CJnrUjc
8LEzUUwfLxhQpwswQIxWXs9XM/AhcInW8wz4SKOJQ/WkPBOu53Kiul4O0xxJgILuXdT2eG9h23uW
h9GDFw2CPyu1/ch3aH5Dal56GD1IwkUqHTJQj+5eELWhwwPOjJ742ojN91xr/04nzsoNSFivzbUr
gDaa2ivmU7/TF7Op2ddyMzqv+k6SnoCLJm9qF5fFyKxoTB8TRUGcy4AWw1MY0vOwItl8AkLZA0CR
U0PrrQLMkIOQBK4sWGU+MOeaL6HTwqOnW7RGE0XD313lAgNRzj9cN96Edu7YIXHk4ymzFX7TJBdZ
jctWRBioytgMnMLPb/Lsdw/pfphkFMpwQsdMCD9vvShzhTfKi4KR1g+ef6+N2LfesXF+DLuMR2Bv
ob23MTSM4MQcpi6XL+omyw2dfY5r870BzFnq3gz7GpEPz89tIOGgYCQa38eDEGWVlSqqDNzSpA8e
HweRBp4ab7LnEbQhXVzjYFsn3pe+YgWr0a7b3mBBNPTHfAtyheLJzpWHHqi04yC8mMPUciVJ3vR4
TGQpSRdhUg+YpuMUkNN6TUMDoN26zn8Nk1JFm6asOQxX4VPqacJigDZ8K9JnW8geoxHpsHuO+ebX
KhK83Y5oHMJVOmPEHsDY+GxCUi8ZyEoSp0S0EuLhmZZLg81+uo1norg9pVdeWJY6boov3wZS611/
5XnF0npFWNOhdnprDUWOWIAGW0iuyFW2HFoZbBLEhgmoEve4cC1olQCmszFFKpIU4pehnr7ozUCn
7M8xvn7H6ehx7btHelq/hIjtVylOlOSn1/fLA+SCnL6Sw169bnt+OCBL/wHRHnnQ0QQnorPmhILV
aYuG8JooW2ljRK9l3yrIwvQ/yHNikzzTnrizRqdZsUJQcDlUZp5MLO4bjLDOVVZTcPk0bRl7lU92
QZ7fWR0A1eb0IjGWvb3tYGJhkSr0H/O/+H6IIYngRuzHeLGZW3/pVI+wxhdaUwHrYIXD/gOnXmxZ
HpicN1wWecZvo9tdhb9zWuUjSWVFPzSFh8RYrJ9YS4+CUv4CmDU+SMihfVDWZti7shXL9AGLTEv4
f6KkwSQ5cFyZHbcRSnlYrbm91YjeC93Q5rhkQl3TvuxcAWHupc2naP2bf1bZvtG9ei+itj7RjGyM
5vBmqLREKlhEm9VuQU2+IDDDavIAn6O5/QVovmEeX8r0N/++lRcJ1j1NBr//hHOKObcGz6LNyvGr
eJHnjjO5+QZHMCL7nbfBlbQwu9xkJN8uP+MByFeUS9yVSFqFG9u1KP3LHK5PqPAuM2M68rEqglwJ
fZl7FrFumpVDhVBHYo67aHfs6CWtb4dSG+z/FdqOwbwvA8dd0deP/87cPpwzRSUif8B4Je3bYEpA
iGti6iT4uzOhZQKARAhMTGKXMiQb+1xB5X/DHEJSyIDNMA/Oh2w5sxx4lpfeg+Sz8S98Scu4uvZR
kQ2685f1txS9NZ8qa5msYyHXh1bIDBzUAeGEvRxg3kUFEam118u9xcF+5xI6dz2jGMyl2vZmg9D3
ljmEWjwFqJL+7pM2YLgDezAq8ZZIStr8Mx4Ymb4BFSUHUe7HWyDfNqRQgA99DRcJjl9Qh3W+LYX/
E8oxHHASQV35vXNPaIcxpm3pqMpshIVFG1KJpPWJRRNjeCdzxmGzo/0CU8I8xlqP84eP1ImTegH6
6jrcswPnLJ1K70rcqxuy3Aj3MJdA12MTrETgUY73aeqmEehddfkVRdbCViCDOsJ03m8BtLr3h/Qw
KhVvlyctKw2wmRuLNj3A0wFKb3B24nHru6A4e8xYwJXh7Yy8L6MyyYXctRXcDR68Xf0d4sVV+VnP
wgOC56fLgFML5kUvzrxEQXWAr225Sg34WfMg8mCDk6/8V1ekZi6o41QMSNYPBpus9LMKTrYQnGcC
BG/o/oCbbbGkuIoWB+kXsOQoq0qLKjXx1CBl+kHmoDaSq1Sa7xuKuRPi4WlWQwETbMRo+PoH45PK
R18x+/LieCn6TQwQ86JCDyRa1tDGVj0Boqo7pvpitFEvgfrD+4pJq1GX23w5iwZanCnyFRjyVGET
Nf/cUcimE9PjEHjoKA7WU82oO7ZWbdOGi6T4j5Z3DSImogjTeqatMd0dbUMrz4D/H40TrEreGQCA
zWNfSmW1YO6vYGQdkgHqINoaU7bCO5kpv7S8c0tc45TeX3FGt++dWNa33YwDxLBrnVRED46XHGQB
JglEhAa5Bzl1HKiJOKlSd99tUPU+ktHSDA83muPoShtp+/XkVGal1fqkLXQadsodq15ZMu4pTfnD
pJ+w7yFFE6/wYci4+eFURyofbqEhL7fBWrEvCIYdzRWnkIU0XbWHHhrXzz/pZ7cU0kC3HSp3u6Ec
rM0strf5P8L4C//GSu3T3I4DZmxGbjhlvO0+iq864b6qbrx4WAojjwv9shWjS2RlGqgHwzLa59ax
Bbg4/qaS0Eq3wkV1CwYUAD/vHBk+bp40zixTC/vaxc0ZUnLKPECyJrHGP9/yEJg8xh6kXse5o+Wz
shs7i3HQ+GMo72m4Y91uMXfd7i9wrBbTnogxkiBzB4qpFj2aYuAAhLSBXMJ3N8SiCsqnxcR/6YqW
Ee8Vu19anIX7dp3D3aiJNsP+UrBdwOkvqqGRYKZrzq0z3TUVuQ4Y5j3Y3HcbhTOnRFkTwm0RPKLe
rdRI3aaumnmNoCIlSmT81eG4nRzzkvlOZ15Od+nl/Faqo13EoTm/qy6tetyulsAJWB95x5jnDUfz
K35eaa1hkuC/ZpOfVFp6pLjb6SnCNEyi2AcktXL1nfNleB2b6FgBOhhlU8huCR11780e42Xub0P8
jnXlOHi1vWdNbzJ0jIK+OG7gW/xgl/jloaVo7OfzZGeoNMM9eEQ/qRFr4zdN+alXBaoe6wyxS4Hb
bsmGeEio2Gqi4S1LbzAJAEfncmtQMGaYb4+F4Pn2Vn85FuzTGrBlDI9Zfbez/eVhBVm3Sue1zNJp
JECA9VK6R1OEvlFopo17iCcdz/FRqqDDVS83op4wxXrlLrit2MltQUVQpUAcwFZ/Zd8o4NpMc2c5
R6Su1bVmafYut6rXIkCPkjf7IzJBmIvUtHqr0C4XUDg3pB0DEZRv0/B2Ml94S1KHGUWp+MDMD+rx
VCpFwKOwiRRI3utENI2S+Hddhiq04eNyIEE7iTXAqDB4S3xllfmDI31Eo4gyO0j1F7SKen6MQ2hC
Ju3ulAPYcxoiwXPG95NuC+ZeERFOAA5+qnw4QWoQfZm2pzgBg5C5M9wGwATAgvmKJlajpwjOerld
wCcpQ4tLGfh0Fm5WXdJjp1G3xrtpyNv1o3H9Tppwjdj59rQKtECxDe/b9odnZ89Z5XCPWF1Ebb1O
+MTOLgXO2HuHxTJTZB8iqhcABfM0hjH0QG4wvFv8y/wTwNJZdLmQUXDf9Kl3LRrG6FOidNMeStGz
2WNhM6dokZHFcg0jmq9O+Mveg0EwzQckFO8mC76Kh7ULiqtza8enqgKlWuQ/mpUYdUn/3d4YyavB
SIz1/qArnuXViZXj1mP7qS7BPb+JHMwN963GV+RqQY5lS3++IUXoUDxhoNuyAZmBBd5ETAQYp1xF
S6cjSSZ1CKUnRdg0zj3UGDnXkRbGee5HzNumSrEp06RN1k+Tgzh77XmpwgX18cBCV2m8a5Vv8e/6
U+EfNkIXQyWcIO1WWB0vlfPo25TcjWFy/Q9H9H2GPjzNSGWeIe+Wd0gQ9ssa626p1Fr9xgL6gU1c
oHNd3NfQ4sV/92xEyTtDW/H3VyQeli1B9ou2cnKdEKPLWaklKdGkuKCh+0MvxvP6w3jQKsEWmLS6
xyCaLUzM3kS9YD3i91bTChSeADymYesR/fWGOr3BFnKjABmzPLjCNW2wBw1copnCOXTSTnQUohpf
hyonoWH+65oYyED7Nacvu0uXnp6NYtYW3UIZl01hjjtcYrqrWxpb6r3Pgm7vuGnaoGWOASC/LSXR
BYwRXTCDQzBj6iECVD3k8Zi+SfOeL4Nf93erbekJhJMltzuqxi8k4WjLejn5iiqLGbIEIQxw754F
7wRVrnuVdt+ovE6d+Djgbjg5ctRDhqDjPh93mQFOks5ueF073erO1Bql0Nsw08rcNNpNcoQ/Gjsb
Oci1+eXcwM9gLI7AxOvNVFfQinBNXp5DRkJ2mKYJqH6BK6W4MOpBgTQaqi1cIEQ3keyiMLpZwaPe
dQTuu+t7iqKDJ6Ua9UxRadgSAx8bFyR73vE1YfTlWw52mvL149vfUTjIIgznjdjGlIDdIW0wT2p5
bDybEJxbkvOZ7YLfjpc4qB4DtxYgHN1SBK0e1aaZgML2MMBneaj754d5lu8SUQzgcuUfZ6B5ChRh
ziIvu2mB4jJx4NRIJabDQKRXCJISlTJEEyW21j8lzEiYQCFLCav0UM5JmmkJvhwTCXGOGw8yeswK
4hM0q+0ZbsZXJ+lWAXT+V14HEDZv3sW98UjuGEsqOKu1yXgDBaUOzHW6mdICwsek8pmE6Q5Y9ToL
UyxV/sgHevNWZ44ZC4YJV2y1fzZVr/8A77XHl9Ut82mdIkS/yDSOELGiFMU47JhEnoEh77cmRmp2
+KMug0IYZqTJgAkPeW5AmfDjCF8nDaZkHimyWpwVQSno5EFZH1IUKezIUvqYCqCUmW6aQ6Orhl5Z
2C3RCDhJ/wLfpupynLw2n6lNS/HIysJYDWjvGYALGagV1RJdZ3X1ZaHtcztALjTmqfX4skHs7m77
hfQZtwhTt4z8vlNbKGbto+qyU80yU5QQWO025U68o27Xx6+R2xAoL1qwCu2vofijSLP0yoUeyCgP
mWBrZR9Qf8HQ7iPK3Xidg1tEBqrN9sf56nNjkFAhx7NMBohYelNzE9ain7h7X3t6jB07lOviXKqn
hfQcb1pfD06QWwZssufdvEXd/M7S+Gisiwb75jIRg+JHMQYoJCj7MsMQzs7PLTOsDXfFgmScdUIG
NXdG4kwa7qpdLBm0xGcYxjFtZus9MpKwiwpFD7C8uKgTaKpJCy+n1sJZbMjlmPWF3Yf3t0i8DDU7
p5xlgABLKFiWlOKDjjc1gkgieIc+UMLQ+SC2ZYsl/1tt4FwfJDZcEEbNS7ee3cY3eY3k+Alvrf3Q
5YwMVuYSgiO0DqQcpX2y6xIDGMZANYda/59dJ+JRNuA3C/SPnmUeYU3PrRl6oGzAxm73MpEJGnaS
VpnmhDGKchgrtvbPybZyslktQNYRjv93CS/KITI1ylIgjWVty/rsuTqOB6BX0+kOmQ/+hUGQanIv
s6h6cNbwLFj/+dA+T+731nEOX5/lLWQ6FgljleBKgCKfarhwytAc5NI8EVsIe1eBEZjqOuLl9xtL
iBO76ELXXWpY3tE8CkjSLcEArKcERvQrEqPo8ZKKFBAk5w+itIW75ibyuf8DE2pTyiHZwoaR82ro
gSv4hy9o/d7kNOKc9lkfRQ/0RSYEcXWfzgZI9nHFeMGnlTa8qKjdeeeyge5Pih3H1ebLDP5NxeFD
QIg8AeowMxotyeWntN0cugt55pWkTRWl/bIB/wUsYySF2pQmGKLHIOLdW6WRCkc4hTugEqN//ZHF
+6AP0B+1hz8US72KH+s2JTQaewmbiQC3JjZO5fBr3UdumWv5z7u3oBrvgi29F3viB2BqIgP/weIM
C+Je+T+IlSIb5tSyWdf2cjIe+mfN6Xrt1lzljVEPY1QIWgR1gTHF0PEusE+hLvQrt4jAP+LTVC80
OZKZBMUcOJ10zL6dtkr4Hfpy5HHsq7SwAyC8dKLf6HcZ47xGHExr1rtvJeCRr2LJuDFOcW+esaGa
OvKh0PucuZEuChDbMiXirRikqKMh/ZXACmoYoPy0R9UYKDRNnzMhD6mDZwGJnuHgfaln9QJnqwhI
/yntzT9laCIIiUspndr2QXjuG8xQH+a4aDkkad8e3lP/+oTofGtw5AP9CZZkZHaQ6UVIzzb9yEcX
aCU9USkBy/zfR0PeeKjGT51txc/CFbCTbvY07qjJhVf2lrnJU6GYr9Ifh0E2/oHwAlf8rwpMJnWm
x71duQh1oaeAKHmPk6UmyB4CATaxUdLB3cUVAMSYdlI4MoTYTp+Y1CIjCKoqfNOoP03DmJVrjViX
YYoxj0jVOuNeh5OE7DeX7LUx0vbK5a/je2781wCZ0mFssGGWr3W4LdSyE6QfxK9aHWpC7mDdcoqg
Ds/Pbyk0yPRYQNiz5jFj1g6jpZCuM47P5khpi8cvIwcpYIDrUlxaR8eH0PYl7ThUirSxO/U96dEk
SuTbixKW4QBXtrvdYKga8IBz+acoF7vAM8M70Fbpnft1+hJVe1WqO0mFbhgNRLLlFeUXLJJ+zL4s
oUuE5Fo9Rtp/NN/dTgkPxX28J1u0tZ1bE27qlufbJ3+J2hXK7bo1jOLMi6DkUDs1kuxJZVP1oWVU
gpd4jaJ5K7JNb6AnT/8XwNfVRj9wLpTPxb9pC2vuT+TApKioDmGQwC5dl/kBKCDQuiG3gJGhPyE/
2q9z3E9MshrtTsT4FvWLxtzLKlpLNeB3JWwXCBWkqDDh/Qtf/dgXZijnb1f8vnqSGEecjIG5BCDA
do+p+3PRNdRRfsVBrxbW6U67JlryviCqNzv80PXv2NMFE+uVLUqpZsoyMQZTKFE3nN0OJ/9uzAi+
8gi176B7TnVONcdwQmX/sAGzW2/CLeVXdtCUPagdefgpuxRxNRtWEhuZlitWhBnLdDmw291ahqCy
BFcqcCRB5uqK28LMgASTyeKAOD3Vv0Hp+lpcdNYknfG/ZVxIyAELEsMQPjqEiNJDbr2LL8fHbekT
l1T3sLu3gRaRSNh+LEH1GQpjtBQuGLnEcOpOQFfxMcqn2BXIAEWLt8I0nNrRND4sN+anfQpvPdDv
MQpiwThlAgGWHuAt7BtwT9n14qf+K1loPvpuIKqwXUOzR44EpkOsYYezy3XpCNVP5XKCMum4ciYr
F6mtEKRZtCZxnzSFD2ph4SqymzKfxTaAlM8m23Jq29OaBjho8Yc6FbOoeAIC3iG/XejDl80j+txk
deoc2KFh97fY2AnFC3zGuzzeHUieeliYMa4+COd/7F5DAsp2XZp1dBepd25qE72yWSnUTfjOOgk2
MS97XRqdECQ1SMPD540llyvVi7m+nlSf0kshM6kfYRxdOwis8HxWGkQlBH+9d4hSBpOMAUmUTJRJ
2wztO7aHRbf2Vv5mEeIAtSWZI6c1cHsCaeKSMp7GWZp8YkKtqKWz1anZp+KJJnSB0+UnRKDY3Nki
NKul3Qye50ODWhue6PFqXlkj+ZDwdGNiFgjsIXlf1f1uelmj5Wl4ABINJU1tegoMqXW/zQbK3d6l
K0FyUr34rFhouv0PuRQSRQM0a6pn6ERpVHu9F9tKKboRgGq4JZwWsq4NNftSeef0qT/KlSSb514t
yOj5rREEZht2ZbuvysODqWmhP1rIdPlOKhcrDpD0xRQ+ZwnhnMgbCY5hW+PPu2TP1kBUbtt9+XuJ
K5q3fq7ea4taHgIwXEhvIKr6bXFXYHO4UUxjGf93rB1COWzIS5muMbqCkx3JLR4omlPrAux0yhzp
J3j41dnKFVzx8BEKlEiqoiDfD9C8BD2+XRkDK+Bn6ji9lJDDMVzHAjZiycUCvrXbwIrbS5E8MRLd
dxz1ujwJTZ2aRatyL0el8XEJivngwaVc73SXgKt0X5k9sGg7Mm+eyGdT6nX60bhyllaTvGvLTjyv
+eDL5MHjqi5TI2XlWmHSu61ELOU0CPY8oKywTf3LAz2wULu5CH24xHPkFdm51Sv44FRYjzjeq7WJ
NUzsBc2aLZspDPNIBqKYXy46UUbNag55vJx+mNs9sWr/gBBc/femhRvikv013qC1wrlNCvCmvP+U
3BV9N6UbcjSrsCbQPvSblVtV3bCpRg/A1N0UnTuFOZ4yvMnxG08N1J9F7fEvbr/f97TA3QF9pItW
lncMhV7j2AhLB26NcT4+21UE5pyN57hf2BaJcnx8vV7io6269CQgEkaM4eMOcY56RcTOzw7gayQB
LOXX+ltG70qQ/aH3Gn6AP/EGqgZWg+GbdztvsqUi5LTMWSDipDz58g1pV60UngsTlJse8j4f0UfI
srQXWo7y9G99x5lq42TRV62wZkvOuI65eK6j1BH/TLXjm4KTG40EI/XEUFCK7gmKcH1PeDPALEQm
JMR2XvkFJW0tlBTk5S6qiSsALKu9+EMkrvXFn40Bk9lv2kl5Dif58o7aVH5lB4wqTvhY4OXxV2GT
asSb1QG/cfM31KuIKG0z+fq92KsTaBF7nN1c7yt1AEYV22SaftngK2Km123EAWu1LPddkTXhHPT0
bYiAhteP8nYrPo3wcozEhdM6kVSV7zjUMvoYHFOyYRQV58lLXMigBschzqBUYJG/GbjU1dV8IpYL
3p5sKu9tMhPeLsPJzwpln6X5mO53jd80VdC9rgk1AJc54eRkMSMGO/38ChZwQAxJd3QfbbSPWT5l
3LeQQ7aG9aiOYRqzoRgLBCd4cBAm2IK/BCDMysF2UtvvhF5ddAjCmKkrG1Qc8OR24ry2AqYp6cQi
+1CZOgRL1ENf/bvxDl7YlJ/X+/6cP/pABErNwfo/WikOpA8eQ1DceBjPqua5H+8wvs5WFLKVLyWz
G43ozQm4H1kEJ1Qk/DetHpTTc+l1Gqm1KGbmzyiXRZqEhNn8NDHqkwW+LOnWekUIxNmtjz0hlU83
T+eRY0N8F8AN5uaiLmJkxXXzmUFacCJSMemWywUuRtDRV2k8K3gw3hYpzTRNNUf4/FfEKkkj+iLN
Lbbt0QjjJwDdftxLHPjfP4ZUtyN/PSKuj2QolBuWJrAVnRDVOBB5T5ptMllitRjQzt9AZzjqMxOF
ZxIbPb20rNGAiGbjHPgUn6vB5O1bw/RzrCgBmkLvyjS+4nQ0wbRC8S50RAVK6cyAcvDUuSl+c/48
vM9yZcV8wT5YqIw6qsu0pb2N1px7UKaGAJwQ94IO2oL6+QXExJDp5XhE66eT8DQHn0AhMU3Pc3ff
i3BYUIPmGhFjuw6ehj5WR5eDdemyNhnlCQtoICUVSaXK4GP7F0ggT18JReMV/iUx87KDItLgOOB5
FcFKEtPdTJMCV4u06uXPTX0AjNplEN/13+GaNjr2nq0GsNqRd0t+fdBTTEUmFJ2u57osOboJlspL
rkpXT7hX3Izypl2kwa1fb1h+XqRhiBj2SQYiNkEUGeMSyH6L6znR921SjfIu6jOXhH4yOY+ecf01
03twWgeIwv4sGDTgx6v6CFr6oagEuYaSbjulMDjLz/e/xmMqYQ78D6P2YA8yPr+3KVdE9ZIkK5q3
K/CzAKrRguEXIzMpuRjHP3GYeYcXnmqTPwIDiVGaSXhge+VMots5U+XnZiq/O+SCk1XdKp2Crgdz
FzO74DEzACD8Abswr49OM0sQy43pgzUQRdTlHrlAXX9rBKqnzLImKx1Z6DvABDO2wOpopUBlQIaH
2Mr+rZxySqzNVJvnTSvHW5EOYaOcHjvy/NiBx3FZe1HS6NKjxVyMbxQoYHyxXq3JMIOK+WlmCVK1
lMoZlSWt5fkgsmRORqFLF/SC16YZQ49Yv0OaFRhK6HQ8wba6lxQdpxlxoKdb8/nkdnBjpPTHCX15
LrACP+IZlYvtDa4CLi2pmMk+E4hIGi3x68rY5FXrMDB1R9bIV5q1im3WRQ6TydLdGJiPUGRwczNb
gvO4oIo+20g4DWs3owVGXWAb7N/DMR4IHDp4jVOekf/046sUrhyKPr5V8VS1c9TGDwJRO05Jm+iG
YCIZLu1oerx9dl1PfO8+FCzBSM2H6uSL66hzAwMiBAQxrv84sx9hlmP2lrunAHBbvQnNg3PHH8VN
KTfKzWUo8N6g2h7XilNLg/WhpZoWZqwJvLV4KvQXb96I4Yp8K2JPKdh4MCc6r55d2aPQn4Zmw615
nmyppDkhsWDEop77RxeUMniRF6+MymqA4dcd8EmLhVJ8LojCxwAB3hCmzbaczqArGBriSHXdv7uR
tc4f3DGh6oZc0j3MSa9BSDKxi/xtQ70NRGLULSohu/ZnoqKFTXpKYjC6ROopsTXjoCnUcyVee+vF
ud0r6wBLr1GvflAX2iOrdDy7a7zEaCdGPLWUi8obY2IJp0/93RzoY7JsG/IRww+4m2hTvKsOGAeT
/d9DJvLdc59aKmh5zyDBWEHKEbbwDU4oBJwfKdwzIzs8UONpdMS+KKImkT1TswsBpW7MInkKq6eZ
xjVmtdCzSvqBDPcmDmGODRQiBQGCf/AmgA9L2xqb/rto/JwP6UJOSylrRS8HTsDap15L5R9chcSI
XCJAK21lyaobG/0Lx3u4qKy+OEoVZaJEXxvAP+MHA10olaVhjm9q5lnhvf0c3mIEhfxKmDJs+D9U
NtcrfCbiBkTdsbe6MxmE9NyZ3/Zav0kpYmEpQzl0hnww0RRGrxDec33fUDWm6ez6kG0Lq3PsNTt8
TuPrNhzu6SmVgmmh9637J8Z14D9AutQAKjHdDireCaxXcZI+HEYNx3Gkp3YbslKj2lIysa9lzE2g
mIP1uljpY+uTEuQH4/4VQ8dikvNIxgXaS+bs4+I4rZkmdaMfSbA9J5Ugn0N/D/AXAUXungB5SptA
4g6LYeHo5L+e6Zzuy+7J5bTY795/yes8QQZnnODTd+Iq4sbTDk/+7kCoI+0DIWyzjQZoTT1pyOMC
NNcxFOVXZZUb0CnO7CEunumchcPlpFlnwkIs/K4GW7h3jzJ13GNPxMxuYOftCssGQRomUpRDGU39
waae9sE9UnlXS+tomze8jFyqN8dHZncTq++abBdy/My8LbaK9Po/FTK/rY0h1x+H6X0RxYgLj6nM
5BUQc8ia02imEOmeCwb8qNlBcJz8QSpfE3PPveikBAgQtxxkKwaT76Y74ut/kr3Zju6wIwR15N6d
ZssGsrUakI5grzJyRFQ8gYFpqEg34qQsrS+HSy5fFqCLg+aSGD56bixiA3B4I5tl9avIpbNy1m8B
p3/GWCm6K5Mlq/GlDZpRQWayVqhUoug3fjgpqrs/XlSfGZNeHZQ/5w8/HJEjiYUahEdkULrYkgUX
z2TQuEmE/oCe9ngENjU4bfqUfJdZkkWqQhNiZJq2sZZY4sPjdI4QNt81icfqLafkaAkj7EBtucSl
fj3hvzdXCma1sdpqa2wcGyzWESRuP2s8o5ESuPBwexEFiipC9sfTcXM6XsQMcudiq+nJ81VVdRHH
Fu2tXeTo0xdS3JObbYEYT7yUOjwBES8JYqh5kATmRJ7tt26jSUfM5hLz7+qZa7D4+og/gwNg1fwa
kCFlrJU7rQxQGuffZtY1Xxl5oB0VTioZXPwIeithi9IJZcXKm8P2KVKZaaYTzJEOe1KMGoF1OJoJ
iMXVFN3VdGhjDjxS1QSAPjVf5FYjNTDV3fXmB7XlPWY4xKZH0TX8T05vK86ncqHBEsJ0DYOFopgQ
DfutMbXNAhilGJhO6crKNBDYF5FvCfVUcHiMJu4l3pXw8lJGsU21QibvGuwJZ65kl+XB8v3yIpzu
2oe2AZTCnJcDJ36u2siThxSDmu1IV3ANwmPXcR8o3XHzfSxyDCaBr7LcCVY5AQiivNfnJ315RlIb
NEcj+USeJwK9R9aZ5a+egfZ0IkVrdNLT+OeprhS2kVSSf+1SMDZbbG8ZMab8DwF99taX4PTNnnqn
XanKpmorugZAgf7HRVPxAJVtCbzyXEf/jqNBMYwJouu9XuxRiaMFRk1LauAahF4uGxW7QF4yjO2m
ehC63Kl2Wk29rUNOp3/TReh5ox85XeMVeuS664kuZHFPax+0cyC372ktMuCq8atYjQMqPSyY8/r5
40/skefSFSW/v8qN4NwP4OyqqxeZoe/uhGLa5kTlkxt2DIYrsZQ5X4c6LE509gN4M6bfrbyjhiPv
8j9I2U/vp4hYz0Lcup13GSD+UBvptpjHgbs5d1QxWC5UQscLp/HyMTAfmUPkpvNZ+/hwyRpCF04K
Mby90EE3/oQaQXul6gCHa5KrSvH32QL+cniNHV46KbzNbNodH4Ak9lVBw9dMZhCAKfHdUENBzURB
bO9heAKWZOktPvxAlTMHr795AYHOwRkePi/MOZTsXkVH1zrJ4Y6mUhl7aiIEaVcBOw90x0glxmB6
B1Sn3lKfCjC6iPAIsKYarLurQGtIoCz6hMQKD4ZeRPNxhupSz2me0d3LAK6x7gDqIbLIsA7VRfak
1C6+bxTc/3W1ZA0YeDwNkhuy1zG19fwJvRq2LZMFzydJV9W+bI3owAY7Jg60DuBlsC1bDKbgjQf5
/yJrcGNdgX430IeuVvhsmMVN8qJqB8hL/6iEkztIisJT235fyFnZSIjg9Yr0UV1dOJhYWd8/EeM6
2gqx5tmwEFR2DZIVwk6NWHvC7ykQWjehxpXaqZlsaRRPPpjDNaosRQk8K2QiuO9ItzXlmyScAbEJ
3DS7VND+FPteE0l3JNPOEIgRuUeL1pTsfW+SqxPTJvR9u7m36iA8Qz23pmCsHUaMl2pWVb4tiVMT
3Y13AvjE2+YC2DKyXKH4jhHM1Np8e4am76O+2//muAGB5xWpLGf99c+DMdjiCWKq/UJgOWhTjypT
CmebhEWzZ5GAd06E5lfCVzKVjok7bJywMdWDpKQvbK0zHO92C0D8tT/87NKGl9Bb3b9hSfhZDdnR
eD7FFYAfCi+gJQiWWsdMjAGcFzwcV+n9CrHYYwjomzbM8TWDuDmr9XteACzSz/bj3Guf1dt5H63E
yKnf86TW67m3bc7C9d7XbYmHhaDKs55+OKW4+3Y+QFfUWdk4q1iSwWXvy9AGwXy6KR90iYD+pHm6
QfDfLuMAANxGVuGgdWhYDXYUZ3QbL01p6Z3yLOZEE3KjkotbmRAsCz2UgWB4WY0ycUrAkPjDQjiW
gjFtueGWsEiQEfZJ1Yd9o4pJSXAZvpSdyNuPwo/PDeERRraxE4eCQ2xdhJqEeVMQjcjHO/9uE1O2
H3V4jATTlyp27R6NeH6Satob7P2qfEZ+Ivf989mTGyhg/2eSwEQ2nuwb9IrXyIKIV9aZB/zAgif2
Id44ujo9eZGo8TOxecI+6w+9hcogeG5cQnAR0nrw2dwX+0QXEOl1CX3atK4ZPko7yZuTmj7BW8zz
xTaBcCg15uBAfWpaKtgDEXGtGJibuh4KbfjhBq1PUYqCf5TmsYbE+M5EniTFJcIey3Q3fJRYC6X3
H5yunGwgBHzhM1OEhG8aUDoV02ygy+sLllQleEH3BvKDBZuO00IlmDEY4TzpBSnxqIrW8H5nx1VY
4Jso6UR+47RsLCT9f1TCNe61AX4eRqdmfef6WkcecKzF41Y0jFADAt2RvdTAr7ddo2bhnpslXpBr
Bih/heddk1FdFlPZUoGBpc0x+VSCxAMa22wjenATNCbQfQustkieU1fQnL8VduHaSbu7+JBbazC3
R+0gvi9fS/bFlkqTzhUhXm7VQyEbRMofJNEXVTC9iNoqCvTo06CopoPEo09/A+d7YT1rcfjafJdd
ZAfOlXn/VR/NSzu9/gXPyJ5Bz3gqMss4M0L9ngz3i+JD3CsSYYETQusCyXrz3ijcmWM/z5yFLaxW
95cScmn3x4mg8trJ0QHGOj39mQcCRgDq8VogB5FIUzviC9qdgz7PRsmaSsIeynqmXWRCjcjVkWY5
6EIU7vaOc2H2pNhzhLEaC2bIxb8AhMZ0WnQSA8DRpttgll06Lw/B/MviUNc9CBiZOglTTgsxI8s/
LVqDxJcwEdlshTTOLFSNmDtUPhfHsPegjLaF+FkQReMEHH6/D/R3kGJFlPARBVg32MSwR2OsiQvH
2AzedEOTQtYHKGRph8DyU9tmRhxKUR1+nFdjTEGzY2pXwUq2wlLXmmlsAgS6Ee9/11oG3569XToz
7Ue6zKCYoj/kJxtmTkhOwV7MuopMfrMUP9rr4mkfQuv+uVRgTK/jpL3vczfcvyS7sFSBbuDIV8cB
puJUen53UAve8CTWOK7U0ui29XAtJKZi3lgjPVxyTs9vLbGXSwaVxFfwUikSnFOVM9isqDYW/w7S
kiL5Qw+lDyg4daRLfOGDEeoGWDhE3bs9dZk/QsEJOhmrsiVXBUljqV7qw2qqoaxue7ANOrRnU9vm
ug+ZLsSbunc5JaRYB7atSRs8QZ2zVliK8R4lejBZdDwcpuRf+Ul3ZVO6WA46Tck/wwmg3FHF7zTM
vqjIQDQtJhD/KQGunM6cLlLun2J2ZjhySx/gPadurdX32r5Unan5FZWd90yVvP2mwOUUBlkIenKJ
ZpkNx9fGoYCqFuRbtrK1quSRJqvWAwbEP6pBswXZFA2GRtz09LD9mpTskqWB9J5Ro9sZlToUXDBm
tsqa6gfnsup8a84gG6zlrc2PuO+R2Sw9dmiQlLegdvo2cXQ2K6dBgCP9Zy+r8Td/A3q96h8anyqi
k6BhHvLnvgLkbdXJE37apyFxdYisuqq3xJ7iV6b+YJQgft4oBRsafVxohtAO6/z8dzdtPMoMy7bY
98Gp4zViSwIkdjHvdhEpknKtXP2l2SUxqJoOME8VFuAm8nrKbo03cSA6KtUbJGYja+yGlkN73HmX
P1Cm5Y0zwaEPOltYaVJXdgj4lo8Ja2Vgal/fo+9vOwtpvACivMPtcs6gcI7crBoLsntWmFqF+1+K
7qsETfeHwlvNpy0q22rGZ9aBnf4qfb2CYwf/Yb+Zl7a7dMD93H56C/kGRKnNjkS6Pa+z7KvB1R22
sh4i1IeXmlxFDyKAwahSyouzMEzruqvgZtGtUYQ3j+gZI0JbtFXTsSysA8b2uMyUnOwdMzYTlLCl
Rr3opkR/0uuYa+6K2vlFAb2vurnOrgfw8PklyQCO/s+XEoLU75Z9Zocrm7Ce5+1xcrFieP5p7bFA
t2HhR8J0v0KLF9/BH9mhOhKJQRpKBHxLGhizbDIG5FRjYq9QMuDYxWyMkiuXxLmq1ip2OkkJ5tOm
dkkGKRy6Om98KNHRkhENaUV+6oQF/8T0tVPkOWKAWKmSVeH4UeJ6ksxQeIeSNTkEaKnbtJFxIDru
7HeBl8uXHW9Et/QZgV+D/zT1L+W8j+F36XNaVeMA3TyHwF31J0YoSYKIkCEhd3PhNI/3TqgQNVlN
SwbkNefCyCBQkaWXy3jc7G8zwFwKFSzPSY2fYv++Jfi1N547VM+VMi736iWaVy2M6maq19EY+u4u
H2r+kXs8CwQIpEngTgWL//LRS7O7fJ1Tn3ertyzUOMS509uABnX5o7JgyC/9119rCPt1V66fCvcL
QFblTjqJbFgE8xMI/o5VSQJYLGjGEhJvtL8PwTFoPmjPY/h6RPMJkFFdJg5JQbL38Bp3KaSuIks8
Faqjy5XU0l3R0PY3ZeJzjolaMwInlvcShmf13Ne63nGrUfRRvphTaOEeVhfcCgUF4ztYjwLkHkqC
C/SsYwpGJc6oJxDV/kAbOrrjPwjnK9nrmZVM8PjEoOT2Dz8J/ozwS1HQkK6McSnE1iKB7M0pHGu/
/ho7NSsslj3r3BXO1lzMqLIIrcIGsX+mBnbIBZgfGWb4rwU365dVCZ5c1QVXpAxM30ZO+RpRcgj6
48RQZbUpnOBWwldsOHAFDycEjUKzt6VOdmv2fKnjf5+MwHN2D65gR6DrCFnMsSbLfLiZudDSaMv7
2zr93TE89CiYIr76syZ2svYcQLyisb7ACBlWDMuUO1GdyFjQeKRz+fVX83xMcdNJjbVe2YfPRPAh
N5Uozumnif0yi88lDDN2m0FLFLiSeBtpNI2N80RaMtwj8CgtoxkozHqM6DQkj3PItdr99KG/z7s9
lygbGUSdDaX84H51gMxuVM6rW3h8UN0Oov6DxFgwEx/SK9z+lh4bL/pmJSq2q7m3Ym0t/5Rtthln
sHEi7XidATusCIis0mHLaDLgAz9CGOBTb766Viql+Jh2Vt8e2clKJ+2DJHQ6PhDrqQovHjOM1L7x
q9S87PeXe/mCgH7ldwB7ADWMa1yIFX57qO5BSOdAP9/Evm3WOWg+lgmFntc8EVjyJdlaZES/ARs4
Q/aDct3QxlFNRl841f94nCP7FYmUY176Jq9ewLxs+BX2WpCi318faaBfB5+VqWenJvADKFCkf8xw
CaRTdjw3/aLtsSD1AvRbMoxkgUHEx5319Ffa+b/uK6Y1xSjCLHrUYz5WgCgBPUhj4a4T2Q+puInz
9Vsnn9onPQMU0xniuON15ILaHqXFZWVPqqP/TC/n+Z+5ZUVRwh1q8WwGNJr+lmCNizwzBuJQkl7a
GiK9ToXtGUUnVT4LpOSjkNobRRvz9RwO29+1qlo564dXqzR4hOJghWjldsUXgfzhRCxUz1uU7jwM
Ol5ZbYodeanIjH1KwtwXwFqjOvocCqT6exDZ4gNPqwu7P2/05TvQTt99OGjVKTC8YQSwJ0Z5/0GE
EJO6VKCdbobW4+uMH2lGe6sqnqAUUKB4zvofVmC9ym7VLh5SDCCoFWOhCZhByfCvobX1zpjKqmAn
fmC56IiIovEhuPPlBCOPKUEY20/qc/swpgx/dW6xH4iprhFkTk0CciTph7BIic5OL1yOsPQzhtyp
nEc75S1JJ+v+oVLD+B4A9ZDjFhyt4cwKf2GnPzdWys2aGRsY6s0h7u6azC1J/tuGmrlLbuAYJfrr
9MdCkVKi+j5G84u6goYljirHMk9ClG40CcfHBrBrde7wy18WSvo+74qaKcPt8i84TPuusgGOR7xa
UAcQeyv4BfNDBxiRRcUyQAhBsoz7HZuNhlqDAUW1NjFbwiK6lJvTXxur/rudRt0XO1UBVhvLZ3yi
vPjx61S0PWosAy0KcZj+UC3IB6YAyLk6hWvr1XnKgQu3lhsyjhNQf0BuH0/Muy0MAP9Ue4zgSV8l
SrT2Zf3giZGvJnLtD43sWJ25cmSRgcZ64SvkQDtRguM4pJRNaMqTRfpKB842Ly+uDau8l5AjTv2T
czQPZ2CSEPoPnntF5hnpysKWdoLD+Nk3Q7bkXzsfYx6RBWgDCS3evOm1ABfPvXtKZC2NN4rXbs3R
rWwBvWKUqv12RA7snJMVjole3d3KdIfzpNytwRSl8gTTSu4gUImUp35wi+rtXiVPe7tIYgnFAPMA
FzMRH0/d8k4katbhYgf0y2IjrzkMEyhGkHgtzjVZvrM5zasfSY0ztsqY+XII69ad5z4PTHWXBsbv
HxWIFvtwzLlbL6P/5HX/P/P1xXNHGuXQrfH7I0qtfAw8rqpQEHIptxeYN0MhFXRBzQ2puya9VNBL
iygWtfnTVmEOV+HVNVGNi19CKag5csbKwtKsCZcg6yUlT2reKEx5ayohYdT6IfLFPVb6LZ7gtqOz
rD79yiHMeLQ9mjR6ASQT8UnxKyIujk8rQaf+fJ2OMczx5sMUglmsuuxTNjakLnneG6ge5OPqUhu+
Z448kF2zBQOPh+kO96hPDIgMMufPVj0lAKdB4HbVlYdASM4C+vzkZIa8fIJjnMFp+co03ZXF3fix
JLEPfYHaisbxpeeix17QKG3sP176EBO+i3JnHVldMnWw3xxitXI5JhzZrtL6qS2ma7Hw9wGVE0jW
Y4sF+fc2YCFKfjcQh/18E0BqKVIzEL9Emfx0s3UDUc++M3PRe/TjPldypFCrLxP3EJnmkzv+DpbZ
gqW4nKGCOkW6oIosgtCpTkhEF6Bex9Dou76IpD/wQ1KsfByHVYa/iJOp4tyGXwfUNpzGF5U+o0Nq
PajNQavndMdW7qOFG2D9WU/MFn9xX/PVVi42xE8BODRC8SzeJNlnziy42D5jf9EZ9yb9LxSGTjCa
Sj3oBmeiP/2c41TkqdNaOYD77IcOAJzXzTy9QQBd4U4g/TqWn26lpD7NyIqrFsbfwUL2YQWGNJBR
xaZrgzVjq1W73UtZs9hp1YKSFWks3uJVVXEIDGHPq1BYSYTVjSVuR0poXJd0eUyw9woPjUMFlrMU
GmXCkssNbNMAza2UeqU7PIHSYreJXge4EaAxdfldG58d2gG2BjTZw8wiLSReiQza5wwmQKmR7zwG
5VlpUbEyHTu8yoqy6TSAjhU5f62hYN8hKqkVmSui5Ub2vLI12CqtB0Hv5r2Xd2/H5uFcsGNc85sN
1YT2qUjxS92r35ijCm3jpeZl/GHDKdAHJv+xmeGUVNIBdXLYpK870usx60H3/fo2NZIXSaUF1pyd
Cc05/qpK5TO0zwXcSgJoB8URm5RAWz6SO9EJCKexlFJxytxGp6Wpcl3ypJDVuGJwBm7Y0fTtwLHz
T5sqv5ltVATg5aysR3JD9sSfdzpIFk77LwCTwxhxGg7d9rm8Lkh12VNGBlZx44r7VGJ7Emc7KdAl
dETysHUTBsXcNImKpcA5UHEnilByeq9xURMexQwufIzdFfLjFkfpFnpxp/oyI/qQqB5L9d2RH2dt
7vs/dz6Lw4gt6nre6b/lj0QPm7g1jLcCZTey+pwny4NzTE8UCK1yxlKEXebS5tmHgBwTN63gUzuO
CvGlXo64Ffs+dNJRltqyGBAPYihu4CmoOGV36Sl0oWMT5c9GgLhZd9Q7VTh1JMedm8cggpJ/hU5M
5M+U/1d+GBwqcf+s5yEuaEwz3GNpOVr7u9NycieXY/GGxR8i2+yt1guM0t46O5t8sM2bf9uLQz1j
YxcGQ20YfO1rvnh1R3KcpfiTVpoc7cu2GTSw4s7hjhJ/4cY2Z9jctW2dpkV6oH9ljjEh57pYWJjG
n68IV1FKy+D3TELHL3iiUkADXAvNhafn5K6+zXVnZJIoza47EWie2KismXP4KsoNMDQsv5t4xQwu
zeaFVejMXhxR3+GQl9lcFFP/NH+L3lYw0FmhTS4xBrhPNjZo3Zxtn0J//hPl70gayg+m+6WGSjTr
AtFHvwDmHJXzb0YxIBtgWakTINqCfhqj/E9kZ+d7r3QU+hIq5b0fqBT4U+Lhc1KTKG1Kqcvx8lIQ
Zw5nUaqMRtacWtT5Nm8JmUUpbzigyJqJldAkpguNlAkYAUaxS7WIRVneRqSpkMBlOO7NrJNda4DH
aBZp51Ho5BA0LMkHwzGTwdk84hQi8keIrcS3lWvwzT3WMAJvFMQiulbiTyoVxN++J/30u6JjeqK0
jsAJCVtrkBhAU70+hHrzNajI0f6epQsT53QfyoQ5yZbplHJSTQV66C6RiE/fG1hweO6DvO6SCBn/
w9tAoBOBnnbEst/4HA00nlo1F1pxLOwEskW88FJVJnqxlxEg14oYB3rlKdOPO/nOxIsXFC3LPzlK
RifHwJp+mYD2mLoafZwBMsOuckXXrONVydoiiDpH5bM6onaY3RbxqRlv4AZx5WjFQYZV6kxT2MVx
efMM/8eu6dxSfNecMEHy0WyAKprOLqrO8cv5qPeWd9qX6vZcCB1vzhlHvIp4dH0InPEowjBAOX9t
uyl+M0AHqLg93IditO2A4I6ILzh40fBDgYQvJQdUoqiQGEqZbhnpGXqCk+V0AKuGGklJsZsysSc8
PCVfe269HAB1xiyJdLty22P70AqUISwlhSeUV0TMQKbitcOXtV+Kw457p59g5zY/K5P7JBXdaR7W
V7QsVpDYQOa2D2S8TCfGYxwfp01gL5t06SoxPfpv+x+NkIPmoXhCA+9y3RLd/4oF+8MWp1Z7UgXN
jUp5iq3WuVl6qde4ParXD3Q8f/g/bEuXtwpJoBtbSfTQve4mC2BltmEBfSIBc7KqycdvyMI4kUtV
OTembt+mqQnPA79WRUW2YPrbsVJBguv3NU2c2sAS6QOs35mgBb01G+zFSHn3n8/9wdsMKZWTLu6v
0KlxkORqFjJnCANRpbphUupg2DZED4x+JioRTt8UXbOW3zXss9BdA6C/1AmhSvavt66aMTvJUopB
Kk97w0xUkK+AzI6u6CRRIATRSlp1FtBVUJqn1+AyfmD1EXXJlA4opLufUMcW7f8Jt3xgEh4WcdkQ
sq9whAXoemD62PJN7eVB85LB62Irgsypd+bTCMyr09Bk2AiogxHEsmDw79+aLk4S/bi/WDtxahnm
FKXfgxo5kz7QH6y1nlb7dKyOYujPYE2SVcglw1ntNrvqFSg3JeyjDeeqqoGgn6OOcZpjJjyhn6iy
Lcr+GN9kRGh2Y8hGqI5/EFlGh7uNJ1Mqv8q7mr6jTVmk0Sp96CBHXuzYbqS8LXjcDvvd7bxc4vPd
bM4gumKv+G/WmcVwd/6B+w+mcbXGvs8OuyMKy6cuiOycjvkoXRupC87fmXi/LsQJJpl8V29PiEFL
sg3xt72Z24rZcjl/0wt5C5peUDYaN0tPRx1NGZjVvCZI8VNUfxTiPORFNdmCeXjvAolsX9LqzOIl
/ev+5YblfJCeoax7XFrztmdGIgHuG5Y0thynRMAK7dwDwfhiwp363cEDbQ1/6kK3znuAP6WUGBII
FcAPXTZknZZG1KbDUg5MZHDNSZuPY1rd27ND1J2OQBaOJM5qHB2HwATbZ/PZjytxLjISFMDmYPxq
3lsR83xEIinY+f9ad3ri7IgzuwYTw+FIQbDmzztYr2nC0tVP97NIi9tTiFXWUps1GYqYNEQX9WoU
VNvEaf3fEZn0vuH6QqbPd35kbpi9ItVIe67A6qLzD8nz7Tfe0JJ1koT8GnRg0ve1QUFvQps4HlP5
4kiCyaUN+ZiSxosfuuQzgvXklDAGyialFnoawHw+/70x8RnUdxZf8pXsXmLn9XpSFOAWwKCTc1ru
/yeRgVu3gJbciOmwZJ/nzUNHC8PIMdUHvCRe0/eWaGyYM9/j+KeTqxMUBSWpnBryUpMT46jq6IfB
B+4u6EnSwdkPVsxNR/cmLTEkhnwL/eWDMSE1Pg7xEqlaP9tsbIBIJ5+0HJoHtIuRvbCbrILGYv5a
aUpnlDLrSabrcZv/mk7d2tyX1MEazB5Sg8CEAlDthKheIcA2huVtiEmuR96JiDQOrqjqCdJkWrPt
59EAsXYGu8zd7jdx1nSKbAPOeWYRszvUMk6u3GbhfoMSwMuxAMUopkUWno1sPDhPOgl2nsDoxSev
elSLrpCr63HmMSTRoxgiLU4HNwuuLH2Z9ow7gmyG3Wivad6XPV4m7qR4XrawXcaivdmgLBdNHt3u
bw94MsL4zV8fTbMycgu/jeOO9vomFhYH+KUdzrxeGmY7Xs8HY0ul0EEJ1rjJGQHlhcDsins7zANk
LM6XMPj3ZbAL9QUaCPRpS8c/rs7YXEbybNB4YVLEHbzRyWZuJepbfMzSk6Bw2OEktPpH2HL4WZsU
JNrzK8DnN3SS0a2DGFqvKw57bTPVHzKIQ9jXGWs2/zeaIj6VKUhyYP4ZQdrdRkfXXX0hW386q7qw
WiNSLM1iGZ8ZgA4Y6jdAvhN18V1sCf0ipAfSvkZ5FpGQA8hPQ+3CoJ/tF3GU+IluFCQ3f8ROK5/S
fPuuv8eL8wximFl2W673Qff0ug7nO1zy/dKfF9NEib/DHo+VlS6vVC4h25/AznC2MQZXnwMzl6XD
BoyWX9FutTnwgsel3O0PuR6pxzOKVie1GRWPF7MzKmsdzqj1jBNVGB7JQVZgCS2L7omuZX+X+siF
6b5NXl7SD3O1DrMul2R0ErDDvkdMRoeryeFHi5o7zj0WiXQVrs2h+0cFTucZkVjf+yYYRwdq6Q04
M9V3TwmJwtnuHUmJ+sTQR0Mw8HxHdSoZpTbyqgfGyBMCKscTOhqnnuCD2PjjRDnk1jRk5USujEwS
yns3q6k0BQyI3E3K4AGaa5utGg9KoPFlPEfO4IOi+ml6ePfjH92o1+xX1O9HfLMP2yg6nL/v0tEq
YKt4/KlHw0k7P6jSHiYU90fOBon2Q8xT6uYrPjazfKLhWQm3640tnNXIasoMKkjRQqeZaK2mMP8u
bGWMP3mpkkiH3CPWz/NcdG1va7NqW+PVS63HXlIkJXqC1kE9CLkrRdGQpuDWz4V5b5Y2RueDs93t
bbDrsjYkaasFNcGt4NVKfHUBCDEqULUb8flys/4krObViWPH6/bFiLrZxN6x+qivqcKCN7m1b4uk
/7g23UTj8l6DIlsqakiUyNbWt9012n0xmWEImMIa4H0r/ICVgBFA1vlZQfkMHDP3WpU4dXaoigGJ
4ZUIkpu/0c/xq71iHA+Q25z33IB9sKWBZFmsf+kE+3Lh9I7nS8Gg9mrZDR+ppOAy5QsH6plJ6lLa
fwKUandrBCkM/1aNEL6Ioc1KQ/mA2JpaTzTfCVI7Z1+WZwv3Pu3RjtnnWKYOZItKaj0BofMKo22M
eVcwyar2e/hvTnGgN2LxEYMEGXc2Vc/WN8qdrn7V1QJEaNVsEhmzV7ldmTBrHFGeDxUA6GTWsAek
6oZq+btSINTGN56e8aaSYwrtTJPloWt0jv7bJveCA+3dGqe8VxPZXn0OKSqHPiju+ubYK4uAKhdk
xWRkByP2NOqodsNeWcfZDgy7HtmAPXu+Np2JXcmfETpCuT29QoxWwfKTJnoDltOHqRIqIQTn+zxg
XE5UXOrhRg+N/iVjnGv/nDpi+JVSXIlTw5cLnJZ6frEuY0NH2Reh3vs5/XJLFZlJqpFyTTV2i446
O6bcoENmzgEoU4CqREmkR8rKnzfh4c2GWJLHNMcjJ7Ogk03189P4f7owfsqPX9pX6dBIRjuPcqVW
fS2Y8qz0OaVCsm8ZHR8Su9gZx4BiXTYU0n+EBoSQNnx3+oFnH3KGHc4rGob85FAxf/yxthJqtPRZ
UnKb8kXEXkhPQdfXxIsgx4+wHu2C7KOZZC/gN0aXpLFmSRjZSF0eQlB05wwkrO3heU7TEknfEfJL
KNhGL70Y9moFeP164MygTswI6CpiJCt+HNjRpZ3Z4EyhamUS9vSWdcSr5+Fymd/HEX/GH4LWankC
8hqRnawYGr/60TdduZ9VIj1gXz0pG2luJkS7kX9OCeUZY8VLU5sKRxJ3kiyhLGbhQ4n86FYJRY5U
A9fHd2p3i+MTbzQWYVUIjQA8S60y+jxEf5fPXbrNWaPOE4Cuu/Z9Mj4RCb7PU+GCRxS2f//lEhUG
v5vNNxW9KvQ/0+JZTEfbIRCHrimPKYqbjpb7cJppPS++JMScxiQah3KwReyMJLrPvuC+91YlaxC6
MC3Qpk1ln+SHxO3jhh36DjxGMfes2c8OWJX0NT+U0pbDar7vQu7E5ppYE2/9CAUV1VLV9zv07ygK
KgXRX5EuomD3oyFJds/nxPdLE2h+xXf6J88BsLeuoqNisU2sjGco87Fy6Xm4LWiUQkNAptHJp5Kx
f2NGaDCdPp2cvOFOHrrkEP3aX62y8qtxN5Mhv8gV9gJxh4LetDa9/f4QsiqsFq+S4B9g8qsxCNN1
3jQjbPuyTz2+W0+LT71Xg+fQ2eGlUxiSEHFwDGVutnsWKxg1lHGCv1uFzM0X9qmvwrl+8B+hvjsH
iPxuarTB7uZpQ2KcVSAPn1TMXomAbTySkIzmVL0wGGQDB4+agHeb798euVD1g817BpRs7GUFi1a2
ztNXOVVzww6kJdpMTQSZ+smtGwUDv5YIWsE+RmEU/B5vReWbe/5IdzIVsvIHp0J6+dQcpOp+nmT5
/GnhUlFrknMEoTjwpVWcU/Quh/N5/AQcc3MEc3ue+gUPmH3/Tv/l85aSbOWqLaGWKQmcB7fY0dLi
ZqYacYXbGZfxoUffxByorFDGg/Fhqzg5PDxYNAKizOEMGHZLhGU659GzgUMPqiJFXQNSVLrS3ZCu
U7yMwTG9TeVySg6n02DUB5iKSMhehZC4oBA7rsUjWDHg/VorHEKY5n7zG2h/x5q+beB63ALKGZ6Y
kAsULlBtG7kcaIEcTw6l7ljjITsyxRkC/a+HqB4V2WoXsyM/4MDcm110gX0qXgJtkie+QkkJTE+d
+8bI7S2NA4fXi29EO68oLu5jQWW7AkIyf7s7++FM319QIL/MoWmtVtVAtQKLGrzHDjoMlyLGKEcp
xR3Fbwdkx7HbVfEjI7U6jaCX3vdZdGMkCQsHvs+qh02FWRQqFl+K6PhDj8yeiecEsYrrLlYin+aL
Ct3RywMXcB0sFzOIPi58Mf+k86B1+senZum+VtQUDsT5g3JtND6LSkTzXOhcv3EgATRdjNw31POz
i/70PT4Y9G4MqdR1sypR4dXf9H0kDHi0FAf01DUAuIC+2ukoNrwFZROz1rigGMWlj9xt8oXqOc4S
ej5phvYeBgDGr7zGEwkSCJuYFqMfCrr1BmQ+slzOzCqHwgPrqNLlBjXsOgr7EAEhY6AXt8mD5xlf
RYli0QpJPDER4CudOUdvlOEmaxLwaEXr5I1e0Nazwkzw/IBg8EHMdypm4ynweKbH9Vag5wTQh/Ia
uxYVd09Rc1HVUPP4XV/f24x0hroOw9YQCj7zK0LJeXnrk6DA9p9JW72jz7O0GFdPV9fqfvIsEV3T
cGpKPYil3fm5QEMabC3gHctArKHZ15wEUMABNFGFR46NMumvRSJsoQ0vVGi6yLuvyAgzQsf78CVZ
bMJXaehWYodUZFMpJWoMhdpKS5bUW7uRSCWcg90Lmr8FJXJJnEpJDJu+9UujbaXWrvS/HSV3NU44
WyVEcqB74qtjKbnvdgi7Ge7AA81ZbB3XIqAGDsFfX+I3hBV5z5pEpKX05VrhwNRwKcjxT0sWrwpQ
ndA5r3sLEWK6HRxfegNY9+/+00KpofWAcpJAdppRKPPvhqRNBMFfEEXhPiIrYfCFxToE2DZ1Vg6Z
hRYtx2o9DpjBIU7ocA4703jWJVnmTsQHVIEoNWPTJbENTJVIoxqmZZhNupeJ+v80wy+OhaFJNYbv
bl4iEuJTgv1xESm1cHDxjbInFQQpTWWT8G6cS4RiZ8hfx9tjgQQCAfFPWG4V3vTHcwq8NCRlEfa1
Ku2I9Pg5XA8V9kSfYWIIQPqmUFgpBwmJIFmdBznLe2IFqybPVHYGYnuIH1Tja0CRBfXoBejaf2+9
cz8mHD2ZCaoVg7kZytafPg+2suNHcfOrYbGTnGtPRflCHDwV0zjXVGb4guC3IurHwpsOwBE1plyG
5//CPq9yBYzF0fpedxG1EAeIv2VRKPh/kpSPJqri6ys6efzruSHjrKBPQCy4JjvaDwMzvabV4QN+
XAPcvDzLd378s2YEv6aNkM4YjLnAtH/iS/h7+14gsgwoxyNLqlMcNAlT8ucuNkaXxdAvk6wCyHMu
fQUdD46s0FhQu3yJlxkiZqt0LZFhfs8O9ocOO1YYmHfDt0COkY7PQySw47Hjw/Tzi3Jj5VjTe2di
gYS5i4oDQUOP93UuQJbDRVKHZ0CmjnEtta67tvhilUUi8DZ4Ug+alcitGjtZom0TuDlYakvPqrqR
2Sw/j3JGiO35kSvZLj7u46/HXoyTk3u8HWj4X7l0UAFjsxrR8e3e8NL4XuRFBGQToKN4dg9QzgIP
VSS/NtuQRm1S4xedw7dU3/Ayv1iTLLfa1GwzQ7ILBadnX0X80ldgEf3ccXtrYvmzbXtIPLAT2IQ1
hgliuQN7V3o2jeP6MrFmeJmkM7vo398K1BkWA+cQHAoUNkLZ16j4To7D6L9giU/RG342mJ2Oj2WK
FJQ7hPtjX9nvMW7MoET4MkOGlcXaJw12MS8/79M4HRllO8mQbbqAAWSnrMull0rcwzE8h3W4Vm6U
uHcw+1gqBYAEKORIEPjJ9Fw6b9/tqJ2l5N/kenZTFIUhd0xFgAT5ovIgQmL6igAJaHNC9gNYKxVL
M/khfjoYMhLvtYHqfi8MzYM42p+MKlFyEvJlvQNeXFk5ewJJaHfYAzEgkRf28nAxhZ/XN49lmNTn
1sozfjDTF2OnZq1s3PhHZ1jB43zOClDeKxZ4IP+gCzwnS86ycKqG1QRQFYp4tzx7z/Spc3IfgQA/
M3NyzdfuIf0ZEwnhYqX5LfU537QVqipGUBpePkamtPCJ7MR0I/rhrAKXMaNlUyyj2T3EZJcTe4Z1
/eUl4Z3DHtFLJ5JaBedLwWXIRraEThQvZq0DZ1UPEZnLlxiZl5mY4Skp3piTST/vO2ttIQN643Fv
exAULjVefqotyeRJ2pW78s2wg1PCTPCsR+eJzpoZfePwm1DlCZHz4KBsftpVJQsg/K0vniSeSa1R
dH2bJsp4l5aYi2BSkyL2gnW1vo32labAN+46fP92qFHOq8ziR7uxRb4nOBvnaEzlh2olN6naa6ys
1Oo7nEqH8FFOBXkydI1QDGVESdHeUUX8I/SglmNTZp1uxKclE4VMVFuZNHH19SCf7qk7Vs2cFq2u
y1WamGlap/1RRYck5pxw3oVI1qIV3kwl4fiUNQYxkKdh1d6nZ9YG0JGlLPkKbiepeeTGP2+TvKz+
2y+vDsSnY17QTYGLAFkLZIU/iUu5YZ5ZP+w4L0EK8vkkxN+BTR+ahKehdRyD9eBSZh4lOIEf27Nn
sOHcAft8ER+dh3Oa7zDepYRa7wknJIwkBzCi/OPTzFJeoj6GlziTZsmZubddOPtskLq21Y0Rh0ui
86KRvL9p/3uLbaRUXjo/NKzHd3WaYBFVMq08Z6Na05psm4ob13UfdCc4JdxQg5lInbeM1fhpSUXb
OQ/8oZBFaEJSKQE+C4F8JIjkU5pUi1cjL+KiMmam2i5SRwx0+qMGlmy8opiIFahp6JKfxjd4P6wb
vpsTnAgRp91bw5h1vBXV1WtC+307vwzbnrJ1uCydZFbMeZiYyCSthWIBcw1g2TNNgcgun4f0qwgB
TH7vygEJs26jZcWO83kxOO+HfoObe4PBlpfP9AYAm/J5S3YCXdaNeADVEWavqHsC4jTYIo4sI59G
ceOPxplUpfmYrRsQOd6m32o0KhKXJzkSi2aAc2ipkOiL0uW3r1RarntzaRIOlflTpkOom/GOtEbw
jLJCCYi7urY5QoUpVWhu1XHOAK7lrhVIXudG/ZJCZp7X/6zOj/tEtD93D+GIjMpCN38cAwU5VDsT
wg86+FzpnnWAM0q/pRCkMLNoyIAJAbRqmC93WwScZM1gUexjisEEIH22BuxeCbRpRyVaaF7z6U3h
K8xHprj2JK6q8AVMXftRONnnzfnaI9+VMIRGCELW7GTeQTpQhZJvtBtytFPZfhRDehy5dconyXse
Gbe1w/jaVoBt1ymNItikmO0dAq+94pwZrNBNMp/GW0aMTAL5Y/PjbYQy/Dm6cEI2SEjwNOoGcK1m
JCLK8gKd5iJ20J/uub9ScLw0F0rUjbvrPXKCpB6PeVy7spwTALPnq3TR17cXICop0tHFSfZRu2IU
7625uI82iMSjfXaKtHVtwDApI2+nRfJfPtubYN2fLlpH3yseuVk0Zqrl/NjcKw6YR7hpZb6u6hN/
FfeTgFkx8DvF61IzzqtdWrMT7QuSPiUUutIftILIn62WSi43yJWZdc0iv8VNXfFDwxCK9PWtuOLM
eBQ5xMwMzynzvbkDH6eGUlQ+rbmmOn6r/FvZEB/3rqflPOFAKHQA9KygciNxO7s/mg3YLM4ruv5Q
cv/nuJAYgIRFc6Sy8x4V6J3QUBHn7G+czs3vlu9wAll7GSSl0O/slV+29QQSEnNgpmco59JsTVuU
JHHYXPlyrm6cvpvT899QrS6f7ADxbQMebbEqeac2GZ3td/sB4vz0H0CJldzipjISX80LclL+Tq1l
IzRz6t7YzSwFBE+dXoTfxLaSsQsCqk4anlEfNI25Ro+jn5RPEgAMJ9LIQxa9/s6RLIesLAHg2bsW
zrUrgvg3Tyw5hyJCZCxDeNoBbIpXM1ce1wJsHPgyYvBppDkXloM3KCz8QP+7I4ZAdw8Y3/hBJ7r2
XRxi7W9QmMigWcbZ6to9BDcfvibjYRZ4NE0L5TkwdrL8Vimu4y5okldQKwt1Nogm/+6+CyMqtTxq
P/wsiaaOggnWQKETMb42eGGabvooLXA0u2g/gVqZ693PzT0+8akeMfVgCD7aXtxifp8c07m4pB5v
wcmYEDOJvFpshYv85DZzo1oiVRpK+IzpF+HUszyqKVI2skpnMbSrwm9MVrICwTLjaSvbTFV/xtOV
6j7P0a2OycGTFih5qd8hhiXH836+IsVhuCK/zWT4MzN5qIM5CSzZoYs/z8N8YNmHNZM6670RQGWS
Y33kHAVpK6NJesGR4S5vZEC94ZqKeaKBzdBX+fFUn3HJYx0wTUwj46HHueHF4b1R1hSPWxH0/9tb
gfi8QqzulnDsCYQRn0gYc1cgdaz3xIIixaNRMr4/YB/NIoKxbCgoUCUqAe7+6gL5jjK9UYRBTZuK
F3dHMuxXvrmy/4fbEz5sWOftfkTMhyOzTQpSNDdyleC4ttFdbDljb1YCVRt4UaiKd/NjqjO5jnnx
O2esiYbycbkgJ9vbv0ByYEXf4DWCrlba/t/0iVX15dVigkr3m0cmLumfAGxBrlc7VxwEquDZRRUd
yHlGxBMEVYqaduu/uHj5wueQzOa8NBoT2YUkcf+/ZQcs324b3Dte7UK6z9lGaJuzoXrBL+WVhsY3
kUNnrbtA5AEoUSraQUOhJXyQFOGiHx5wT9nNwQS41iVN6ALSMvSjo2DpOq+yYW5XF+jtsd6oMfkP
xSu40Qc2m4Kdv9lBO1XaHQkKrF9JBKxGfL6L5ovcby/NerngYUB8oMN7mamx4iyzdB15LoHEG4lP
MZwW37HL5PuHzWln+I1+eape+cxmP7ErwNxJ7Y+K53I+JNUQCrjL9MDdPMxyd9sEbUSP0jslXy8E
EeduozPSFtdCRwzL/kHhKCsKh6CRv6GO1SPBB1pwBy6wOPJ7qc64amAfEOruDXGCLJ5/Ep2+32ft
9i+xYO+yDy3neeDnswCdDfmPAMimu3zpBROyGc/rJExkAVajNQc+j2Y246j1FVMpP6rhDggt4m4B
Bc6858qNHd4U/hfNU23vjIj9QLSn2qUWC0+rZ7h1LWmXA0QHgUXncl/uxTmWPKJVg7w9eUGxKqT8
aEHpmu8WoBYjAhRCSXwfrJvh0DFwQf5zJ2e8Q3EMQY6Nm3OYhIhA0BQP1QrFeB92XErCcqMbqy5R
WoDCcp2aJ4nXQqLdnH4sF3SYPOJgUHva0OjOhYtBSz2uE5qIm2hs1N2XXu6MAyeHYFh2+LPTHMCc
phe5+9/l8Pu3G2YAObuJYyzYecmZTNx1HMf2ko8hjVV4ZnCKEsRYE5W6QWDkSZWSgBtbeVXbndFO
A2iqcJlvxL//m0b5nMpodAERNsC0qbJKNLhB+EvX/zo3/VVA55Mk2kAPziP9KeRKOGHFUoQPLzp2
UrRmczW4ZNRrjvu2AtxhPOowMUQBgjpTOi1H+UmA0cpdin82ZrwQVK0bbjhJJnqj5XJwRQOHVxjM
XjT7frJy6y0aynQAK4B0d+162b8r97aP1Eld2647OrgWSyKYSjaebOeVit5Obu5VtIHyj3/EuIDI
xzkG0El4O07bp/oUm4+hGOVKkSievnkcU9ecM9Krbx3HEqQEu80MEF+N6yquR7gSm1tXcQ7Gk3xp
IK7kPAyfINJpP7oy0lAH8FoeLU2BnncK62mf8cuA0REWCKTi8UBPCw+JyUrZe9CYCUBgD9QI89s2
jV5saelf7AHSHw9x8CquFzrwOynB/X4Z5PEDG6vwWl7L9kuvj5VkgZSYArT520PP4XMFBr+sifFc
3QjdqV/3YwJg/vnI15/iXo/paPpZ066HsE1GJHEgRjy/0hZp7VFpxi5qdCcT6AE3pWmKs4Yaavqv
AMB554Pm9doSmIx35zorbXnz5nkLV1HsA8fnBKS+DrG2vZmR8tuI4oYMipIeQrt3Fe/Q45ZlmZj7
jBgS4rPryX1LZT9x4slK2oQoNK26hLFoMoSbX1+uoWDUDEnrdtSLmKUGOLHD+Kw1ZK9yZXgLruOl
CKQNxsoP2R5mhFRwIXmL5RsVuZxrFATtrERk47Jlg8KQhZbqdLiONBVWwrnmW8V3LkzzoOpGOhH/
AKuo0An3NEU7PB+kM3QyNXNPk5cbQc0K2O+IaHpCwIlLQklhAx7JbjP+3dHeq3bf+nFNOwp1Xh1T
KHxfrHm3IyPe+rm5BpAQj9MGBVqi5HI80t1XT13dyJlaAVOUMG9AgXwYm3AMDTuSu8+O73IaOK9x
x0Kqs5D5dGujxQBR6CAs7jtKkFcV91AY1ynaU/dW4QvO3XXOte0rdxucPwjjSowhlj2c6y3Hod4O
3KlNCwVLzxP7PGdvSLT4x8lJhvQodiTCUva20z9JDj5xua6b47AUErkVSD+GIMCFetSu7IRuB7jq
3f7C32+58TqT8oMFLF4UgMGy45qcSgCX7TpBxjmVmoZDIYNUxg7wrTy9HBgheWEnroHzTIbP13CD
7ACTykexY8oTseHiT34610HYqPcPD+ct/XtaSrjFJe7DlVCrBsEsL0WEnc1iccrtIWbaNUYvqLNM
t7UIY9gBm3ALXTp5X4nqZ+UrA78Ra9o4e34K3B24KuOCV8d3arMgGE5CT0biNb2dze4SIsd9Um48
VwuNLi0TDS/3mf599rUoNzp0xetVuSb1PpOzuJbn+TJDog/gPdMSD2q4K7HmximRL9vKZNHmBj3h
UVglOKSldV72toMmG8MFD4FYvV5cRc2de4MPrXEIAQcLLHkzBM2R1LzdkZS7gz1+7uOUTxNdrgob
wLLwuL92HWqig5qyrstQypnSKDb+OaJyGiBMm1a6RoDesqe7iXytgImOcSuNJKGLigGeQtBx++95
HLCddpFjlJiPdaKumcfhqvQWSdyD1qeP9vHlxKcU2wmUBfWErm16WL6FduYXTyGkOdRKr4Dwzohy
HstyPnpkMI9iUMcXEG7TpclQOk7LFeozLwAh9AOJZ/PyikWcZOe+68zrIarp9KOapmDmcjIzSZzA
VfqJtmuA12VNTU0y1aljRteJkbL2TFgDozfG+v4iOFo1UMYvW61bAfXQAL7r1fLtwpOCzq3v0f15
FI06A5MnHF32ryrizpfW4PjS7FSpri3CnZPWaCgkJncuZyNoAXyZLUBV5oA0Ms7Qw5LNCHjb9f2Q
FTtp1lDv5viwcrRtwXIEB6vSgd0dVSmG7yoLsY5OkVV1KYoCKIAM3Enjz2XY0cVQPGrL5/IvzLXo
ijy62MzKcpaeCxEGSaW88/qIqAHfoDFuljiv4TemWfuF4APeKwuiEK5T7bMTyb/dr/Hhx2awPatD
aJnPMPr8w0VfxVSAHWxRvbH7TOB9gSuEMMzSK9uKknbHXuF+jK5iXB9BNs3kHCjwyoFtx3ZssPvz
rPRx7DOw+jUnScyeB9dkLB8XhNpSOx6FKUxkqmjXpKtwHtgvsX1afhPDX7TPSLI7NYmFt7F4WmCz
4f39TxHy3SQAt/hcrCNLcJWJ6BgGmYPg/PwWjRkAnAXNtFx7m/FFDkG/ttvC+7ff0ifaNWu6elAJ
vXvutcluoZr0pYwDFfTDcRJFUMRvvU/AoB727fXOdIVL6smPjdh5YR9cDvPw8dO6rFBncqhw/f6/
sjIc6fzdWjJqqF/CzMdAkHQ+TL0HcPF3YnCm00G0kfAzAVmVL9+tjScPod9oAbXicPo+C9JlRhEo
XbNJ6KzNWXKPIrPhV81AW1ow8k+QD5coT5Uv7j+VW6Ycv2X7uIYhiAi9/XceURcqpYUmIRURjcDu
klr+j9r/ANRWxzdNr/dx6yBk5IrCpfaRlw+hw0WDfiyohkknMTPHcy78870W56CTZYEhOjIklkwh
mefQnRnYmqhEftpaGQBSiB2ekAXz8Xnu8drQGxZGjtGSs3OMNOIfY8fF2hOK3s8VSq96cthyxnT8
YWelCn57GuTxEhqf7QiL0u6d+aH96QR80SBLo0LK7Tw0iMeELLugNQnV6OnFxa+2VpeAM7tAsJ7J
wNtDNDvMzg0kLU6cXT65MkovM0V4IGRxA0ZqdL3ooQ731eFNF1srQbM0FROakwUEHTDH0FiDr8wP
VEQApeLrS4J39//dMYtkJtxKD9QLaXa3EzYhK34mweyri4OWtoVi7uvFAELalEL+ad1k7U3cRsrW
lnhpwtvg7LVCOmwjfwr2SavncNuDdExLVuU1de76Nw0rc15GZukqH8uaYS5LBnhIx7+Mg+MyHqzx
H599A0XSCh1kKesdAWHW/SMxTinDe3t/uMhLPCxJtbx7Q6cSBQA7+mItElPVUOU3C9p+J3Oa986H
U+cJcaZH4YMoHkg1vhPCuj5E3RWIqiDW3v4ZErIw3RLMc8hXUe64B9f8VFCo/EGYkWqPwMNEO3lR
xwOucjXgVp5G/q/ZmknoJuGjQEILC7eTXWaYJ1wVx9aAAdpoJgRn1Q3jhVEUi6MhVrZ181KGtNbs
cT7cLb0xzhymu4JtpEsHBZ50ItlGTuCM2UHr8sdzdAkAtZ/ch915zUyC9AOihmavN89r642NhTKF
9PpWf8yGpSmDTAKlaEumxBPVMIDVnzNd33vndfb2qgQfy+K/M2ahmDV9NqAfQb5LStdldWr9htc9
Xg0U4Ih26/YAneBJ7h+D1PxWwfvFi0/dLABpHCbxtl2OQJnRQY27ds38XuoIT22VHgsvj+i+x/ph
SUS+AnaBXRlV518yYYFZJlmh/WAP9aSSlGBSHVC9Nk77vxNd4J+jP2L2WqGm5zzD4U3hHwpR6pKE
n3XZINlfoyms4I3xrI4RM1sChQ2SEBOweFgJzIgmQGrDvo/Q9K1onQWpeAia1VtQdd1AmncoGSOv
GLo2UOv5EI/RIm51JrnQuYXj8ZviQELLSCMIG2y9M/sEp9BUXnrsf+MMG3dekI0gBXqasIU+MYoV
H8bxI+qG3KqRsqiwY18jMk8lGETa62sbiDZojkns1bcWsTzqDtuc0FuE8pg46LcRAq67lUozVxlQ
5dzL8MhWZIXFF5fG/KHvGIk0iSGjgqz+A5RnpGa0mHJnNpxel7TWMAicjhvnPSlUj0LSZKUSOnLW
6E6Pz+/FkuQVFnvIuw+/DmNbguZQAwR1/zPwd0jg1lufcS4MwgGk6abvs0A5u2lyQq19ev7nRlp1
/Ek3LUtGwHkH9wQoKgwg+DJBHgGBKjMluPxAm9xSsCjUNk1Lu2m6XperN2BqKu+/idPJtHnQHAIA
+cfPxCaEDhSa2rh/lmcIU+LKHZ312zheE+E6tW5rHG4CJoQBYCBDTg4N+jWW+Z3DmIcLLXgF23bL
EWMVETJzcN+9D5YMQx8hrnj7rpHKrVTGSJoOErVpTO5GqK2xRmQBvLQt2K63HFAuM8tHKSM2AxJr
Imn8cgJhecm7o2D/azrwTN2Rjc716fyIc20nyx/FR8h8diB5nBPa7AAyaELkoXCMni1OJrKuKF0v
wGQpCZIw49xDdSdMtdPYkzvM1BSIFUMdLW4TVntridT9z2LMEql4uM8Vzq5ThnwIAZ/24OSKqvmv
XVLcr0DA/uNRICnAzyLOfvSXcr9QHhntLhALpe98GpOB4c+nOia4WmeX+M1zhI8cOMhc7z53f3Pg
6T2I3PxXgHhO67VR70Wv2VCCa099g4v/grhYl2U32IYoBNy+71UA2KTy3Md7wnXKUX8rdPUPCxhk
YxPbAomD7vbIss/SS65uMbQrzQOzfQRgyyuZK3tGDNhSWD6WmUogO+8aj6UoDRZN24XPIWh0wp2j
M2EbYHJZbU8VzapMkdNyGL9x5NO5X3EtPIMBQZOBQofzAmCAP+tqfULpJTkDKG+/NYFLX3KxI+F9
rPPZX0afaIrNpZLNTlZSUjgFDcXnM0KRiIYwu1pVZLXRZGUQKpZ+F70D69ts9rDBM6qItczXJ61Y
r3pHuRj99L1nFtCJFdi//Pa1/gSH0CuJCnl/dclT3tiX5K9/1fWb9QWxOLNooAVnTn9FHGAvxW+f
unUT1aLqeTxXKuJiZeOcq20la+VOBVcsleNB9+aJA9o7cKTmBNGFWcwPe/TKiuYd6pjP4dVhC1TD
4wEGzcdXQEdyxxXo7iEs1etVYs6nhs6FiRQbALP/AQnVmuIWQ2yxlroDgISh1yrJSbm2AK/dhegj
ra6dIEC51jiJIzmuAdfHikxbuAFegSVBRYONUr25NmGmHucGXwtsj9I1I4TznYkJivK1Pxkz512v
+ZHFALLG5zNh+vQp7zEd2BNlBUQicj9WCR/f6cwrk+8X5LjYK5hF74suIu9BXMdVci7XKybvxUyx
fOhixHhTpsSQyOAO3pTJGvwNRqulFRmikUTvIplSQycSlxeXLFj+bvJRpi31I6rjrTHWxvcvfG1A
yXNQsVQbA4YyTn94YGZHTL/SwUEzhvSz5WZS63zGHpxpYPS4h48P0UgKD4JYk3W+ayEOXMJnh4mG
0sSqxqVu3u/qT755ZYtn3c1CRL48ecUPFSrpcxi1dBqsoEzVh2Jq9SVX2cmA01cT0VkXSdCGS8aF
NH0raBqbK0mrY+wfEC/0QGaUXotdjm8VUtaFfhicHpQHTmpjLTy+8+oTLi1kTSR3Gb1St/8Pza/l
MShz26K/Eov+hqOdZycZV+vUE3xGpe2Bssq/lzbOo3dFBoYj8PnpRWRS1BS89O/rlIKg0NUGoz1s
lluOk30E3ZymEp3OUCrsAWjl2Hz0NT98ti4/SOfsg4p5ns8Jqbuq8AkW0PNLRKu11bK/ikeHgr1j
qx7OdkuIriVC5PWfsYA9WTFJHhQspZN5nADlKKm9q5zzBUJ4tbNNy1NqOrH+fPNUj2sOarGpw8r0
UYgN4DY5lbetSu/J94etwNvGwXu9b3v2RMySn37Xbknrc8oXduFit23IhxSbbfjLURqkub0wzZTS
D8KEYrQphOAb/a6P+gRzPwJEuK6R1mK30f1AvosBYm+PYBvuF3Z6yNjH8s1m7Vg9r4PyjjcFDCb9
RsV+jQQsgzHElxzkrEbUhtyZYUE+EHEsjBtc3mV0Io2maJs78OqqauVJdWnrPp2Ulkom1lcrGGL4
izaoLNXQL9EZwoCN0JAKbqWFuIWkP1Chc6Bw6YuQxiqJY2XcTMMJa76RO3kKaxibqVm20ET9JJhx
0Cys0eHb7Kid24acbV38QKsCkQhPTpTQMqhvVWr8SAebVjKRlm0VYOktC87bXsT9fNxSFbOSteCF
j/zbwr5vEpV8cWE1VFPmHExmxl8/ggY2jOOV7XKZcgZIfauKg5VyyxUbBJNjUdSalRYxQshNhzqm
fpFO+uhNN44Som5uj12jqohGmichwnjREW53hY/lt1/i8k6UlAw9/nPE4EX4r6xuZRqwfpBmLIy4
AP8WDepVIUDegEtFsWVGw8bw2XDEYYmDFFyYt7iAf6Hpj3FNakqFms1xcsZ4hJN9z+sPzGpEPt2v
8aPjKujHTEQKa9gBCDc1l87k/Zj7Vu+lfuzVidkVdxyp7GlXAhw7lLU8gJ4oqGVmhP9VNwMmGN6o
PdANADfyI9NG/AsSzzgGsf28X4W66X6tRVDpR7v2k6jV7v4UXvWK2+N3O+z/EpaNQuKLc2oM2k+E
cgIXiAIMFioia2G7Zz9BbOok872s0zA3QHQE5//8c6xBLHbwtkg8kbvtJD+qPcmzZSViJLNT7LrQ
YZbJuerpmygiQXy95Ly6MzQUG691AN2/RtrDAhUyGQdNg7uW8AOLx7TwUmfN4hDeYM6Pu3bY7B80
848mS0HuNROdcDUaBSZxT5ulu/0YYfrwnsOi+BKDjFWvZpoz49LzihpdpEzORuPip1N9y66H7Aex
rZpRWqq8J6rsFAbg00BCqTuql1w4kLn4W/FQg0BpleL0xchrqOY62gHs5qP/7+hWA9NO04y2jTaT
sGgzCnURVs4k9XOWmXRPY7ddTDyy9qlgr3Re3aozzHxdznee83dF58gG3RSdtMroZtYQugVNSxYd
8zfSCac7LxgNPDPl6XYbZtFFjUsbSt6uOykTRYaqWHn598BGlPpT7dEhejjQKjl2ICyFnMW66kij
YwhahmI+SkgGeFrIyyLHNKzpqmsA1McOs6tTY/OpG+b0Zn41w5JDw1/wRRvYk99x/MObbL1c0zXo
zsUpIEM2kVAHOYMO37m7rfBLjdlN7EQYOxyRVQ3NxGaZbKMIvSCVROQCVbm08abtZh0p61D1NwHo
rf3Rpb58GG2XJsVC4qDODWac5Ep0G+I+BXO78O7dF/CLBQE6GDU0WSbd/GRYZSgU2xxEbWQOvVDp
Ey2R7uw3Gu06qOT2rL2A1V6IrhW1qq2EXdxf/EiCAg1E9Ac0zubisl5ZklngsBzGxBM8gcQPWQBL
hoojj3s4Q6lQmrj2QTqbU69m0QK0nu9+xO3vtnxyF+hh5g1M/FQC8O/yyjspfXHKGnezq1ajXjra
8w//IH+E5q56KGxcfZk50VQuSV4/MSref+2yZPY9eN8ybIYOcbxo2aFjykptUfTVFYfzdsNevxVn
6NEX8YrLs7BDC3ryeHAG4dAKUTjx0pXlYDEibbIckFlX6hvpSuq4BASb5MKUg0aYOguCXNgnqfRS
hlXI9xgnJSZKvOZZYT8Y8r2EXwzwFCkx0mGFgtOb9rXGK02/OAPZSe9Ar4Yi7u6vsdZIA/CDRZ0m
OYX4kVIWYhzWGmFCTDMvGwJ4Dd/TGUy/kYX9P+k4eoEw/ODbhh5Ew28f9j6U/MOks9tSV19MKlYl
sKPitSTwSJHzypTEOOXYIn2iGwX82vBzpNECBLx5UOclXiJzGCoHNvRbvngij9Cw44HqgC2Ed6AH
1zhQyu1/8d/zLRhMQzZMPgvqug2jLfOuMDctif+FF4DFbuZV968eFhGlU7L5dcERkhmam1Eicwoc
7Ga/jZQICchV8riJjEiJ/WiviwZYMPkELDXij+IzHvcMkNn5cWlzKxCV92z7K2KVXXAEzfTMI/7j
CG1Ka2uhsNHFNSR+/k1MLN0BUHGJnGHxanLMWIY3kwORNr3yOSTqojPPVIYjHXTp2doin4dFrqDC
R93liZ4hzLl6WEXfDkLBXMrtOcXA4oDoRn82efRXNm36ChUVkU8SGfZMS/fOR++MGBooXFNfebtg
7+GyGu0I55VG17Ojk1kHU02sXtjMQhGuksmWnxzklde5RS/nGtpwV5bsLuqK7iMFudmhUFpDVXyQ
JTFYjFVXgHkLcSfxaSVhG9suLA0x9JhEch5h8tqhRr5Vqdpl5v/exOTHI8QYMrsliuFsWeBV7q1C
hor3lO/wWRjvChTJBIY5jj8CFzpisHXjkdoQSWmmar9KxGQB3k7RziHoU7jpLOX7FS6WzVy1fKSY
/7nUqwUr3fPYhOFgO1qJdSXkNqfyM7bwVSwloXcEUHK2Py1zF8TQtdjuve0EaLGFYNIKdhmu5qcd
wxrSo3oWG89Yk1muugMie/LsUKtUQwvt/CiqzeEN71+jDpJ5YfQt4spL32q+d4gg1p2/Vtb2eNd8
FAiy89LG00Crhx3a2X4oChRGKqEOpTT1siHfz9cy2Y3L13Cm5wEtTDWTsonqhz3Q0b47wH7vk1vo
JAVjulVYQcfc3lOMg3GMtU9yhiQMXoJUPwohEzBQVWtImIQD+9WgsUWk3u7BBXFydLtulQOfJE2f
o/QQwbVzOS1cfokur4FGUzyEceI7CAOGfrB8igjEgxBbB6HDPK7qiI8+Ah444U3aTnP/4UouSRpM
vdJdj8c3LPm+FpBIAr+VQqUhW1TWTZ6Voo8MDUGtsba0y+L4HlBKqQVJjLgW/lAAtJyk+DtX5+JF
Y+7GTY6eXktQBc5hyisAijJM4vZzSk3Tq8gZyGgx09ExgRc8wHefwLSmJ+XCS1stR5ODdR+lal6k
Xw4lhBbotEF5kadK8aHagd0HNBsNL0xsiwOQmTwSasQcdFALSkYPPUMLKZbP/nPcHMxO8tIT2wpA
qIZzx33SzbkMEWBqN/d/WAFDnJKM559v3u3RFP1nVlWIMg1md5puvNus2yrFaag2GXdkoSbfph0h
Kbkm3WdWH2VjMonIncRYl5vqO3vIxJLro1zuI1l+Av4kQyOU5FcRGzIj+sv9Bh7VF9tZqhccxAPs
Gx6IIHozS2fUjxWBeQvlJUTFEWSOAVXHerCBPUydar6ltPYsf9hmBil+E4FRvE8djrRmYjkRHNr2
n5mZ2K44UmD7AGmVNawtbdADCT9lVtoCLMQGBr0sg3gQcOAl4vYoRYy6dBBJbZZlaRqZtaEanOVE
ZbrIs07bAHqNiWAHnqPP20UNNHTpwnkjyYOIG0qirKVDVfURiDifvq+FB6mdmiKOE3qtuxAZPV6Q
tNL4M7YglmWJLzf3T+1p9j+JCgu0FoxHRN3V9sHWjhrT6CaiG+c/SRXFap7C08Tgotd1AsMLtrio
8mtD8igqVS6u2/xKqec0z4jMCSTfbJl8q1ve5A/54zEG2pDc7oi5ZlxwEcVCyaiizPY32Ue+nZLC
xrRgAyNqoFmlUr484FZ5lXvP45Z86iTRkr07imCPiVzieA7pTmfga9x7yHDFbrMx1OYSIa4fFKGh
VFv8yDjA9BDZ1odOTktiCaR2I6u0liqxoqvDVTLQA91ghJEzCsXgCd/o63C3/TPPiouvVg48cgV5
881/q5zIt8SNQGvHLE0s0hekNpvdcSiDF5tZQOnpuovlxVO22Q16jANvI3icLKSsnK24WJOpTbt6
D7T7LsJIl7ULdSe6+e1F3tg8XQeH4zFvjL67VrufzvYWLbuIrkb0ffG/1w/GI2OM7qntuX44y8fZ
l9YY93OKU5WsjVkuN4LVz2Iz7yQVCsvrOA3YABXLAOvVP9wZfiIQJky4lGGyvKNHZhPIOcNjxysO
n0Q2zHVCv1U4E7RObt7Yn9Gv8b1Gditxoje+a3OroQIs0JjM7YafzLfomyhbA1MMlVs8K+BmOUBq
lDyqiJwQ/ntWJ9jp7d5BpKnUyXbHXQy9kEdcqOmLzBFFVmdmd4RB6rY613dO9SJM2copPPrlKfmy
t4YBBu0Km5Dj1eF8Q0cqQ/qVcefLZBQ5cIjuDEZtoXc7b87cdY7SBpjKF0XrkRrl37pJO/uhqA3H
ETju3aNah7YgiGd8P1V+eO8p6u9q09nofT4DMragaPiORe7ZZ8CTNZndJ/mrnV/xO/xSe34jSZlH
ELSQS3z+kYUPJqA5o6KFhYP5e33Ob1ikETtZ7HeMeNSJBcNO9llUW8eD/n4vXYBE4rmWq41b0gnv
BPABK2QIfFf8h+/ei4BkuHm0pz1/tS4CknK5HN4T6hkkhp/GK8asJoyhcK0XKfQ42tZtIjN0tyBy
pqXLKS7fqUf7CuGgWuRvFfEPLXiiMNUmJKvoadphGbqPqWaPk6L2rrq9ZL5A/Ajan/7iO9IEMvtW
IL/s6M3zQSGllS/fEXFYcSv3VcncMrOeCKmUnUk3RgKo/iwfgS286+369wPwh07elHFqL+zJKnMB
RWMSoOEzfyJJzdAh7WcXQZFdaMOgWj4LN41ZPx7wOY8vBxR0v5cwTwxZx6iMl10OPt5tHfXIhpoL
4x2afCZZDexZXVLoqpPcun7/oQqmKRrRPmlDCrml0xhPJNRknhcMQuSp7PDcRScvPh5/CJM8Nh8J
INJUiOYK6Gqnc/H0AzvRLmks6WEj6aLuVWGEaM1ShiCVAcRk16lkJgPadb3OG7fmX5IB/C7Fav+V
dlAZSGTI7bsdCpqQQPvvrbsclk9uJnW/b9ETvP7n6BGOpyHRZxiReqeR5i+JQq3D+jpksEjQEbft
+xy0gPJdcTjGJWs4ppXx8u/AJva1RayEZsvhw8q6Ws1dW86dDBGrgKsfFCAL10CWDz4upoBt4dJe
QAK4OQ5SJ41DpUTu9QwR85nooCwBec2n0y6hSIbRoxj76o1oX+R6f1zYCwy56oFmQKfQPDy19KyW
uGtYx1ts3PminiRzBymr6Q1u2Yy7sQKpHxayLX1R3YhB6/OdT90Y+gnyGkY+x1AMb/bC1vA5agKi
CDHO1WQxk6l6i33s2TA3JrniotbTRXrvdSgQEIJO9dFVpO7LXbYVWDUZem9dzM9hu5r4bJHotyZr
Mu5B63Q5qH8TmSXec0i0i5VnjruNlFQ1VeyrIeYsCs0Hhdiwl8+SrI/RAO9z6ANRfgyxfqhm8qEq
Ehe/2fEp4gnSPE6Y72rp1klzAcMLnzl98RzlbXnl4xB6CNOfacVyolygTI0glKfXPeRRz9qMQmN5
Ljp//yP2jS+drIAriLacJXiPELsaK0hm7xJMH8KSb1VaCqxABavCqRDzcCEFVSGQmhbaOrrIPTHD
cIAXKoEdVf+Kj7DMwsV1dawclRaBsNe5wHxR/BPOrVhkTeV7D9lJEFMCUbEIxB1katMWLmhwWhqM
DYNv+tfMJRDXhTxGmA/GB9EQoUw3RhlNi6t92Mb7s4FPp3uwAZTTljHd5gI+DD7YRhCHKWGT0pwT
rEs1S0JIdPd2DiNIkjkIMo3Xz2rywtKYJZbT2DI2PprTMBEHgaFF8y39kgciDH0WWi6Xl40wg6YI
KZkD/B60Ur6qn/1wJixKwKZgZhRNgTwIDncQOpIJya6vRz3/KpVJMNKfThjiPAcYzOHIHJF1Y7tZ
o+ZbrqBYo0QalmZQfQjB5d1VyRFz2UzOh19hMH1x9Y2zM9lWeKCDRG5vJRXED4SngIqyhtTsH0M1
MHJFDFTBy4c0yIjPBG+4pUsOuFAmwZa6teialUOuZ+S/oy6+UJcwR4FFhA7ORojyrrO7HjlepCUn
niSu7GsWhgx8llIqYno3WtSbYmWVl8j2HAZDOgWA+xANFybKePpOkMIaLx9qS5w8dPwKK2CoQWDN
+zYltKpkzMHYCbOXb2Ob3b6IVlbv1hxrIoMOw67wjmnCGbtKJBYMsliwCoAW+jML54UoBbA3QFAW
JkBxoVvMAuqxzawaCAcAUJUD+8Ea+ufTDAcTjhvm4Mu2vP5Btra11+1gnGyade+wo7NSyWiDFanx
87RMWHyfFaG2L5P/gBV36lRyOYFmcoy2johUFUqCgGIvlIIwQIe9QQy5nfRsa5oaHjmQKp5/oUNd
7/KIFIEpr+Lw8W9GUUW3upe2fJvc6xp0cQVSC5KH7Bhw6Nnpn689h65Xp4azSQ5Y4swgjlgpxHTN
rgjcZW6Zg5bsL8/+gLOl5izlBb8h+hm4AlpXyh+OqKNsxXqFyLzxJYcEOeJqKYtYQ9GGlg4VgFDZ
e0gONztSPHvs3meWH2WSCYPWxMm3QSI/hlA3rbf58e3ftkg4xxnB3N19srBGdgvkfnBLIErUKKh+
MaQxyedXNG9TE0Hr1/EjhNMUIpAMBfTjphfj9Xl88+QYef0fS1VbF5szl+gZ+XttK9ALjvBmsR5T
/jI7wmesDlEGCaG+3DlVb+pMwIPD35UJN077O+8q7Nmpd13TcHqV64UAZDG0R8Lh5FI1kE4kBoTh
6GkBXITo390DgVkFJ3fRE5kDlPWuuP+llnORocq/y1nXAmaJ/AZ6/5KrQq2D39nneSe1PsnkHW+u
BSdrdGuheB9CKeuhv9zg7mnmX0+VmpsiI8L42QnUhUxUUsXPGPt6/zYCyshTGhTaINVHgGXZysmb
GiOBIu3XM4YDLCp7u4OcDqX9p78bKXGRLa3ioUOKC21NxxLrAd/8iwNGMTGNReEchRXebuLGslSZ
8pcUMWG+f4tMWFAuz3Lop2/ME/t0+kJjh38C7XPPZJGaB6WUP8XN6xOraTbXSzkptsQ/8m8LgM0J
uGW6ED4WnjGImx35LTxEVktnzsAry/8hObiussn5UHe6ukH0u6dePWCYajKdl/SShDrpcY1yYG3o
uEf41xXXyaCFW9imqKY6ssbqlAFY79npLePCfCOHvz7spanY3v+vBW2Vr4rxkl55gL6DHSQJxNjr
EuAvIMOH/r6+cN68fty9Sm8LTN6QadF0z8hxb8pXW509CO7fN58BxC5fAPa62TeFZSDnmdlmsOEv
QseRY3hhDq/zBOEtKnwnRAV4es4tP+y+H0L2fDaBcSR7PsjEXyeaFcuczhKkla4ArNHSb6NVsE9k
L3mzFb6JVEzDgITxdDWyPvxAK9dMKPdRzgaPgVyZDXlA3ORHrOVtlTj6KjpgoM14x699N5KQTTo+
TXU2SvrCGh82GpwWXfeezSu2rH6a1vWVeHNDmjs6rO1Tv7MH2jxSplUJ6vf7In3Bbr5n31IrwQH+
xPuohmmjQqF0cFlgslMng7/OxFpKoaPHYLCZj7RTJ5+ty6FRdgIFFx+EF0IxDWwZ75Hmp2e7N3Qf
JlmMI/D3HUf8e/FsxRXOemyMJFv7OwbEaZdj3GHcmVj+VnpA1dGumxwDQVOatfOiGWFtHQg0uOu9
m+iqaoaC5lJqi3a4Zeat73gfvuE/AJq/cWJNMajSEzHgVrP/ET18XAlMhZM8irBiqnGlOgZOCePt
EDKnauGbXMAAWum84wDMCmayClXUTzkc8KWamNFkXm6YPY31i0hwOmgmct4ko1o3/a4lrchf+jWF
oKGE/8VB8d7rqDwATuVAMcy+fBlIJTrB/5klkXzSBx8RNBVIb2E5N3koSizuXrQhM3ILlILQJTFp
1aHE/joQd2rrIcfr5yV7ydo/NiRbz6okxvhUpjRdGQNkVw1qJlrkm06xc+y33XKr7cDMsUO+EPTD
CszrE9S2nk6oLRWrEovwjhdt+lXzEN1DKHOFMVXqGsNf2jZI+10Rz+qOga9L+5rzG/RGxQNR8/Q2
MX38CQij9sL/9Lz5MZmFd4mGTqKZg3nzhyUw7PMiZXng2qIQO6NT/PMsZ+PAnrstzWPUvhGGpM7P
QwtTyb09QgBNrSrFEQzJUyCGJbB4zQG1hueHe+0yhlfU2Oo9ZBH8CON+yTQudXiIG/OIYbpfZUYI
aBRpsAPVU6H06hFBTrPCLiS/sDDW9HrFYqAlJ98/3JrrIkyiIpOrwgFSQ4WbdN5M1eBvmDXc2yTk
Z1OxcFOSe+e5M0mwR4yd76Plnfllx/7B0gkCN2Jk/WT6aIms1fRlT5xwKdD6oj1yerd6lLWtnc1X
axor6+QAy0jMvBYNg5cKeS82QMLTb5y6JKngCbgpBtHDMD9HrP0ikl50+xLuTRz5duVYbSMwyeAJ
Czbfo+otxGlznrWVlftyHeh9x8fkxSRlJlIKe167fSNGTai5LOlGiaEfRSIiMynbUuhbmVfGRkqE
0lr0Va0YMVCSwBkLK6fxXbdawrsKud9lgZPSRYs48w9IOtjbFN6BPyJ01J9ZhiREVFPCcxL7na6e
rwIb7bw5BK1jDCgPADmSP7C8R2hjkq8M9OTgUNd8Xk5sHoYw2+2nAFbKKUfXb1VNiE7MohVG8L9l
xnZs5/wsrQ94ic/BrtZ6CKDWQQBzCsXTOZqsLPH1ysF5Sm8uwkULxfrwVVVpl46e9ZkYD0gJPxd+
HAYRAqQFJe36oNFGedwl+OK14NgksB69jT2tNY+3jEG7gRCPSe2DV+iMxuD9gXstKurOPcZFIbwA
5Cbr1RI2DI3T6NweWD0OyMvCYqiTQr2F/Yy23hwu3btATsmOmzGD/axL1cYExN+eIK1JObKa5YXy
XxClgz24dK/MQfwu98JRyF7NAuIznjG2jDphHQx1/3fzzdAJzluxcirmJ8zBUzHwS5EmProlnkbx
pgvDGQXdQCemh9N9wSjw29L4YH0wPzbemOOX9i71nd1O4/7NUwyBhevbHfo1+NwStEMKFlTYLHGN
EOcWVyKWrRRDRW8lBhnsTga71uwwYKjgpRBMW7FTPoK0SgzZflkNj69a/Cd3xjCgdVCGEOw7F8jI
8wkm8vuYP8cvTHDVY0Q94/RFrCNvik3mi80Yfb8y5Lyswsu8UuPVQvvlgx2ANLfcIBuCI63JPutA
S+6UDeK8T3j0MWNlMEwhpciWedNQxdvS6CjlTr2nt7hsVMt/x7+khba8qBiRAfPzhRfiJLgomBts
gkkTzZrUAocsa9hN63VbzOsDFkyhUirpY9aYL8dUKmkSdwcEutNuaNQw9IP5p0VM8Vmmoy/4yOE+
GmJgIwMG7i0U62UXD+S90PxNz8Zc5NwZGLVyveqqAjMUoGUr/acWaN40JsvrhjuHBvpfX35XtPv9
/aLHWrdRFcM6OWVuEv62A0DpqZcgnBeesdiM7nx1l2nu9dpemEuPmjqg3kD1yVaz78heyhTKgS+4
VvkcTHz418YLK4PBNoABegKSiSWFB9V/viZQmfDl20209iSOAj59YssPFkeSG4hUIDbk9vuACV3H
OOzAFtLcjjserPo3udxVXpZ4ptS7AnOKPwa4TGiOSSYMW8sgEfPKVXvwtMxT8W0wA7LNqW54Cop4
yCAW2C3i2bFKtSUpVx1YBniMt+7NRyUJQ1MS1NTKMTId4Yr8KBWwNOlze03EuVH4Awa6MQRcgXzH
K2Yj+nIZsMNyEaFTecimeFuONQB1xYp2WOB9i3zGblAJOflkSvhobK8loAcAIuC29hIGaXP5wqyh
E+enc7BU8wrpJk2PDjTjAclzEo6IZ+9Kaof8iY4q1xOjXdwaHhtFhhK/jBQkj1B+ylV0Zys3q2OT
ZjfuAvkdNNb8SBkqXsJBolTnoxWuRhHn4nRs4i+wDSlmHUnk6YAN+0nBtpMBS/vDJ4MmAhb/YkiO
Rqc7k43uL8z/kj9X8q9l55DaH7wwEg1lD9Kk9w42MBLG6yDAbuhYyMZBiLS3iqGbghjmrgetTP3r
oVxZKVKubmuBomHvk1cKPVmZbDCqcLPRU/fm4e0d/u83uNtUVmz3l5h1t+CZ724hU+Z4pyrAlI4z
yDk1alkSVfYz1pHHBv33L3EO3QSez/Chfe25xP8aLtPT5fzNWv5ehN9AkeV+qBQVtOic6vKTfwIb
MtQwgCf6eC2Ws1NSkOY43uHU7hFPjL6sCvobrC9SFAQnDiUU4H+xo1ifQiMdy+z+aaysQgOpr8Yf
r6LLi1+Qctd12H36leEhUe9gT7sbKus79jtQSBCnK/wSWErlLR1on0tCmGsfmVoxLAAYkbqspqVS
63tlnXTMNjprOT5W451R87jHr2q6+X3Zp3k3Cj5ot0fzCZtJnwk+d8WfL5i8bntSSb+0HMWA+rsm
ReWLpRu/YmUrwnBp/wr/f66jV6Ai90WLTrnU2dXHTKTNhaJOhSoRtuMH9/tUZX2zAH28kdN/dpGM
TE18sZlHOuHb1uPgOKAYXGhgiRuZ/2jh7gBXMeYQHUojSMsDdpR0pUJwZieI1D8sZRNSVudDYYPR
F2ckhAeOnYb0rtnoOXs9smZ5P/4UUvNR4tzltCbHXHfiKTaZkSemC1yIq4l0HUZlQRUpPO2w93pF
FuuCJIswo/uOj8FEJeTW4hkrLpt+XVdLwbhPK7jINCk8DTKOMIVkdceFs4PTy4WWONUvup2t3Scu
m9A8yCxUEzog3kjJRlpPNemzAAAdjRz1RGXMmO//6goKrWe+uJ2u9ZiaE0FHRbnOgedOIuEf+Ya3
L77ukD4YHGAmHtnJqy+aZMPRCMNdwfTkzZhjG9KlybU/UBadK7F9Wam+vyTLqWeYiai7UBn+Bf8L
tm518peAntiw4T6PRZMOqakYjwPV+Uh6+7k2XDz/haWrc73hH6yRdygKMH1IfXqI5jzQPippOWNT
1wtojQmT8hLvJ/99X+xD7y/qEejeJbZfcZLL4cVe0DTTsWhj4u7GA//wWL4OuiSrboaNMDK9Rcu+
ayd0EvnOfgGfhfiB+/5xloAK1avtytNxnSKEKIct9fMbeUY/iaJmlJyWYGaDBYCq0iLHnzRglV+8
r90PAtugMtRb8Ohl1s9W+SrqeNzj9GZ0RbumqzfTjgS5CpK6xQqQpvyCYO67Cqt7Ymoh6GCmo/QF
RBTH14QGC65gh0c9VZ9x17iLrDPeQMlz0/m6XTePrRdRCMyOb+61VZVp/gofnYR6pITGsacbqpmi
zWQiz1ABkmMXxG6ox6qcBbmIQu+IpkqygJOY5Vn1kjgAIzQqrowm3FTel/fuhI1IJdITnNXkrNw7
eQDHoTxfZMSGb8zoC7FDWhDmzOctyzJ6DmdtQtkWMsKtg85phhnmJgBoL45bQsilagxAG0472e/2
ZFT+t/nRhjR59/b2/F3OWKH9Hz5jcHiXcWwpnnbiMahuiRkdiC+Lzfi8tiIQ2kiFEjM/CmZ5tKFx
GoG+Y0y/c8sxQt2544PQooAA1w5OoddJFZbsVkZLIqxfn+sSegerwjWuoz+Rz6AXj4Lyu/xGyvo6
9WFLwffjzi/Ko7kjg8xitRaqwVjE0k9sxTFhSN2q9n8Vuqysjsh7EkRwt/lz3sci143x5gpukEg1
KeJ2+Zjn/+ApdwVGa2W4YX3aEBd2fWZGbFDc0nCcO4o665vj5TuVT/zAUyRbSo9X6zXy8A7pDvCU
yXi+WYo7+4B/QukDIDesEkhpfoBLOmbVzxPE/oeBhK7WG/NJKQvC8AA0nk2OAbzxwfFcBAPWbLpW
pg8k1KWchOCsWO7xaaoUsllJ6GeiAsKBSrrcLRaHigCmRiK3vtYKfGhi+aq+ipYZRRx6a3nYNczB
ExNUsVX57/GAGk4233+6g1XO+Gt61Wgox5sc2yUeD/fVfZcbmaSkY3JQEh7FU6HPCH+wFJmwkDS5
1NW3FBwobhQIBtlaPWU37EqB2yu8nM9m2fgUXlCGVYrGhnLaRYxr7qP8GqxSB5HHxHL2z6jDDM1V
4hrU75MN3y1Db+Ntc+PKqXZHIlN33sqn60kKOyQbuhbyOlC70WwFs/NDsx4fl9rNPQUQ6H/mR93v
ZxuneDYYBwjwBZZjSEZN8sEXevwE0DCB4IB5TfB9iFz+lEzWnHJcHU6uMm2B/Q68akACjh9ppglH
d9CLJ6kFPh1fsNHtHu1IlVz/MMMoSJjCeuuUxh3hYDpZBsEBHtR/fg+Si5oPve1D+ARMbhUvv5/x
5WcecZFNfFkECuzRWHrVSzx2nJsmVm13LV59TUB/j/YKNkPIdOvV6m6dQCsYbaG9ajq/nkcyw3BK
9MZGFpV9klNYGSJN1OOoVTgH3rF3OEklRHyOFFtnEqSKBUqLwski6npG+UiONUoUkIzmzJMcGmqm
nLSPykVx8uqZJYHa6y+Upyf0jSxZo5wyRzYiqqiQzxdmyICCCMVcwkxl+ibgotvKekQjqzfaMhBC
rIVUaoysnkhn76cbmhE0I0+QrYD7O0bdy+JGZWCch8KPOKl+CufyI7anLZOP1AOEuTWkPfADbZN/
+MKHjXRALOEBqCHrLjHSCIaPg0JbbKJZbKCJrWKQuUIHLV97JZIpiAZDuxcWmI60LulkTMxRPfqn
FOFKGkZxGkI+UaW310Eew2cfK92CLX5q7psQSOdk/UoxZR2WKAQppO0DY7c/bBipYcaTmvJgp9L5
TNe6I9JHo5VOSPZdOcBPPPP/pMP/CiOqeXqqWN86CNIFFTk9HPuMctJYOvy9kWk39jKkaJtTmVf/
cVefnJprs1ZsSMBAiwHbCkRggAz94jBYdaidEH9O+SHR0SZtBQHgEl9AJxADtFo7bE0gbeJxkDgb
v7VO3MImeL78u5wOxBLFHC0sR19NIrPDX0K9ue5bXDY6wb+z4QxliTd45+RGQekY42PPW8T40bwq
WxjdVnRMEgGFRwl0uYh4KbvTMtccPZV3kaEX2aI05/xCSCm+89xUpzWyz8Lr0WoJd4D3zA3XOwhl
8EJgO648zGBj2QCLuYbRwZ91HimVtLazOzzWPNxD2JqG1xurGBEg5rQvs0RoQ7ngVI2Aa+O1Ng+B
aOKkg6t9ndoixGy82lfMSlvgFxIUZlPbgRpXpP36Sf+CtMqU18K9M06YmD69iqlFl3CNk8JSFxHt
Xwlb3ULcbZn1ADK0Ul70oX+o30PjhqwnFi9O9CirJ80QOYRs3Uze+M//YZ+6+GkWaocXJznUpwMg
Bb8ww4TIMyf9uvSjtH4PdGRwOfu2yWSS1gHMJV1ll9V9sW6ZbiHrzmGsJPwto+VzgvYqNH2GGY4x
Wk524rd+wztNGZFC/OLLXAAzCEQ7xmEB80AbpE2kgikBmZdCia5OeXrXXkOzKif+tb5MqoOfW+vr
RQ5vm/MItLvy2/R680ZY6wwk4PCsOKB+JyxwxwdHhIOVTiUxtD04XrqZvc/HHxabYEqqBbDB1JVj
wP8YJlTUkDUGplfpzvtFbXsc0lEE34CHqwpLFc/rLFT5HeL7jRHZa1B5VuAo8o1560MKXeGHeorh
L6T3TrcsgRhkOA5mCVbwMZrvLzTyHD6e9Wd/LFVdixwWaEZ7uaE3Nb7Bx009fvJIhNSuASdUfA5W
vytFuwni/vDkTh4spfN1W8vB8COmtn8C2L1EEgZcffiPTwpyJxJfrG1rIH5MXmpW63WwnrCj8Sb3
3Lv/zluDbnaC6YynAs8tdwfanxNvlqb4yJmAcvWjSKx9fyGb29M99OnuLKIRFN/jl9KxyIQkz/uM
swkpqP2fO5yfKUgJwVSyWBB2AsAwOc9YIrisZwqEea3vQiODEftC4zCEmqBGEwTfK+QzaIRjW5dA
ObOzEtflq2Oet/kSbC/BoyddXM5KPe4dOvXPC2aleJImDYY9Zo9yANrlpXw8DoTXfWKjTx7MvQDY
TmmVHJ62BUqZDsm1Z3XwTJmpJNVWmv//DOJMJSm9X4TTfgT4gzDRHLIbTOgupemwKx4UPKjVXukN
i/K95OWNtOKsBaUWYryLJsmjzt+bt+YDYeMXpveMwbf8ahj53b2gbmpJs/1ZSTBT4yCHWWWZW1r/
LSPK7fIRdwkKMTkj9YBbyoMehQ64VyG+TwjiEeW4lxFbi34rroSbSP9Utrkb2xy0mR36HU0OuEr0
q4KIqg85Yu5bVSq6CyqYiGZ+qxZxj/MJfGcXdRKQTCoucIfcLJ+EfMYq6BtHCGhLJtuhI4IwgFCW
xGEK0Xe35BB8zy044cl5jZpH+qrm9Xw7JgYHhbPuqdoePlEfpJVnpcNRlHxvBnH+Y32kxj/OLsH0
YGE/fc7xGoeqRz1u2z3pTkBQX1C+p2KDvQ8NRXjdP2alKDAqf03Igk/vEt5grHhCR8nttY9qu3q2
JPlcheIwUObvBMd6KL4eC1tKnrj6Vt7aaF3luMZdRj5ELiB2IDpm8/l3eA7lyM9m4DtVsolnmCbF
C+hXBuL+N+0J/2ZTaF3D7ZE2Qo8TSh/jBPAwFcQOy7BSQY1BuP3LbdvtMv3//mSWTN+7Y7nN0rYB
tt6K/Q3Hkv9kvXn5j+5N8AYQZXLm4vHx7SFDSrOeuN64/dYpsqlfGmsgc0Ssyy6DF/6+SxPJInG1
2X6MEC0GiUt5RECEi90rf+VN85C7bbUZc50HjbXcj1jH+yAoCzgv88f7r4X9TDkfKdDGGZbhLVdY
Cgb+BVsKnc6qRWL9DqMFxP1Kx+pwzpAj+GSQsDa5D9r2m89sgzjQKUYmw/42mlnaJYdIKEti1Nci
oq/csbK0E7voD4pxrYnXnY7c+38izu1Org9/e1qJKKUW9G35NPLaop2NtWrB9lufT5HjqDw9WgUq
B+b4Mbskk/ut70TLdc1nhTaiaB2TrMNUflQheAcufFj4GEnpBn2E7qJXBdG/U75YBeeCdj20l999
1jWJL++x9Ae0EOHA6MC9KGPThtVqv57uiCNTgheMry6zOInJtLoADTmrAUX39x8cNiuklRWG8wtY
VoC+Q7SJSjc8y4Z3Fm7o4lCi0rV9aXREncx6bJh0K3ALsPq6sOFn5EnRo1aOg09UocvZvAPryluA
DRTQU8uBrCKtjDXWbi2/jEGxFWzr0qavLYYknPUG0TolWggImYQct9Q1mStTpQb822hK9niUK8Zh
ya5XSRsZcjeZulHrWEuJEZrz2TWX2hWMR0+DBd6lSpjQqmQ9Gk3zPfUrQP/lOBQYMwb5rv31cNXZ
n0afooSaq7oqoJWnjAfU4BfDdN0UDH2ZnBZTdkyY82ve/PRcqvx6GBnkaRmMRVdC6MXTqvTuYK9v
wJLOF99pewWTll1CLn3QBc/Dlx1Rsi0mljwH499eGBELClNtbbdFNoplkyQMpoLq3C3ifL+AqoiJ
vFcAGJDvpQ60pQY8rHY351ykAM0DHNX8ip6NsDxDg67mNZDbL8PcgqYobY9zQWFfxcs4OHuWGx/V
hTuhPzZhZfnViY37OeeUfuowqIx+j4poZXvviY3CEuK3mFnFmBSnvgzElbIRMT+1nUtSCXSWl0Jl
1YsMhuc+Jxv6Z6dUnM4cOOnRVYjb8cgZ/A6y04c7AfThlNROzB8udOMGgXUYKpuBB7uNgX1hxUTZ
TfsyqbTwJJ4nfHHfGf1Ot2dP0iscvRCUhosvLCeVHOPp66RzDX5q+MkOxqL4k+Nov9yOCjnHolie
X2L2cFh8+bfd3Wgbg8G6IlLVmwt7DcIOb36jr3BlpOb5VehEXmFDroDKohGynf5f96fvgwgK1rwp
MTRsHd3xyxSeqibdB8Ci+e7JXO6bCu2LAeT9SP25BST3fvI4Wd0t7HYmMovW9qj3u+ZTcRedMIMl
u8T/LBnGnI1pWqbhJ909LyKucoB+VutWQX1XDkduUwY8bG9dgdpUDfGdnDxCDc9COf5YpzbD2MRz
1cyasGSg8ezaqDPJuzxl2TtdNscRpn5ltYqxN5OEkCy3vz0x/Vyp01JaHXXGSRtX8fttgJqFAKIT
OglZwNa+6HGJ4r2qt1Awa0JQYZB0MhOpW/6ysd0yFeVuSU7x3ts3AZWUGgOvkYBAUjNeUzIwfp5U
EFPk1fXwAPuu7u1cqp+DoMa2IJlOspsz+9WUfkTsTK5cGi0EKmOQTmgWtHEHFiD8ImHeboKfr8hD
1f8Ld4BJRL+snLUJhY37GobkI8Npar9JC0r0m8O0qtTDSOO/zJcRvP9tAaA675KINSN0XNA5SOLh
mloXTipKmXl/VJdyDm1H490f1tksQfdByjWr6Y+9HM7M9cY9ligPNaG6VZzjTXYw7h0uiZdFMyIY
WVBQSQU14r7wNe1YepGU+KjDoz130ZWxdxRvBW0uOWB60qP9dyeHurJN2KLND2l59qTq4FCauxXe
/z/BjCCKOc61HlZL/qHLizsUA7/0tJRvjtq9pEF1kkiajrCihrLNAkaOmRPU5SisG8B9Fcl3eyy6
DZMeRbTkkURoVhn8vAu64srtJ1Til8KItwUEgsbKeNrPfEPSoO1P6lAoy3pzqz1wk/TYcsbCz/LY
oQcb8doScqmeLHylmnD3YreR4fwyoi4n/FkyiV+XPjG6BP8pJkGBQA6RyjqDjDpHiRmROtL/fVxM
x0V3qLVxQCuXUVuacobj/S+u6QrVWa1Yx7EeIC8lZCsmOn9L+lmJlrvalzbqwWWZ+zVBn62BXBX4
poioYfAfmt1hs0JwzCSvgJTVILrgbyJcr0tfHF+8Ix4E9ze2oSvq/ZLCn7OOZzj/iGP44XjMMS0R
hsRgW/eP9pkOqZ6ydj1PNwPZoe3k+VkedQb7AzRoyPHysBEnQmoNIOdRff758j7lKxgsVtMwRa1m
4QulohGXXSk6dxSg89w745BQiSITEnDYBwz+uOm+zxGqh4q4IAxOBefqq9/bpiQVsIWPSX37dTyn
k3neItWENYaMTxo0vVAjqetu847whuV1q86mWVhdPgne+ozME6CVnQwjKjCpvm+CnMaIUoB5cY+k
H69M4G7Hqdud2RKX9NaxU/R9Ird27UslvLtZd2yGB6H/leKyKnCuKUyKF5+DcNH6Sdc0cXzbAIRz
ETeKVHEsO2/tnVHVjab7P8lKVt1XWu5siXiv2zwoT7fa8KzqeTwimWGoRbfRT7pZWQOmP9TM8FgU
34JgkTIkmuSz+u9rqEhyuJeBI5SplxS1q1YEpJb1rRTCNDJH6j93jF7niGLQkKt5cxQVEf1rebv5
HOfeQHyCDPFCk5KKykhnVk8T2LUJ/dp0dWQmpKGsZEFp420TL1ohIOQckTv3KCTSjhXw8IMSfbOp
L3rRw9bnl5fpnM5/9EirInemJgsZZ7Qie/Yij+SQkC1mi0Npa5p0nYg40/+bPFYy1AJTurfXVCcf
UEPYhk/NjePl/9Qe7PsV4HuFltlkEhSOFNhLUUbS20yXQgXH7kj6zRdpxrxVCOPt1+C66TjY6nX3
c7OxXIf7mpOGxKQV1fOdNjmwHWFjbitkDhbtr1W4tMVOMeAF3EELrceZ0L0i5RwMecwy4EVx3J1V
9cw1bput7OMlXGWYqjFfPgOnox+OLBNeoON0ocPZd+b7CUTCgjyaxx4jrtBN20R+v2HZUa+lqF3H
EQLdNo1pTq/IvP4MLXbbsXfVZNLBpdzEK/aMtfFOkXYj8epSFc2NjAudkyx4Fo2cdDJ/6CCFCCix
CWgZhM9O4U36VS8K2VdOtszRloKXGH3G2O6sHIBJWsPnWWImqP/rAHfByagbzyIXqj2lngc6xGPG
JOa4Ox5nf8szcqAjxWjz7Yuw7CKN+pbcXA5XOtk3FCqOwOyRxr49MF58nSZUdPIJed4JswsBmpHw
yxEPXW4KCEa4054ChfWZBoKbctxpZWn53FtHM7Huxc02aI/Hs+yP1D9qXxG5YZ4/4kdVbh76E69x
Ufg6EJ4E9kvdBd4pnCRvl0kShZFECW6vjTgAQxn+WbsklOQh3b/33nGzjzR3RvxgbzgQvyqDv0I+
k0Zgx8oO9vPRfQeK0o00UQHaa5R85OLN+lbbT1HHkko3jIPxP6EHMJhUGrDjp5Bg1KTn3wj/7Q5B
TL2H5VihLSNtuDYi4K7y+SAFUYdbFPL0J2HZwxp1b5OsG5Uz99cKh4U8QXP+aGKEHXnjc6I0og9E
SqVCrZ6e10xA3oDYqcZg+cchIZ4T5Jcs0JYenAOeLbFajpiEH5BQW18nGHAu8VDXr5yoxQuA0fgE
/O9RgsIx3HR9kMhnsKoXL8ABQ862WMb7Zg2kAcTlIzTOsV+ccfPDjZHDGSecnHYkLmb39xmnU0UF
s03P2pb1yua2vms7eEs5u2m4jDHKKgVDVCD8f+O6cHe+o3excuCeaqbd4SNDONiY5FVMrL4izJ36
xe5Iob8Pfq/o2zFTzow+SzIXUooEo3QuMf7sK1hNsdPERKVzI1sfogPw4VljCD8ry9fu5C358Fs6
ElLqoBEZtFY0MnfBTaLd3k/985SVekG8ocPHJgafE7JS0aOHk4UpGZqPQddHLyml+lMiRRDTMzm8
m1UH+8/JXBbWMqZnQCJ0ul0bdi7ztgWH5PgTXEfBLCIBCPtK/WQ9FhkCRkIIssxEVSV2ieK6c7FU
1B76CHr0g7sh4vWfGWX3ECE+soSgmXerVAZcjOGZDVe0DPzuqtLsDgpB4rlcoZghquZeqmHpfA1b
yFxlHngSLJgdIc58O/UtRdxiTA7D3IrX/3os95TVmdBPU+2ymPNhQJtm3NECZ2Mn9Q2k3dIdOlN6
CWsYUDiE67/eHElYUn7QnmWewavhtumGPSMeMWMcEHSWfYOY2fHaORuKmgkJXo/Ky1cwNBUTw4RB
wxCXrf3/y9vrti3kw+AX4PdG+eChli3BmHHn3Fmwtvd9V4+iCvOOxg0qA/mncz/b/BNt5WphtufM
y3qmtqJ8huMA2yfTfmjAKiFJLK4ES2h3yYGUkMmQJLw+9OgokOMTddA/HlVcaCDZ2nScHwGtGQwZ
y5oRYTpEBH0Q+0x2kjLdfJmb7bYDlG7AI6fv58x5FyPe9NQKe5CahYOCmXzIQ466SPh3YCv1gEfw
EjoAraSFkJe6Pr6GRHJdQP5EXdSmVmNC6jx2WVfszjxnEFyEqK1P00Y1DL1b5D1A52EBj0pKE8W+
or1Xak1BLGuSRXApjEi34yfRxx8jrfn5Yh2Z5iz2/p/ddatwV9tdvstCfcvJgLYBaKCtNOY9cswJ
+YzJMw0nFVlvYhk8lKCIGf64AwU149xoGpckcOmbxuMZGLavg650vWmEW8SvF/kHl271bKOCm24+
Lb6a1brn5qHalAKHnCZJ/pINvnrA4Y3wRwTWzOmfZZf/Xg0nzhnZGrS7gIIliXUOsP3ozVJSlIjh
EgTWe6X0jtnJqH6uzJxZhAwu77lbeDkBYP2Fnowko0QO401U/Y6JT0c8uUbVPVviSiPAiEGhZzR1
NnyKMguTfZ0rDatFJ1LFXZkA7vbT2f3SDX6OZ70sm2lFNznqQQAR7Q3uetpsBL+HdYzFhAJbJDHh
YLLaUhVusEmhrPa5Y90lPhlPZyNDnvwD9HuprwCfHLQW+oMC2IsheP4u5liLgrZz26Phzg8JJZNz
VU2NGruS5XNFg0sZdQmTnzUdAhGroAqk2J8XVThF9b5lUp/Na0li0UstHQyAuYOVoli4fUh4ikmw
c8zTC6vHCN8sL0QcmpUZba6PAhiaFry6VbIPklwplcTb+IDkBuUtFGpF9vkVl2MBeu2w5OB/GYZE
FB6NLNDuFTf4WsUhdVATN9thyGiHPHXqesaFzU2dPGXjbrDLfSYDhEEw9XzlpTBYsx5RoXijHn5P
mgn+Tyx7ep+/Li6d+7DRjh2PncMvfi1EkiyZdKTRetfV0YE1TjLtjRWUP41ZhOLg9oCavQWYftpc
g9tgSoxKqjOicCU8N5l8+EAGzNHUr0RCn0oJFn+r7vNpyhCbtAA11wUZtEC65TJY8GNWCnkN+/kI
kyWyw5tAEuuEpGxFQn1OlQnuHddS1iPRz87rrBy0fJiDZM/F0vfo7Og50Nl4vgREC5P0ul1qozJe
5Y1qqSa5Xau9NKB+odIpZ7+0HzQ9cl/lAngrUk9jSOriwrVBkVCmRNRI07yz2Z6b1ZMTtPxTxWXo
vQNDS0XVjX4M2FVo+U128b2738xxgyK1QSarAlGsKi1fjtTYDGXkLqyZKlwSu93OhbzjAbFCtL+R
4pqqJLbZc+3JlagwW/XenAHaiWk9LI5qi11Q/BLs1GZL68+xHSAt9mcNoAYSTtEkoYWsQ+EP7PnN
M5PLJvfxE8MZ0AXW/vpOecGjPsbUL6cxWzaLsRETV3xC88lLh64gXKzgBMRykBBBEGbemNKfiDZZ
9oOm4trjgqRFlwCkgyMZwhxht15lRfg3F1XZh2qneAUAUO01cnZJQOfAbSubV7pJODoeFhr3Pg1a
y5QZPJbkdnOcQ35g+pftZQKA2kXhf5B4mcfjiXM/wwFmTqLHWmyAdPwZAuk27tpkmzDhcJDbfGwO
cqAynNV55q03ma4LgkGMugNsSmdWUmBesP+sY6/dwXnFusHe1FZy6Oj0K+bq0XmbVqHuJLpYDEBl
UPD219uoAmtIFjuxIWekMt24Aui/kgWd6DRLT/Rjv5IQg59lm2nUWOFShywtpO+//z6nq7L+QPe5
Z7g5Mp5B6CFdKlbcqEd9bT/3u8dPjBQW6rJCjOnzCqzBA+ILHF/Nap/Jz421IDW5xpfRKvIjXz9a
TYcs72/CCNombJ3Jz0lDhSFttBCoPTSagrSmwI6k60Ivy7gI50No6kAlD7+y02S4fnODo3bxd432
aCImuzsLxcOnSWmi1fSv/OG4lHDVojHgNE9YhqlNiKN1h9Czi8LsHYeyftZHDdxmLTnIzxXWR9ba
99XJoHxYzzeIuKX37vI58sldtvFbngyOGWkpuYMf8hMVQ7wCXK/Eu7yiDWhm115u5X3fuXdwJeSZ
aoBH48U97VmTANRe5lzyrhdZBIfV/pS5D/bk9YuCVA/XuI6LtmSvi+f9VK2LLyg0J+iEha1GzAwt
ub60wIX/xflGva2HBAxMGsLGBFVa5n6XhxkiRd2oUf2CCmJBZ0c7u7SJui0vvJeqsQNXmtL4xtrb
bso2V6rjFpjxbiFlVz8MfnEKbtXZrTZ8ZE9fmuVxNNwPRswwcH6y5Y+fnWGx0B01AdIKqKmLcghZ
dcluDSMu5E/RUeW/Ak0BlxrmAPaFibvhSreszWYfqRoomVCKdne5+XxAQSL5tCrxV2ovODLhUkNH
/FAsNUOJv07Y5xTGFBMJ2cmUvb8iZ3YLqk6k4iMBs6B+EnL5ubUlx+T7Fop97bDm5H0/A0/Of/Yz
T6QzbnfEIwUW1wLEkk3x7Cf768AGve2U2tgb5WejmYR7YfGvsiOHmDGmmuzNxx1ZJcpmXompWCoj
2lvGmzLU7/Lp3XYvvIyLXtn/2abPI7nB1X1SXkkbpEGuPSjPuwY8XH6lzsFQuCp508dyy3i2lbKk
W/kVpQEEg5AexuAduXJ3Mjq3z0LqqAugMCFt7rpWZ58PXC/1nA9cu7bElFKI52M0bJKEM7cqFrwc
+fXjwMF8MeqwgoT38hjs7CqI2dtHRnaqLof2vgEZlbvGHPZgQ1q5nVyTN28Rc8UDYdwamBq34BDp
/2yBeKXhlv2GYQ+EgqWm5efzu2mT6SuFxUVj/fD77NmhGEyGPDrZ8AitRXz2/di2NRs96YY/fdWX
1ZW2Bdn9xmtnrEJ7xeDo5o1OGmsKaomeSgUPDobpIJkEu3KEsMULeGdPsey28+kSyTV6lLuT2KaE
OC/RpwlI1F2M1id2mdkSdjhLcjlvnYzjJod5IjIluqqogx2dbd5ALxXmfTUMpMCpuFp+dQlrhzhS
1r+BKCik0b4YqmSgQBlhEDfQibbRt+jQ3y2QcwT6o+oT3lxKstGZcsBrXOuUky5zNcgZZr7Hjnbk
tJPrM3kQwS5DJn/NIm4VvGbN6YVeJb939suRc7vaHTUdUvrNuA7IF5wjnI2TaNVuUUCtyO9kag+T
d57h74gVWR9LAxKlpdAm5FE5LB7bqpCLp6YuLh1Adk6h6Pt+0GbzIvHtukc+ntfBOpKUjdDoeUVY
fH4qVd9DfP8AuQky1+g2+fEHsBYp3Hs5D5rHCMl2EQdUgkXMAnplxz2nl1jjztgOXjMjUjbD9Vzv
IpUqSJG/HpWPwvPJEzLwQ0k5nJt967P8rXUURFkriLbssYn1DXUqMHmpBqj9VuFbLShWI59DpEw5
sfpbM6nEPPxSGNVymexOJsg6EauhewhXzYr3A/XzbxhIGY/qUNzTzgnigcnVK3vVoZ4nMX07RqHN
VF2wRWmUyvWPG7Dzm/6n83OUzf6LJeSNP9aMAj3CbAvAZXz6fgNWzehLtbX1RNY99WXTzGTrOEMX
2t1j3ttLRB/8C7xzOohigF+2XCli1yqvH4MTQrt1xWrhMAR4QQiqJZi+f9Ri74IMZS3qNsLs4APs
H8oKY4lqEPjMH4ZS/kZiUnaEiG/UAozDFXjwyjN/aJ/hX/5vR/GwrYvFiIHPi6YhpxSOp2oHeP11
RAtP8YKTSZqG2hz6rqtBC2WMdcBYQrzYLzQq6O0MrAnQ7NdEF9orM5U07RTwnH17VazzaoCIo8gk
FUySXL2oDNpQ8HctPbu3Anql4u0ZwLMcPSgREOzSxgbRBHKhveUhwfYmwFz3iVuzzZuC0dUc4ck2
8sO2ROrea+GyQD2tEbxNo0c9Vw+0SPZ1z98LBU9NEp5jyZD33pJ60pqdsQys3rrYHBi3LxBDjX7K
lNIWK+jMPRWyl+SKODVq6TRwUBGtHwnCklqkF+c3fAAZE0+BEfUPGsRzrTLtsVr8260HQv60Mp14
ukMsAdahvY3swDu649GpA5KO3tTltrydcor3ITlqxaffwX8UXVtoaZ3FhiYrjV/yPsaY3rU+A+Q7
Nu5+aW09n/NicDFn7xEXMwa2f9NbupZl3fRYAa+sAD/21krPPKfjfc+QM06MShktXi1HyeUBIkUN
i7rrnHYVC6gIZ+WV7DU9v6PlfU17FIjsgWqX0JP8KftaqJnUfj6xtpRuci0LaAAdPJY+0C+hy74X
3rdYtHo9QKrT0r98+7+Z6RPQ4P3jcielbYEiIxzyEWKTCVSDyIeDe/6G0+FIhd77IHngi92qP5Yr
WTp5vRQ5NfXmx6WuG1mkF+iGJqsK0hcwq1Ykd/e4QdpO17OuOKqit7IxegX3WdCLlqZ2tC07WejN
XQd7g11fRp+grWY9NyilNwY/ot/verTy/DM1u4HgKL2uHS1RuDbBS5fgAfAll2DHuhP65mMmF/8+
yRTZCcaFx+kaP9o0lgC171DYrAAtqsP8LqHSKyLmjErRSiShlr6uRO/mI1XGVZ2TofYfipG6MMgb
EXb5sdfeyQu2YQwuBAeCV5W6zW91WrA/rxpg1/FioKXFX9zoXohFkt72VXAHnrG0d8vPnccyI7Kp
rIMuXU6MYpNy1CB05yQ3ldhgJBC5RRY/FUENGSBqkZDA+/WA3ctPwFoQiq9bGHDzxN4WPpJTvYRR
iXpUIapTu+KbItWtEvEviYxoQbU/W7WxHV0G589nbcvxXmyaQavcEGujp76spUXE8j2t0/9NW6wY
W3iKH3ow297kEQa6EdWxFej0Nr8zj+/nol2jvkCQ1p3xul4Oj2BOssEqpwB0iSzH4ca5vDNLQyqF
iDIySetRZQwX+DpgB7cbfRvS5WxfjSHTJIPFNxLgiDsw9dtGP4uinWHj51ppvZl3TG7M6BDSUK9e
oAsnVrTpboUckkqv+7s5OBZQO4STKDqzeLejAsjy/stlAYGu6aQh4RRkpMgvEva3vH5BGfF0lBw5
+MXnp3L1BfxYm+sdXwiXmdYtWmhNye483MF6e1R1SS1nwuf2BsTC+G2H8HRolWNpzqHhKEYGasGA
P/A1WM/F0jdr6d5kK2YGg/wfajazD5RM2d6vHikRBtyBLQ85e1LvuBf8JFwTtyQTJYoD1qhG8ql6
H1AgNjoobrmuzpVbg9wq+JUnjnR1porIEbkr4TxrEexeLADpgLhTZIgmI6y8FTsFrY7QdIyvlvrL
q4JCS0PeYHSHqTfPJp00oHXg0/7bt1+o7NKlXd9wNoVUfXLhXYdEFZVwHxSp10ZiTF2w0Pwd+/6t
IdWYBHqPdZlEqhjUOxmQZICotlMrTWvAv+orEdbuyKVutjry/go0CFXUT0a83sSb1nInFsduZGDF
1SM1Bo0jv7psWnBEeViyMqhGM/Rvv9PXQhMwNEj510sdQindrSrfe9ACLw9uvIlaC7xby2HJA8VL
yKIu+qWJUEe/ih2/+V/+EL06/Q743dSAGpjijTvL32WawLZrFFSw4nxfX/ytD+uevAXzdp9ai9rM
JNQGRX10gy/OLGDQOfLQQTE2eWRSkCEd8m/9grnNbzvmL6jStbNj/XBYRa3TOul5I0Py/qA0eEM3
tvN0D8RtE0VZtWMjNagWf2BNEcCluXon5FX7E1fz2pkwtH91QUcDZGB0tB629U8aOni5Ib370U97
JMqlUQ5ogO6GT7MkRPVnbD0k4SWOunVrcVVKCKRNeWWu4Dj8MGVlbNzUoueUH97vO6ENbpA7Wym1
5fIvbipkqh4JrO4ioQ+BQ3Zjz+EjXV5I3b6GvHb/lPumi8aQWNs4dHthYUVdh1xpYVavq2/7FyS4
v+TKi+1/soD/QJs40wUY01RALC2I5gNUVCUAvmFd8LMjwoWXvJ6oTs43nmVwSbVQH2Ng2534WAJJ
NLxCCjegtXMaTJjkIWQUjgxNRXpqIRJtmTS71dpF+ylZqaiD2Q7UKDiHyP1iu/0DOLHTDLyQuxue
5JDznf7olBMxAkqcPwYYB1S/JGoMpmaQScKRZG4gxPN992gXqNt8s1/mLQymsPjfUV06i2rGc/TB
NM61hz7m+R+mzU/bjhmHbwnAXFUUFsQQKOOrhG+CU6sP6icKZ+v5g+ZvgS9zSy8u7v9iFlTdKotf
YO3x8upMPizGseSx2oxGqFSxLxwOBYBoUqm3OxXKhaUMw1BC1N/SISWymKiGu/Dm+bKzK8JTnNg3
CQpl2xQ4JZV19TrLudbWKRcRlJ2IRK4L+uIX1hraFwo7mIvEwMhLk8Z7ejuoEl565O37za/rwZ9T
7rEpIux0FJl1GZ1e+9fLUDxHLUa9wpDOKkPWyCBJa62TYhANLCzy75R7rTcJ0roPXV5/eUAjq6f5
5my0EBV929/zFwBn2P9VFj3h8KdvbeS87Qo/m+YsNQQEs4XSZtHDr28tUXiJ0UiumkEGgY/kwtTC
UEREKuhqDqa4J5Vf6JCtY6WQz6k1+ODENMzfbdqSj3SpDTdNfe+oNg78xS2OvcE+S0rtucY8iWNi
Unu/GMSGBWUHArw8Xki+ANnu8a91DHrO1OjQWoAAxOnh0MvTJFnAnwyC0PSeSIkH4Z7F7Po8Gd3I
pPOAfv/1CKrhgWwQ0OPm+T+awzqvhbCEccOdBOKdW1e0gg3lMpt/Db3SbUDgv7zihnw+v5nM+evk
OsN8U/F8DTTS3ltxaEJdgP28p5ymT/6i/zERes4rr1ow7/+QtpQSbFnYH6wamnuu6lxpy82/a7Ej
eztXUPWup+8aBlVN1pRfB+k9HbmHAAt0UcO5Uf8vYhCkA6xMIAtHRuobIUyNJLM8uwVjkaGGfc5P
luNkJTwR2VtNYKtwZUu8UQ96asTMbxvucsYoMX9iDF3bTEU63nevSDwz1CrW1njhqEbzQzncTgzY
RJBZs3+oNZELf4tAuudN2zTYNzBbrvMzLHQ7PXj4U8Cm6vgYLf8SWd3kt0bXto5p4zdURrxUZvfZ
7mW4KK7sD3zNuAsrFuuwKlOfgcpaqYL6PRzgPt00V1Pc5KEbinKdWWWOxEtszMacdTHiAgp9KApH
K9eWVedxNFUeDFPCz0wt6iBeP5Hn1V6ex30mHZXxetN7OKnar6vm8ftYEKX8mOibz/6QpibqB+kW
W2cZtpc/+OV/hubuS13gK496Pki+2yd7Axo8+gE1iNdGWzJ8xkJCH1Iy7VhgCpG0o/LsU0hM0EQY
QbHCj6tjMnbnxigVF3nxhl1rH5MhWjIhLarUSP7XPpShy30CTgOHUBF1ELXobz2XvpatDaZHs21z
R3WGE0Hk30P8sNY68pHpQdCOj6ox5w7IYLAFOD0kjoVxKKGeE8LSHQAzHWz8LPtv8h5jAtQfRQRA
byYzR9ItzAhY+NlSDdH7VGzplhOfCVcvmZYaXmlVpomCnmN8aq0nG/4WU7oQ8gIfHE1bqdoGzqZ6
Nn6iKjZOEaNzQxonD0fxx1vCOclScgwmVFaWty+jNm2JbeTHtDFKZ+rWhQOJ174vj5sqYIYyPhbI
kWvm8KUSAlq5Z07E4TCIcLD86I4kVgUS6RUZGecS4yyZSNwyBbE83jR455c8a7rK7dJ40eyS5ljF
xpxbEqlDtosHQY2Q4R3fd3NO1SJjrBPJm1VcunjBdgx46pjig+d9bkCtH+qQ1l+KaN1iKANJZ1hV
RPm3l7zwDt/38eRsv2M7YK47ZL448UHVax9GCrZYzMLIhkBTzg59wdsSuS7CTWFE1WOmF+etQhaV
XMt8EKlL7cJpu6jkmLUo/C95hR3PqVdFX5EOZ63oVUrjVJo3P+6rSYANsIgL+qE3JGFNU2/bupn2
/Ct5p4IkP+PI4khLeapON8bM5xAwVJydcz75nNZ3nH/J4RzJ8D4T0uABCOB0dEibOOY/o0NNP2Ea
tpIrkHlhuOxk7Ww9h9rNl8R6oPdSRna8hc13L4n667ZhLmLVa8NIjdED2friXAz2FX6fDG/NZmV/
xWSFDDF0L8ntFFY2jRHYD5+p6S5pgUUG8fXvQ+rmHfoke8ZnZQjHlJch7HtgSiQstFN0ChtbPE83
JLPE1c3IE37pdHD6oaHvvzbaH+8NOz6kXQQeS7k8XtoK997bkiSfzEqeS/WbsvSwATeII9919Vi7
NQTPYo3PtyKzf82bOljTUd+tSyZjJ1BnCzai6ImGkkCEDnM9EsN4x/zCPutYdiIbyZ1qIynA0hC8
e0ZGR6m2tR5uGXcoG/AozCA+dsjnXxU2bFxmn/KkCwDqA1MiEjEw0DfNGVDVDPdO/Ra/0o7ZztKT
gd+jSpOUkpt9ucJaW2Geyl0QY9Z5SC9PIcI0sRfrOTGjOQiEhCQE6YybGOiPUb3eCUI17O7ZXtPA
2LuO5f0xRKMOBy8l+HZo55tWsJG0nv7DJcgsyPm6xIY4ySJQKQgM2f1TtgDIhcLkyLo3apDxwFJ8
1B/RjClG633nCXy/A2pwlCqba7vSgM7erqKnXjGed5UpoTJ6f6xfEIrqdozindYckvnNXzAVawik
Ip1WTiEqc0LCxIzJbh/NOi6D+yRuSSs3hPL2VAkW01pMGo7lybHqdnmCXJah/290M8RSsbnNi4C+
USx/lNv5/T3WO8xhHr592HKjsDBD4ORn2z87oWrZEViMXYcA9d9scmIomGQcgNqljrCCMelQRtY7
bUpWVLrR3Z2xAvLtx2WrplIp3Ow9f77Px+mlQZYtDikAkFZQHPgDOoDTaUIn9O0mI6luLQ8/4tPk
GUKzj8tvUv7DkC/vfzDbTqiOwJBqLo1PGVn+8ook2iqQzb9d9B/95OHivAD41MJZZiTMNX76AxGx
cb4mXO1tASvOuMO/F9UYXPC7L+3q9SDF+PmtFxmwS/BBGsF1lPExIWYFp7qHwSnLbw02UzunM+5s
QMvRAjCQ6i3htNxajVhB3BnXu5VmwAEm3cn6QuUdTP5PiXFsiiLKP9jTSRB0L0xksd7c6btO5yxv
EuUNJs+XKFW1dfxpghjk2+DBVku4fmWS2FOYz/jD4IXMyRx9lzot0D+lpIqN3AjotA5JY5YmdreI
P0iKoQNnkFiqXTjPfKJApNZqvpelhKmB+7roQFxPCgApsULLdPcecg7J5I58zQEpihUKXWFzjtuq
jgjUnZULEE1nAA1ixLDtUo0zkeSLImgZ1yFtKteV0xudwLo4lDgqgi3x81f7qLZ1JyeIcJK0Di4A
JF3JEOMpdqh2B1jXiJf9uMrzEOL8Xh8fXCY7IsgvKD/54MAS0IIFAp1yKieJ+hBkCqsWhZnwVZfB
5Z2t01VLrISVkq6iKtEGSe6goVlQVvI2nc5SXxPmv3YZVfTaLRNEBABZ5qZp6eeGDYVZ4eupm66i
5lFeCCZLjQClmuMMnYyoYCCDCgO2G1eMwjmWyi9LW5v4EOCQUOY/iaolyVZY1U4SqHljY8JQb2ZR
6f9Ku9DJ0eWhULBZBvmPHJXpKqG2FhgTBlUZ6aMciFGan1OF3i0/pJj8oOr8npeiVlsXmVA8QblQ
/Zcikf4RFd5L+3ZBZWixSQ3gx8+78WTcVmA8ENYLs19O2l11qAXbMHC0u21+tLVgCiyWNY614H6S
NEsh/D6KQSXsS8tM5x4gKjTZ4EvWsmrh+loqNv6UXbj5fsKDvhalU0QCsKP2/QEnCANyp1I/TK3y
syZW5VEOSwacv3O2SWtxIfMK4O/5h702efM1Y6JU9tJe3lPt/RXLtsrjyZKgmrcPNv6UUYk22Ggn
cDsSF8MKt6NVHmnLtcuHHV8kxmHyMqOmWQHa3JMAiRMMUVpaMST5bPuhaNwONefcSu5VTHdqXalO
fcEnwWxyDogtH1QpuekoPr8/by63iOnxnrRtVhdyIPsatzsUFuyhtLY08EyWl4QBg+sFZbmYOQq3
ixYwNnuLIDaN0f1tqQVYDflj8tvkSNsD/dB6yyTYDNSWWIZerUYGj3o9FJ+hIFCLcRMEspT82Y/T
pgwLNY3tzQRfpDNvyEwR9vlM0E99xT+Z7KzIvDM1MIzCjpW2Dr7g0A9PyQazsS0iq0PWfEKkaa8K
yJAEUH1jT7F4bhrwrIWxhaeivvVBxwK95giYKvRhzBlw95l8KXxGUEklfc3i3w49RJYq3k33HFed
oT9aSEzoaMK21iPDlq2DIA8pPeOTfi6zdmBK3DfW/6xjdWz3VoZokaROBEapt15P0KFxpxVXMhUd
OylQRyusdt8MZno62ckNW4QymtqcvtVP3MA2T9V7P4CcxiW/SaF2ubpeEgzHhwnoYy/wn42gGgaF
Z8NwZsF81KzIsQ9ETBbIAMyetm0zOFpBH1jhWG4O+xx73OExEIuMiBEtnuxnMP4Ni/cGIzo9dPl/
cUj8LkQRF0c2vXiJVwaxFqnIhE9kZpkfv3lnb3caN5BDR4r7dsEsJWy/aqET5m9i7iRzX8NsiRQE
g8lSc1ORCO0yGEDJ9QLRy946POIJJ47+3fwlKGTkgdwGfJnLvt7GY8bDq/KkDWH7HErFgxA0M/D6
5A4tW2nZ1HJG71f8EbtcTAbxOhf2YrfZXsdiZ91tfEFBCXdUt3LYtku0FTYAQKfhJY7GwF8fAVGI
Z0nuwiIrivqfv77Yz7tk2VWm+uGOM1/0n3fZF0MvLyV8CVSHoiFV0QZyyT9VUrlypT3Sd7jmnQkd
HSRBbVfAhnlkylidy/soebImYDYgS5k0LG444pvRk987VuZB3Fxgpy5PepenT06wExZFr/AxfV4Y
ejhQnbuod2601c6HjB+Cja5sekmDaJsht7fwFRQSfr+1ujRFMysN/T6iRQvjKawakiGlACFhCW3c
ltgdtpv01pv6nM+4mAJyl8CayTqvHGCe6yoexGCw2PI52hUob4+MpHzj+tF90PPKC+azfeRN7VUp
8eNJEMVjnr/hh70Jm1EHOLKq+daaJFXE76DrCujv/PEOFbwAWXxCaRfWcpx9je+pb0FfWAFdIOc+
JEJKLyfuxQfp3cCckAsHhN+jqugNPvsbqp9Z5UIilo4sxJ2eI870alVHUkP6rcOF97Xameh8apsB
QfIQ1OMgvuFJzaTzETpwWzgPxhEP14eSHf8Yo6pZqxW+CDQpuwCtv4J6Rx8Hvcjc6M+45x+qsTIs
0ert9836xxADxJPvYduLSHy1T8G49ed3imsvOqAhjAzK9ff7712ie4LYidLhmwX/BJ+wIP2m2t1k
VeWRksaGbfM4E1G5MKmlz80ULUBJIQtUuSwhd9iVo5ZbHUT+MVWG+Xlmf8bBMp5whIf/xhC7mAOS
aXEs2BaAqcJj4H7p2JkMLW0cTO0dt5HhOvyfh66Z7m/BsO0GH2GIccIRKw76vEE2NhoUdF8laM2X
0zGe3af/yQ/eEK1+Ar02ORNOl7fzNXlbWW2WsOW8t9lMXyYUMj6wlJmebO9ztQeisLEgGhJU4aZ5
hVn5/Fo9zQRqIIWxYVO2VEVPR3EeqY6EYYBnM+9fYs2FlwEafAjijUF+Jtm7cC4TN+vncbIIGwi7
vrM0jhGnGl4Vqy68AuLlzX+PMKdTLbBCKVCwUeoT/DHXpt88at+4hQA7XwyoR5kkd3s80VMOTmtS
tBZYGcadzp27FY/Vf9ERyEsiWNIiIobmSE4nJ7pWaGcoAFjV+noOVNkqRPgMhrzotiZJqeiBSYZX
D8eLLqAKoXwKIc9bUR9CKEyWB1oBJ6V5E5CZOMhC8ecsAxZODYob9IiU3Ke/PD4iSVvw6w2kROOj
/4chB0GjTmDD/gFLHONwQYEy65lGz69UK30U0JYYE6/o/etTMH0r+7IAleJEIT57nxVtZVQhixba
lMXjof8SfzRUlo69m6d8HBST7BVfBs4WvU7ZK5VQ3Q8VQKZVHdfdCyi4Bv3Ic7Y4PXCnqsvH3kiz
76Jvh3FH57vmFJRFnF+brnphDHEaYbKSIZkd4+d5qwTc6VpGRIHpLIR9rbRY5OPGkuKoldnOQYFV
QIuyO6uU79a9WN7QNnJigMveeiN24ixMaL+I8AxKW1hzbeRrzOrtR7A5HNWXdmEm2aiXJoLN4tqz
n6nOCnNf5RsDp4n4bvQjxjswUy3N/pohb71oN7BErtqczLUhsdgAxS/Sf9Kb2qTkwMcRMM4ri3t4
eDxc2h7TTY5h3wIRUe1lOrWLAL9S65Em/C0VEGKelS3hBH7OVLY+hVZM3kMA/VOQUGByH0awhlnw
G2ChnYHKB6mhMItO4EcQiwKppkCgVpg8vYjD1eHDwc4FNJDBioWKjcKR/FR/4jwhHxwJ7+uZIyzO
8YTA0sfKDvkm7NlDK4LcN4EVDwNBNKvT4ajGCVxVZL0qgz2BhwcSb/PIFMcxC0Ri1YdQRoqNItRq
sC080Rg6K1+lttfuXFlCgxMRj0+4L6eTzWJm0esZ7jG6Dybk0yO4K8AMlo0nQ0nXNDQlW9oIGKbn
v1QJhz3cjqqX2AUXgjjp/Q+icrjPmK+g4InxIGf7Qt6o2qjoB3dfYneMZ3UKeidCWQOvw7fRgee6
4ZAipc9A9QX0SkcM54g8mmv9WbbCxPtC3Mg0N8aNLgrqMRczKSzXgoZ3QWwbQ/CNKV9Bs+TDfQMk
l46XmCib6A3tq8gY1irrvBISnMcxtLODuetsU0Cw3DlDrVkqhC8bZx1d+RtTC34Jkh99kLP+sG6f
gybNT5p5KVcdbuIrbTHTQ7LcywUAmtwok0DPCGwe2r6/2ItriTIgsDAwkvN3KRNyMvjz15ZT16AQ
7Ny0OGsE0B9+tMiQ84D6WiP8sESbkVEwsnZSj6tlRW3Mi5k5UBlxnEohxBh4Vtcn60DW4A4aYinp
4zySf2aHrN/dAhuRyxSoq94vSE00c7yu5HmsmDINEQT2NHQWroMN14Myv0sidUmU3YujVM7GCHrN
/qX5u/NH1FNpCmSXtzManGOQZwoXJX11bgZMRiRH0RZ4+HDQuZqC2x8f43Ul0P7BA5AD8SdJAquW
x7kEaKHg2WhDyIgkqOrJu2v+g9EHWGmHo1NhKrkrNim+XiTMVeh3/Fyw4FU3Pm9RMtCRRbAXh89s
1KkvCguRmfwkSQVv8PfwtLJ6V/feSlIC6zHvaRzhIUV6Sj2dZrT2m43QVLg03z/oTnrhHO6O8h9C
OIo5UTY5CoEIN4UzXfBQVFJHkpFHRTppO23ygOB/dLgT2aOoTZDEwR8BXiWrVRnOBAChPcY9Ipj4
sY4XQxcp/yMVUCgvzTEUi4tHltoW/jzztn69gJ7sh+k5q/tcMkxHybUZhf7dHfZoM3in3UDuYhu5
TG0JtA3y6fUCl8tsIggtKJR+eiLZ5KaCbBHQhxkRpml8JvpOVc4D5d3f1QPLakLZB+IYo4RVVVHH
FKRLKtqP1GTelIbcfN18ljb5fdBCYj4UHXqGBtA/XG07VLTxwcSCkunehNdoSD6q7FL353MfzrbY
QLvH80YJxmI0f7i73JySBkYbf2E+mTU/f2If84Y8zvh6kvTbbv1jL1sL/0zutIoFlakzcxSadZmr
niw0dMiuJyvVzSKDznv7kFloHg3XdxXYtdXVDMwbqWGm91AayW6oilPuV2ZR9VEI/GgvTXhW9W7L
li1e8qjEAGB49xmHJhQ6weN9Euqul4D4I6B23cmZY/i2ByjCKNZNlbBOV5S51qKnG9AKl7niSDAq
Fh0C1WzSO9mFNuBt8JkHh+fsn+I02CHO5socZvbduaLdYj3bT0gWq8CXEBCkY/QVxXYGzbLYBvMv
5r0G1rUtA/KrUC8spdDnZygKSkpUWlKT0mzMfU4ioqJZW7R+Ekx0wgFtqHNmDmW8bfPhJA/IxUrC
7pk8oBULUAvrJSXfhHnfqNX9nwaWMqU9so9Mq1PGMIqzYyNBfpeFByFw0AheGWWCW4iYQmt/zIQb
49htivuphMzxCZchEWpGTMI+Po1q1E2+U5+rkmpUlzoU05jJdOyHPxx37A5CREQdfpldGgXwPr9M
7KeHiEK2tmTdndQlGdYtMPF4Ln/wrl++m6eXCYDaeQBEQ2I8jWkEqhLzF0VcwWfzCQmggoIkEVhY
pozi/2824hU2qDfVpPSIMP6sJodhuxK9J9S/n9wrp9CCVJG3+LSFTIGTnYU4ETZqtNE8zeleZ492
ZkupyYEsiVqdrekeBARGbGJG88MtEeTWnEp62BgxRzh2vs6lbiKR70yjdBQX4ewyyfIyPdX8VhG9
/zW6rnR4q7WUJm6GYY6SUXFZQdhuyY/RuTqYh96U1Hx3FBjlrOjtgmQU/FjeMJRMFN3OXBDXpWWz
UWSO3SDsTiAYP/YuShdxfzham5LbTelvUF2/MJZJswpC3U2NzuBU6GvS7l7+d9KFp3mRK3AhJyZf
Fc1/P7q+tE+fg0ySrMnQtvOjlxaWDAYtvKV7AipklnT8zrZMIB1Iiy6mOVkT0ltsXsZibmlrF8OW
pl4QcuBoazZLmqLK6xyg1fCp4Xd7TE9GKCQyThj8sGIfRyMPzXUuo71bzAqhtOOugeHRkFXr4oR6
MJCEZvrv6dDRi0twCl4EO4S2Fr3S/YySQmNtIWuELOR086DaCSgVr3d4HqGQNcDB+CiJ8HeBUPPM
+Sbgku7e/viVSt9VoFJkxco24Dld7sHkzIlQjGvqmsfGyr4wQYviDBTz+GrCM3PTMpjHXErTye/9
HJ7APSXFPloTxRT+n94tsGvPQPjsD8NOQcLHirGTNOrb5fk61PekMYhu3qHjtbanroZJ0Etq8D6F
rL2mdmBMkG6pfUWLrzFBsLE02jifq0S9oFzsZ1sVpKIuz3qOnNr4mt/R7jHL1X2+D/1+tFDFrHw7
MVaIojYv9BF+MQ+owNs7vCiPVy2VwW05U5KTInGmdRugQD/hkXrif+TMD3FGD7pcYq50FtJmiUK1
eRze3agqqJKUZtdDaK0STJsiXzt2yenI+C5oqjKhdp4mpfim024gwCxN/79NDTIcjFqGN8o6Rqvw
VCj25COieroMe6oTJUv9QtpU9xUizr6DKjZPF02sa80411jy6qDkhIAPS8amnOGDxeAjlZlIQARp
86EAI7lu2ootK4lDFiMKAYHXkV3BC0KC1qZ/BmZbto9DpJgE7m+4wjnoiPV+tSw3Pj4yRyEL9Kde
uaF/T2zc9u8cuSwGFD7yxvSwSZBFNU4/QvnpntOn4s8f3Js3xF4xLGBSqxNzY8jKvpNbf07FDKMj
CTvTqK0Dixu9ccH2LDrmOm/noB3hAmjY4F/gelinPaVKa37DXE+Q8NplB5ofzSl6wz3tV4vA9UMb
kpJbYaaMavRame7a9RGQfEqaAzyyZD/AIX5MGCeO+0OYItBrgGHoMvIls6vaRk+g3yJD+VcB7Yy2
V5aY9khRvw13XuH3/IUb/Mp+/Gk2Qiw1ZlRt2af8uvWp+LCmHCUZeOSMVedlSht8FNTd3pnbm7zO
WEyt64gou2vo7iXAZ6+I37tJmUez2RszhIMVmfHvUzv69c7xa1MgULLMjIzUT3nmgZgxi7RumyuX
OJ61ub3Dtu2FgmnSohwfgiHfY4N+jULlortJej/ODcKZpZB6Mr1QVzmSHBPdVoDmCxdFQ7PEcC35
krcIR63SefUsWK9rp+BFUyIwZxNyXJpHpzaoTLV/Gzi0Y0xwuvpGb+XOyYi/qGZoxvNtnKFwVEnK
oMSBgLlPsyNCLHL4/BmCtuWE1UoeBiIo+5XSvvjy35q309GwA8jPkTXPG+3/jsRscxrFpiHMWbpo
EwIxAfdjCGoHj91i70nyP6e4i6CYojwh9uMXwX7fYRx5S7VZLtqJSlGv+9v9PFn3Oh+I3JPZ7oq+
9bFoc2HBy4xTgrVMlgTBCjB1aUhUt1tV/N7nmEfFjZYJ5zA+U7WsSGa3KFSBHD2p/iJbBlYJusZ5
JOXjYnK8lJ4VnXgo+Rn4AkKGZ+EiAFB9LwPIIqnv5Vap2hu6h81LkBfCneNmiW+WBHBp7U65Ht4T
tsNlqRxdbxSb1pTpytWQnKJs6lnXYGDZ4JHGX6sj4TW67L/uCIRRsxMd3CIRZl2zCsxOvXbWbrsf
Njb+YULGh2PEnSZr8Zhy0ipY5ADqW6+77Tpr04kDby6VNiEJFIb2E6iY4SiVXnf7mHZBya8f4oba
pkNEQN+VzqcRXHudgKkIKImcDheWIdJmVEz0zEnMLcYA8WY3U+bK5/4hHjDr+woBxpX8JTs80l/e
QPp9aKTzDFfWZaoTe7vzWUUv6hWORGlUkCNIMvMWALQhF5vDDzNqjsozeD2Pzf2NOPEes8Kk8G6X
tlM2acUDmw7rrgRlx2NFoAi/wfr/dBw9g7dHKDuuWdhtHAM4C46gZqd20dz4Xc4q63o3MoZzVyow
+XlhOlsJnAnbztI/YybeSmOYHAbJYhrJFc5/j/q9+7BWYMnxahiTGPHAQVLwO9VA+25521ybHiYN
MComBd7R2O6EIhQJ7pmRxWY4fME6RFZHv3ZCKCdVuiOPALMsukkIxcswjlW9WeDhYAJvBS1m72Kd
77htaCf785lB8kFm22ZwiCq7+3z1fWDr+HuCardbpyrZrEvYDnr0Myaoqv8w7kZpc8Py3Q76KIz1
j+3KVtEDiDM+A7bcPBKGRCr6mbrldWpCtAfCakZkDafbVdCfH/a//BSzlbzR7avslbgC8aXCrusv
KNKeTe2LPfoFF0PZA+GqC23Q99fLNavoSGbjvb044JpHpa1aVXpy7gKVFDWG+bKkvO8U0FkkNzq3
koq6TprslHM8tLGhSUzvmsSDmp9ht7OLs3prK5vEyoqrAskvU4YmK0ogHifxzhGh0QP6MnglDvx/
fUixC8T14pBAwhJEuKDUNhIm1DNoDeIytJLK+tjF/VROz4rMcnEEmihToMMbDrMu9mo0REgOP51f
T8YdX5Qg81o8vo3zH69SJOwk+FJmMqI6QJR01whfbUBgU313Kve4KfAtPeBPUmUrSRy65y7eW29a
XjjjXiNrcEbVGtYudBuf3N4J8hZqY/nsK+82hsbk1a8eUJVRdEBPQruYq0FcConS0pGtbY6l/8nX
AZBUxLi+odTog3RS2REfNX1Dg9rOCtqffhJCmIV7auEvYEbonNteppO4Vt4Uo7FyEf4+SIMmvAjs
PW1FO+sd9ZxrILiX1OsfJTkJHHoXBa/Qg9+2Tk0i8sr7KSVG0JF0IIfPIlsWpQnoIWUmhLrx3DP3
wD1A5w8QSv4Gg9wTVxB3iDkeIQXWCOz7DaPWPOQG/qyYHMGiPoBzrlsj8ndEgIIifc4+T91OFlf0
IKuXpLF2tQaprP1Mtw/oPFWycKnxZ/i6o3y/SL2Dgl+0e9n6iNYrX1lzkrisyuo5jdiMSYeOEpWe
it/QaNxu2sfeTGT/SVxSVn3sYlA5Zgmq4nNHCDdhPNTBoY1onS+EpuCxC1yWp8gJjKnpSL+gbH3x
Qr/o/zRXAkZi4GEr1VYNoOVNYPFijQ3YeQUrI+lKbZJFJ+leeJtYAI8s+qrRcK6BE4VacdMvvljV
MqJZE+HCVhpaw8TFrbLdyUGS3zmNnWZgESu07JR9i1SmMecj+f8pQzYAfjrxjmuf5TU0rl36136E
jwJVIfWGK/1NaQjA6j6MxkzbOB1UOA7ONAzwJEfAiFh6QBkQpGMQjUNzk3tDsGXPuJikTYGrpFSs
dhejiqOLWn5oxR0y6XgoHNimi/V3ZaBPmTo1zQ5pEoZ6bDK45bxxNSrWOWk36r0U9n3NveHTaoby
18xsCzfQnuOo8QMzdRE28eAqGEi1D0Wu6oi2/iPWSUUjAw/rW2Ks9Z/KlOslSfaHbqyKQfczrExE
UbbHJzVADFRUJ/OReKqVMtwJarA0qAuFURGMVbYzYNa9a4qZ+2jz/pHbOLA7J8Sz41AOWMXyAU1k
RL0sQc0QCrH4lq+2jVnTZRBwqrZzglRF7sLGUhR8E0KCNr1vhO3SROAVEsFP0C+CsCnoIANzzJ9o
iSJKOvS6hq0C85fILBiScF86MuQ2Nqul4fxEaBo8zHmjSkhn2JQQTFF8S9oOA9R9PlbG0rGX5oUz
ujxyrw8oL73DTjKLN0Tbc3lSTfeucucQCu6OmahqZ20Opxk2a7CX8BDYRzNf7G10D24pVMdq8yJh
eI86PxpcWSdjFwwRQ0lluTQJPIDBid8Y+0F4dAL6I79MobZAic1Y3Fr7gGMsawGWezV9iga5Q1nl
c87aGM5SGuEOtSc+m6PqNyeBnb++a55VoGfeofSiHrEpds1w6VhoWVAR9bi83eoXysqgURc12Wcg
hdgzrMmbl0SdQjJlMvAkSiUYAMi/y55TWr/fgcbWVyBSuwMu2p95BvznC/Wbp5vn6dDInvJ18D3C
neC877oukpRM+wGN7E7vPRQIgBIuoZpNGl/n5Z4ONpuzVXSgqHnxNIlRiyv4+omEZY7KUu4TmU68
pQolGPAvZ5H9N5LZXZFLyn+MBXALTMxwDj0Q32eIqJWfQXo1acI9frsAVZRo1f7Wqh/PCiKLK5QS
jTzeSslD7Er5oQP34AKzr2yDJoGe6UYzP0nZrGQJxR45CFks2PwXmoyMJH3U4Plsys/Z1GRBB0n/
NjNrXXVFTwc9Fhr1jVfKQ7Pi1yiFgdRguMbSFN613ebSeKnaiqciZZh0D2w1Q+PiiJQAJvDG457w
vImbOq636pB6k0z8NMmw1H24O5/rtIL/PH3V/7XKL2pASRnPbfSdwj8YsLqk/JvKfyG1ERaCe24V
z3Q7zRCDFGlgoNWbeNuQbX/No9T+fNzlH8xZ6sEDfXI/VY/Heywj10LZBeyr8UHQOqy550Hpis1v
eTiFnX7p5VLH6CfHCkk1l2Fp+Rd/XF1YZrvbA0wz1k44TuuLyhufHn4BzRuup5qkLgj8IBUxA2W+
WXYfud5Pe6CZ6jGz0I4WlOOo/mhlejSf0i9lXbDV5+sMo2U8pPB2ekoU6BNgxsHo24xlzDOGux4H
3GRGzPPJI9dq7/94S/pH8AAcNLPXd04gwuVCA68OwCmvEaSgxdSY2J/WaS3GsAgXL/e6eFntADvK
z7cfPSJdACDxdiKDOXGgnOLg37EpshbIdE+Ex/Hl0L1hH3kTV6i5AJsRL/6Nyj828Rpca2slBaOX
xxcSnx6iEzHQ51yzB2eyrLZ9ZfwmZ2kuoMneRDAMRJGyOk/6D3EcQNf7w2xkeDSCGZsmowBOTAEL
j7AM6Cpvn1aHJfRCa5GKusoYJweSRvGl4xZ3TzAeoNiHIL4NkUoMAxi26JnAVPrhvbmGaufAqLgP
rcTH+cyE4mF06NZIqYM3zyLO8sEXaTNfDVP5Tm+5Lvqp1H37LIJyxiqcWGMznunr1qxDTWbe4oWx
VKk7aK3rQuApaNPdDZG5cry97jJofji0iBZRmrXE6iaJibpzsgYUK/gbqZbrzk9V8hhsBZU5QBf2
lIE7QIQNMj9RDoMLyWLleEGybokzhj7Uz8dCXub9e+tYo4abyH0oINZYr5FQ/qFCzXY5ZVwSRUco
/caKHxLSvv5Q6lOEcC2tecURxDriPt4e0hu4BqXdCYLkBRCNYNSj4WmN+zUrr8bppnD8D9ixXjbK
ABIMo220x+KoKQP+T2cFypftipBz9htuel0rkwycnDzr2oGp5QTlystlfi6zB36i3k9HwEFzVoap
xmOjA8imOZwERj3VlyYLU61ue/zWqFHn5xEdNGSsqxcRuNK9sed92Ct2BW63EhhxcilgPjrDS7VG
7nsOyUXBIyhPYlwGSsJOCQaApLHShxrG6PtEs2KHVu9Smb8UibMdvVhp9k2sjSui+vbkO4/k3zKn
SJ3fbTIZrtxw9jOzHysT04M41RthPTTHubHRAWwX+GbdDeQqE7d0f1SE/o5s3RjRcj4f7nO1myL5
VWC++BUj44C2ws7kIF+jwYSFClnwPOvRtVEi0NoKWxFdTazWzdTuPhD7aGrrjFsHfV7tU31w+rj1
YEFHUKzCbMNyQC1a5QGFztt3KeM5bgApOnNlCxA+ULNpYg609AOMPk/XRfg/xWhaFaK144RMiSP2
A0HnO7SS7dDe/87N3e1Vlz1X/zWJnZA14w2d/CRasELZVy6iiwXYB1pZWZYm1DIVBvO4sI6tpG+b
5vOiZMJbPzZLLpPGx+zI7VUDrzjhY1xuNL8tNMnVU7tpsYH1GGH0cuFO75pS5y/D/F5axQFqEg4I
Ann5PH7EnlosOrou93YdlefMHxXpA5fbKmNkotlvWPT4KV8rJ+3cdmw6MjiaENCjV/vGmDWtyyEk
hXieIC60mt6UVlmO1IxHQPKfy4QODr5QSH9BKsIZrfc74O1VwMNdzkcLHhXOO7/jZBsP0/54qMKo
aFr2TQ2P9s8h+mpk7pPpy/pCz3yDsKIy6GdNRgNUyG3AhBgO8Zx9sRuYmHGA3o8loNjs46ERffm8
WhqUKGRu8/DqxA6Sq8wheVinApSnewIYSMuM5bElc30JOvRKrEAml0SqxVJKflcZ8E9jQ5pQJaOs
vGeqCpLUJHj+/F0PB5iu4d4d2DDCAhcdKFfELBJNU/0YK3lIOHco7lIbNAP9EscY6sZSc1myUUWx
swkt05HovJzRkGZyl6VxSBBvNu3fpD7KztjL9Riu7oNj4g/U7KAz5qm/PN/cM91AodXCtjM/FLy+
BWnsjtobNmp1l5wjccpoZVxHWXdxZVTtODOBLcv3Nh9RZWI7NlMui1bDLy3KHYcGG+kONniAh+cH
1X/YuZSUeYOU+DNdbI2B2j7XKDflTXyOic/nIPh+e83NG4I5zlvbS4nmOjBLAoe35XFq9SoMVkfl
PwHmXl8bHdc1Di6IOV8vzzrDIPx781UHhu2TD+n7Aq5JEdK0ld4Kj41hVgrIh+eo+EFJsJ+feVwW
cWaZeiWnjpXM8LofsObw6ul1R1y9yUoofB2vL6rEFCTUOtP065h4oOygZ+T6mlLTbfWXlgjea1q5
VcNizC42fJjLtVG1atjyr+wfgdEAR5OS/hz29mM+P5bQ4SjM98zwcO22XKHDlI+1In3j0mm3ZAJ4
4VCZ9QlVtJp82E4fM5ieqv0gihJDA/zAcu7OtuKo8HEkcKz1BTO2rT0N/yR53pxqGAFPQIDAW5Jq
k+DcHYLGZM+I4CMGnObCBJTLf2m1iZLBANbs3dQa31ocTPmyGxmWWnAKRswOfk0zu71fouMAHYLk
hEBlGsI+EpCdBe51KmMkZWJoDa5HCLgiTJ8kJJ4xNJO6DcvjFUKXY6FHGota04G3pvo12rAD5y3j
iqo0YKJWfVNv/J64F1mC6L1SBzMZqqE5rKHcmU0/GdxMHeFFZbvOzoWyXb3tQ1W98JE4Y1YDf0eO
I4nTC8d+YlmUO1dfWavcnCPwDOc5Qa+hHqNPmPxRZZbuCADcpVuxFuhTJ8940xP23rCjgRCeJgRc
18QCSlJ9jSIyAQLOaSFA9hNae3O0oV9cfuK/raW8vnybvCoQKG4iu3hE+5vJfkWxkfrSwJzWz85U
pdhTZCTvO4h7d5L7Yr6PfJh2Ge3ToC7UQqSnkBR0zbxLtO878Jg0EDTWFvZbR3gX9JKt/aiPyME1
+RzgTBpsEldjP2mLWUk9r2DEOOCnQkT5gveWwdubttLQmsHXQtYAlv8Z+VLgPqlqyie/BDTigDEY
wc6v4sMmTyRo7eVRW2v4698me2Z8AJVRlD/ZlQwaxdcrp+qMQSJi2lE9d5RtervRQVIcR0UHW8Ed
02JP4ltBNTaTwBT5mVb31PG6inLcguR8IXrPIRvpmSSdfjNKgZT/yfVR/8XVmLWOYYwXwpHrp9vy
nt0BdrRmQurNs6dqyYhFE9C0k6sLMJuu5b7gxcwRiyoC/Tr3aQYXIwgFjJQyRUCYMOCKNJ6LsmOH
5uf7AGScewvjprLJ7DhjZOblpU8ldm0V+HIZDaJi+oadEsgHGMig2pr8xsXiYQ2sGVnnqri2KSP1
4oaxc8Fs/AzSqGVSPFJFPKJOwLDoiPT8O8HuEctZ63qI7pup8ZYAn2G/lEjZrQtgIG7fcN/I0jc8
mm7IpiUsstcabhhgzx8eRZzi+JZSy3I847DkGpv5jj+puXVAM00Exxnc8+qd4LzNK+QI8meR48Uw
DDyEvaOsZs9NiIxgJ2l5x9fb/seWbAfHBeTXDD+D/JdznmOtxGA5dUA7oQ5G+8pWnGcpraCYguxe
9XMkCcCixv8Py301jOmjv4kRCr4w52gEV3BDiEqJLD5w3MIy6ydCmTy1eMMX4zTuP0EqKYAEwO0K
i/2k/lrTyEPwMOt9WwHlN97cktw/3P4snZgiAoC6oJJu/eksGbZwJH8u5wf1rqFz+fPpXGVj7ydf
8OcoUSWDFQObzX/KlXLQwbSD5T+ii7eDQ4+qg/uAMQjqbnOt1k2ITCsRZ+tatwoZEXZ0tb5i4Uau
GXZbU1ZBWR8OiefK0Gkxq/Y1dPwRiYtTVssCMOx10gDL8oNxd6YbIGwYc1xsfPqZtff4z3ayicoO
N66DOPg8A8ARVFNQCuf+pYEj857lQ0UhMzROv5GfoavUWPMMdod34G8EoRBJ2/52MrDz3DoR/xVT
6dY/zR2z7Tu/EVj5gJRApl8MCWZFxUWXE1LzIYPf+Eq2bi5lhV2hjEpRrYSUN9ZYd/3cUPAZIaW5
n8yIaetDPK7TAo4pHN6QbcbXWq11x61U3vg15RhtoPFMbflcc1RG5bQkNXyxW9kcV5bvviuYWqA6
/I7aQXF/73jlHVWRSLqyHYP+yvCPxf7JCD1hUWoflAhEjbyBScsAQ6gWSiydjyWS0bs3qcckj3Fy
ZiTSoDIQtB/Nm5Z2C3d4EH7CRFUlHiLflm+pRHm5v1Fdofrnlu/PXLBdCTCsz5Ii8SQ8yu33/Pzj
t+peDXuRzBOMg2HwHhRE9acz/u76eOx2wCzk/4/H2KQcwLNbtjxYhsKX6FY/RjHlJVm1vuMcIm7G
GRRDhxLlqBQK2N+XvAlv5NwpkKX1XWxrX/c/nRFJv6rXWstOGnesHo0qhyr7r67GY9gveZI2wgsS
EUECxqK9wh9QPbuw0al+PHP3OCzK1nF8DN94AVQo90n8z19vqqtiZEu4koAOZiazwvFJRF7y87mZ
gX/RcoppIem07HIwUHjWCDdB1PjF0UiSP/eVGKIKVNiE08rmrHn/gfDyY7RWUnd4gWPRHborZVSa
3g/qW8dQU/wHfghmPLEyXQk+BUx6PNKCMStFRNMdLUMut0rSDQAibIKslLlTs/CaaDTQJbLQK7jM
QEOHpouNoBFEzYhbBfrbFSdPFoDkyemYq4i8o2XMi7ffNMqfBeJ8CA6sa8fQrFIbZFrHTeIApgLg
xJqh4hMKoQv5dR4h29HjQ6cTawgjWDZvRLPseikWKUizJuZnlh9JeuWi5eGbOwLWpRHBqF+a6LOS
TR7H5O/0vCgjVZYAallES1J6DnTFHYqcK0B5sYeFjEJaY/Hum77O+XrSrJ2jFknR2tB4r/Q5fBtQ
cGTeb4ll3m3xQg+ZHntn3yMa/9bcXyWWVN6/ZA0L0G2M1WTjqeL1XYMTkLgetyAyy5PqoM+ydx8m
OU6lgcmMCTtsE+XSQnTmmp5cOWsGtYIT+KYKlkZghkzlapPcLVzw90hBl6gcw5eLYDmRBG4JOJBy
+3JWBWxdrRfByHdu9rVxDrLkNRTsttIJrmxQLq/qrt3iyn/v8FtmT3hptUz7BXyjjnRws8sutAoW
lnz3/a5wiUj/bYIyQWQi7Lfgg7cWCcQx/ecNuxg5jRpFVPM7JC2s+gIY0OyuTnkCJRIFUHFVcQlM
N2vqBbQPkcRHWDS2alNBaaEO705bPNYbocSndB6eU/JZH9hoiAA1I1UcYsPgo4q5jMMYU8eNf4G7
8QfMxnkfWmd/PYMLQAtLsAO9fSfy/gZYS0aqMudLFR7NeoVgCwAPlB0NN9L51fdk0wxfe7xKXPB7
3WmDr5O/oNggChugJ8PE1Os09XOX3Pu2fe30OcCs4Wdp43fkcKGHS/+BBxc4TVgz/JsV9sqe44/5
2wOuTJ2kSJxhYVXULKlVgQ2gd2kWzE5LmNlIeOVujAYgm/0avk8CWuhZ4kHG5uPZfydxDNrzKQcN
ap4FMEFN2P3X8kIxqIt306s7xV3r8w+gA4+cyr4zSkbr/2rsoZn6rCx42x+DqTF3l/02wdUdmBX2
bfkCoVDxfw0/jnd6MVsg6kWzEzhMFJ/6HJHvS+oLMuHY/kizWyCtnDnoUA5fVHSY2Eqkq9lhysLi
xo/fld5yJmTsLtpna6eJvnDrEPBxlRSVPPRXU6loo10FceNxrO8+jC1VMz6+DhgxritPOQtBp1GN
hpLK1fdiYS7K4DPJx6rLPN9jhjrOwi2YLLvBnPtL7ycCD8OpKABSJxFmekIhtYO0jTV5oUlrh2F/
KjeggLoyvzq/hNaYCNdFIgOOwETSvUO7WvBLWEfUVzAAxR4327nPRaItxFPXYDJ8rTujI4GrcF4i
BBfa2uqJlqxUD+9OqegyqzJ98sCeloKVq3D9Cf2eEDEprfvQpGUCTHv/9cDXGKYV7rfr9Bpt5DiJ
CRsadtdq5qRjaeYptWWcCDpEDBgXZsC14Mh2vU66yyBsBFmy8mKkSKIORmAOZ+WryAwWo/U39+W+
9cRHmkBYrWw9gi2acGuynw3ATH9uJwZzlhzuekFXfSBE3xF3wicHeG6Slh8wqa7wOorDwbmjz2hD
/MTVJpQg+f+pQ3GUx5bLwFg42Z26KkfuTFPvX1MTnjMU+eE7YMDVxBCbKZD2F1U3CagoSfwmBk3d
MU2gDDx1xC2sODxCk/K1gNOZKqUvfHCf0lEN2Au4HTW5r0Ur+fkWjMSgDBmKTNd/x+R5ckAoDh1i
nK/3xPpXNoNCI6CVyMxw7m1Aj9PVhBuIrcNTrGGBnKZLqcFGegoNdqfwNTnAZ3XD3r79H+f4K9t/
cJ7EIGjCOf0qlyT6gZhvlRUuIXb9WnRCFZWIHVqBJtfMlspcq9Rjnax84XlCQnDEKXiowz0hiuj2
//LBmonysPwyAV2pbaaFDV1pxgYrRT3BjlciT4vJhwL6Qqdk9Rkw0V8Dq+/VHvjl0t5bev84XIyt
N+mQt1s1iwVp0V79guyD9C2WvOZmgwWL3s3ccTARJ0hmp5XHONk9ZOyRCQPDhavBOHFB3M5iPUdZ
PJLzz0mYoGR3j29baXhMZoBCUU0AfVuCtC5xzPbe9Knl0pnSdJEYTEQaNj1OBmKFc3/wRwuw08c6
RCCV9fDnWhGUleL96FAkAhQtyo4jsVp2pjd7S29W7zKU/YPHe73tsNi8f87PbWO+RN5iM9KamJYa
2qaun0C27MCdkGeRilkLIJMk4QiE4hhRAZEll0ekcoaIqIrmc2IwW7KR53+P+uBsex/gI6nOxqWr
dCel8XAaKpikv73lQy+MujQPj0QlL5rj9nmJHwTyu4x3LSfnIxkbIHOJ9jBYWywYYISHxkFOFf8N
SEnXyBJw1q3jWRRo6D9b5bmX54NnKZh1bEss/YmzSbgJ4EgNfouRFObA9B0IaeMEup6pK3Xfd4Bu
AvknjjHQe8253hf9atX1ynx8X84U8svMfMsHwOBafSoBcbo6f1uNCrvlCw/v0HqcXDyXZAgYWjCN
XZpIrsu6wOnufnXOhnObolxQvnex70QYdZA+hJgxddUwazaqH5Sl+QuN9AdDsLTkfcoqO2cXYBWn
zow4uR0zTSVmEWXKFgwvtqkMCNG3S8UOTRxJWH+rd1QRjLLykyjG6JCjF2yZ8PgAvcLwY6IFrvKI
pOzfu+WL/5T4u/uFjDrkIMOYD0usNemVbsxOlJFBLmj3dh5kq633vsi+BCjbafG99KzzJEzkkijY
q6KtPbh7Hp4fMgw2wv/Z84v+5V8+lGOAXBhYBlJexYxENFMUMyPoCsxsMlg1GTZ0BS2kdt8obNh6
p7Xwn67XFwkyxfOx32KNBtFSrz5TeartMGZXz+4PkvC66AugVwyieBG5X1fYXnWlA5DzUZxEFZnd
TQsu6Z/syqlU+61sU186lLbp0UinHHZLm5F6n2rrLzPQwDd9euFbB7GIAMamBzLoMXwSdIo6wpom
NYcnowOsu0eiikDy/YAilsVWAGkObCSwsCw+goTIxq0Zy+WF7jaPylyyV+kqlW5KMxkDMi/KSXFJ
QDNW51xnoNUuyfP/UPXyx9gHBJJkNls6uVmucnRthVVq8LpOiUDHfoE7pjlMCVPSnvz5MTp0xCnz
rumMmBfbVTCQqfOqTIqYq2wBW2nhRhYCiBg8Nj/TIWX4/RXN9w1ZRhrdK+SpXEanqof0NU6STyaH
yUufRZJqXlRcyFSzSjBNfVWHkBNCwpPzhg7mjLr0mFGLEj33xZx9khhU8Z5+EUBujIK5Ci/m5HP7
3WzY6xK5limEKSqpyFXPc8lIsYCksWjSZNFRHxFNh5xCSZbZTUvuijKgEWLY57e7mLSc4TZwrF3g
oNJdeYP8YQf8vgTwJyFfuN2zc3x7UiVsIv5lENW+Tj6vjTmDMk7IkmTowpO/cDYX3Q9Bs5gTS1Qr
0HdNJc/ONZu3CNY7D8rqk4zQBmrpuv1T5MoG6kQvZ4YqKARf1YebgxYPoIiB8xGAF/LU5eWqoL5b
UIsOneteZtmX6Dsshd92/dlAZ51Eg2Su+1HSIgwpWdU7F9C3gSMd+ExbPiqClgEfP5yry0Z/qD8B
jPSBY5AmjaAsbuYDv9lPBmWsplyJtQFLKixlsNPC32mH6E6lsgNvEGBGjQy5OVKU6Pmeobwfoh5B
lyuWApFsdJtHrbIvdhMiRD+W1r+/8xXO6FJZpcK6wDgdOesVLo5dtrGTh8yaagKmNqYhb2wIqKSa
I0lKtkrru32eP27XXyw2cSqSR7Uc1sXkhg7KQfmTPZcxzfKaGMc5B2YGeg0MHaoHZ2h+Ey5mU0Qb
x8av4fP6hItVPQm4Sp+GXFoF3a2XvGiQ3phDnjBrXWxw4L1tVOTsog4MF23hsp7qsSpqwGFbTq0n
zxXhsEOT9ftyI2p0b+pPTfySCypXzMDxyy4WSTxc4X6k5iIIX7Z3eZJRQOpOOAW4XdNOS2JSitQq
HC9v4k4o7QY0IhT5QFQ5SDa0gsSaOqQsNHu2A/4TtQUmYnbaLCX6m7mhooOEDnDf7FqkMHOfOSwJ
QwW8LdrO1L5SVpkBwc85+t+4sAFnbJBjLROXafVU6DB72N8iFJ4iMf/XTH5eHShqv8JNdg6SSVR7
OONKSC2HXxouKNY7AMtNCI60O3onOxjc1cNah5dactkPSnmvP5+2GcqAvakmFy/QZMOirsccPa1t
5FeZOtLUZn4MFo8UaRic1gONGNM1miUcNNezwgh+mjBsSHBD+7UQbvOY4NpYtT6sB634GKzgKpPD
P5rOc+uLnoGzlRYX+YsIodkff/PiDBjoWEG95bC9kzr8cwwvYYocW2NCFpmkdU1f7yXKBE4oQyKT
YjM7EzE6l+80Ae+6I5yspXYibVbwrgu9+sEOBKKEnByHY2VZFT71eY+/kf8/C3OUhwNMYE9rrRiH
Rl1AUkK3pXisR9uPHaj6eZ+K8kwDmUAhaFDYZAABxqY9nfrYB0Crs0Mr0kWttRdxlM5V8VEAmV0Z
bT+dlNAFe13PK/Q928KPRXPNCJPU4z2pJjw2u3iuq/ydwnBjewsN9UOES07Xos+HdGZlijiVEqjs
qWVkuJ5dIQvVeHKgrcLu/FrY5zrVD9sdp9rJA52e5T52Wi5nF++hVKkquL+/rUilPF3P7f+uos42
D10JLk5uuu/qwjPiCctHkHTInz34J8xH/Ge+tpb4SBP/JrzSscxxT6ydaH6s51UNVPBQX1vrInTK
8f4a6XD2gWbJIVohDbwnu56+2DOf5t11ezBXcaT5HdeSUmbKJrDyrJwRgTrfQFhCT13ql40JaLPN
VxL6HswM36lCt2DTYFjyciZ9fqEByyIyOQeL+7Wk89HpSNQeUjb5MKd0EgCC6F+8JKbXVtY1y5Z+
qExFU9AHVjSnvDbmwZUlV941K0c8NEij+Q7QP1FIV/qTqZIO7I8+IiI+qtFugX4d+/TRXuAjzXan
TH1NBPxjIZdUPSb2fvD3Um7PsBXj3YA+VDineO0VQg63MrXvxtPlPGLST22tdku3+izwJh2JTvo1
aC5ftrM8exraL5LpzBKs867FQiYFADXekX+pS5QVCHw4tzgnAd1jN/ZNXYaEdLzd4IY4k//7TUpV
7LWpEASadWk+fF+v1Evzk3v5YZ2lWNwR1Du9Kjtye7Et3PobrnydkOVxAnK5mFlOvgkoSlDm5nEz
8h8pEHTbUnZguz8x4DyBoprjYtryhb75J4s6AGalZ4yj4tVSygsRUq/TyqTobVEeEdhc7rNGWKub
gwVYLSe1nw/Ieaor0ZEuG3t7Bx7rctV4AT5ZwP6vTA/JpZtgCg3zfzG7LvNCubVW2096xVUqx3ij
Fs4R7zHhguVNgVyljYU2SC0FcLQXJtyc0d9eocoSXDEKYem2wdo8iMjq0QzvEwEYEzHoJPvmgKgB
yR3FspjLbx29Pimeaf/GqUCA2xX+vl9GvmiQY4YJjfVajrTVpIQWJzngNF58Qng9kNRRMd8N0vLQ
80T/3+CIPXDVfcC21rSRW6biVDnXgfwcwgjGh4u44GDxIGkeaGgxo9fca1X2ybKUsYH4/sLOzPU3
faNKFuxmMn+5zopVvBmP/EJlZPxMBfauh2RTs1PK8OT+ot/HyaOakg029EdWe2lqXK5GzvBQYXUQ
VE2o4JPYk8QnCIhymYq45yx+1DghJd1QoDO2euwMawjVFMBieFyvOAtbCYUyknDF8Gbxob5lG4VK
OVRnU/1BvX7XmP2MNqdl8mGRTjPZFi0ttG2z9lqNJ+spEgQi//qbVKCz4WwR84lw0Uosdydn3ai4
c86BeNDp/uT6z6Cq+vxBaz9/n6mG1xA6QuKzgocqijsf3LFDbxPFh43qDD87aeX92SMiTjRLqQ0B
cKouOlcJNFVgDOtsI39kUZI3cUDLNV+d+KcxAQTeMpLzM9FbsOjFvsQXx+s8l24sYQ/uA3dMf8n9
4zT0CECLcmM1v2n5KRbAChLVYGL/ao9DGnBeIx219zYkl/df8PG2BM10NVMbmhLzOjjBDs5gU/8r
gsIJ4BfNGYmofhfSaWE32laLR9BOrP6nbI/wPJMcmkfrhRFg4+FKofcT/6hmThvSrUFAqOSawRwa
a7ooZsIAg+QL2o1MPR2n0iAvm/UpAuyANtXKKiqo0VQomlQY8+Uc4f/d/X03K6R2zMSuUDsdd4kM
3+6c4bPKzSeOmzD5zamJvOTeg8HVlELoEDu89wRj6S7PV2GQ14/LbGzzcK179CMcwMKagT1ZOQEB
ZwNZmWmIyeiFXC6lNFCi4qdPM4UK+mQBZhBdhp8FusWpPOItwhvbV2wwPEt+L9Gwven6pdgbE+GU
cLVtUjHVaXwfbXV0q44x38cbJEK9X4p/oJscGSYhgvrKHxtqiEPl8aa0epeOyZ7KVD0gNvJL2b5G
E80YEH+0N8XpxhWgXh/t8sOd0r9tOgpgyvnsyRo/0KHDI6o481bLfccfjMNWvPDwhWPgk5hA3zSE
gTSUN0Fm3NvQYYO3BVV+3jN1Bb0p5TyZOfNjZLVAR9utzcYMDaPS+rUKy+W5TmiAwAlnWV9t3lxi
0TXUSsl+yO8F24B7CsPwKq1aDMAkx+3owaIOfdnrjOFJCKBLE7Mxhu7gpsM4RKxBvWj2puovmjUK
8Njp/o0IgePFGH1mkQLWpZhN8CjrLsC4jDOygaoy7SP6ojLo2hCnd9WWko3DJ28hqNsvCCbfVApS
S35DPXtHUSrox3/bXbqAPCmr9YsskJgvbHZ7nHQB77XUXVYKzGFCPt6I2pTqpZrmp2LH2jkqsTXU
YDPjc3NWzGfZc4HBsnrWfBvvwjQm5AwDw4R6UG9TCOglWoJ4KIB1NZr/ULUDl0kUWKkebq75LI0E
HbxsWG/K9SE4ZkaRhGtGdoc22/Us7jtAQXBq/7ftoWsMzCfxL5ZQBv2j5uJ/zq2BidEMmUOzvlyJ
IzpfHxLC+RzK5P9WtFFUJHuBtZjN3wIsPB4pYuNDHVjqAVrKf/QpwTO+l5jd71nSY8AOmYroJwFC
cDycHf+wHBfnl3Ttgx42cISbrTcwYgcPwrqGJ356xyasOHJYsmmcWfjgtKGeMn1ZYeoe/Gund+B5
YKw+Jvm+v+rEFZa/YEeoXj8XfMVFY7H8UtCDhvjNuGt2aOjX388kds1sFCN0EiBB6sn+tYqiRNfJ
BHuKC7tE+jomKQgFICS9U8E9/2EnOConUZtu9v2FTT5+OJpcfr83ul3aatzEYjb4aawiXSvamk4v
AzHwid3wdwp6/7mctl2TMqwXWeTOmlnUtkxSSX5KbhssIi1G2V0q0Vosp12PXSJkZm5jVV5uB+iL
TjC5ucJqfgjQLCToESigpZ3EZZ9EOtdd2O9mhPuwLJa5vrVxkNjtp6aRdqhYe9P0R/BJ/HyB8B4X
Xx3FXTfqUMutrdPfjYE8JFwliRL8TISc/+qfOnIA1BqrSPRQDYnnusUmTzCNcBWnQJOH2KTKk/mW
JnsnU8JZigOm6thToUW6t2Y1+vUzTaoOE6wvD7Cil8k4iDo10St9LpOFn2meIDZUSESBAZNNajDJ
lbupd7wKWGCd8fTVt+emBY8goDHjJwZfCwCR0GdMTcCvto6WQv6R+hZ7K+e7pFJQb/EyfBBJzpDP
O0KSLTYgvk4mfoJOsVOG404eTltK/Jzkb0zXuSvfZALp2zLLcXgrj3Fb2qp6lH5OAyygIGPTaeWh
ljAh9CFJUbVhCSL1kXfLcbssaNBfUeoU2nV1HfedEOlil8gswUyfm55lp4zeSbTa8PGT2OHSUEVH
eGlwaNJvDKgBb04WfAExjgRW8gws8Xyr81eB0i7QMdwuE61mmrdoBWPu0KQ/ItXW04mzdHGF9GyS
QUnvS5A8+EOilFQjLFVGPgDUMu6wQTeO2e6g8MjCLiaU8m2uqdBYWlVJJsiT8UNcNiKAlJdTYOCE
u57E1FtpcpuD/gsyVumN7wEEqPvW3btwpgUEC3xvmk6nyZ89vig+h+l/7abPIhcofXlUwexd+P1X
Bhf2GtocgUliqTDV+YH6bRaUnKZNAyQHtgZddba4v39mNng44JZk82XA1sO4kX9EvmR2eLv2P7rB
rk/KsbXyraM0SHVyKn7VKodZRV8cvU9oCzA7jAjl3FRj7Dk2AhtSqlk0Ax1B9g59qMTbzj71l9m4
1VUrS57pQ4QLNtBPb/HGyI55l/BunSiU/i6yKhJwYjQ7cCt04A6PDqdP/V3Q0FIYwzsOD/++8OVr
4Cy/P5hNH2qkeis6HGD4ufCwb0yXcNmmgsyudrxl4iTz+w5M+sOGevLVyo3UKkaUUDK0QoHYZc8s
i+wlUorHxSqwh8DIqopGFrKDihjIL3En3axuR6VKWMa60aHAqmaIevW0Jo4wmX65Y+inTc7LzLz6
QRhOo0s5Nevk1JY62i6Vlg6QjjX/gd08COPMIW4egC1lxtiQ8+Tp4vX/yXBxox0ei9ad6Pp5s5lm
Y+mSMLdDzzhJas405oh0iugUSSM1rHd6fGPG8O/3clUTq3lfiJoz+bWjtz4PdXsGTlkFEuJLScBx
92atOgM31q7opFOfcdDGZyEzYki4Lo6lRYrpuUNb8nBgZb6MPigeykMnwbpszeLVrKq9lZ8IIH+j
byLTlJb0FVcB2ARhMV3I3hZAJHgQ5OFRF52pAROVXuOnrodHL9Bcu9XHPGYu38uCk/MqTgbeW27M
Q1/3zPG6XBI82etQqULkn640srTr9aFh4X6CX9s7U8wk1BxiM+Jrz7gSH2z9w8dibq1qQDVxKwtV
lVQdz+acarAonnUlU2n6zwro75A3dwXFROLs1nsrKu4LcEDRJz4g6uidVmrPXELKr9Ux6plfOes0
gLdFb0bBPKZowiNgzlOWn1877emQ8WcBtRDtCWCLulaUzByrEyWfoXX2FF+2Upv1/Q+DW8kPf/4F
NPxAA5riNfD6gKx4AIA8N1bOq7jJUlJ6TsnM/8CLiZOppvo3SFRdTA6ArXv/4ms6EA5b5vFjsScQ
sLki7bVOzZmPPqlKc9bcJTBgSCyhJs/oMZkglRwKPEKiwYtwgTpilSmuCNuTkKay0KEBWnJUBEIr
XjN7eb7PUwfPt1s4KmIWYwQC0mvea77y+h30CLw3+rncpvhq1pBVqP72LBZyeigeKvqKZNTkKowz
3se7jrqcfCd1lMRGbYFlzzhChb9VFw9pC9iWrzfAamWGViUsgmPg91SyOYejrZGFzVP4Bl1Yqd5K
7Py+6+waFEHDQ9mKPWFJazabjdzTiYCFVkaGSkvBNPhHMn5PeZUSqk6baFxA1TyOKbOtG5LI0KKI
7Fv1kpzcSSChzrU40P0qbxYqNg7e6dARRCnBMDR9mkV9YwY7cggakkrJ6fNiXcEgD3pyPno1G+Ep
KBTyhH6m805tDPUYFPc2eKQmpNQy2NXvIP1Xq2Y7mN6XhNwja70yGt0pu4QfKT7SVvetsXJIPCCh
dYqWzN+pgINiUxt51mwLKaPVLDsFv6+NEOBliolBe6lopFkxbPTRvNBZgvJ8nPTb43JWT8/u7MdC
WiHUtgb4z7zt3e0xgJ/hty/hSdOe7VNeXpv552RZWXfa9t6Jb965ZwjAuOsbXARgtIhE9BQKoSuL
abYXjWsemtadeCk8WxLtDhHUVt6d+gYovxSlgz3XJfMZyp31TkmsH1L6y83m1hPWNqtin4lGMY44
r+tBrsG03wLwYaki0V9ZUHcjf719NGHOle2ae2ZNs7e57Eh0MtZflaoxmqQAkLbz0vmZpJzG+Lkh
B6r+Up0NFrLs6zxj9fZpotN0YPpZgsZnBQu9Qjb+BLE4sMqtpy0ReVvYPbSRUGQCiBlilT5PWS5g
/KD8zVB3coK3zk8L/WnNJRVWk4itckiJpHoYLHd2AZcjhmAgMVV5iKuu13QDrBWSU0CbqPQrgKcP
sXlDK58Y1m0I910MiwmKZefOKcnMiI+JR60F1rDh3fmNRxWXdEu2wMDeKWfCCgSBR9ydXawVSjfC
AiOZSw84kkB3mY5CLMjMk02bICMo4YTS5GGf7mTnyPRkL7lI2NRfnosiF1yNQY/xkj+9RMiHYhOO
cCAyW/zdlOWhKaN/zO0LwVSVXTEE/BZwwEY3H3zns+ATgAQS2RxKCEiS20xk390+53gNksD0et0W
/2g+JYE0NYX1cP2EX5lvZRc2tWRrHYCo79Z3aI+2g4g1DTn0bvfRPhsJJuSt4pjBDPcEay/5bGbA
P/gHJHloOPw6vuaYsSRl0HhJSs6fIHyhvS2efGTAeJ0okXlJ/pJDbOd6h8lBVrOh1sqaHXdgUloC
/8TPfDr3/HG7RXCNjy5pXVAkEldBdJ91edsGD71Dhx6rQiOEitAbr8iqtRCY4jhD1g+MNdAw5Fv9
jxvBSQpWWRN/WtRmjWKabYyvQLQBpWIH4ZQyfzTCBBlU/0evWJVOpnu+fQ6qQPjOWlR+UNGnXQXw
ZLWvgtoxwb1+J8eEaR3Ga+kYvafE+lX8qSa/bzUfOeU79f1MmgixuhUaqnpBU4srJgcDwAMkvoie
9LI+lfl4KmFtS4ImiDwkjZ4F4IqKTpF4RWqnHzlIiNe7w0e2W70lVKP+0VjYF49qqZtcpGRfefmb
8ggohhq7scIDh9coWuKRSTFYocKAiw212z50qEJTLw4x9iqC4RblK17rzRn3gvkpY1cNAI8qYTpH
UrKFawqMkSBoudOLtIB9zFV1iylVLeE89jDlCkpdC1nfSMa6jmJPxEAcjIksRJNxgZxn5CHBNhto
x8fFPidsHbSe8PU5amfs3ZPCvXFkgGwDzryvxI9Hd+Fo5/eEMLEZJPAcxhqilZ3Q9EhGEtBm/K6c
dNL6mefh76euP2cXz0jmBQED0N5+bTxuZCxDYAkvGajOzAziNDzqOo7ilF3/dXveEqBcQejl5SiM
Ih9exC4cfbt8pklV7WmfzrG+B1A6VzRX4DCWzxq5aZhyUGydCuHeJs+E+B1ezBzaMCqDlmGso7lv
8sCLLKaorLTk38WIZaP7FvLdaXp0raZJgKKZgJa7+psXMkiszqeevDlXoMuVlc5ov+QQKDKkb/Lv
R3xTC2uqcITcD7cQh7lEFPCMJnFlReuqBfQB2eMrCP3d+8HuCQ6kyWTi5u3nJpjKyiNK52JWpNXr
r+2K60kX/vnAeP7zw25KfXs1c/3/XfPIn20vJEatLWt3DrJli/ZQg/OvRt+APRyziJotkANLj3q2
0xKuMaRF67lHeKdAQzsvQkw9yNO9caJIRdJJOyZt2Eafj6V3D8UXDdBjcYf1Y+zZfLSwqWMBKVip
PVpLgBvz/pq59jNsiXYAtqSvFpYEDJr02tb7oZQq9NOdhKTe/Gm6hdZ3guy/x37cgEgg/yuZdyTt
097fWdq2t1sY/nkMwiyNa116mJYskpSBIJmqteSoXSaNXerfah7d5X0375PjCDBsckXF12KuXGf8
OCrkj13z0LpJxey8H7i9svEFAspueYjD9/iEH/bMaogVyEh9G7f5IMT0W2mA9+n5ScEKyFaY5Jcx
5MQ8TPvLKM5c3KlfXzSXLHq10eDYf+EKhU3OZ776U8slfw+bwEz71YYqltq2qJ+/DeBbM4q1u92r
sTTM5XB0I5319VEVHu1VoE/2XJl/6mpNUh1o0Xbm397bWrQhbeD8fjxWngzZCO0LhiJxKZTL+tb5
7iRuDak1Cegms6wu9cOCTXvaZ5LCmTkmnpGHwrBggce/lCMvhPkPaqDQAZ8T+kgZYmdoI/q0J38B
tYTV0lINqwEHDXzR5EwLdtUdebogCaetxikf2rt74fmiaiTUjKVbGv2Gq95aV1HszRascGO1EoiW
u/ifmZ3Kn88whHIlwX4bxGapuGY0bPRxOpEei2uJ5k2i4uEplqUp16+eiIi7sVC2YfOgIFgW5PI3
pg8jQe8j2TR+mX2pQqE9/SPPShDgLH2C78mcLw7uFYYgCF3xgBPMZPBIc0B1xaRH/lZoEcXDSrQK
UU7wocVw6ytiRevAmBmoqtgCZWo2WwTcv+D0crM4fjVW1At4bHQuRCNSfcQYL7jhkxeAkDQKHDjG
z7sIGWFVH4KyC/r9PvsSKNoz/FjOogc3fLN1X0VBim4u9MR+kYUQKSIjKKHnyJFRMlCm077hvWSU
09/vOg+DQIuIn+Ibv1Kvmy+UwAUvO9IeiOHxZHWsDbDgJ+J6fm3PNPC5l9BIZsAyfxLNDZ+r0Drf
jrU6maxwqQGo0YiPGyofNv+raDEKQ8CP3kLlDAFhDwfKykSjWesg3baa2N10EFdgQugBVnXs2v9p
xBnnZAnl02Cdccb7r2IBbUi40OAh4YZl8BtRZPtfWD5tTfjr6o0vw/7DxiMmRQDkRus67q9F/5Z5
JOlem6z66qz5pfeULNmzTsZgX7ErPNuJQQpByqZzaLw8WR1hwf2pz8yRw49LSY87USTDHXf4NcmP
hnhB8WfL9lBZC77lhWTsA4Agi7W9d9kyaIiDIWLILzbJnHPPfqeTYxq28gXHOtE2lwoCRRYeMJot
h5ESD3veW76F1CEeM/Z0hHJMyJSgHPKnBJk3pdiq3JMNA4EjI4fGWBSxgepnmHPJyOcI0Y0qvnqK
ev9RwJ3ua0RtDlqJM5giDvJCCvBAfJl+wpU2k40z4L8dqiL7csNgg89NWahj3a4msaG86nUHvv6d
BQ7N7oXndCobueWPUT15nVppsabc5WBvESzSk99DRH+iN6d/Erb68fwirArFhWbzEiPK0ns6drDV
+/95XPeh7WhTOYqtwX1LRRBb7jJMa2ZkBfd7GeK4Y7CczGOyOMtb+Mwu8r5CmbF1u/fBZFeTJhm4
X4hg+8hyNp9+i4b1NwypjUoBMQPwjiPsdQ92uOc1Es5HkOuMa/58d1DvRbXOgJnQ31SuD5/z8OCc
8g9tXq4tT73zeiB5z0u0OaEzIlX4u/kMsd8W/+l2yfEt9jj2znLKhhYzGVEaaCheUr6U3GmU1+zZ
c4HYWPT90j2hItu6PG+uV8eTDVMSimWbeSHW+4Yok6GR2rpzlE3ckRcxlKcGl0M/vS3Iw5ffgoY/
CUqS/VoCKTjJDILFvmnZImm4A6Y2Itc+hXwzIN4fazElhNQYuppCtuR+O39DhiXPWw/nxKOwKDBQ
i1QRdliYXJREJigvfxQObyuRmoLsE61RGZ6zQ8JEZUAoDqgx8hWU/qlySkzFDyF6d/dpTfl4z7rN
3cTCfIWxwmhgZDysQQrEAghHqY0GyV+/nobd7hNZOlnd7Km/fQewhVz1juuItHL2JTf9cZJhpOHM
0zbbcBEdhN7s3VAPwSUzi1El2ep6EyrUXzjMi2WXqRmrdQSeDSdRBGFnTjEY0fAIo7OHVhinByud
6ZmBPRtaPTHZNykmvn3pUTXXkNn69Uhag0toyIR/Fxc1jGBEhruyfZR6ALA1XVbsA+p9U7XDZ6rJ
hJEN2KnJTsbNq4S/SeFG6RhuQQgXNJSPD+8jDWShoytIIevCsvZjYhCJB+LscusJMParW7tK6Fxz
QSzH/cqPEXJZ9/bDTccwfQ1dEpy2ZoPFY7t0EzdOu/NGRiQlGe5lsVyHL3igKWRbD/NykBRd6YsK
vU+yB78DHoYMF2GYSFUH+mR1Kq6KeptNhWuIlFEkE6jcJJZJ8eSrk0GrfgWyJFEdFCPOt50pXvX+
79KuDUesGa3CbTnRx07FZqYT8S2WZnX3FA33N5UJp9guvnQLIjSRtlht2IHF5aqGlauUpzYjh0jC
LjMiBMM6HJHSi0zVvauhOCJF445QbammN0cd3yjpDoRTqguVAcqsBtqZntZwFSXwYebZaMaINI7I
m+BWZnzjw1B+dREA9h3cuxJqacW5TFQcVTTQVfXnvVqnRITMty/h35de2bF1JcoteSA/CbbTvQ/5
hpWTrHJh4XipMW9w9qRRCnBJm93syswtqxl9mMBJZzAa2NOrMgjnSqe1PlUdn5WOPIU9R4tqxfmK
NDVUfaCDEvPNQ2AJuJutIoWewtCF+Nt4uXq+l5cfv4DxWYEHLkqPFv537vcYhsRfhHrCENckeqst
4c3kQwYKYIuGxJ76V3r6ag5borDYKi91zXMlTcZKqBt0rX3yEGaIBb87d+hN41LQzRrVMcQ6jPzw
Qn3xxehBJkH6Sf5Fd2eviS83Ld62SLrvRWsCqVDl6DWXNCS7GSfRLqjGRq4uV9a97DnjLBWUPa65
t0E6qZzdPkwADXe1shTlJt2Gn7rZQzUbOC7keJCGcmRIYbOYJHE1Ia16aaAQtCf7gfVBcHEjcPbR
7r7kIS+O1XiNoj//13morhcePESiFpF0+qWlXxFfKa/m3Y9/lMCOVm3sBQemx5CtKKrfLaIMTZBs
ppy6dSCS1BgZuDovrnzTMIEeIILGZxdSVwv6IipHQ0Co+wcywd+4I+agbgfFHaEe6LRU+wGNmZze
yfVg4h9QVZaJYVW5yt3Q1cZW9lqPjuEvgIfL4J6TGN9gVWWs3HOX6uFdMPsVJiHkRsgogtysKDGl
/Go9OsUsNu09iYUY52trRWa+zZP4AIFlEAFUMZi9x2P9VcGbIYpKSOD9/Ir/EY+bwmU/hI4EXIQ5
asVtozx6gW//XGqd49csZW/ouKPeHbhgYK1NiBXjhBSV8vzWkOuixNqCCv1k3PZk5y/mK1l+O7W9
lzljlqn5u+6iawpnkGNCJpalFTTqzG3AEXKiUo8734MwzIJHK+iwUrhqUuDOLgPx1Z2N+fu3xn7o
uJGrJ/XxFXJEy4rSl818xeLqnU8SAgE2BXJ3IuD6EC13pLMhuEYlqvYBkq3jEuQZvxrpC9phF2l6
6jhCk+8sF21YwHIxGk6jCtPO+I406ai3lCirQ424pYh63ciQ9PHv7mSphx0XMgZ24XtKglWy8YvN
XHmbprfgtzmlK+2iNhM0iMSCQjgbWbZd1NMgbjPGJBMigRCqaLkFssmMX0kOR7VTiYSUcjoMdVw1
D8qtEeaF5rVDIgUqsxaeDA53CWwMxSYOIB89o4sksmorkUBSgR6r5S6yX5rqlqaLLlajiTYNlnvV
E4n99+z0DAtXucj0sXhDZlXMJ1DSffF9nU/wVmjp/KgfTU9GmHY79xEW+pwssgBth1V70R1k4DlU
+bJDsWwdkW5hVnKT/J6orQOF9rsiSHK1aJKBOzfX/dHP4940b5rUn5bJWnygaxhGc6mYJf2qFK7k
HQRUrD8TcQGhihlRtolL2UXHemAifnTREJ3cKNT3x/VM/Hndrd7HQsYwpfewIRcLX+hzCW/pvjtC
zmssHWtGTXyy8bHYz0s6Y0OJ1GnbIMp+hQvm8nEZP6M/vL758TAFT0OLlWG3fopBmrIjfiZqnSa+
5xmB318jayWi3zy9xrDpslX8DiObFp4igzTmYYnxPcGsTNDkN584oC/JRX62ovSCCGT10ePrBeoH
RZL05kNJIZ45/a9THlgabKD9n0wgOSX/XSlX8sS+W34OrPgCfa0M4YKaw00/IzErXdteinjMO2jp
ElyjBkb79HbbFSu5R9wynkqnqhCnnsvp05eXgznzSIBeUZFBfL9sobka2iM/0BpIX3ADjx8K+N8o
31tLYUXV6DDUPj+m5wanNxkRzxYN/xpwJ4VEbc+/1wavzy7tJvXE8rlg7wohCQJKVML7bxYkIL6j
mDbxjmoXdkr3+pKD3MjNzFzLCeJrDK6dQZOL1pMki/PGgIAs12Qdne6CC/aopZHshGxKvB1PftiQ
MRf5YrXEv8nBg1fclU4dgb/rLEnqX9TWxLfpMjoO1uwm355uxovn7juarancJq5SSm26cq8H2PTK
rj6yZ2r9TOtNRYfP4ITXnzHGTT4y2OowELpv4JEwnS84dksYRwTDW1hnjCJ8jKUDHSztIrRAH09y
JEwXT5GN7dgfjYyUTwfMR/IMxLh8HN9/Jkmw5FUVfg4X0wmLQ3J9a3HfSfzBmlNZpg6Nfheyn4CM
bitaROig33ZgBGmiKAfX4avAhpnaF8NAjz0ldN6dorYNxjTQK5c3D6SAnq+DkgH/VDZ1YVL7G4m+
pW7evURVMvV/YXmkHDet37H4rvfq2LvIPaLfseVMNlL4bD42fwn5uE3LfwoVIgjfKSnuu5QbXygZ
AV2G9pYElFOcCo6xr+1JmboGHidnP95Qho3fjff2QdZcwbV5sQKXPF/GaaNdBn4xjn0df+rHux2B
4yZZx8gJYSWvuLE0ahJ43/9E5kybhCR9LHy+xQzZb3QY7D6DYg6zNGJLCVm2TSwiVGfG+q/BgitG
avyJXsvGBXyyuBoY7JG9Hu7tBNHRMuLeW/cunn67pGC6K/CFxWF2bCrnsQW5PJQ6cCE4r4/mua8J
tHIhfQXdMvsoWPKFxEE+SokGS1q950/RX8VXFXDHtRqwFJtD9dwx3j5aygnnP8iKhwNN70yMIP2X
fCnojJEu1gtjU4KZ0EdEuCU6rXyllbHeSIojlADeJZmhOnjCK8bROf9kfLP/qUHEscxPFKnUn4/h
HCC0d47AVxLqqX2lfX6Kx/IcyTUfmelBUjdROAWMYqD3FZ0AYPvNo48ofwAf5BITef9FDC0Q/STG
qjvrbVwRuRs40CUQa+0AZcNzM/oa2pBg5itm6gczzFpe4KeCQW4H6AZEJr7iaAhS4zOxvlS5Dk6g
b2BuybYhH60hVMJr9zvu13WlEaW4tvDY2h7wpLa64KtdDwThhK7Oz3EJ9/4ckFqKNZmoam/Td5w/
85yNJGDirRe9MZsaT/gBsCVTU5/njL0HrSlCkC5OpoQ6X3tHuctlnk4u1ouIZb0SMnXBdm++3WC2
kIWgAzXQYWA1TbDxAUo8NN+uQogtjVOA6egFOZXZTHyaItjE1XjMLqFmNOI0LzYcdARgnhRglFJW
MlTm4Y2TZtuZrFl/YTPRyJOLoKNMiuT8VaIO/3kX/3z/Q+qcNIuGRwQu+h2krBhi9elrsSOaH3a5
75qtdmrCjqjZMlSpwhN4TNbEk+/yzrLtW0DesQ1LRnq0dynrH2YADNqI2kEEPtyQLKCYAzHuWClb
EM2uFutfbnqoS7/1XTxrHr0y3T8k7khwGqHnd3jtTLQTYsL36693QoksZpPEP/gbqPGwJYksEsPx
mU9dQUWtRYA7O0oSjY5d1nNggfjKSiniDuITN8YPSDCy/XKBcFcTSDiMYPv5uMmto9GyH7B1vMRc
Rl+5ig+jFctR3mvQH3skEzZdhwGGJrro4TZKhoBrXAkMOXyFk3Pf8KBXxvWQX40j6aAiMCcIS/Mk
ukNYfEYeHaBbKcLCtOq1AUKmc3gfcm218feVaojfsXg5msQaZM7f54cismlJcCCbjqstbS3ZR9OP
Ufy0YhDw/m/DLGXyo/eHt3eBCaGvfCcW6aQ8cyr3cSa9D3IpCTWM1RVClVqEbsvyW/qJpOXvvmXT
mJ+2W68P10Rahe08fkAm2Xjjq+ib3HCQ+WX0NIbPYqlCt9JB1ETKIqKLs6GpW49Em4Y23iid4VE2
+OJKeB6rGMrOtGxc1tGbNa3zVwpHiE9egfk7heFrmc+HgbYduEjnG7gZakF1doESsI9yuuWzC6iZ
4WwgmM7il3OZzdCfW5lIpRi8NE1vDQaIoGcTPaNJAxWVt50y2VJwfU6R3B1SF4mmmapUbelXZz/E
PddkgaVQOGGGO0PjidKXJ4QZYK98BdCvdxz+ifa7K8t6sWfJAwPDTo3cT99FllmlrTWYRyDB85oX
AjpmFetr2X1pMKWbM1Q6a9NQ6TfwVhaxPsaeDxfTzIFCqkABPgghcB3Uv429QCvWu4Sw8su1fSBl
AdNW6y6/5l4QMrjfadUyTVPtMbsa3blZnHSWcmzKE3/pkJIWZLVCv/jtB6S5bnzwDFfmznOb4h2u
ib0WZrnvYpN9ZucTDkYASvTkpBvKiLIvc5VDt8m1VbkTjI6atCzfhHwqc7jgnMBOUPZ4eISbs6H/
Qnv6DqIiPmerW2U6s6RK9y7Y58rGyJNCr0lcSnt9VgAnXVlPHAVfxudtkUtTwNjyzvIh/rv15V4/
7RJ6eTtc/cmy5z5sHQsxt8A1SX9k8IFIEi/sYYDKbmB4lsDPRqdN97n7D5bL8GJkQbCoazgvL2PH
7/U+DOegwRwX+L7VGSI0Jd7G4CXngwju4ScEscRUpTlBqdH+8B7tJp2puIcjp7/eQy6Cx9sejPTQ
st+WjV5hy5Iu42nvykdRPXqEzf0PWMQFpTWPwVBgIBbZMmJE+G7q17jxd6JxroDXbZkbcmA0JHtM
78Jj7OYYDJtaagsBMEtn/Dz6egQo2toJ0vyVSFqSyWTOcdL1Qkn/gUI2lGum7NDQd2/F3VbeRAnv
Y/9O8h6RbELzqvLfJDsg8t+4JE206whi4bXwN50alixVkMGjra+4VsxgqTF+xsIJDIomxaNfwnnC
v6VsyhLxe6CTUW60xIGsLX+MPWhMmp0EtgdXyxPJo3qwA3OFCunv2dX99wqhlUKe+4EQ+FVBO2ji
TX7AClf/aXLooYe1nXQXwvmVIbpk5X/o6CoFzrGQBNZwQQLv+2G/ODu1R6UWpTqcqDkXiENwZfoB
w5/qucIbN+xGeCXOjvGu8lXc9SZWSn44JcOFwWNoi89AyjEPb6nWNNA5mvg8fMu6cPHSahwy+8le
V1Mvdg2RW7TZadciDeHvlDI7JelMZvnpS7dl9G9Vah4R2FOrbX7hMp91CbduGhQqHLTvHdmLr0A9
6KfjP9LXGGuVhvbWhkMTfKhYKm2JWXO/oOA7LeDHU7TmfD2xWhRx24qboIxRQUZv8R2RRuLOocZF
rYGZH0LXCBrAr5CBPtqOEBDWBSZVruia6OgUTlhMNPWosh0Zg3TCMPyIeNI1uiIQDzI1ic3TuAEy
Mk4zxy3HOXOr1xRmVdNNHQ2s5GX691Z5saGz3sAKww3EBKTJiE8FUzXDY2Ibn5WR0nKZp+aQlej9
uudYEnl0UJ2yM5yDtWcsUKLxSRJg2IWtJYZ12eXJdaewQMJ13KwgjZO6U4cr2AsnawGzlmqcDl+f
l1PG+RFImQ9afI3tOr7D6oBzYCUrrbO4EpRaziozZHpW5eozCcJxDq1rPIKer3CrFqjrhXn9825E
R/xyetxEOB0dhdNX0aaWj45iqIoVchaz/lcGh2yX5eCbY0nt7Lg9eAEJpmcKa0kyFQ7A7A2hprMB
kINIKefZmt1H4wo0Gi1g7fE/3ei/RATobkPK5hJZluyCqEustSjtwQ5dU1pC+qOrcyoRbY2A6xKM
sk42nBJVQI6ULoJ2cEQqIMo+nEfihvDwF6ukp6HAJ96z8khXlj206u+QSdPb7ui6J1m1iKdCoXHT
H+RBcUgNDtmrmvpxiDtiWgFNs8NUnKtkEWXaEXYknvPVsU7ctGgv7Fc2WrqPsAWto3ePVyMNuzE2
srE+/PxdpDY73ON6dPcu7ZGtwUx0FEX0aphRm8qfLLU2MUVlNmqrSFZYDA7MZTSUfUFF0062EDie
WQQ04VFIOnYA9kRzJhtfTDZVFdMhohZj7l/+XGeKCHRea2OKEdjiWcR0kZtrsyBn8jemrFytOwFG
sxIRl3RA4K6aV1skQqSIGZSh8CYUorvXB72QE3tKSdU2h63Kv4555nGlu5HPR5K0Uky3QxpnAStK
nMvHkIRmJUJ1eAD2r+h//RItWDJPy/lMTfexTJrgcMU09DQvxW9ErOUa0JW6DwYNrcrrSFaCMvcY
oN7Rb3H+q67Brxq+hw0Ow0aldzAQOZYY27s82fKVx/CujHmSH0oLuHWnmOBsfuBhFMs65vt4uzOH
Wx0L90YTNfzOiCaez7XtA+u11SygtnA5RHyLLIMf+16ZkM61yDF3MY3zHygPQXeQjmtUoOqOKVAp
kV1KvheHM0FM2r461A8BzHwBdinsduLqAX2u718jXx+cEiGVera+xStUR0hHIvx2TjPa+30ckd/K
5nzp6T4ag2C2BcPigS5Bl9Py9TPHt3lJ+/x/cGLsLPaVFoxqxQwX/QoVyNlf4c2OcypOiNUYs54G
1bJKQHOYXuj5aqlt+wDaHYy1hRLydXQzW97+5RZGreSn7RiCHcneU7SlTqXLw/u6BLw8eBguKLv0
JbwbT/aVpNel9CZgJPBtD6d4uiCET1Rn5IPm2zwYwynR0i8hBKBHHuRquIIGeiL4nyDwPehruGGI
Z+t0a1aeNL8zJC/DBFlIK/61YiH9YB9njukswXVWS4vHnRBnszsWm/yAs09e+jIg9KE6naccRWIQ
d5PXom2ODhtDUxX+gt+aGGjZh7+Lh07Si13c19gTTst9uCu+Szh9i9/ClYN3P775THrZVLKxEVDk
oGVcePShwS0uEakr78bE74azU9JUpWIa/Yd1Zntvyj4aC45mLL3z56b7SvLxlB05crMe1uYUG2+b
A0qQ1NP/4nEaNs1ELRTVEicoGRw39ifsbVfgUp+zLt/YxGqS18LfWPI9bxbmH3e5StIRQaiQ3RO/
LBJtUi480HxoV22+ZeRiMjz7viHMC2cQ0bKUoaT/7UStTpzU7/SomakvoF0zUyRjlPagk78nFssn
ZdbMah7xze8r/YY/XxEaJL0SVYkhOq7EjBG8eQ61Q1RHepKY42sEYihisCfhabn98fm2mUjP2Ahj
d6XkVz2YcAgldq+gsavoubHBPw+4h7YGnJrw0RecGZZMDtLso6HPeqB+lGW91STFVOrvAMoVxqa3
gejpzqCFzeCgkeJVTXXkwaFaC/JF/s4toMOt5zV4qnCuHyeHAp8RD9/VoxJ9ljgDfc0yoHprYCDK
gYKQXRGQqRbb+9uBW1GarXIr+eVgcQYKYhHvGEoXQAUoC/9chazWhB3bGNGifD3DmyAj/6VAwdxv
vecJ8QyMY3w1aPP4pMEwRqOdWjAsvTs64ilLXGEB2tlGVJsacuRORweMy4fqKHl53ftMpLwY90+6
FqiASEUnY7bPz1ff6bzWbg28f6+hKwQPhqu3TDcxItrAFExg1cnrxxViMDA7WeCckHk8h2ZudnCp
jppREk1TkbGwh2MZOqyPx/sUwjJXEt4meTF08hcFs8e84in0m86JbYuNYFKCbNFiiin2nv6tFB9X
mv334IOkjK1PdnKH0150PgW3AweWnj9EXKqooUHzzznfgJ0HZfsk0vaRzoi7uYmv32uedZzt8utF
5zDw8R1LJHL1giKxt20EmJebC3t/Uu3Q7hzfeDVrPaHq3Ve4yqlppOCuGquBVIsZDEzWQtEokkMg
ThvGBAQ93ynz+xMSsjJsB9ry7lBoWnmwrTeYUt9sJz4eOn9bG4xF1JaGC3Hu+TfAthpE1VfX0Mnu
QW5gWSU9z8oF7KSLU41p9cVw49BMecFQSYziA4HiePypcID/oOTwGdQ9I10g/KuiMMKKF1pdU71d
gX2+fZVmVtSipEXD7WWn/OPN7AGpxelREdCaNqArtSQg1q+j4wYv9f1Us9kTiKlw8DllaaSNny2l
d9ihIxY0lmMTY+HsQcM/SphLhYyqQ0Tx2AQDFOETvwMj7Q9rHcylH59poYVtreeLMN/r22VeY3T0
TI1FzV4Lkm/7UW9T63nuTK8DyBV+a4VLtNcdsn8CgJPqShXGTKFgDFqXfFL3m1+IYIQTRZmHKEW4
SLPl/v7Mb5GUwhuvBtxgbTg6jRvtZI9ZsgywGNTqvGS6xykV4YDfhZoL+ATPQ+hoaXDinUjECojS
qwEEfDJsr9luwYyrtcrRlpdZ81HkcWfRR98otQ0nlxGfEWPLLPhVL1UGEawJ+lXLNq/oiTF1P2Yd
+PXVEALMP3eZFFKrz0Q+oT/XcktEVNXSz+pCoU7PvCk6HyLlNiRxl2Uj/BqC6RE8Odq0F7blit3p
5Bb4Vi5MvZAAgue82hr+TuF1oL0NUvCaPYDx5r1ONTbo0tFdgdyV1MnL+5NRfr+wth1MQY9zsntm
PYALwOwZXawYunc4QAMgXlOLdQY4DPM8HbSSnAWwQ1u/O6+ys/iiq1sD4gZoMeq6/yqwcLtu2sJP
juC73GEXJSU8nvafPS15diGNtFSKbZ73KyMn65w9qQF3ZgHWnDoWcS5TnOKeGRw0toFba8oXsZ9V
CE6efLsuFkTiBHaIDlMwoh6fdl4Z3XWc6qCAbcdNHBgJ6D9DF8psLDXA35a671+szVEfjOJOsRu8
6oORa+JELL5PT60v4/snFQNz7DVJVXeUw2B1yKTU6AwHyQM38/9SJMU7iSxWN5Y+9S242h/c+f+p
FpXPdjoyX8D5KxUqrl2lEDcErc+oBO4pFAOZEwV4mUR36BEclBnKKNVmqx18qWxKqaAiN5msWPfJ
BVI7Xo5Lk/90mCbph6/GpvjVukFJ52LpAD65zraskGhw4EN20x81jFVUZoWPHyPKPMilvfEGIvi4
ZDu/tNkW7X2M0IHcD41H2dEBdi7sQZejxV8WZx4iKRjv/Jn5c+ios1zUuCNuFmCYcoS6HAwCcRlD
4+eL26OHhROGnRAK+t1FGSdNvZmc1eupMSmmDKjvBeULUl2D2C2tCvDMSrleZM0LCWA+cNQ5jsSw
Lw5CUdeGYCYzCQp/Wh8QDooXN30zfR6f8qXPZBpJMo/xYG55GxEwad1LiOrvjIzpkFMUIYHTc6uw
50+SFdHaUUtcqR4dIsecSZ+J2wTNaaXAbCWK+5mJW9mjjbxAeiBz8UU7YKlhnMhu3vmC8RB77WO/
DcN+flDvB3eEQTAsLnWBpJwBU5SEbq5v5Ugk5cdQ2erzK5p6ICxhmTklYNUU7NuJ0E9yE5HzNxT2
7b2rDCaeCQnUsU5Tw0L1nLSHvqQXHopiDmB0oM1xyZn/gPxEfE/6eM0cIMDQiZPJlv+ijOWtBtQC
fkiXpY7iefDhcfGhaYMZ5XP5WfOtdkqxttA/SjgK450SJm/1sjdKtLrX8HmJXZbacgaxpWatI1Vq
8Skomn7V2x/5Gg9/RuidYCfl72ivtuyslj4W1ib0lUa9ODN2/8+KeqRjX6mmokhxzApxyoeG25e8
srGnbIiyax+ot3mynF4ClpD4NgiSIumsxp6FDQ05A9duT7DYi33znnJ1BgMnb7o3CD1SWSYihypJ
VoAMjftAo+ge8+QanMUrmx1jlPbPvAjeNusYUB4Myi4GVeopSPpNvu/GhmFYnZpQta7RvvL4gOMY
O2L00z2/GHtoORvP6p8KN6CNFcFAbLc+Qf6542FSUdGExtKkx8AbVGSO5YFL/9/ILx1g2BNHY603
VKwlQw6FoEKyQqQGvzptNZUzZa0Rp9AC8puPYbHF9VEad+E7TxzQ9mGXsKMGYySMiV6vl2NI6JGo
/IVlaWUkemU7iHVW0nVkkBWEuL6tZI56zjlh8W5D1tReEzWJB/W1VeTVdVF8sKt4t1jntCXsxH+3
3qnjsMXJe7LVqIpXJA/KN5oNxToPNVmXa9Wr0FHNrrlnaaj6Du7iU1vBBiae0JpuEx8Ar46J0LbZ
dMyyfq6lj4/NNkQl2PmSsHpvSMrujWv0PqSVFThWPMVVXqO21M10J/kYjZTzYGn2J7fuHQfmq28z
cwoXtVJViNsQ6rdx/Cbh4nzQz1tfK3hW4havMDTq+1/qf+OKZ5QAcfMc6Vkc/6Cau+bEXW+fucOV
ktR8z3Vxc/oI8lTM/vTQrFa3HV1wQTBMI21U7KWjsSbULyphCoim4J3U0pPq+aRaSTLjjRdxDOiA
D8acvTEvcFwOnoQPTYI4FAGKaeCOmZKuSYYZo+lTyeHSw19aCqfrzHxncZZ68fa27nlbLAm4zm2h
UwWUwOCmhstNEYPvaWs5cFos7L4bdZp2heZkcT1QUoRXYgCNcogO40I/5ZM1048x6aIXB7ODOKoe
/+VjyT38pd+EN3byt4SMp4H7Z3HgxfMrjJ4RJsRPcyJA7xpb54yExxPgVHDId03dpNVXMTkDGIU2
OW6YA9RhoI6nSlhnrRaBf9ZsAD9m+DetMFft/ZZCD7ImlML8YyW/rM7wZuNVmA5ozTIVHGeLfHss
agEM0y266T4sj4ol3js8Xj8MpVrLFWpIPclKWYOTmEgMEBVfkZTGSgXemCv7BSvxfL4TnDSAtD1S
JxB6Di5hZ/UkvrvlMDt8xHLKS4NzzHmmA4nlG2MKf9Un9xdzSILDFzt4m3uJmj+kJR3GaBt/JoZG
Ok4n2IEEWtDFShiM064cjjWRIc6ADz9poxDVuVJjuMxBzIc2oOvLWs4L2hRRh1uIQME70uWQCb6t
lfoyZu5V8U/eE/INIpKUXUXSvPg5zBbgU3kCQoTrmvGnsvVo6lV2qsqZ/JXZL9Rz33kgrhmzI+Rt
SstoQ1EgUpOMl3ZbOLzXu6UGkRI38nOaH7R7XwgczdeJ7lf2ExNDW6yp+Qa8oUmk+VZ9XALnImVA
lbwTb1I7xWuL/fsw0X49gg2p3477IT4ks1q6SjFUBKHGJSiHlec2F+8mYlFOZ3Nj+B2AX5ysEj/C
lKa3jttpABRYdUkgXTyXB7Hw1EpbTSTrVc0epmOIT8s9AARwTn5YOgST7BqnOSL7IlGLD9T9PiLR
yXu6SmXv2nuOQ7DEW8ce6yijSJmi2DokIzVbGeIzrSc0yALNpXtXLqWU6Bwr/2rxlL3gbYAFEVwY
QTIzNtC2+NzcmZUPD9mquxkpLs+i5u11Dsv4RZ2GiUn1VCL8vZtTWwerHH1sQDS1VWVCMO7ehn+I
dRCOtvlkbS2Mb+HGfE4rD0RVqYhvrj23O0q5frBAf+Yj/k+DgqS+N+yUQ34jtsJxbkbjnDb7vRKx
tGZHhtzPPjbUq8NgHBlI56kUMeeoaj08pUCZmM5JhzBOYcB6ZNZRtTLCxpKZduxouTzbpXwtQYAK
MsdKjaXdskq29mEcQlrQJPlwbN9t+zIQigS2xAygpqRxqTeFvSE6PGgZACBblXCKdEBKMjjS/1df
SlKKWY/5YvpWG9r24IlkVh7q/23d0uabZR8UFCbN8p/HFKlRPnEo5FHtEdp+purw56X2EQVz6Nax
3rM8IhTIDWSy6pDFKTJT6h2JtKx2NstoEKxQp1LQU40zx2b35XaqpVxVsLd3SCuDJ5b5TRQaPw9S
kTYa/BW2oz0WzkvJIc0ASef7cD3YToRG2nWdrR8sAEQyMGk4JatNy9RQRFc69GVn2bHBtFdXf2U6
vNvTiuog3z7sCF9RSRXTiK+tMJuIGha9HImnBAOMAuoHudXVbrpVxDzKTFMsvf8oynWbDsYG+WfV
Vrs1hgSuA48B4I2jEq8fsbIIsmIb/paXL5K54ef9mupXIYMRfJ1APtdW7r4b9VsRHbPB8qWdr9+J
uoTN75stmAIJzpQT5plA7FciC+Fu9X2nitQ8hF3xEoplvTN7gR8qSR2oEjXza5MyeFhNmxjMpvw8
PuWwJo6GbXuW774vYrrdGRqsV48ti5Wpl6JYIDkn8/GMyLsi+RcLj3vtJJOoJoUgYqQos/EeNNAC
VhZlY0gjzgegMkOpp3I03AFWn9mwYeT8btTzDWRWoB1xMFeAupjV4ZIofZ/BcTWH+u4Dv+IoqjN4
sbJiHPaxNCvUCEzAAOrokSAQ2ZWFXVcNh1padLsT2tfJ83rD6JR3Wx6FWKpHGxbiwCoGtrDXdu9x
FhV4+RLGKGCeat5sXG/CPE3gWaUinwi3RabNQjLM6Kq7gQK4TC6eQmrHhytzJzBnSXHacRRe0wig
s0Pefa2VZ/s3cxLo+BCJCr5AzodevIFmiUiQgfZocQFyHWOqZqGRCRkueFrpOs5Ou2Yi1axNAB0U
UBmOmxxIli3SCzUxtkwUAINU4vNhbN4pyRtDatxM15h3+ZDTlM9BIptRSUufKlGjNPRy8+77Bmti
Lf77bDoCdFvgK8+sBPs+j9nG4A+H9RFSQqU1Sx81sLganpB73/Bu+NrV+YKjG8rDSzqRa9tnMM/j
XJ2J/Z201MMH7PtJqKtAEMDgs060SZWlLFUrlYQuyjKmotlBRZS5jIHRJ8P6zVbL7ZEr6+X9Z4th
DlJN3k/54xTzxI49Fh3O+Lyu+i2QuaBuQuEZ+yil/W/+29LQK+bkTgy6s+Y93soRSYmSnNuVNIBB
vsGI/MkO1EXOYs15Xi2DyzAaWjGjg17VJIEXJ3BQmc+uNQPzxrq3X9bCHo13cz8LwF6xqEU++/iW
q22NFIBHKGWTr5+ITJXHlHUJQQEZ/mZRq1yyHA4KETR81Kj81zL2cDpCwtQU/pQM+OOho/AaLVq3
j4EHhDuMnLlV9A1k+tosQwx62BYWc+3Tc282aFowY3ERiHdZ8ArBa2KxgQPVvJJ2BU7ME1A7oNVs
IbGZItJ1SV1HHZCR/wgYzPENkAY7rS9dG5Z6pY/S46sAebq1+C/dQqrFZcCljwjAxBWFhhasEwdC
i1MNdV5lx0JiSbtBs17+mPdJn4MdLgdHt/wJUiIgYWJP8bhhxZOqlI5U+j3boUtWkYgrsF8KQ/af
f/Hwq0Gk++gjWQwd5H0880BEIBkHZLO6gC4K9BoW82NlrwRJtWAqfrKSsDk0jSyPFqxjKdSTUalK
kBBW0X1sZaA4pexWAmYgSUYHPEg7cBgvjo747coyI2IsMtmExrML2b5mAkthNDBM3ocLWpam8nn9
C6FrpOKNkGRqqt4PkcNdO7CtUl8M84spJv58zIorII+AJBgT6cByI8qoiCaFyipZd7KV25xXYbUL
pU6L34yr2jSKYpu3sPuiNe0VDIZJJLAfe6bjZzRPFIJY06e8A2ewBsGGR8LuzqhCDglQtiscxatH
dhOKPTiuLtrZU4J2Lltmk94G+tuWw8Fx3Bi4EbhRo9cPAcOg6CZbA4I0avEhyejiAvutCpLq42ky
8gjRLwy48NfVyvizrNvgOEsQRvWpncwhIEGxRAM4bfRMUX6d6I40TM7Y96UPGooaq4VW0YFy+OTm
dHQbWz5I3zzRBLPVIgr8LIE/Oxsp78/GO3KbpOW4/834tlknxeXM4hbOxWGSkfjpZsRBIGh7OxqS
jQSFSj0Z/eh70iv3OFF3Rya7R01sbYCda4LeAFBn9y5vFFltMbyJKj5++uOh276TG6Qgc0ZEpEhK
RndCw/e9y2oU7DUDyALuBB9Y8qmR5L1j29BOeGCcKbGE5qKzsc7nm9sosALmze8SFRq/ByCpql04
ytrYcs7+TkqCihyjt0QpUc4imiSrI0YdxPExeRyCqTZN4MVyZCWcUWT2VQ6R1k10SknxuNJMjyil
0ffY/csnl8xNZ624QgVDKylkVdRwHHXWe6VlLwX0OO3z4p/kMcPHrb6AtF2ieFjoldvBHAhz0PAa
HY7ysAMs2cAFRLjvfYPtmLEKqm0ZxmvBQ90253xhr82Lo+8e7JHHdGAnvaK8hemSFoFh9ere1LfC
ALrbDSAwp4F/grNBfQfqrmP5qY3NlN4dLa3dyYwlkq5n9KJh2iEp14BhpdBzBe2ZzT2FcSQQ7pXZ
Psn9S7SCNTUQCiFXi1q9IgpnWr5a2YIAlRMgOiK/mtUWcxMHlii8AmDiX70NO2oSVMX8Kom0Hhhg
tA2ei3lc8q9oEM4aWXs4QgNulDloG1+4CIBzJFZqqFZq2TnpS0bxDBEimOZQegNRcGUwm0wVAFoy
jZkizSFocvJUVcxCtdDghRgiJn0OuQ4dyqarEFGwjHJvb4C76L1R7JZExLMlnSaSIUDfJI56lLcc
1BMQ/BwNXHhunLRSK0hXGIRPZjIWOVrlKE7Ee2KMiabte334IqqBIr4TiE+rklPUK/PdpGkqIhAI
VxNDBSORGQbXwVDRkIgpl8CjMFSs/jUpbRvhiFXhqV/L0V3EtNE9S9W6QUb9yOphxmHEIAT85JgD
fcnKC8R+tt+kuxOfPfF6RyTDjIH3Ig/PuWa2s4KFV8ovzTpg0ytBA1dpZ/a+MMvd9RRsCEI2Y9IW
ywdmshkxw3G/r9MdQ5PbWIRbMPKQdD3dN+Yjt2F0EOwXitFF68JlBtfhLIV1f9Q144qy9vc9fG5Y
LOfP7EbYoc3R1QHOGv8zlTHYPmh6WjTHNfrHQk6rU54+ixv8Qyy8rMPFEP1tveKF+wFOlGCuPE4N
vxysP4KVuV/w04G5zscK9raGEg3OIp/RklfzRWxdjFzBCtfJSFZT+Luh9mIeiTwxwDimAVFNmYOT
oWi9JBGDE3/zkB20fEDVLO8Ji47D8lQvZZuk0b/dtoOI2Ls/54FKm604cVD0NuzJp2B5GLWHWRth
e56wrO3UoXGbb0VJsQx6v1c8x/qId9SGqjJcMaYL9F9FeY+Ndr9vEhCArmMXAem1ab2UbuwCGh5O
5KUPByC7iMfipV2PuVteKR8sOu9skPMyr7FGzvdNVJoOB+yuhcbQz83VH7r9E0qCpv/oL1glJdSZ
8SnfIyCY/+5F00C+SRnhTzWkHtxX5fl64T0LDVE6B0BBDhskApruAyb8jvceYElJ2nWcvelV7HIx
ZZFfDg8EtIzfUAC1YzzTdyDDxrQXWgwl256jcN0bpHWWu15YmWBv03vDEBlJYi9ag8XG2TMM6Uv8
UFMd1PXr4Wzl+oCCO5tmbyCZONf8Lok+ml4mOAkJp7UhZHts+SjuvBupQoQwHekTuGLeYOYs3MdY
bT7/bLZGyK7mDhZSxcY4KedKZaY3yI3Eatmn479FonIS4stVo1kaojHdwAfHNPgQ64ptzMp8AU0A
duerqGchBH0dLtRvCdjpmUdyUUECS4NFx95wiqWRnjhSqcblPFWqLMKOGCdRlxe2LfVDU07tybjV
lFAzfCcX2z8aZpSlZ/mlhX8beWCvdgOt9oZsYLrXtesEpFpgX0Maf8J4HRcOd2Nzm8yIRMHh0NcW
FlGJUkck4PQ6n1ohsB6oUnviFRMAmykmM1PTR3ZGn/y8mgZgJtPzxzZcfaGaYx70Uc642xZ4P7IL
SkkoIfLhiWImfUTOrfp/fecWqPD7+QeSIxZtAaIVNMICeB6FySPZUG910WXkzLvNF/xDtaFl0Qyh
rnJVe1K/ELlM//HDArsrnpW3rnDWnCzUTHxiI5s1DJH7k2AN5aJrTT+LxSf3X7d8fl307MAxs6/U
tHyeN7HSA1eWyhSGdbEfqcgeT5zzhsilTfuc4ZvqxfC1z8jIWVZ7Q9+mfAu3j0tHPYw4Qsb2+uZl
bvZ6GXeyOdQQDKgAJa+F8xuPuia7xwL3TPbp9TbeON5mjbo2t46gVwOZwzEanVzO1HeQsBWBBL+M
0Wn9v1oG5+L3Tg0ux1uiEPhlIN/iK2ZcoduKuMvIqnlRV4WsJRq4Y0lN2d8/ycCm1PXHMSbOG5tN
qscaXpBNWyW6JbzwqR3+tPk5Th+JzR3kvAKv80RJB1qSkzs5up5ZzSwFwaJnJ9U2RWrn/8FnfSOF
XMa4ANKKqHWkl+k9/XH7w/A699bsu9L9I782Awy+tFq3V1WtLTvMxC7z9cKtImu1urLVa+9PAUG2
aHZ/qBIT4YqxuRoMEVIi0zq3EJ1XLxmN2uCePogEgNbq0ULuQHO4+i5wJJWaCejnOmui2yp08AzB
iCyUwRrG6IKmthBkwQLOnMWftLA0PR1ulknW881xqMmqqwJbEIXwBRgucWcRm2WtPsWjWPPBQOPi
HgMGwKo9B/82JnH6PtBwE6N2w+TgNhaxLZ2e8wgfWUkOz9kUb9WW0YFrRfIkaxgDbZ45biTX+hoK
dYUwPESlkTuU9ZUK7UcvNTlw1NZJuRr0CYOpsZiCAKP4PFNFXx4PgkdBTj8BltiKzpN2wHPHxRME
ovqb/Ac556HA4hbLfqYiwMdFQAq83eUrj3ztdCdO200W1KzHTTuymRF/Ia64C3jPzn35jx06f5uJ
gJ7qzoW5RI9pP6vxtjK+MDUjEX7YzkvMvBD2W4V2YDhe6TEFIE1EURBar2ggqC1KN9jS4kNopxsH
r4RUZzHwi2r5J4vkfkA8bHmTZeVqsu4JASujgQSvPf9JVf6Dku2m4vJLp3S3rFNfmNi7QWu25zf3
WChFgLNv8aSRTMPqFMqwwunMdKwKllunmODazYns7xyvcdwd/fMfCPzO5l0B4tKe4nRuEaq0b1KZ
iHObxWO0xYHPeum6NhXL8mkTpSUpQZh8R2kHniuHBiu7NkQipUU0OZkBOZQRj00IOCP/FxjBZ4l7
heS6wE3g8vVzTMBrq/wMwImBLKZSp98fEu2SOk13JMQjCL1AZTGsvvhuKlZKKAa46rldx3QiaJzP
Du4ZPwOlc5FKgqBHqF4apjOa3xJha7jK0eM5aC2M6ugcGliYHtVk/Ujb72G4sK9cj7NqgetsLNqJ
amzsOomYdtM4LyC/78YyhCgss1cs8I2Z/JqNKy/+kOfBhkBngXyZ/hPqt6GzXngbImGjdgZULrMu
tFzH3kKMWllnSd1dROj60KWIJoh0sAeYVyHtgp+IU3sKA7pKrykq0hbfIv/jJ8IWY2LCi27p0h2M
bkFZfCSlyNXRYwNIF37/FEBgRs4vx9VcUlHXP0sQN6rww0cQO7Y/e7x4+PQMfUIP6f3nG5tcqewM
rGR2SrjtFeUL8+2ShuWDNq6FCf4fCX6qqhdUsWAx21NiUzs3RPdnxb6dFxLFOxxOqrn/cIAHO/J+
wEn2FMj4wWOwgk3y9pHYk/KhVAd92tQbg4csp68GykZtlSxIKRJQILK3gEcXReWj/yM0MmSJbkc2
/pP5aiQ/4pHIsHzMs8dIrD8pKNzdgjo5er+2vXZZpHTCdyDIgMNysi/vLpSQ/qx1APZ044TWGWcM
6JvynhQevirAZ+vC6PcBFysrC/JmXd78jaiphkuy1DgBtcCqzJf7qs37FKmOZRJY/2DOKB1yvhb1
191F2Ev/uE98tGqtLp8+SeqAVMb6OXvgQmjRIYKUxBDJ7tY3RVDopNXRwqWShBEHVLrOFMBFHm7w
F36A85ZOy/e5kgYgEYMYU7G5+MHPTcX/zoXk+TOQdfdxvVor6GBOle2CaFBw4D6c/5G3DxqVwqHi
P77qDEPnB7ezEuiZk8/5O//7YXwN+1a/xhpi1z+6UvMuIAAbvmAWv1UbWvLLcQ+EfWMMW+TA2IFD
XQZpe070ywzQloyadScSIcppIfBMRxl1aouD5bpiyoz4XaiNWmjffiuju3RQcj6ZnoGqV3kFkbak
5m4sPXVyDeU4LxSc85iNaMNOUMlKjNJA+61gdv+Xw+4aYJWDUgQh9F94gRyEpQmY4Qv4iKcYhhJ4
ufUfpBq+Ii8IgsHaiD33MJAmKIJs0QMmxlZJUWwZf5XX1ebGQgPevEsbvYdy8aH33yuk2zsqWgip
K5fTe2nG3V7XMziX+zo3Ymdsqr0jWwsqzRYAgM7EyOhUFF4vwVtrne7E2EUftjpwf92v0ZTshbmq
W56PJy6KVlFppWTEzc5qH+gWNAIr/r1lkyRRzcv4of+V0I0wQQXu4+t+VPm4gGK0GruE5Hanvxkz
V1Hgr5+2V6ZYX5VoPQjb+pblru2k82j6Kk4vVHI8EjEeaF65JpCW1R7lqQiVHU0wE8cbJPs7IzD4
/KAJatpVUbOc/ic2wzJ3BffHEzAaJ9A8Vi5vD0q4tups/ZLZ9r1bG0K0MWO+iEUcSsgWqmOITYV6
eJaZr/hDlgR2xfKUrgQHKRanjd6HZL6YCUmF7Qd0EPOX7yLriCytlf4jsu6ez1A06wHVz0jTOZbh
5oMD5vVrOQX+3pB2NfCznbzL80kDxjRC/wfC1msvPY9xmUzY9WoTue0y/JTCp9VG4BLKiV5H2/Yn
CQ8+Z1ZFvdidKIA3Rchw77UZO4Mouz4+D7d6BR1aEMqq8zRpx2v6LdN1HM+06TMQgz+5nwW07NlD
+F3NTmSy4tlPU7jDWeed7PJ40JMRDXWn6Z70e10WT8qZNK2FlrU7kRUDMOgYt5iyIyk1+uhV4qCd
a17enaD2f6NLWjbMl26CyOEMKS+gnNN3QUKFxMqYvwy/Bq5mEQkwsMkqnwGf5DYR8iz35cxVCv+e
8x1iguIbV3bJ8X8Oial0LqtDtUO53rxmSMMG8mHqIHCyOxMn+neBKLvMzNhQyVHcs4Pj7D90ddoU
6TX8/C6r2JslCwRFgnm5sqzyb2H0jzTS7zBYe5DvOGs1Ng4jxvCZOiXlADJXfq0nu4qvF/NJD7UO
ZC+uIAqzFSwWHDyWpZ+n6ovgOxm83QQa8UwQQKty5VnjkcdPg/HvCsk344t1VLxP8nwWU52GEghW
NckWVT1M8On3g9LTXYswiYSkE1mu6+EPOncbawK8j/cfrWSRgBTRvf69DNEXoZv9X8ulZio60nFq
mtqRmYnpGBXGy9gA7ELsXXZATCA8gU/jCw3OHjeY3JfrFq2MifuQQ2rGkBgHLMSM2GH9WVXC+voT
L6KVXmCtXv338f05OCdBB8jGa3tmfZnc5hwDPuKHLgEC+lSUTam0XQW9gG7faq5dzWT8U7ZzVvTq
1Kns5NZULyNqU2a1DfUOFZHLdSYPNNmmK+jek5JkktBUv6qvbzPYfun7jgMTL2vWXyJypt+wTAKB
8WkleF77jIUvqU4CdBFZRnJKt78tbDLurdLR0xz3c8+y4Q6FnCeGZzQkbhMei0dCoHa+c1+qF4uz
BCyc8WmHwV3cXCddx0J7ABgPaXIsb+pgixi9M1bSTv0PKk7Z62W7Ou5F0PxM+AR27t/l67jFFu8t
ZK08TXWRNh6BdcJ+nPtMmGMDm5iYM7+0uT2Yeu67AC+LQGc+HHXqXNWxLbkNid66yYytyqo7Yrsf
HHbZ7K6S9OOHKfMajM4s4d65Yd0oamO7N3rYWHbh/oLxLr8UitVTInoZcjJFoG2Pnc0sjUJbY+lF
Gkcsl6QJp4L3IEt12VIOrTMF8H190p+4n7Zp3xRfoNe8wDoUDzde5ErYNlbrfZDRnfoIsBtEgZjA
T4OTy2XiHb3u6ZPLL79uEZLT00b+hniyYxw9FW9JFV57ZJiAeL4C0mSDBQh/gDJ/y8bzzosZ8VAr
VLNPEPuVjvDWYwv0cU5R+rGXZaY1NO8yC1TySePuNroxpQcfJnFjk5/q1ZW05sp9eI0y93EUGN15
xw5ofKTF2hKw/A6kGB2y3K0qsfGDe0GpnsAioX1hV7uwMq1e6YhNHnLXgXH1X2sju+IvjXKBljCh
VeUoU4l4KBQ33sd00KHp5FuQqXbgteo6jO8uGFbHCSo2HMYZc4fFAaEBrWVdaJ19UDmQOvXlUqwR
n0p/spTYZxFL9FgYulfuRgDBmPeEdXL2YzoeZdoLvc5eD/NMeyS94VX9LvdMkCEM7XVBhh1Ri+Bs
61BimvBjpeqn+2CHzAYUggvYg3IMHKv9z9Enoahdz3n8hf71V6TnmTaVTKaQa9FhNMZOaRORVqju
H1oYO4g9Kpbss5ZnFeu3ytu2n73Z9O57kJ+shic6SVVwJIFS+AR7yYIaDQhlqymvipr8xTGUba7s
Uxdw2FWszGY95Y/+QXG8Tk7Qlwd/ZLP04QkvQf36x6vLf6Um0QrtMh89fJHrlcteSitFPoLIgpU/
d84w2+/2TK6tm+RXsq5GwlxFQCMlBxQzSGpGLR6UqCCGKBeGUK5OGpz8guudxZai7aHoM52m9Q0T
ZrCcbqqIsPGhaxT0Hmjec05MPuc7+BLX34b3TGlpLZe492b6Gb+9LU0/LHvLMO0NLPaTcw0k4Jbt
Du5fzM6lMNAyoB4K5gtLAGha3B4GAHIg+BAAP/okobFp29JfnFFgPESqNdaDXFaIouaDx41fjPcv
0v2uC09FcAYKm6wlsaUciMPKFBdtEZLKWaGludUGXxJlEe1qj9sjiLkRa+VB59bDxlwaUUhbiVJA
ykWJmzTDvJWPTFPXqBc+1D5FwOdMxUj+35rgKF2deLztk4TBKgwRAnc6GickhGL/yEo1Bxs2IJd8
PCDjSjB98sUwhm0bxkvFVlVTPEmHLKHf0s8Oyq0vHHjaIGarvjjCqKDbdpV9jiLWQRZslfEVQTj3
VxrEwUogrzEjlprnj3OymS92yi6UQ/nC9jSmivR/pXdTYML71itCaOfKypg7p/miiW9/+DFMYlNN
JaHtZV0EQrjmKN/gMHhkEq11/DOg/aUuiQW40iGt8Vo1bjJeCV1GW57ToSS00X1GAwapP3mqSs5b
txHAnwQpFQMlUG0j1felUP3C2eg8cOaeDQXMvB0XJx3YEsfFSQ/NbEVuilPa2HDOLbWKks4zkgzP
g1/Ad1PsLyG6K9ZBvNw2nbvtQR+cLxr3piHXE8xI+yk+LzXF0kg46NKKuDS2+OR1gTloAPhX07pe
EtIFNIBF8bQRHMNpck0TDWoSv5UFC//dfa1FFkPJoQQRhCWh2Vz9KRAU44rONfMga9es+R80ROJy
traxE7CAaK1HnYeX1V6s2vncOuAaQNGh5ZNb1uKGxiwR1NhxZpdL3WCZoeoi2PnzvWTJ2vIJG09C
0ij2SvXLJe038Bdcb0+3ADFrgq9qVvGL53eUW+0JF+zc1XlyvUY76nkCUlrXr00ItNFmpw6pYP6V
PMGfAlvOINo+2Yyd1g24CS6yyJfiG609rOgyJ+2ZdZFLgYnCytzFKOq9J7hS2FxTsqzkaFUBQaYw
1KuZyY99ffgC9QZx3uvkVkKfQu5GKCD4wGr7OLHKT3Qv1etPAJkpa2iTZ70AJHqfbRLOGViyLTzP
kjF8xYltsvGsbYKhyfX8re/sWg7Z6caltfig8MU0XsIIlj6xxG9BcuhlP4z+/sUAxiIi7WUqbcpg
rxnED9fgt3L71F/rYCA3oTNE6dD++gRTRWVxdvyzmsYBY3FfK0ojTFhsEGfX8kxpyr1dObBT8f6w
Vo0cCqm37B/eFYCxnr2BMuajC29FU/VT1dcc++E9UO2h6eFGa74rmwiGLUGLdFFO8hJ+fwy0WgGa
R/KhpRn6jkcALNyTAb9HA/wOIoNtIiypR0tDYlxDfwmrGdErub8BzV8o7/iCNJcr8BH9ZgtWnwhA
X8x8p3V0Z/yXQZNu1ORSyknBfQt66GFS/6I/bp03cOJ1ysKlyfhSXqx8y4rSTAsU851vp4+j/ghE
I5veM5Fc0lOyJux5b7wHw+2bU0UnstU3zkBNBHfBysgRV9Lo05It+B0PlB0DK2j3bjwK7a7B6xVT
tTTvwlwNPszHA7aFdi148WCQ+ZkW6CWZmDZb5qaRKTbqmz3O2bwiOGarkK9aqzjj10U5s9H7LxXT
lo+XroHUSpl7O3bYh9silqJXkJ+cU6DSMZORa6QmdlxyGkhHTl5wuzIb6/KKLO4iFI4WsyfZUauY
rvRLj1Fux8F2wU8Yv+0SLv49J6rXtqsojLKIk6f/2ISd/OwD59nYKfqW0Z4wlO6Ffn5n5ouQPWOY
5Iul8U9qfo+mm57BpG2RhZ4jJeLAcEpAcj8aQOiDByIISB0K6Kaqq/ln1kkaBhoYifevdiWYdaos
RyDbzEzd3P6n6e3wRNR2ycfSevUJmUZPPRAu39tcWq+nYqt8+Gz+T2X81Ba2N1PEFMtE5jz1JL9N
SBGbMPU8yKArHob7O4IZ/LLX8CV9N6j5gU1fqovw3MElHppww2FwrCwytc4XaHAYwiYHl7MHYojx
q4JEHgMlgGt/Yaxv1Xh8glY4UO73DAFg3CDGDfWLeVE/Bv2G9tfi6+mWD3ozp5a42mYzHsmoaJ8U
rD+/DjL3sZj2iGUGJ45l7ArI53PvAZrQtoVXk2LFk6hBN9hKVvD+qqupsnL9STOwNIgPegKJLdGb
XzKFq5p1238l/+gNka+m9GnV+RvHez/oru3vNjd0rEMIruoh3v+gW7VO4X8WU1to1+TfjdcRMpU6
2577aMvzR7JDuwyGW1NLR4S6SXJ4t4RbHutBWenHoEM56UxPjqHy/umbp/qhE0FtQTsixaEB/1ur
pGNyS1xp72iuvM2U/w9YN3dmNqxJ7MhSQpHtZ2Q3d8wh6CzJ4eHOiGHqaTwxprLA7nUEaUE4WwOy
qFMk3XHbjKxtuak7YhJ+kgWZgfPBO1sQKpNx2EeRy/nciy4K/rPgyEMVl04LozA2fj4vhoKD6mdS
hXEkVehtNGO+4Ck6gjzzyQlbgPtcUcjhwm4O9mpYBoxZe47PpTeA/PzLhUVKAGU/duGWFFge8Cbn
WtnCxCmhiMti3cxZLi8MbUtybDBp3AxPlFuAFDeiWIko4AIXHleTyQ9qNsDRovALbiY8I4HGpVsp
VuJyCKsEGIpfo7P8P8yLvbohCbASHzz9ALEjYXCcwz5KTZq7EHpNlEfXzrYY02Zao0cwX9fT38k6
PertDIhyXvZVgEvgkiPXJjCVAIE3hwDzJUZ/KDYTuXAaC3AIyLROaEzFyKRu9cH9bFzKtHwQrTcs
O7f26DL5ceIlS0P4WluGev0X/wqTcHM8074WuYa7xvamDS2AKTDaQu0eDTAcYKi/OhfSN5ZEZfto
xuO8QgLl91BQeT/QCY+jgPj/7ijIUOnjEJnWEKq4jEbCy+GNpt89OIz6Bkx9ktMbvWCAXhqazQEA
tr7IgBtjYOFR4MNM/VHypkkW0VJ8JtA4NF2d9IO+9TX8+sQ0xjUMoTVve/YKG5YjgYtuKNCYAjGt
DoAEFfQsHhmUgpzDLvVQQr9TdmsWpzOQPKrsuI+phYhsVlqhwZqK90LhizMfQdK3opVnjWpVOjOk
/QGcuWmluxSNFTRr9hbP5F2P55Q5rNl8cNtgCyxKeNWtAeOrznSMVyWu466yOxb733wwrmw1Hzmc
gltv4EBiPrdBBtrwVeGBnPUZgybeFkK3HnTp5nuN7BurjrnFbsAtbnAMg2CL8v/GU9555DaVNrh3
26BTAu+jw45lP5i9ewUjNj4LtDBCH2Hx92AUQ1LkfNVuFpgl/0H2FKyUluz9bVq87zQRb5s8TgB5
P3IQAgLC+/DMTzHK+K4Ep1uJoAxbujXs9KfTl4CH4nguHpeYSgHWORane1N6jExZegw59Gdy6+qF
Bsk5w6Z0YdaAcUk7e8Pdyx+riTE5CFUOHiNIPpqyvKPtrRlU/h10/dhpNyGyvB9CLdDaYSsCxdyO
FPVu7x8sX5ChBq2cgE93XZQSS3xG7w6C2MtXpwbHj3PuhJE3mZ+IC7w4z9uycG6sEYAodMSK2C0I
1DZuhsRCTJ7hf0XzKse1OHq/MKF4eULiHoY2RTv7B11ZK8eny0OAjfTDMcZi07czqOxRzLk0zKLn
6xD/OY2GohqmtbyGoP6I90gK266ErNN4n67T3ntA1xKy3qhCywYrfvuzb2beKaaTvGjdHdcbvF1f
ySe4Qx7lhakdcjTQWSbf/+73JFv672bQXML4Z9HBcxzG+kIg1wF/6FH0FhD4lRnWJGPEm0nLaFbc
iVnJ6viCODCb3mMYYdGEaV8+Vk1nQrmKH6/FWuJgHDPK70zIbsYlaEPPM2lyvIJPxKffUZ8rmvsL
V1AORZ905UAlsqRcGsEfgkbHaGLUpdSY63+9to7ydTYU3XWkDtULvhNpPftBMwxoxOVxaXDqdMZe
BJQCQpV2TgjeFES2xZI4l1mnfcjxSRtFI0xeutayHzTzYzL9ZLcWMuguYlIvdusZC7Rw1JTCScYm
N55mqxgR+qVR4Y11UEI+9CHJ1knMV+Xcra60cJYlNI5V16zUuAkXT8OMA7o52uxw/ZeWd4zw5H60
glRLw8Z3iXs4YQ6wrH7+clUQsM9+LU9HkAD8Gmj3jf2yGHToIO3LDZhHKVWKZFusYMG4kRDpe/ia
5oE/kZ/8CO/+94gCWa9DXT1i7Q55r9dBLgkpBtYvdWgzgbKAWq0RB+i9rgYJqwPMHx6cH6Rt6v0T
HMGNvzUszu+9Xsf5OgWnRR48lM1c2eJhDYGL/C5WfGl8bD5TAJ5E2ATMprPihi1a4ZwaIPxiuLgM
Gc8NkdcY0rpLuJr3C4Ylddd8g7vHsOQ984tZEcxMt63DwxlFWX3G6Ss62pJ7drzrsZJL8Nr0UH2c
wDMX7LgOau+QYKKSZTZHolr6mHpkGaSzfZgYk51cd+MrKfmobjRIrDjqDeKCrVsw16BRycZAwng0
MexIj28UBTlo1Q7owYJU3qjnebn/RnOvaRuEwifUEX6W4NC0wNCdlY1Te3o4jsF9omPAjkk9fWEn
c3d1O6JAtJFGvJDPZFq0rdFGAXJwzMHtYw1nx+P3LLCtgfQ8h4FwQ83kvxXYy/44+Hbq4pXFe3oM
EgPBJZUj4I9o5My317N79jsnc5LU4RnwGFXn1g8GyrHfNQH7ptsaP7JK8BwNTYvgHzH+Gpb/Uy+7
BgDB3AsD35g4tLwHwpgX2rBR5e93tI2UyLFisVVHIGQeQlzvMmii9nHhkTshJSlSx8lCRwmaPjR5
1Z7GV6lc7s5ido5aauGTXXHoppnluC7Qm3DfBlXd0g4RmNwRHH0rFG7jhx3oHS2c5G2YONwL4Rjo
EEHfMf4BnXaueIZ6SJi25NMgN6x4FZE0/sasotH2yuVKlv/B8KSKjMsgPHpeFCJoXQfLkKZMa24Z
GcltX4WDIG2K+IwFrdWDUAnzujEQlCzpn7rDPqDtXbV9E/2s2m7gGMugvKh9JUpit6+Yk062WqVz
rk/de0KaBaYyUo5UVOTPdok6mNzdRatgbedirbxt+I8TICmRlZWyLgTBUbjEesWTVVKjc/QkIDAM
bS705Q6M5jDuNp+4Z5dOaUakBnLIglRfUsl1zk7z+4Y/SHLC6ysOiGQZcVAelXBHRxj0BeWvKuY7
bpziXoSFk3tzlKh7yNnJD/yHWRUZgqKYPuRqE5LWjVRJHy9LgcH33244QZVpScL6crQzaRh6Pb1Y
TlBHSBQjVDdcJmiTSzZFhVj85w93YuKgql0QKqlzp2yGMS6ZR1GtNBL4dTgc8i38UC9RwsXvNPcJ
ifSjIyQogysjpOWTXPgKQXiFukUX3os2PtCGeG/31BSYYNw+bWgxO3ZgyQX4dav/152Q9wjazqV5
LAMq4HUo6V6MCIMjd0OhEVkHg1logOinsEPpVY8lLYQVtQaetEc0EFw/4XoHnMWc1IoJ/VmcZiFk
ub1WijnxSeKgzgG43CSSP1NPmbzq3AJwG2KuNLH0eQZ5128/dlknLl8wHmQZNsL1XGHYpNLCUa7m
WK5YeBy03sOFnp6O0rwC5v/VEOra6azqw6Rocr5pWygsbm3sluKKeEcpUlmJu5vMZlNKVj2TtAXg
lv6xSRSabuSHcaH09G1EziJr14bHIoKgudKo5Y43hH9Q639CQdsyAPB0Yu6STisfCt7uG5jev3kq
KpFlypjziAzKXO60yNSPNuik10ontR2xg1XDWpszlYNwopRfNQMX02+q8QCZMTMhzSp/whtJ33w4
4cI2A3NfcfKmYd5CaaWGsi+6Eo0/6vgyVGryArGFsG0S6+DLO2/rk42TVJOh8V5XHQx+xPMWYdDB
k/ZDQIw8D21nB4y3num+wE94ZLvmcJU/A81cOHWad4bS5HVRGynkL4ihD+VzXuRTNGCL10hGKC52
MCahoU6ozFskiuAdvUWhaweptQAcn26oCPG/q13tPKckbBTBi0DFoNxAsvKPicBs2pBH7R7T3mPq
VCkEmVhkYYvPzM1FEfct01ZhPLbypR4itnbWpkICPXcs1ShIA+Ylltyxo5aWhCslw1Djfjjck3OG
34kEbtkYiUehXYCI/jK5du5wBj9DwszdfK3wXotK+oTaV9TnnmWbVvBKIkJ0VPmPLqhKySYxM6Zb
5NKHepdi6eDH5nqYCUIAm3YJ67e9RWWO4j6WyoJN0gURhOfNio2SkaRZDa1GiBS2kAxEZ6/Fjjyi
X7vUisVS5EBUp78aGSgz+Pmj54N60ZUbCHJzCbpoheGQbsYwcOcXkoFfFWG00Jg1uPvEK7U1nirt
RLYTq0uwt3Qz+N9Wo1ud51X/pl77XgrBS9mgm8saMqg97DnucIRgSwt1uTXbM3RX5Ud8rNuhvtGa
f3DPlKtg2Oh58IDGJn+GONSFwsxOjuVQz9IA2tzzBNVcrq53SYz13TJa6wgkQRMXk59JB4W56e5g
kEgurvAebg+kWLH7Eyng4rJGl2+fDcXOSddsr1QYJIr+c0jps1eQOKQMmtGhXxlbY9L7iSsTsIQw
KfLevEB0WMnV3/DoZ8LtK3QqrkX0b5nw9N6Wcy5w0bE4SG0d2NnizqjpMtD613+MAiblzLcW2OKN
iOYrChCYotCD1zRyObdmoFNtQEcYSZaqxugfrSnIA766TfMfI7wj58AvpO8ulb+xbXmNT4r+JuDg
kTN7khqcQQmAWybQAz4vYwSe9pCBcRN7bK1++r44+WylDz45SgMTR+R+Xb9BTwRwwlDWuU5TL/Tg
5eFtUAtLny4evKtG4FG1Ls4Suvb/ytgi3wIwwTVz6Ezd4kYjkJkFbNv0v1+AxRa58Yg+slpRWZPU
eW1ZtqO6WEj8BiZDBKX8d+aoF1lpR80qZMRHJaBYUEs9EjDlO+sGMsBzQko5Xfc7DCRTFh/xh1iZ
z9qdws9m4BlaMOFAoVx/ef0lTQ+0I4kTDi+W0d8G16ZWCzFzcof6KpUiy+7HfggDW8OHPJX7x0aw
Pay1xj+7FBugXmIZSuzpm8kiIS7v2BH12wMcfq6bNacxfwFiACY2JMMA1ckOU0VopCC3zriKyRn/
DS6LZ6D1cGVteYepQXWh5c7RGvWShvbyCJD2EoXzKk3I4KvXJnEuJ1R7hy7mSu6wkyuIno0jl/Lg
EpKg4pVdHC5602+5/mQF0SqJMoaaILAVNSxJTdNWbF95YFFYUhJjtH6AdLl2CeGC31lyVlxexHsS
gSuOooz9rLvhLcqk+zFmL9H6dJV9/lmNrp6N3IjYAr6EuF/b7ruHlGOS57PqGxv8rAeGpv7uA7q0
3l5qS2V3dQzxPS2Q9YqE/n7ZnQf3xLZIzaVh0eVNmfEW3kd+KFgeEleIqQ9HMms+dxGQiHeL3825
zIpsnnb4t9Ty6jrgBlhY7MF20oUlgUarhhM4Wxz/WSoJ5yRlOFfcgtJVdq3L8cx0Y0YyzC7TXw3C
qdiDv36633jyJonuGj5GsSYUBjFMtMFkmWmADfkrASoPLujnes4jlFbrukva9T/61Ym4QyUjDJqu
mOIuGGBKDv5zub/34NLpW7Q1m2gaACdUyEVeRmULRy54s4ioG3qFna3vP5ALfND9DX9uGyxr7Nt+
LPhnvfmpwdEnT/ATdQJP39NlC0u6FGFc7TimO2s+nkzJO6IHq6EyCRIZlSLNYXFHfpTyBPehmMZL
iDkmJ8dfvWyp2lt8DK/l6O0hmkQMEM5jNztlWC4WHjzSiVR7Mslj9JkwCFjXhfIPDdOnwAymCiXf
7RZrS8jUti7970xlZ+hFa2yFvjMtEd+T8pLvkZuUhoZvjIT0pmjud3lId2D91QYupHCsOqWTrLjP
AXaTMZO+1EQdI6zjIC3wkpYW1iVeYolplRK3oTvOkfw42EbPESTd4kv1yuzI6hZ4KJWP4BlnMsHn
iE6KmYlIJtePRcqzZMs6og43pQPRi7biAUxlTLJk8PG9GJ6OX4sWyDF3ZdbkxvRW1GdAjS3TWYs/
WqNdMWMB1wqAIDVqkW3g2rs+5OWFfK+owbAn6wgPEg43u5+BfItVa9c5UnuR61wlFMFcD20mknCS
UJSiryligZn936B2dm12LXjO3fFC/89PnpI5vvu6GG7GSmgemoIXMaY6EBeiCaECN7D58GS503Rp
A3htXzOEDPhhE4ux4p1SOvso9+45shsVFBLEcC8E0zpgzI+CaPUEk0RuQ3uanv9tgSxlFZwLLbZB
FxS+VTUjyst4CX2lcFmGj/WHAo3bwMLevFYYW2zGsylk7ZYdoBvCoj5Ld7lEflHOsd3hQhlBAdOY
ZD2/Za/QJUu2lS2xZd+hymsE1NvqVB7bHRlPTHKxjVaPIZK3NXABwxFthJJ/6McfrWQmo6Km1vXm
nY8uiZwPbMFvre0hlbhuZL3oCKrhqZyBHWDZIv44tRDW+kiidirQkdWLxcjAichKG+Yg6s9x+5CC
Ew8yQwAWQ1wG60fs7N1oZV/OHzRxnEcMRgPU1LrGPqYbFSeIh8Rv/74Yym32XbAX+NRKOVP50Xf6
edYAHXTO1AEnfH1X52RhdoovrnzQ3I/5++Wu6u4y/vbIizNGencrRzn6KN0SoimSggBZ3Z2SRHo3
9g4TvIotNzNi7/Qs/V2NVY8F1eSf7sWAugoDm7DF0gzzvlsMqRCkboVzR6t0k5e4Ay4nILzdrRJ2
r8695n1B9nkOTYHmR8JeyqMIAMSym7UIZPhW7z7Itydo5Bm5VG4pjxl1+7QHGtzChYfqrVnEjgce
+OlNJse/hZ9fAiLwUlUGDXzf8Key8Z6a4ZlOMCpr89KqiPDguomr1bfjtc2JI/O208jHEegCoRVL
rXj8HODOhcK+Hp4movRQPxywJIuElFZmunltbCVpO99oCE0u8oWqDECEuj51V7Z7XV/JOtDUrBtv
7cbH/3Pu2R42fu9sVUa2woiOCDhf6AeMqTTcvso8sI/4kz9P1E7hn7i96+pAnSHekjcIzrvjLgWA
3Bhe1DNfKiPJoF9A36z5NbucGOmDgEZ6IFJmOF9Rn656HPvyvBDK3qOryCnucmSsgpOaxyxm+ons
5bRFf07PpOTvG2aiKeNTiaXsyXVMZM/5ReQ3+c5em1quj8zWU5xyLOUoG87O2Z018ELNTE6Qr7j+
A+MAoGiVZe9/cJMehIpvp/M5zh4RgBvEHKc8tlcedMnAt2oljxMaPBGox5UAytbyCPYJ3DvAkoEE
f2wVjWFjTFex2TqjrmkOGyAOympUidF9enCTABmMwJfCYQuCTErp9006K1Y7dnF8C8z2rucIf1kS
J95K/JuGPGt2XsPdzfaikoDq6cI97ol4mASmADWi37iaq4cQ5fJtQZyv+gLHfTkN9k7u+ANOd/OG
vL5A9byHh2OnYkjMUXTWIbNqhz9IGsCufZiw7Tpze5M5+2MfIVxXTgksP2/V5aYcLRk2NuZepsur
GuShs1R5PsrUoOT3rG6205bvVsn3/sgwN0mzjH1QeAo+Wo9G8RCUZo8IzJceiaJzofy61E0jp9aN
pxX9/jfQE8+SFN1vgRmW+B1dRlL5yJAcpGIpOtofgMZ4wz7suhzPnmO5qSSPPbARf0LVnDfZU2kY
l8nZ5Orq7HgTGSVfLPQ7orktjkcMgLVXf96fbel/KbW7dShm7RRehSe8br2S6jjJdy6Xb5i4005+
dO3pon1liKIzcFqGZkn8fVnL0JpmhDXQToNLWS4LthdDFz9JT759UR0oiqHX7SurEBupKPKWk5B4
GXM//5daYHa2eCnYswtk7JCf0+amfu5AhBHsqO2Aa1s4Zmfxtk/+Lq2a+wBf/0oxfjbJVaao6+mE
nq1UuAy+ZZi2+xBW8XKsqNteo5RJ/QV4kpk9oJtEasav9ybOgaWfxaveIl072iCIN9ldauDLQ2cr
zdkeQp8cqAFOGmxZbrYZJcKf1CH9h6BB4uOjw3yJ74x05z4CD4re8v/fIUK41tQc+9fegcIopbok
qjX64o9a5IKhVtngKdAtPM5VKrCKx+rWwKhDlCgqHCerVXdSJ6flJyU4522qoOagThRat3kXmMvj
HEoudRNwLAqwbOcNJ6yKl4PZ5BwVKTGUsaTmafaz1e21tublL5bBIL/z0wMAyiGD+MUfummr3VgI
GfUv3klpjPDBeSXLLDc7mxs/K1zuMFUF7iR2YpOD17HsLI/8viFsNFcZBLhBIrD2CXCgBdebP+q4
73wLLnuBvgqA9hrZvJWPr2efFOWyLx89G80DLhTeMTHpwy9rGBoxfXgIgPKMTJlS6YB4xafg/4K9
x/98n5hDT/m01H/rCOZkZE+P1eHKx4ybzHG55Uuf+xA04mfSOUL6euBEJdpiuAPENfwZvYI3r0Pw
Bybk/b/y8j/wFVyqJ7II4ym9km5B3IfPBHrLsEx+Ywn6RuFIFgbbqnVuRZRSKLK/yW2Jlg3PYUXk
1oOnyznD6GQTyp/bP7KhgVqxJTnBUEp0BDSrEzYB7t+5fnKXs+NiTGr71jWUQBoz9LV7eQahGdJA
Kx4SU91Rb/wz3DO5KLd2YSny4Cy4pdunCiZuMKqbyrDbm7r51Wa5LLQa8fli/37XMvRnT7dPAjIN
Iwe8E1uQ7lj2BNZ2THHXB9zuw6dbJp4jhhlQ/JZGvZpFKy9d2PbOOro9me/YGdMoeRDOk2IoNdHr
iuJEourV+1slCEbUnDZLBFt2IdCmVXsOdkkyBdLZBAJEphoWsgymVX84jg4N2rYt5vC3mIYbqbvm
aygsvIcv99sdswILsXwJt3S56KclEUjpAirB9CJlZZ37U6YmMrXiOKIrdRH1aGmqy0fElnTpcDcP
ih0gVSLEW7rbQ7M+LhkURYuPou6o9vb08eBHiWJjE0zVvNsO/hjxYKDBz87T07/fpl6aCL3Ztev5
5E8POo3Fq+A9KlLPbeRUtPHDbKpgjNgLsgqqUXX/540feT7WJz0+nLGY2JmihW9aR+BibF1O3LAJ
BLZ4Vh5xoa32e5IeJxE1Y/uhZ/vzaefykYlukHtEb3ZRvuFBpuhyfAjyhBp/GXSOp7wCn92AfWyp
HdUyVFMt7suPZQrhYEQiqMBhh1i7/K+ty9tNnhd3RvSmpswWD6efI7lgLZx/wKxQvz7vcGdZjsP6
yZCDTj/cQ8ta36q6eK2foQK/gb2+3dGVgeukgf+Z1Gy3rJcLKEK37xBKaigcgqDsWwVYcwnaiPXM
8c+62R8kJ7yBI5CbfzM8WVeIxRFuSkfk6l38tdxtbTMSZoUSGsxM0lhDsiUhp0WzCYvmNAo3m1Ls
qv/NYk3LcxuNc7UHfCS/ORJ2UogJqtEDBx4zZnNKXwzxx4KnNQpZXkMRmHOnATtRIkyRdyuCTuuL
iPby+s0TF4CnGUeMLiJgJfezGqRTiWyPLUhFb8WnA58x+gdL/nGYNgoC5JBQpyGUZYHkp7PRR1Ko
ixn6iaQ8IoB4UPwnLRfe++e+ltz4HazV6P0Y7Fb253iB/53iP7B0kx+MWGku6tpjkg1G5FVKczeM
mES8QFzwcKxkmsLZ0yWDfWOSJY3jRvVwuexGYzbizg7jUS4sK6FpFIaCge7yRWUX8DwGwVZd/yGi
iDpj1w3s9XckV7RI+I7vQb1c/tGZAZ9rvZzqQTGRoPGg/+9oKbwh0ggY7hDnYbVivhca3jyBh1or
q3ekWTt3sNeIOPgkP3S62nJJ/rQoUXybNPK7xhE77dEoBcBTPWfKjaQPQDmWeHM6ltQ+mkg9Lnko
3J7fj51C/4uPhs9Zf1map159F3/CqzCQwaam1yhyrW17T7Exq8bWCJ5wPNRCbunlJz/iP3rhA3RK
YuKcLnjHCgPitJJrFVjgvoqwGeJQ8K5kMPwsxVAhuYl0tf2W0htYNX4QZbIyfn3O6MYELc9A+uWP
3Ufj094pJNyzGDQrkWVYv4yhuLxylYAeIySmUbtvtZ3jFxMhHHi3xuFGrY6O1XY99rhVI3eVVxVu
sMhAr4swzaKHPIl+bF70NKlj/oXqdWPjk+mdSBMWZFp8jGazS1ZrqWL82gI3wAzPWCXrLxM4b1L/
qywefPbIs8fJ7iSwEVDmtAh2qqBWzDRXENzC0lHybvTTY9KYJFzdpZjXZRZrjHzJbsIim+G05dZs
E/4MaIStF9wxk3jKcFIhb9ESGFhnJdgSgW4JzS7XoXDV95sUWAG+AQB0wS1lc4a9Efd3PXTWQbKr
GezeYd2Oc9gLIS6Km8OJwn6em4mi/WyQbOM7WpBR4X3KjUeuUfpCTC05BQ0AWwoPqYQf7PSP8YbG
ntd+80lXPiC/m4cznB/puL6CcrspztYvnS4FWya+eNrfqMaN9q1HNFMeMIbs159lnxDFLZ/z11SR
DRnVuhxU0BIl+1ovpSRkmo2Uc+NVwLBVL7fHEBAkWORKgZr79Kd7nfPIgMRJTIX9inw1Bw0Z217b
zuFMPOYXcagJIMrVe/RL1C/AgMl3ZszHobpbspHbttqCaSA+KTucdXcv1Odmwv8xQ8gpbsjBogSc
Xr+CseahwE1QQUzZN3zVw3vIuDlisr0bVvtlf1QZWW45TOYmrbSZQjurZO8myhz1zz14e8DY+e10
FnsCg0nZa4i8NtH+cNuMGD715733Xr0KURqQXbXVGROEFwGePQIoaG/WEvfB86UXGN6toUZCUUY2
aldVVZOzPZ1Ejr8u24ZP+xbDrxKB2FycxQihu/eVWZwLGB/aPdtKsA/37eWnK96/EMpdUS39DCLM
gUtCwsoeXWtaQ8Rn3YQgjyItl13oKjbrm3IUPkvSG+lBhXEYrefhCDmBxkcZEa/vA8NXE4kMVAF0
SX2MiJ97UodgcCBcJl5D5EbSROenF0EB7z6IYiCyBSUBkJ0x9eiWVHgh3+tdVYNvKX17vrf9vV90
aosJ+vLNZC01KWPzjKBljyf7YSFSKWDTaoKmweqk78lbWCu3UzbfNPReENkqGcFIprkNhSOMWdcg
7d7Cl/CxxifecCwDMBHthK5zW1rIbxkboP9EdguCcJy8CeFF9BAunWXGO3ICby+3sCCrhRRRvoXJ
m+qyHgZ/K7Il2bwB2uVEbMfPYG/oyA1WkhRXP1rMyp2V0xDb8hGtJ4EuOCMabiuRxp0L4bCWzBFR
RhDFd3UU+kaBZwdpVAK3ipjyoOv12USdOfPxsOoVYsNBy04+728US9tkkydNK5El+qCegw4LKAno
hqF83sGhlDdppkG0EaRToN9mN3NGnOWZlaFDuxoegGRUTjglvLh3Engm3iXkDEwRDaG7jfAoX5wy
K1rWrNyIRn64TdNiyhiy25WRXoed3tx1mR1JK2YcyfCM18ex7vQfR0xmMQDV+LCfW1g/kM0l/QbB
OQcXnjoDyX/i0HL3ndRsMHQv0Xf6bqhlr3871oj4Xdlv+x834sZnJBQzANayqDtN2mtafqrrREGB
yTOUj9ecMgsMU/FS60TF7bIAvsm04mkS9OjtcOfrLlMkO/ha9Sw/5lUZYC6PNdQ3bTV2KDMdD4DQ
Nyni/N3cyyxOU0J317VdmfGo7jV6rnHQxxbpWrxJABh5zRObcrRwrumnnpc/29YOq+e8KHhKcXLp
CQvteVb9yIRc9OkKp9qcQ+i9ENtxuviZ/xzw6VH2qneKaV37/yCe3Cf7lCbKV2B2AgCCtDoaFhu1
5T5CNDdCBVFLxTUhZSzpLYPfVAEszqqfdXGDKg/1Ke32lz+kO3Dvs/NihLmMZxcAGNMIuu9y8QZk
+M/WeKeyOXrw43zSrXC5nyB66TIl7v/aDn5kDvwOnu56B7F8iMQYN2mJHCVi2DII6XNwddXuw/Y4
cXyI8mBkOIvGl5677wnT2o87GJ3XGcEMt6d6F12snBSv22iDZflKqERxdhJLhp8cQPbr5zQeG0fs
oh96kVD6bppSlDy68vyUwidYto09YqJWG84IMxDm2BpI5Vl4Uj5f/husUX7qfo1ZykEujK8FGXZd
+u3po7f9ZBzmSe6+GoLblllRry1Z6G1wW4eQjaRbkgLZgrbv03K9z5uNi8opY3DHUvTm3TjyYZ5S
U4l65xcJ9854pj09USLmCuNRR5fIhbMUQcG4WKeGNaUlYTrwjcC+CDmQ5ESVCekIXIjFceiEx9DU
OP6g2GQfkX77tbJpMq7GBVZID2mFi08OzNH39cCSrninO7FxLJQsCzP2WztDJUO76zRNRQ6ovFkb
fXdVsUv/PbhLFrKv0qFxVCEDXoLfxsoHqHMWdo+JzsnAh4FtDZv5IAt2qrITpinewaervGGGAMnH
NiFxaagLxeAtbsJx70VSVt/QOSn97YvMhodliP8vdBdQZIMiys8KHnvP+2m6NYyCSNhZBsz7+wYa
AWn9Z/4UQqiiQFn2zP4aHLr6TZBDzY8GTguJwM9q1KvmU+PnHyXo5LTGXH2CGdJ5W/WfiLSJenY9
FPpjzyTlzmbnGf4HoaJmNGaxZelX7eROWYqFu/KrO/55zzCAcZgXGZsJJvcnFheDk7vcoRjuSTIO
F8lH9VZwvii3Auc1LtQmNBrqz1+lztP+nIjiZSOQoesBQF1LmTCw5W1JAoaZp13Y1q4lwQkGIGA2
VwLpet60tDAWdK+59w5uqi33OZV2ZVNWqcvF3JMKU0D0FV70SyjSC31Ww5zS0eIkeASDM3jh+Ilw
ELhSeHSvTjfpota7/s1K7RtLAcdXd/uGe832OKkv+Hih2v14dvpPcBKnVyEFLRoTm5Vnf6iZyPYc
BbKCapGCwnH2Es05kfZH52v7BE3E+7Vz1tJULAtxmELMMgwIMWEM8uDKHPrHAqpSgW5V2Ek9ZSzI
tXPmPTY2GGhpQoKYgYG1WTBxtbTDGzCYQqhFr0ddt7r2IkLk6Irjsminw1YqLbSFLx4K+nZEej+X
rSDcFBlC+Xcsmt9dk7CHzC/98E83Yjygvc6HuWhQXd4xoW1jJ6O2l7pC4Yb4rVh/EnPiYoeMkrnY
lkD2WPvq8rvPxdStRY4C3z4cq858DlyQ4lMjvPGdCVAXAyrGajC+rKGAPvSAX7mWX6kYLketNL6S
7iEqpagHgiMKMXqW6y62VSfqDnnczQGO6fruqWEAw++XHTmBzX9cmkaRfzv7mEBjvBZu0mIVO/26
pxj/z9SBhL2KgIOKV240hfZB7H9dQmCXkJEXQrj6qmu/FPdd50XrP0puHI3DGyXekkXWNMxQXTJq
C0rV4anskcJx0/NyFpu+9UhgSrkPBqYRe41iH2Bo4jKlDbFoN3gab+eSKYbr90cZtvJvOA918QdX
gdADbXQHx51Hf6C7YsMF7+cBicsqn2FBQXRqifu48L8QDfV6+KRuXl1SlrWJeSTJErA9bVeqRtXJ
iDXTTIVKL9atd5sZ9g85avEt2M5jhky1QotiWXkoXb+9FT9dVnvhHoFSGtHj/Ij9WPnXz4kz30ag
yGDuFZjxrC6QLWBV8hcDgnauXn1cNCISlm70NshtnxEj6627T6aUh+Weki3byqzhTW99phDi6vgS
t8kaIdfKWrf25SQtpPv4vL9bOTOaWA0Vc/lh874quZKiieqXcEtGem5eApJafuYrqHmSilhyUY/u
46YQgTDIa+dW0PHtbmISZkHoEsNZ8Wn5AcM72IOqmCYgnREjmKEVrkTNWIjsiEGL47hOvVvVmJCM
RUOkUHreE822Ob7ceyFsmidDKGVXrHFSz4/MdWFxjQt2myqchl7UyMP1KBrKez+ykX7r2vN9PMYP
4tcWtLot7J/y4daau1UdSPzVuvN2Qu9i98CvcxtUoASBkPzwz3yb0EqcuM+KYy+wXhNDlbzVbpje
Or3ASuGp2V5Qk+ur9C2RmQL3E5z8rZjvdR5k5j2NzObRksr+4VtRjS7agXu5AvKuBBR1T1Zs+cqm
v26cMIDNvELMUMdqbwPVYobmSRzVXVmtsZ50UO1DcgQejC7AQFd6ZQDyHpGlw6ae8KIxHXAMuvD+
zG0+pyjPciU9gBCci/bwdrXF3bajg/cBxJmMK04JhqJDn0vTT6EHahF8gFRT5pl26jmAOn8vV9zW
Bo8eM8TQu8HsvFJG0GTTYvOmWpm1RsQY8L73Hb/Kq/fa1NbzZkxF4ZiqujcncDcdEXY5Nss6xcg+
oWpkQ+Eb6djhE1D/jGX267DaQ78hmQjGuOtl5hIZQKf6CjWuiR/2SdRW0wpeAisTe60vDFgtUHhq
SPFf6oy7M2Qoa//x7/aluA2dqKA6xqlWMYjoOcG1JXkfQwpBBv6sZ1QZeef8kaef/xYOEnKNZZXF
G86vGLGrS5E885dlZGsnGUXBfdVIgzeRJK6E4hvSsUQ8U4mDK5z6N9SsVanv2xZIVym+rlHnP6u1
WJH28WJZJUHcqxRy45p3CeIMuMN7Tv2IAcxpTjcnSaVOZVHdNTPUalA37AZUZM4+fJk8UwKVLuN2
SkSghZHIrC/fS0oNtgULSZ9PFrjvSpitp9D8deeoKpxDIof1FxWZb3lkPzbUwmdTqdT/zPiCNUvg
T1G5obfxFi14wpCcUzp4g/t6nTOMObCAsZRdp3V8kNfMKO4qvjgOGAzGCnoGr3fXI1xPH8DXnOF+
YKXUHDcFf3RAu4EHRNgxfzWrPAAxuXbPIZg3MTTi5e48uUBdMRAgpU2no9iNEcraytEbXUHLbMZw
Hx+XO3M7yqYnt/YI5RGk+3BG/clBfGefhm6tMYy+w0TRkQiB+VG8frjrp7b4JVMAHm+d1Y8UF5cd
IC8PZQJZrfd/oJGJ2DnHjqOx92p4RwYb8+BBQDjfG22hHwIM83CeBhYuwnU+s5sRi571PKvMrqXe
xpzUpE2f86QNuvGkCtQstxLorwRCdYzUAN5hI9WwP6P9c7M4ySQyWhGuX8nL6pqXaSamLXF/F1Su
mfn2sXnMON1sQ1Lwgm7ySDdbqyfvq9M46kNSKIi8q5I5etN74blqN7tP5rrWWeN2yjttQkbUI2lT
6SNQATCCXSKC2w3z4LwqcZTQOQX7HjqC7Lx8qMVPSdcdQiWgfA5YRpy+m95Sl2SB7rdm6n4jvp5c
tL8WPgzMuDGAq+h2Ty+fsA5lYbFUdt/8p/d1jyRaM/VMrB1tAIfOGYc7z5MDt8Jc7m1rpHl81X9b
C8U6Zs8Zan66vtji7b2SKTXeXclcpH5XlYPN8YEH/vIbHqoxKO/2jEYbGJaZAjtvfl7oroKzcBq0
EhZ9a0A2DQiXtsiN5/SVwdHkiNEDtZaDYd4YGSycD/s1jm+tHxlPxmEzAlZpTNqfn31p9zU8TMHD
vWsEiKQ36gqBi/gNFfQGyqjKqwHnlmgRC2tyvJ2Gr7qd+EppqsDpFXYV8TucGQwU9BvNIJPP4AYg
2HOsc7qhg0GNKkTGuRYKNF/o9RkGIDxS24i3Bn/CVbXGCNpqs2KeJ0Uu8St/auxkISlGTVlIPfSU
+Mzyvxp4sHZZ5/L668+pTODE2iXGO2QxWmCs9z4grzG6U72BC30XBDiU7/3vjIXwaCskP1gF66d5
oB3TMo3AByi6+x63trUJjuLQsZXRo8yfsQyyYT+CfmiEKaVua0HYCRPHelQVO2HEwHmtTwhJdYTT
mHlx50C/Z1J4EySrxDLQgGTvouHX1WT+IApScWtTFge4CA0LC7XfZrPxTxBhXOxguoZemkqJD6Zk
o7dAOYZo2V5W5XV5UCi1pJLAS6aInHbeJ/Uy/ne+kI0Ny9xZYB2HKbRTqKEzzGWAHaVnlMYSJlCo
SLA34U2uk0lyO0pFjDw3q1bzw1mgSjbnZAAWbKMTwpvESHMWTqn99WcJ0P540sAbyMbrZLlTjs4S
A//SKEfPFxYIcRs5LXIYNW+GVhDfpJyNi0l1BwoQGLxTG0UQBeOB6VtNCwxemA3ce0dTSC4dQpzQ
m2BiWAz9bMVhMsfAWU/SxAxL98IJcQF0STJ8tXDWl3DPIflQz8RyhZtgHV3FG7mc6Y9w8qC5/iIs
Sx5V9X8xImsuDOw7bBS6YX4sPqd9G7FH7ugl42tBkYIbOCEcMwP0ZlDaLkAOkSXdG/Zd+71i7/j7
sv7FnQrbCMK2/wtNtbjpf6eSaiVQKRkIc9LOq4SHexNWBuHzjauSWmvQmSLXPeing7uMaue/5eA1
knyzGoAMCFiUIVT9OKnB3hVOBDukV+cvEirxQskij9eU2KhbKYUyeq/b8WI6N+H7quDFy3nuE4bY
SasEeK5NmtsKXaZnyZfH6kZw4gKKGiv88ajqveucky8QxSPxKFAqfaivnJ1dqONifMWBiIp65zf2
xf/+4zViTi7S0yDViIyJSJuO0dtpRQ7rxaKmb7FyX57NRFevVWT6jEB82vrL3hwN2VK/xNYZfYxP
Y4xp+GS0k6Zuzrro4AqVwyv36t22mwkvAQJOVXSkvvC2vfx8CZfAPQkZofmitBqNrux9VIOvpdz4
gslL8KOlWK9fLGJAnZ/C+vDlbpyPn9bDAa616kPK05BMGM7vtcqPojnOkbzsd9ORlcU8wA1lROtT
QWKAXXRuxobvaW2RONfbTGEgImgC9Ry8DLU3iL7sPJ5R8JOB01EbB3il6W92qJwFu4gjBc86z3g8
L5Oeu75JUF6Bmd6m3C9k4ViqpOFHAs8D71qMlHrHStXtNCJgKYNzb4bA9I2b5DwjWWNf/0i10oZT
4280qCRukgJ7lNJ+iGaYN0akgGgHXskYE7xhU7YEhiGCJAmqDLXE3dygkZlt1tgBdCr7IDdliPfS
fXZfHP4VT+J8R25aI9A5B1FpWJK3iTX5CAQZgmIcWT2KQYLAR0bKLYeSA3iihWxWP+jOSmY1dyvj
cCTIKC9frgsadIOeOfzoBRlO9oDODnIQB7ctzE+LkBW32rCM1ZYQx1K/X72kbYayowvhdJnTO15V
XO5D0V7PZ7sIVQYot6av/T2KldQ5fimUB/6lIimWiFElhZROK3EDmgIRnMY/Tkg/euGTZ1IsDZMW
WQ4MXK9mpIrJNyhSqR+oH0zUQwOdT3rwwCz27rR9bJuLibxt7Opp59dGidvmiJ1lDfjyDIG4eENG
24p5ewMu64diLP/pKtxZN+Or53K18Zk1tDHTTaebMjMXgAqmpVD7CEp5a/x1Wd1jwXnIk7NNG6g/
XGyT9m8Wte2F8BpijPvzEBCHK++PYv4VZ7bv0egN20M8a/I54zvxtG05ddRUX9WlUUPKk1Xe5C2m
N5lR0ygM4+6DRRf2AOvla1scFtdi8sFIowBOWCamqBfLRu9LgBgoDyCErLrBA3P4nD1yn4qibENm
dQ9ZBKM6aNUeAcdpzmX46JC44tp1D238I1SLeRW5sk5cPpyfY3dQB88gmbvi9o9uISH+L+3oLGHd
zNEu4mOeEqRaJ7ZMe20GZAhDNW8AlDWNhGiulN82Eesc5AYMV41KZbRVPXiCrSM+Rbtlkjolpz0y
VzUUdaFbkRQtgM1myAw2dCniOzptjfd5QHvUGkbqEwzQFL5rqYRUNYtuGBkTkVPh2u1DTm5/gMQG
9PPER/pFeb1+qK8BXP5UZbyqgZeCwOFWXcGaJvAiAGC19g3spbwFWv08QEMkEQOTHloULVxnGnqv
sdM78VSSRWdxOqbbDFBPmLD/M8HlmGt4Wm3wDu001BhzX01kUMNnKldnT1PiLrY43grdtr20zZOq
i1WHK2teoIexXQw2YjuNx14yZ+qBpDCDMm97rENraWCNJOoKsN0ZOkDTYjVliAzq4Hc5qbU+QyCm
be6vmnUh5LezViwFc571rT1vxtRYDr3oPUtDhiEBWLN7h2rB5Mgy95ncts5lLnzuTTcXxUGAl/My
PWspRKDYWmLEMqNnJpsJTobIjIbQ5AJ61aiS48dLcy3D6Ank5buFv8C55w0RjxnH3kPUibRmrFe/
qV4qlsorjRIjs0F6XjGfYxHS/ht9AS6LU/d+4TGRA9HwRS5yKOzRakL42WwRHqyPuQX26PEykIvf
mMCpJ5vmyy4bt04ywGiBNP+GlCF8pixAG1dtDPWDKrAfZnm300+P3UO/17dF/PRsvSQlTeQ42xO4
Nt5mw66rcZzK9mnxfvCd7bz19gtNgPnfdmO/iSOkEdQdjdEYpJ5Tmpp4KwEh/jro+wlgoc6daOj1
P5HGD0/qM9EfCn8TfzR5/bgrS4x05yiLidgCJyo5E6BPmAyiUGBlUekflDgleFnZm+zEtF2LEFtj
/1Tp+talMgm7XgKglsdDrVZQD26EBu6J8gXSyywEo/WLyXNzXuvzbLMliuJ8JjJrj4tLH7cmkwK3
TcRUouHe6EsVR1633EAiGOJv8RPKDgw9hGibmApR+dR09FZfSXJkSDGtnokZLgImAmzKkRBMiTfl
6zVZHI8+zOAV2rpJtkrhMJw+r747mr9GGs9h7BaMUMwr4C5YkKrzwjhh+V8FHYkySRn8vfWQ6Fqh
iNcZmMvHYS0BmKINkIoCx82BQOMNjteDu16RXQUrewTWFJqmkK8q8ubq+hrwpL3fWa83n1jIg+3t
gYvtCcfl29n7XgkeJwij92GNQmEYQsRgVld/Ma1/b8BlSsb9i1+oE4f4OGbSMlYEv8XXfkJ1Lvjc
S3LZqg+btJgf8NfZ7e8cxnKsFoMY+dGFvD/HXz+y92sCSryNzhuQwJkVDfzfvZJbXxKuW8UILnMD
FTDqlRgLgCDtc54jeTotZGY/we82cd1RW7S2iX4NjIz10jjxB0x3AfETeOeohL7Peb5AbSqtMlaH
Qffgf+gUGk0EbbLwsNfqr5wLqHyE5JB5q+84g0BhIRJcn0jLCyrsOyw4r+lztWb3uSeMA4RZ9UEF
BJIEs9/pzqXkcM0eudl7nJrZdq6QBpgDM8xSSTsz1P7puWTaOvweu8YKSXDb3BDKzzVqLJssS1jz
Dtxqb6ip+5FtBru3njLIU8/EIRP1OOziNi1Ydnv6GYtm+Abx4AxY9ShQw+F0pOR/oTC4bu8nIVDg
xgA9QvX2jrr/OkhlP/mm/GoUnbTW5Mg1z6LYVdEFRYvCs59kAse3m1Fi47fmpn9Sxy2CQsUzOv+l
SjUc1ygQ3pQQTRyTZ1anqxKbvu60FYmtXrXx3sSOt+XeOgXULH+CXPl4lUMOlnIK/JZE/iirJqRf
3pRilt1TCT7q6iZY12IIebA/O1krEkNNjNPjn2gNhiJ1rusccI7KXiz2TeHFjdLs8sP3M79X0rWG
yYABtf8ToNk3lr6lwo42XNlouVVMO/UanEdDv+GTkmWMv70bDMSCDhlR5VxndaIDI7FtEK1lMUng
MuZ9OSj8FC3yWb6IcC6uUxfTiQOonwcgGDZ6ZszRopgFp/e9KvpzDpMmjtbJ6d9ZMfhIfDrI8R6R
YyknfZvtRC5Ln2KnQmGboBkH3XSWgpsLtPJehjPTT8XTTiqR2q207I0mfg5ub4tTiJ9LbV8h/DWN
JhC3gDtljY/UrDF+Uh5dX7WvvJWvfp/COmjMvCr+1q4fU7eYKKZaAQnfhsKHKuMl/8B0fai4broa
rU4PDL9x6rq/LUfw6VweVFXd+yEtQXNe+Xw9J0DVnvJqrIg1D0BhwwZ7/rbqHhtdDov1b88uJwDM
Ne60gG147zY/DQ4W85JWVrSdUCta4p91eNEeA9Ec8yLvQUDDvDN5Xr7XwtR73IRC6XE33IzO1S2/
4D9zAYVjWYC6CYdy0DiHG45iE8cV4a4H7COSB3SDGblgFmSO4j0t5GP/BVwtNaTssmrhrbjMdCJs
UCemp8P6swKAaVo49FVsjOD0DRWakuiyxmiT6snHrpPJbLphQBaX1KAWimkqDfBjI7JWcg5MS7Ud
ngEKzZvMFudtxEp/AB75JZKNcrC1qyu472Q4qvfktP2GDn66Dy7wXkhwUmsTpuZRb2fj7bgd8WaZ
k5OwtM7JhJG77jqEE3JmGycdX3ot5r9fYkrJN9SIGOQHaWnuhVNVFYfyHxc/xjAVd42Z3Go0ejca
CCjJXQ1obTSYIyvtkqM0WLnZT7Ip45HI0zXKN15KbU4QBDXbvErzypY63HRBLaTn0SJy27HduGYI
Hh+tVtOXq2/heU+9w7m52ugvZugRdpVQxrFrPfL7CKZPqZDOwTqPeSVRJqK6pF2GVdxTCQp/i1F4
ihD/FTzYSzDxqevKTSC4PVc3LQd879sBO1eLrMMMkb0eD+TsBhU1tCLQXgKpz70qmwRPm03nsoZG
6Eel2glYv/G17ruhGYZ2EykUoXzVphxTi7HUSMWFFG2pwbUgcf3hytQlmbPDexmb3lTrohcW3qMP
RylPDmS6sGSeKXc3ZA7bQ+Vsyx8r+sssRjN6IU7cNjSI78zAkafAyw0rz0gUWqbbSx94RaFezx5+
BwzxgMS7Xi/as5OmPiQ0VIKsj3XQROgCGgEQyhgSjy7QWHLGjDiDJFr+h6A8QggbMNsQVnEc+Qz1
sa54ME/TglsaInpiKdyDmi2F/oCuNx1roruhFeixD4cg/d/0WER6BfcVqG/K4q/BMtgR7GvTJdee
ZWxeEUl/gIOSEgdDrlLOJrApiXBgrZ1lVwH7GzK/u0ofGgoKaKsMeIW/uc7oA9H7xUYmdJwpkJvb
FAKsPOnFU9PiTx9/7waR93OSQmgrHZdltTg8aD5CfvcFpfW0HWaUPJYYRXGKwR2lUotFTAZpZLwP
NdMBiYSQJ7lcB9gH+tgWMASGAJPZ6ehKK4efH8MSbitcakqJnlqB91mAhsguYYZhqMX8UK5kYz5D
3rXUwG6korSgM/e3G83sXyM7CFk6i/YveY5tN2ynz9ciYRTGnUE6qQFpJEMwkc5P2L2UJbpOD3Dx
Ul2DeZVxem16u5NBi2Q8Rj9egzq3S0k7p9ZW2A44LbbwjxP6DCNJ0RFhVvimFY0Pu3Xkgyon+1Yg
pBBBqcijeJG1wXyUJ4soGrJDpDnV5t6zyWDP3Ph9xD07KKCSsd0I/LKd6NRC36nAGdGUCbHo02op
iCqLHsMzPBydczQ0T6ehc2v29Dg9ebAxXrhJ8CsZJ2N3bJ0leS6X4rMrbi2h+pTgaoy4eEI0rCYH
BmY0xsJL3GnU53tdcsDGeLNPB8cCUVTNYNQDyKs5LCwSlT0YVwxkutZ/V+jpURYYN+MLUocl4T21
fZSvyFkFe0ZLbKNWWmAqPyT6/H/qpUUs/J0anhJ36f8xoiC0XEhC/dFxYDUWC2VStAOiSE588Qyo
eoo8+ZuvXRB8FnG2qmm7neOfbuVG0ORq/qe0FXrYzfaPGzuVYunzXl58yNz4p+iVSer+1KgLHhH6
z3gPwRmtHHqDpRNEX5xRBbeO6MeAhKmavksVsHHHjewue7xaueMbIc+iaPcd4WQwvUpMPIjknfvr
C0IxGdY9q+E7eOXOIhAesiFGYEGe24nghd/mJnHj3YDRth2J/VMX/hW3nv0ycv7yvkojQE+MV2PT
v+TgPYDRGtgcU2Sju7GxSmiJ3BDkRn4rD9nMBsvZ8ZJ5AnIFYXCurxD5P/1i3uPvZQ4pqBWwZeSi
fHqVze+o+IyJvAx3iXLh7rmM2/Eo/2E6X6AVd6ga1Ksj4exgv2Bl6Bzr509zO53kzl1SwmRoeAyI
V4wTEmfo0wat0MolgI4eWgnFUjzPCL7OqaVKeZj1i2x4pL4h2N7fWbdVf3k4uzq3Z9JozjAiHhvC
PHqdpu1WIdS/wk2oDpE3CfsDptN2oSV4pkbHM1Hl7v3J0VByBq/Y/wZ9bBKR2VV2fL1QRdNkgiRO
5GIwmfexFqKC4uMzTzPzPxshijIco6cK3AxERwG1RtRcovHfiXRJMzp4spUbdEDuVBxGYiqaIBFt
xNcDyFhY8zKG4AumrBk8XRLpXLmy9eFYLi4xMoyBTRwbbpFFhWwBMRcEpJGwV9HKfiEYZMnNE133
/nsS0C3VEk5F1V2Dscegbq02ak7T+Hch2JTrZlx+hdKXhLwU2hy3XgazydX9wAaCMDLPTaTFo0bp
+HqB8KFGznIBDiCUQKPQNxlx7q646bvy9sGNVCof6YnMtIaRKTyp37hu0klKLkvXMBFqLxHmIOUl
iBjF0YCoyaWnnOHX+ENI7qHSbXWekGwyF0HHVLb4JlUohkA0Qf4YbyMjy6ZvRQxfDCHW+Ayz6c65
BrMWl2BIl0Ey0jxN+AE03bfjhPMAI+9cf2bPpd17fzdPjncP+iyNB1YG2GRI/HlzSkdbuDWPEAjH
r/6ZaLjvbZH/1COqp73mtovc7KQ7resDcfFiWEQr5pS/hRl/8k5MHXIDWRAtF0dYt75aRhOUzYr7
9ZZysYE3r6o1FDD0fbrQD5yNmg/U344TxNz1xi482wTxUs+pdkbClmgJd5FvN14WFZgFA3i2mvBe
89I2DODMJzoXL3ZCqQxpNJyHS27HHnMmu1WGwiGO+4tGq0cx58grXivgiCYJHb3i2g80wwOvfshd
p2EHDEO4H+Paaj0rQ2ClLruhEFjm5TUTZBXpPIV62iqUJyvosungh+vgTR2hrzFrDAWVZZ0XlDAL
XaywWwPQPO8+v58IhEG2+y0FmUymb6kfSqFwBGutPCt0Buci28zwLKlAhEy/WmeN1ibmtUjKBYAC
td/TCc/ziiOf4RWv6lawbaYpjD9eyuvSo9Z0PlEEEVHEOhfROmA6Y2PtaikZ61KShT37NQfzuWLc
XBzcajpwxrvdV+DAwhRjp9xYz+QqtMz3eiewh6rGCvWrxE2JExHequg0Ov51RJF78q5ehbCzAWPR
7LnxzjFGniTScv8aaC/a/fvND3FHtNnSy8PknHFw/cyqUN9EzJoag9fZFbfMwiyEVrXx7sWzuwMN
x9PPX0Z7askicaGlH5J9uHI77jaDF48RKelIS0r6fC4y1KRhvq02fhvdli9S7OCcDcJa6308odXR
uZRq5N5HxVOP0e5Y6d1oyf+nEVvD9b3egoyrRDTy29anK4NK8SkB9M9T1tc3479IeAYH0wLvXAzS
buRdFhmFJNAoFadGETp36TYLhFLG2T4MyfB6HO/kf+jrKW4MhLcsZlZXvTc/CNTO/2wLBF+ZfUMA
7JVp3bM2oGAcodn4C39k+IaU6IZ09m0lYXLZNEKyXtGGBsAv5yVGK5Ml/bG0ED6RyM89UzIYM4QI
+/xEixr2rRKqM1DlWd+23LvPSmDpsXeuZZX8ryVsgDQoPQ3VLaBaO3Le2V3ED6A1gsCz3pEocb7u
JJF/yxsIz4EmdrceQnJhYe0xGQLiKRxymtKNJY4AIyfW6DWsLMPP/Y9uMypwPHqn1OnL65NRsv5m
ZavQWCYVIA/9b19kB4zHvfUXlCRHgDWjovfLS4lRwFF3jrDnRlSiEVU8I+Ce1hlBXuyw+2gQQjml
GJhbjqcpEJq22ahJnWCzOKqYCYAIjbGgjD3B5R5SAU98Cxp9PhNK627PYQ2GBNpy84kqebcMS3n8
js7vBib2/dedZWxc+WjStcbnwERWshMic5AAWeEkCqUaIrBj9d6navJlOZQTNSlarGezlGekymuC
V9lh8cN44qEOGy+f6ls+qzq0JFsvo/KjNcBq8NSf9VkiSn6EMtGdE2YFxY6Se+w4gm74ZV0+0XcM
nuTIq9wfEnxiV5GGnUEOQiySTnEFTuPCT9Ybcdxm/8nSDpTyLwk0ld+bKcHlhUiYqOObNT5ziDEZ
jGFXbDs5OSj/H7nl8V9t2Y/eHmise65mP5mqn0PbovBFVmMuBQFj36WwMazNKx4huJYRvAhoPw4c
NTIbLZsWtnpUtayCZfrdaUAcxML6P62e6gJBJXgVNC+CXkhLSZzXr+Atu0DtmyrFVmc+MZldDgr6
Py5kx7K01aaADd2FEloTbASfv17yN+lK5gaI90vPOShgs+ZQcHFovN74bnSGsgtU1w2MumMyPIXw
r/zz7U4X/OOaURX0eibJ5KSWgAIkMvcMAjhbiSTjyHTYGZbX/yNDrZheRnit7fB7vEPbTLDnRFYy
p0lpyq6dcon9u6Zzai/p4BWZRKbpv3luodfab/uK3k6HSSqQaJQ8zSCh0TnQ5r5zgBUTuE/ZTwhK
W+RwcEwxJFQ/7dJKgpCTBUYpBmnfcwXKCK5c7ucTP7B5UUVW3NJWiAiD9RgplBxYt4nAEtuPwF7y
ILBJRnwA8nlkpV8T5XBjd07VaBsHaBkBBYHwxSPk/bH+IvsGZqXi+ur2Pj9kBrTgsCQKlqnjNKQT
WxuX30g83K41CElta8xu3VDs+fwGvGF3MovnkQiT+9FC+nEnOwRVtXzNeAOe/moS8SEPiJjsRLf5
242jByTJWRD+iLP5sP+CdP/DdzTUZMMuk9Gqkb13W70L6kZq5XV5m5uipDmt5Qms5/d5I7kisUiX
rqITU45kPZ7JAp7E/QnK+4h12Xmh2uq1X7RTE+XVPa0iO6sv3kM38GlYyyI89M49IqVbxevfGto6
wAHj7f5Guu2B+MYMkMpX+1Yc1h7o6sAvWuKPvqwxWxrRRq8QadTVwUz4lqLyZgykANwKo4WACuFu
MfKuHmxNW3wZtnpCd0RSAltz8fTCOzmsg+L6tQWiZpDdeNSL8NYA7+j1x5Q13y9Q491ehzpwQGQR
5p51KLug2rTLRkRzAm4cBjWSX9OzFnQRxUfv+Xp6qJuz05DZlQ21/mR8kQ6yHlYDPrwdv8lacC6d
ejM3hRY36uUjBfaaJAF+911YnyRj47NcQ+V+NwVuYEAXoQi/6PAuhwldqNpuxzzQF9DgGQSfbfoB
lyCQtJAe8bRApyd20GWlkC+Ocj7tTIsTfeGn0rFk7MpgEO2Xt6yVIO7erTJbe1sKE9NzuqPVvg+u
j7F61ZRRxEbC7AGkm8GsHtOgsrfJHJdB2zbONFRAKxgYmiWfTjkjlUK9+hffOQ+bNVzaRHc6is4q
BltvCnrvqTZ1isQseHJ0RcvevvbqEJYN1jfjr6ZEuyop1NfVVr0Gb0tvoOxy0fE4Gn4d+WR5jgA+
wW33HLIywTcJMugfzVaciIPNHc/TWCKROfwCMyYLAnXZO8wx6CAk/NlNxyjyLp6ed5sIp8zI0mCq
uE+cVYt/5fgV5iw2lnMQP6PoLyZFmu32Ij2JVuH+K5j6Z2RES/nh9r1Ph/PorpLLBAqvQyo92Pv4
FuBkZjcDdxw1p8cMMs39niKY7CnQpETsbf9Uelo0aJGkFJMKZrpof64m4D/nWBcSjWWVA98iLAjn
kK64XEOGla8QIZfsxItk+S9wubQLtm671EZS5SZeffqfK22D0WxCPyz/qleBVP6Ij9ntY0FidzH7
TeuHGF0THsFSz381C8VPCX9vtIQT6E26p0oNnYlFX5A8Sghe/pAvQYOPUblNQ9FvUPUyMBlYqWHH
xbxUeGq/EQfq9/Cuu8JTiJvque4ty5DWQwuIo3/9oW5aQ77MfPKrDfA8Wb3tCxK/W3x78SScUw3r
YPUqTTfeLggdSe/x/ANahH/HwY8RJ+WDhfWbrsiCo6/nlBQJGNeL11Q33SS27bFCq6XGaF04Od9v
YxqTPRGLyhuvf/p7COvqIYRSF4NFAwdpV5/8kcBhDvI3UAdEEDK0MtUznpprtdBS26FcF9uFIW0z
OfArrDgDyvYFlzW13zGws0tb/qMzk7GIaNKVMffOgogn9yBNxrxG+emkHg4cjQMB2If5Yz/vIst8
0cIZOFtOXwBvbnC7Ynw5jZKQwsm6kx8eFzInh3r/uJReFsMbl5Lb1wAM30ANkKG3ALbtLoGiNw4X
Yn9acLOO4ztfyEHkAwjveY0wqaXd3dj+pab9UFVXKy2zYEz2ziwIubQb0Ko7tDukUH84OB5pvKBj
0FubEoYZ306QbdUeyEt//SxgxVjcdi75wPfzVopny8l/OeRSTlJZfhpyVYilsk2n81TlT9j+bbV+
wA+BfS2+305/qihOYw6PWeuiankwPNt8D1++Kq2orf9IgLqDOBhDJpVoA0oNSypZ6b3sTAAXM6YJ
mVy4fglxIm92E/zQ/ZjUaMovvmWVf88hThaq5HwA4nyiPXLyEU6AYvYkyQFKEss90TalWhf/GVMs
IR5VJobDbo5oZ2wLWC9uaBBITxtywSHAHlECVBq7JfWizJ3iKzpmSShkCnu2hvTjyU+Dc4WaHgPc
6rx1W/ttIUFzERr4+DzB46W0Be6i5C5CZJpPMPON0uZ3TS35QIug6sQu/MbdOqBiMzID5iNiBnmp
B8QB7Sz7Hk1ygJbfqU9QOsh4Q4qXEgqRy/d3dcURnIotWy7arUmkXqHGX4MOdURLhGieoBcy/ckH
zMUCFy+/3ChqNYdH5qQCB+5Xuv0JTHKLmYykZWiK+OyDdd/daPn/lBebQH7uiRiz5QxP3ud/4vWu
Rgbw5173Nm8TPkrD1UApNFqSpu4ylGSRLgQ6M7GWOdPYPCHzSEGxjw5tNGb0YxmXU40ZaA6XTAKL
ZAG5yBd6bm6R5p8ZCZI2WzzULNoyILFBvaIzIFTBXFaw0gVZCF9itoJjbgbOfeFG6lI8uiE2lvDo
QSQNhhCbalr93xLVQ4t7qKP7/BSjcPWPnOAggG0fo/rIAToUotb8Jhk6XHcOaRkd8LAjJeggvmXi
RydytcJljeWzEGLcZAD6qBr2evADMLNQKjTVm1O01iiKd3q9caeupMJyciSjEcBSZ0j08vljYVmk
b8meel4jTLU81de2spqPwoicqKNtQFiF6TN2m8fgchLXvyDmPAOZ013eBL4xPK7tIMC/wgWgllcf
yhGQEp3FPelYfBLRsZL5EOlJjI9QZPIW58g9ZGBeDcQtmQCdJbuv3dC/jYQnfO2Y+5qzqBw8qmBV
OekyZ5O6i5ssBIpdMinx44q60eQMSGK00pwH74SOWBVlsyA6tpPrzWj6tuGvFusOY6itR3eq2fOX
p9tfwI8taOgC9VQVsYd4AZmXB4O5yXonwpKIYZovAGrED2yAkT0BXROSDWsP8LU/KF7CPl0sh7pK
cWlaKintYQWBVq67HZyEwdGN5fOZCqu8j46DSJZb37h+qHH9Ipu4snzyVdMvBWYwKGT1GJBdRUxp
jTBt/l+NFaqAasbdy4fTw9/3743avjMnBRKorc+NbAbz1nb2YkvaNAa05o0U/upH9hk2XjuV83eQ
KXfiRFoxHM8MnPOet2bZLhPHtkiK4rAbZiTx44b6M9iWR9PDunRWvoIlSDSG+WXmqiqLG1dtdjbD
vPT7g9Ep0cFpDbqTIFY483XJKPsrB/4xy8tNuBCzxsZEcQP3Uu/jrN7Hiem3bCiboQ853Vdasti9
Mb/Tugy7dvHyLT1g/nM4jdJSstLe4fL3YRI9a2DG6dU6S9Lq5mYmlrtsUzEMppcWdzGZJFhPagmO
/4g/3nZqoFURJHAJMpNeoAMQatP4cauk0zL1gthQZsqMHIrZPjZgiDw0oLJkLSTCgoTbi2qEAwM2
XEJtgqRfxYOH14aYHE+O+4V2zG6f35OkkApPWNfA1DsndIyzSO/E2zsBNrDhZ4sYkplsiUiiONXJ
1Ma0ujjJpZ4d6FaGhXD02Uy+KM7tVM1Q4i+SqUB7xGRPxIVziLiv28vGIXayQxI1aRu5aMNA57fC
gKyuqm0qxrGVYiTjPt4IGTvQWczL/ZM30/dwt6j+sioUYr7mrjwMkiIKt+5tWyxF8CD217ig9uP3
TSMUv8NO2o7kS71s96J5oD9nK2O3CV+7ouOV31OkkR3sUosMPiXx49TS5Bq/h+iuHLfPVaOlyNHb
X41yYZQYI7007vlOZ0Q120H0p1XahsinwMOOVILUYwQzZ6ZHoUH1lat3v1qmfABPbmr9c3Lk1HOL
Y52aTn3UKbZWuqNgk3mYhhmChjHZM+Sbyp1QF8vvZbomDnvRgN3RxCT6jAIgOG8gXcTuvzx0LW8C
4E+f66lB/XvdbU9ZfESzuZMnzGhQQOszl2GB0GhAkeJX6bTSMb4vcZT+O3FFPRN3zPXMQ9mvwWxJ
9bgWEGiv9Ei3igqUf8hjta8o/0ZOcHXQr4+ZwCg2ZHVYNBFRegHjprLuUS/7UihkVIGeBuLYkOLi
o/naw8a8k1iqaDVa6XNOu8A1Ge/3yNxIzY2FT0sIEdAnyr7p4mRPWoVYMF60B3T54dYAXNrHeKS9
dUYIDqOrAbz+cXkwJPSRBY33S3jYnk/FHXehCRFu1x5hvcCUUqURyZTXrN2PUS7/KOyJDkNWM0mq
UqEi0CFdP+CB4ge4QlLUcEsinP+yGRKmn1Y/k5NITplFRx5dWLTKDsxuWUL0r+yoz8M0zPAK0Cch
q9cFSAFVQDNNMmPBTX9VsTjOt0MtElNMr1bmnoj33SUea7n6MsibqmnI5hou+H4JkKWL16DBIho4
DUduanU4viPlV0IqtpZVSJ/goSvkFr78D8b/zn+wtb6jw9Sr4GvxOmu6RkCiYF/HmPZ0PAHEfrAt
XUdTSOsfMdr0MocQm1EJIWacG1Uy9AR5uOFoq0IWCY/RpuxNBdQMB5N/3X8uE90dW7B8yNewRlvF
B4prSTic97hahVqnjj7WfagIl1AoZjAEzLMEtuM9lDFxf6RdTWx3f082OF17QBXaztNkw057iJdn
vdTGbeQHUdMhbi8sVGEo4w6jpH+5ypbR4noEcDkFUuC83GJBGY4oqZhvIvmnbG5Wd4Fu5SQgKqXO
jZMHFO3suAlBQPSI/OeoPFSYdOFGESrEw7oyI1eZLUTnYdJiiy6NNXn8GfBkjOGtebiOKCX7usO6
NG6r98kxCxkExkSmzdA97NKVmcaYGNfYlzwC4XjAAlYuVw6Z60PFI1Q1SacYbraZA6XGtbl7Kl8J
0oF8zdZt+7i0s0PLiUYvSMpFFk6CdmCKIR3DsNm9db5vI2G0GxGaDR4oomHSUeLoHQV8RwJB9i4v
+Tqoz33va/z3KIwx6d+g8/UKYxTli5bQmt+KM/+HY1ECmmAF5x/XMuXVlL6L2STUTWrkRWgK/nUN
u2qyezD9VKafJcc3hIdEayk1XdSleEJM1WQyoqa4gp/PAPK/Jf2L+bJpEvb32CTLXy49J9R0nc5o
/PE1s4rH/7ws/EpjpoYoG/QO8YUfFWel4eh3A/k8YL2It2pU1E4/oxCJvjqEQkn1PnuTvwSzMjB7
BOJUN1ajg573XXzCGluwXHG0GHCH0HnYPkKvQoQJYrNy/Cgmf+LUB1saaHRjQ+CDVvJPG/RmH5yT
/lzWeo2dn6EGg4GpuHu/f1fcN0o8Nimw7KqhvvBVzMEElakUDCaDD1R3C54CrwWxvTn9QZOk2O5k
qx1pKDGVOIdfvHu0OOqe36llNvq3BY0kP99iaEHNCA5qISYIcJTGQj2RRHU9U1ENAIZNBObNtMhA
NmyJd9iiQx7RKf4j8eFTlwHLP6ov3zd7wg8p64QIa3kcW+vDoOp4l1CEO+pR5HJbeDXLUj8ENCAk
SWohwkzVY9oolEC8HoiEsBSQdAbJ6Ic5CB4jXPRKCerZl2hAyxcMqyASl1C9udDC3c2s5o0J2oZ1
ExMGXGnaK62yDWRp0IlSV1hVX6M+pWugajF619/N9u7JFkKeRJNiSLyY8/TW+8UzT/Ipfe+dVO51
jTXJ/LsuabjVHmXntCg3QEasGAwNcpsWW8fUaXXHYGq1/dvmvv/wcG0qP9zr6G5R6AOyJ3q1wlu2
6hSn61ZXKsmKVJzllKkHl0jyshXGV58Jq5e/Uw9qdwYRghMsCqDxIOyX7+oczzX82Y2aVcj+9ltN
FZ/3jGYSZCE1NWBjMMyqZ/o9f5m9Rhuw/eoJENq0XuF8qclrHJ4Wysd9ybPBovorE+rbC6GtaGmv
4uiiFg3jPI6xFUZZE1fir2esY00kd1pll0O3dPlnjOOei69WcG8jughg6UqPYIzGer3vE7ZV/deS
xR2mpAjkk1OgqZIuVXMZE3NV6uX+3R60uxBxtL/OQTCEUyt73zFMKElW74D/rFkfImT+Y7OqVhzv
NVDfeU6IkNk1T8pxnumydD2/+BJjJu8E2P0O3KQZ4XG9FStuj2LHGA1bZEOtWhYu/VJtF9uTw6wG
WTr1dzKU+KWUEFcOsMIMgqXjqxzMkRWjLtfLgstUuPTPrTCfO4jxsi4mY+BBPv4wIRyqIY7WR7lF
7+HY8xECEUvJa7JlXsCta9RgVPSYzYKqdzNwq08BkQWTPEq/RhUgDArUyBubY3ep6kKYXN1EmSPS
iXBaf0qz9aTOk+qr242xQVp+IIrUbf+NfvEJ6BmXysHZvUBl0dI//FmP+7SQZK9MxqL/WcOshCxm
aR4wGBthYQ5zMUegAm7BQCKiUuT56Ik8VasBO0PIK5HEMK7YmslbeatGShWB5StrXZjPdqAVemNA
fSKo3h9y7IfJB6kDwbomQ15pUCyn4Jep3Mb10m38qCddFhkNmFFeK2zJ88F1vT97I3Ym3RpMN+7Y
clwWoqEbFCgMXFGcp+4hK/gnA4xTomEg8hPLIUMN06zksVccl/6l0A5JBzSbeSewuqGPGUnh4Tu0
tnFKpTL+zlqFjyWy4FnCLFFA/L+uP/0g5+9ebCU9RmsecfwgQBYTTCYQG6BHtls8uYV6T3iduq58
FbVGLIJwh/Bwe5lwFxuyFOb7AmzAgPpDzB34oH0XjvsEtDLM3HZM6KnNX7YEh2d9Lq58vLTAvLnY
ie3CgkJae8NCsAZPvbQ3CQh06QjNG8z2ehPog96Tz1caodVs4Ag4Ssosy2kPw/whP0iddwjUKJPc
iWJhnd/ObryNEegVfSEJ+X20LHS7UucK9xNbsArnANBIzbLofR9qdTBdmh4VXYPa76CQkNt2gIng
mh6eF+MeKKeLAVLceGq4qq3GJj09conU/T6izEybXtQxKM/PIDJThfHXT2kpean8KzJmOkkIn2gn
G4bfW8u8LELuvt0cgV0vWQ87DfGzAhBH4IMPOTamlUCmtjpWajjMTkJyNcF8kisqw63tsT8uPiNt
g2Ou3CI1hYr8VFPwQeJA/Jufd0oI0MLsnQUm1SSwo58rNuhJ9IUcEDjz5LX2wsdNtzMqU35AbTxK
atcDreDLzV9IaY4b7HijSb5Gzh39JTZRVkVGExiRu4azgeXwean7pFPRMJ9WN3ij7QPU/zSAnR3u
/pTOlWzioCTkwkWNDq9Za0D/EOF3PENXTWPHr7IDVVsQ8rOimH/o6YjNK4bT8DGRMGdpS5VZ8GF3
Yk6AWKaohrIia+xKl0R2BosWDzeULhl1Txwvy9VL4Ez9p616/STk6A3cJL4IgPGRZpz5r/CUBeKR
m6UOqdW5IDZM9zwA6WYi0eyBKBqjO9X+T9mZ+j+ZnRaL0grl3j+QwMEDDEdpNLDZCRj66d4BGMHy
q9wmKCovdgQCyLOq3bxKTqp+IcM9FdeU2szbRIPRTDkHnizRcalX73pemtcgM6lIXMDZivYCbDoq
dLjQwzFPPk1KosJax4E2a9cFQ31KJ/GTrcQMEqVoGlV85n4K8oo3QzdjY7g5Mzk8VHIy+ZR7Kuse
Cb7ttKIUIvwlaw8jkvysMwCmT1tx+Ryj32nCnJwcFV5aSKpVx+x22qzXtBj8AmkxZy+zcPIMODAH
GEOvf1MA79910yUpk+kjpZ0RROZ1q3quP2EWXTZR7L7eGQ3IDdg8RGfCc/l5pwV3knLoP4TJm3gL
GHTgbIfJeFuo0lryFg9STMxbqiVCHf3/oXQLx1qkJE2W3QHy+HP9JRq3XtB5VkvJWlON6uMhuS8r
ygbwlCSt1+Em6PxaC7AG6sBofEmsS3o6h5XSTayfz+oqLfu6KJfqUqs1Qb+htSu1odz1ikXGXczs
sJUtLy0dqjI1q2+J6uAZwPytNJr4KFg9g/Rp2iGlyZWM6tuhgbN7D+lhDtoTCX1ZmCQFZ8XqyFqm
4IHB0HwylkL4m2aiq4cAUuVs8C1cjjCWbycZWYVlEob9T4oEUJY9v83F/YFyeS7thxOh4C5LC2aA
HRk70Sks5CmOD0I+KlYZiUkUuPqXaiuNpkCQDTaCgZrWlLIBEqNT8/3+l6v1o++Q98+kOyHHVXtR
2Dqrxnfk7bUZfKDNqf0l6jwzoV8af4jQ3LPQjng72IYlk3VGMuibVosthj9qfXB5OVBt9rFrtljO
l0n6aViiNFLMqtyzWjq/Jvp/uu0LHSTvCsACn6OrUvbw0O0HsUvMFHl0TMrsFIS+jsWOvPpd5cE1
36rnGcs65Bl6jaezCXjhlQfDjmxZ0K5N8dUJY2gIhqHvomaBQaYquHwSldRanQ7/XSfWmHWTpyJy
8RO0rOk7fVe6eGayH6OFHzS0pHaSNZeiwmOZRcNV4DeJ6OwoCtVqdAPNmDIHQvNhJOBjMiMxBX3+
ekkOIVoy+P+mvd7VhzW50dHzoQRIo8P/dJ8BGkhwt6JYW7oFA57LAy4Ad+ePCZdhMQ6+DY7L96C2
/bkGp9XGOrVSMUoI+PXpG9qm1VOLAkF4WlrGw+gMw64/bqTeYxxBTDh6Fb7ZjMJyta1ZgEigpyey
0luRGysZ8z7nyal1SvvavftblJCo0Iz2G+uoYuGVLwszistZ8raWi2sgRZjC6NyomSZb517cGR/K
S6HogmImB1WqEhlZgyAPlFB+rlngIpVeBc5kXqb0GDzOHxt57LFzDG7FfnYWcrnRlZRYAaoqwSET
5PPBbmuxARtFHFPCrThGL6j1lRoH1iIhGaOurEvEnrO5b4tuNtIlHHzrQ3A0Y7D0udcNdJY9mn/I
2QXtMr7kJjbJ4AUeK+4wZuAUdMAy/b6Jp4zlw8tx00GqWiculY/Uiart5Hnj6ADw29tVlWNNKFmX
NUCoMWXEB+HoIaE5ULRA0KEdTxj/waFz37BinMeUEguhPyPJpA/RNC3trTUKOnRqTf8R6HIAO+cM
f35s8DS/ZQMT/PLlA/fIMcfxR651Q5xPmJkgiikAK2zVJDmTLChTzVmbpKfO46wih4Re7bteTL+g
ErCc5vh9Ts8UkCzDSV5B5PWmqiLhJtb/2zLw9kEi/7qieBEWAkx1BgiSmoTLXHh/c/5rwi1IgN7J
nRXxwL6HBGTnjcZnmZs6GkvyAD3Nkwgafh20dKfkWbnx1QRvPhCD0+AamGtskzm56R+5zHvVDI8i
eLIcw2NOLAY8V1UcaQw3FM7S+t7JxFuHxXJ4aUXslrv5SB0mkRJkgj+D2+A6/CJ8vAVh0maOc6i1
5d2N6e5yFn8pSCl1K4IzGR6d9SPIwCTqH4Muiz/eogUvylnSCAHun660eVGSJxCldEzB4W/CXh8A
m/rhHYxF0zwstup3j6OF9ajJzPLM46/NWQZ7+L8TopVXQqJMfsJxMjeQYvSZTHeQOrVRoC1SWWQY
tq14oBohV08EH6pCKMaPJKlRHR+0Pxi1qD0C2W5lxrPfBrgpe18kWNHDM/WJytJQQy3o82RU7llJ
G+CexBQu2zf7wGno5dBNea2iDtUdsP+R9/E9LMHwEQS7DaSyuTS1iTb+krc44fAWEXDb283O0FVP
mmQQiDn3PtAvTP1/6D8TuW26mQE8UiC5C+dVxgK6YUPuWhv/zvrsNKxWCrljylMW3kDEgjILQwse
Lrb4vjN1eZIolCKhbRqbg2fDmSxPVYF5zN3bLYtKmYw8A/5PCjsq/6aQjXjh7dihkVW23yBAS1AD
DwJt+9UDHPgghQa6ewif3wvTFxyvYkGjE7ZfvptCvmL1cct4ujrgu52j1OHQruvBYH3NdsaXVrlY
g0fDrPv0sl/VMpTm3+8jSNEpv9wkVVKo4T0XzBvPURhia19cDHkocu1OvShzSCMPqPzCHsSPSjOQ
+2IFmUaDXtSs7A/kYisios1SKfNcxABnbi/mDVvJeQ1/hHWjj+OULnGL2kcI1l9E6FgIfsrGXox/
ET9tHuRazsyeB/zfyYDbsbmZ06p+gDx6mFuUnwAjMT3QtlEE3rjxa+j8kbIvaZaXMIBd75aXno4D
7WKqSNdOC6OyEqyorVNibNSWpYtPlDLN+HybOMQ585pk8ZedYQtFzr1sf3FMbOZ4+7XHLlqi8QoT
ObHDknZuEbnabD324KcBVYScKlc6ni7Envr2b7jwb4kx0dC/Y8/xffxDpM4cmgV7FE0pRpYrqe1V
1u0KhUrSwWERurhFkuizuFMO34iVORsVxGyJIPdtACSg2Oggi6Vs9JOW9KYAqkZTqWAfPz0MRVgk
ODHgJ8X3Mu9OJB3LOMbqaXu8WCQ2B9Zi8dAYqGjnke9BLiFn1FByzYtqPNQLdL+p6c1N0Xe5J6jR
hnh/xd9OF8Cm+TfKVfhtdldnlZ18njrGxUIhtOP9PwYu/YamDkjQogcyhRDqayqwRa70o2LGJtpB
ITBmRhtbMlztobRekSGTdLcE10qhSlVhyeo/ieKQ99QzrUDJoMQiXIoHgBpPWNdK7hBimmbXmDFC
TV1TBBYgCaFAiMqAzZ2RmcRW9qx/JonP6QKfscOudmwYKxe3uw1PXunTOB2k1Us+dGw9lBW8KZdW
v6+SsX3v7RpE0L9KRPsYxaJOhdbwfU1vu7HT/5+Q++3M1J43+Um7rrujI6pvnLh/t2rsFBCs8hlS
1tL52jaHAEM5BAL0RQkka4KwQbQniEodp4/k6vxvLCKeFjx9OMKdMP2mJMgcWElJTFR/1raezXBS
ftewcty7b1tKGUrGe+HmbDQWpKUpWrbXA/6hhwyWJIb5T4IEvy8PP6Uu/jPclyK6/ZkRsueVKP3Z
eX5JTiKlKike5EBQ6qrSnumXeJ6wMPjPN79SqqZMPlmY5JIqXDttgiMvR7NXzPk/IKiTMTz2znrS
ctffx6oUByV1lNbI8Ukz1knMWIlOSPsQKorr745HJl6lTUSqNVKV3I5AtZGL+rBxC3Izp1nH7hHV
ucIWtIUa/YIyZ6sQsSKmdartBjU7gP+guMPi3r7La0HHZWpGwIw/Q/1p/5XVOqLL3PVLbJmXz6Mu
tuT1bxrP3eLD2HZP02q/Om4+dnAdOdxY8gygk4JddKp7YaATPG5RPAGjzVnzODxK64C2VUQyqdqx
tZR2lxcUk4J8kV967VtMb3Kx3B1Rt0N3TP+eOjchrr9qztoRZgD+xhuwKdq9SbYDqjBoZ8LPtwLV
nkJexvvnHAs+0g6n3EYICnhrQJim+z85Da3/oRWpMNRE/Xztn2h9ZhBmfRx1CCzA/ZTMdcg+eXx3
B+heXgu22Esbjrcd0pvu8InLHvCdWOvfRLT/ojDWMs7EBIAgM14eA7uMWrwWPVDZI1ZaewIeV96u
xAbd28VfmYpKQ66C+l8VAaGcnnmfTkKUVSVo6SNXg/iPvPkMBevKpc4yrkrG5p0A9Yp+9nIbPm1k
C24Gmcnvf3SfYZn+LXBRRGF0eandsJbR81lJIQ6J9RCVssjDW3hVNVz0SwhB/vCuztTBydxyjH1R
XFKklsDuTPURxFbtbFeytFhu9qAu7NZPQgr5bprS/P2fTgSWQbfB/Dv4Kpxq3CEMzTUrbMf0nYtd
cg7ut22G+6REjxmQ+6dWqk76t08SnzQyPYacyj3kWU1pcbvaONH+Tn+m8I/+A6V8Es3DvYhD9wui
Kcbcx64I36FRNvZBLE2vAgHKr0zt4tZquGSjdEyhN1euGJIdW9fuYJkRp2VvaqgRLMAOKCcIEsD/
l38lOhMzLdCKCxl+MDcusDDMLglz6ILj2y9AFdhfitrLoae/DSATXfHs7Wmn1qTvVinfaBd8CE3W
H29slOHHN3zX3zAO70zqrFazn43jv2jNWiv12KNT9eY0RKviM6C7v/R1CFxMxqWguK0VWd5NXcgb
msrFdegHqTSxGOhlaqOL4ymqT2YPnG9sNtrr7MpcZyb5fMrgqe+7Icv6cwcgqfBul/a9ElRs2aW+
oMHiP3gtVw+Vgi8WaunfZ9u+/FwXsieqtZnsiw8ctlMvMbFkp/pKD9y+PluENK5KooOsZSL7dR6X
LO8cnZxrQzZo0MNgkz9HUO5uMydulvI3soFFKZFK9NAq28ZG+P7RR4MNhkTZHAHYNSh8Eu/lOw3a
eKAmikO4jaXoAtu2ol8p8pICf1+l934Lsai+wpyU0x01omjHqGtJGLioPMwRVVDh24Q32LD7G8zn
6LUsRsqsIJgLIMOY0sOLqgOI43gxEjdGXGtzb6HmZG5/bC+AGagqLfbHUl9fTFuN6vi1VdP8dr6U
08N7MkUmKXiRNEFwi94h63Rfdu4mlbg9guqOzeS0Bjbn9vzOBliNQKpSLTskcVQb3xTltXBqkvLI
VwWy4X0U0k2CVb2A3uFHBxJvuOlvOvuJDZBbG85tuEA7Q84frVW6LVGZhp6DQWW5XMG0xUeNj7Ph
lM5TIQ8dn5QLK6M7bhefbkvRr41u0uLZg6iIqZ/OlUEAJqcDDOaFzymsLQWKEQyR6xOoaDyZNzHd
A0lBrGb/Di6LaZPHvM6q38ukA3RXhi8lYxgUDFyRxDtBUp0/ooptufujYWijgKiC0s7gLrR0jjtz
8wWjdzGXYwT56NAUoNlI0ZdqWwMBcL7c7S8mSURYuhXtOR3bwQ0ttgMZs2VLxByp02r1IfZR7+Jc
LIcxoZmWCDBlmEbRw82qFv785KicJvO8sVl06fFTVlGF1mj3dn5fEmcFWq0kVC/Qbmuya/jx7+lv
JD1yr2+v8rr/y0eDHAFKUchh9Shx9+rjn2FQT+sRaHmF86jRMWvpXjytSc3PmEA8NT/FKH8pWBHi
Xbeb9DDXVLjm1b18QIqfiB0A2CBTKPtj5MMl5kABrEbuKxoYw2lTnRunzyHFHcZs5Hua3iEK3DCM
qxDKndjK0pUiUbUYIoePiyY7llg1li+pJOzKrN9l/g+gGqNeUF31+xF1BsaO82M6d/gqtZfTk2+H
oJjLq0NVE/WTzgNEPpfTeKLmRmmPJ/0WnoVF7r2feJhfk8CAMwT1h6ot/+ReLR8bGot4BSbbVOQp
2EY5YC/LNjM5/WRF1fNabmqFEiFbSg2G4wEi65I9L4MngmoTWBbtlc5wSIq7fBOVECvBtMjg0d1l
HaA/POeoC2PsS8N8f9gARKMb9ErLHBBSDfl85+yF17zKFKbppvFa8QE3QGS5ravfetcOR+Cg6zdE
n/92qjO1V3+WTbVunxEQ87c26tRt9EVOXchoOXhzxEWAEy7Ha9EXa6NEFcf4syrmUJEfApBm9YVu
GD6HlFlkbr4uanGEbuHoTOiNKxdXoD5X+wsc8t5pShDxPHNZb9REW95gRaavHAIiIprHZBVfDEcN
gEZltZ3mFTRWeVD0ENRvmmC8hKkhUnXK/nQsy0ikILGDhgTQ2ZvkM/8U/vXex+Stc7vdbuF94L8H
ACNqc7w5MSoemNt61fPZy+v67smr/ELr0c9ncjfBK7rPELwDp8kKorXZc6BkIgaV8X35voeWuDg4
XEmasWPk0v5xoaCzECBa+hM6U7Oq+B79bFzn3RRQ117dGhW4wFfhkVzLS6DBlHb+IBbP2IBWq0gv
oma9sU0y9P4rOKXuetOKHIgVpdtlogFQrf6THkhDaVICqDMD4avwThEuynQNl92dSCC7ZrTPmxWy
PlQAQB+HSvtKmc+LDmo6lZhf8ZB05YgomCZhRfwXgPxC3JT3PjwzMyzd5RdlQvqDIxFpVfoWUujo
397zWiYWuPIIpGJNvdQvEK+WfXTTqImSeoeus/Y/7zd+UYfoYMqk5vdfeRd+fzqAGhXh8hBnSa3D
h3Euv0AvuiAjV9ACVjU+ckv3zefecSWhuCryzQxBrcZQ8LBCRyucCB6L1Pdji5lR+oTe3SRUlGJo
Lhq31G62xWsKaSGkEtdbEgiRO0FjG5dRUUU5PvtHU/a3We2YnftLL5oouAcjKOB2vIE0U3rkHRXL
bE/ikVWGxnt1Xvzb7Vjy1USvw7r5c+h4GCPNh2V+MV49JxNruiyHW7w//Gy3gm7/bPkY3gZmha5g
sdN0WedrBsVK+G2fsmMn2k7dSSJv6dMchak/ul45kJD3IbIWJtAlSRNyPsS0pE4fFzUTX94r5U5N
cxkGLe8/PfZPp8+j0Q06AK5veJlF55wod1GidEuE+ig7tapM0ciatFU/oPYgQbGGKrYEW/6irjrK
MWF5gy5zvOR6VVqLWlkK7f1x2A4Ry5YdaRgW7/f9FYdXJVop4NYWhytVno9S/rNMldAU8UZQfBKR
mxyJMMvW58ESb/rFc/eTbYCGs5V+jthOybpR4qhwqu+qGGNIxdubv2OZjY7TQTpsjuVdEmKJmQVk
gZBCH8ZMykHzk0sUm4e8zmgnnnEaaIaV/DwLGTf67EW7qs8svAYZJsiPxStekQ8qk1IEKVGGAfii
zidvksAlicru+dFCWiB5n7qhveffRlnnDImk8QFZHqTa+5lrTDWlIG8EpcvtJxxTnKZIfBTNnut2
2zXX5XSwcbaJTDjr1XcD0Al6Uiyqo/JeNjnCnX7IdOgjSpJg6Gh6HZlPxGQKNB7SyM7MZyZ19wa2
4VzhvJiCaZ7UY3EU+DM27p8gj2suGU+stAv1YE3rQX6EkNmHwlnmagxg7MuzxM63XMUEMnqbKrZD
eYvsed1HKiY1L52c4B/PlGBT3aK9dbF9O7NGee7MXjhZ8E6GjwkP+1ijVCvWvLFt8ZvNLVSXAWMz
Mm+vBk6nDfcqlVle8JZmvaZowxZoDR62W9X41+Gk9yPXzpeAQJq1tqyOvv5+Up5oFHdnk6hNZcTM
rdAGNlu1rforQYXyv4Qfbv/R0JuW85sILBbPAor4xVLQ29BZKsxTfSZ+gkiH2FYMwM04CRkMOMop
jaoeJRSc7pQt0FSj3BBfioDtbCtw9R49ZUKwyctivHVGQhAwmKDoQsYmJ03qekBxzthPK9hPmCSE
sjRPylFlQ5jwtLiAOENuzbA3DBOhRXA9XgdfetOhowSd1GL1mRdn1hW68OZ8J53WGg59pO8SO+OQ
3vA3bmWuTJfiWCbe4+XfWIK9hQlQ0PobjJ3sVA735YdV5ecoXIBXCrnhBzA/YViuYLi/pwBEi5T6
VuwproHzVVc6iG1myOEnSzjk7USDufTYTeEF6clANPdOa/P43qWQvTT9++ElNt/uFE3oEIvSzHeo
A5VU4Xqts2jSsoJdEuZZWmMxo40Z5zIPgn8NbhDeVhapHvsUa7Aq4zQenwPuPV6/1fr9PRpe9O7R
yC7xVlP25M4d2SRziRnzOmbYsH4TAGph/WSKhPo5BGAZ+IT9/MN8HUcjHqAgV8/MleLwdw0Pxvp6
A+zKT/fnXm8xru4m9Rd3l0/9kCJMJvnU/KtGirHqnka9dpUfT3sWkwwGQ6sogffhayjqln5ZCSu1
ZaWF5qy3kQFB0bwjxflhqQpB7RjMRdMnXakUfButTgIEiJ0WSunl40sro72aut+PBPNH3zYcnRWp
QRBKg1pgxGf7FW2D33Eo7obCywBglifqHWS9eN2mcqZiuoslDP0XPzHtcBpurmJge9UEU+RTr7I5
8s5NjyZlyrR6U9FKi3onyR4Mf9pBxWLJIyGettOQ40YsDi1812W8/UEvabZ7Erua63g3DZAEHmHR
ObZYKCU3G05ADgm+W1xWVepspPCoKci3G3QcXmnRJfdbPBozy7fsL5+Sj+hxUA2/d/P3jEuSM9R4
NmkGZhMRvCluKKc2AkaSaqwZVWvCSLMbt8jI+zxUz21p836dW6PNFiAQwqJVM2GahM1jjRj6cmiM
wUPJCOekc81RTW2oTL8CLksmbp1w69AEbOOuEVzjQPrci+D6xeiDt4FSOOlIx87abwgVySJesc0i
+vdl2TdSnpytXHnkyQD6YBqTSEi0dbwNslB01gAES5UPOttgWHrS4q1Kb2t5WKIsMw1CcmZQKDXN
MjX0YZ1HgTP05/fcE7GU9pmu8qE7SMfOXB8DEBq3vDaInbU+bQL+ght16JFbhZ4w8iUyto674li2
C6zTL3ZrSs+051zwycgCh6bmhLdgprdW0zHS3aGBpjMC3VoimvuPygI8j7tLZ0VHeJJhezEe1B10
koXzQdpEj+ISaz87shZP3SC1l7ZtosgNXg0VqzEAVCy8q5UGmIT6ms/MyDtTxoLdBHHABMWMjl85
UjNPvb2kRRyXkuD2tLymC0OEAhfKp8rsXp4AbVTihRilHc8ngosZ8hMX/tuUn+jSyI7hpGbDyRri
cENptVC5F234CKDOEtL4gpJ/7VFZforCogWdWWMRb8JQGTXPo75bK4g5IycUUwWf1bYdfs2i+3NP
TgXJdKrae23uorh/Ei8F9hB8N07dm8IP+WfcK2gqs6ZqbaD8zgTxhzzuogpuqqNFTjjQfW77fSRI
CcYOfBjcwpEUC6iI11fXpgBW/gf82B+1INY4n+3zT7cLnTUKUGmh+P9x/vEQ6daObgKVlgsYd7sP
OlLWZPc2xdI7Zo1oPwrZkHH6iVhzzmGUXraaYm2fe4VzjmuwGixNp0MFnTngLr4wiCKVHuzsW1Z0
nX0qzbbltpZjMzvXIgfZ8QVW3SeIqgIgrFt6yEg267qHEGJVZPsenSvD8Ihh2wU0WvQNXOU2L5AH
aX6RKVR4/BQUgZ7DYAoS78ujp4X0SjI48Pz0jEv6dQAjmr6+w/wjzEyi884mFa44vUoNUBHkUVH+
rKmWQW5uCAROsLwAtpsauxhiuiIWUkkiG84iW4x2l0LNBVaiEXN2r/6WSqe14V0+clN3+PiXhOK/
i5Qv3qSqnwtux702E4qrQoTqRaHAlycof2XAK3oLG0qkf8fkyEBZNMkCp88rVwSp2eyvwesJ2B9o
T+KMcIFe3TpVda1QCZAs6BSVuj0lGhmIhdqGq++cD//jFU3b+jOy8R7XNoTu92zVf3ilhbCH15Np
ym2MXTveIRZZWWQY/YYvRVGr2kfOPalBZ/STSMchFLwYPaK6pHhg/eF8m+guj3M13UFab5NuMT2x
4h4DyBG5AIzp74hN/NOPD7VaUTxl7xpcutw/R8UAYDNNgom80K5rA0T8LcaAmU0A7jl9duOWXGuv
z3E9rCIeH6HPy6IxakCpARubv9sg906Ag8SC0pLYBNP0jGmsSDZopZFQqBBFQdpf/AaIwf93G1IV
pUA4Je2x1ILYykrSnI1pWHJg+uYOP/kPBMnDhWe6yqpLGNIk9di3suUzXhQRuZ7Wlx9EFImKI4SS
7dGNIbUgOB6k2H4NZRhPZETsq4Vq4y+TAkUHiLDz71JnQgX4AsiDCIvugopAm3jaaHOmdh65qOoM
WlYrt/IAcArXzBj/dSFL+y6eaW2LX9RbJmkz0ygtDpnIPGwvuXXKAN94vVMzYw1fGwNVcnu4ZF8t
+SKpsGF43t/WL9/XjKCveD88UWBMsaGjs1phdMvYD2qbUMSKCw7LiLaxACtZGjOXEa559io/bbK5
fuyfAn728Vb/0MzBhrkoSwLoGJV+1CgRxFqdrdM0ugZTnO9bk+ZCZx5WoLsK/YvxvZbZx3sxBMdK
m1zerwQEGV9BsovDK/54TzrsnjTnkCZagSmk8FZ1T5ZkoedDwW9eRfOt3Tpn4W2BNjU/Y4TqBeHx
gF2K+fneYp3vRTPH+6r0sjz/nDmBz9rz34XnoTgdr6Qof9VtUyseSoJgg77SXlRVT7EYFfeCJktq
XAb2Oe7Kk4B7Fj5X3vzPqTZ6Jvr4bThL4hiuDbUrr3D5aHsRluL5gJluYIlV/vGu1hUGYWHlRfOu
i2zwlkBlV4LKrvO6Rf1i0OraxohDjtpJjzJIq03ooeQL5iClEAfcHY9QZKJ8DlpY0NfAh0axhefk
Q/yI1F871nAaZDOIpHMCEyJphSgqweZ6NOASzk2Gr1h4Ov2YgRGaZFtXhSathiJl2CiOGvxSZWdR
+9bU4OW3Jeq4paRiWkJGqA4BcNaz0x9DEdlTDxMqkGK9uCmXYlqScR/FgZ+WJRynCgPTIlyU+Vzq
wnSL8ND2x6mOX5F0V+OcDIgj5a0TPkKDQCVzFUryAd4jWEZ8OsYpL4H2WPCTxBo5wzBX3L5g7y8n
yFssoSp8egHremmYNBIxOY/10PkXQuvCpT3tq7eC1XBMvEQKxfHE+Hi+alxEVn3bcPunMRDvomvI
GIyGG7F/B7s781rj2Gr8qvFVJ+lEbcQmvVTMkY68f618wDmUl+bo49/hj4/dslPztAtWqKgIAbwq
QxKKzfDDAjemeX8knzwWVmZ3bP8IhzayIlNk+95a/7lNPcjKsQqjWU7AP02EScWTVXownGxJ0MJ9
GAiPlJi29Ptp22ynv+1xukdSqo8pog04w+m7En0T2jm1LI+Yf+AT2zrq67mDkicV8XcZExt/P6lR
mRpaFkZKD6KTHROr50EOxrVHOGIC/KUY/QjJyGcLXFhQOPO2fG0YtA6Ur19C+VE2ils3cmGC+oUn
oaasZgc7DBlOQiQmrACWw7O+q3QCIv+boc5A/Ah9yWjxjh7OCQBP5TNlrpW6FPTP2cShNGvY5UJf
6uW242R1NAlZYDsCFbLmxLp7/Bxt/w34ugrDWXVpkcpJuw/labffor7umXhn302dADcYvSwmRHvU
4fA6ZIsRRPI1DG8CHl0l6T81Q+cO3n0iWGWi5qeInOkpFFRlCMzKUjYXxuwIGWxs9fm5MscdLtuT
ZY1wxbHRcBwmvCYtNrzbfVlMfjdEGT891Uk4jLfi3f3NT6K+0LrKGsTZNgI/2m7CwePuMULrgVwZ
f4ZL5a/jc9Zi97+8K48eXRa1fIJzQym9jPQyJE2PAHD/xolbG4wsXKsy5ptlLIJ770xHvrFgsvUt
3Gxlu2RbOA/Rmq3+6wwnp/BDq9zn4xLW8Pk8RqodIfnog4JzvCoXiueMFnZUQCe5rY+ljcD980tw
ksD9NpAfPkPDwxFl7sEC+8SY5w9yKjMVNcagPyZRIfr9xEsL603DDzbOlgTPo+pSR94i1JkP5nCE
GK8TAOpIMV9IIcJnmHUfPGFTHgbaklGtnh0/HutYqXCSnVZDsMvxosNn0LZ26BkEcgJEIDB+t45Y
d7sWRJW/0fZyCfdPBCJrOlKFzkPEoKeV++v0rJYGF5KWkPz6X22al/bYzcYWoTq79YITz5pxD5hc
DjRL8TvExoCewnMtYaDJTHwzcNODMLny1TbZqtCKSH+6Zi1sSizS2WUiEzeg7tErLZM0m6ys6kSk
nrJbgG8HGl2PSBrlTqan1gXKDsGh7J4qLD0Ef/qAEEhgGC14eK9biPRDWOsWHLRSYjvbJjcKj5+R
XyKr+NTLatroFXB7Feim1J2hH1NPTMsnRCq31fHOm1BQO+HzVZXjm3gTZRpyvmHBCiH4noi8ikGz
o8pYu6Vr41ek/zdhG6QgwFGk6pF4kJZ8NFUGKnTV4Nck9wUET9f7kYINbzjG0L2XNo8YRGK/EN2n
/Kwj9EHcz9CqX1qsuAvOd9qXn42ZHfrmlQZLq5lgKDO/jZs0p1KyrwYGuMssWxEnHx+J7v1i7tjF
qbS4Vz7wlqiZ94ZUJ1KHEH20ppKg2gG6Uy1AlDEDhs7dr1Rgjqrv8HrqYtqceUqGcMFq6cSp/2SO
vtQ9R2DeRIe/pur/Ic92BENw98QNmBd3EcWOS6OcgVHBzd21D76uA3E2ofGDTeKbND0yrQ1pHURJ
iF5RCWTTSFJB1Cb0fO2HRPY/sIoxbmSGmv2OsDyxFyrpRBwS/a2kLCXyKSQJK3GqOIKZeGfyM5eX
z2bVlXIPcetAIsVmXt+O6CnHAOnxXo9qMMb5X1hU47oz2AlVDsDzPvozySUA1XjxX6KhDYS8nPFt
3PdSxjaX5GMJPU4SvYuTcaLaIEFrrqGKzaYYJTelUpr52Z6o/OcM2ewYIc+6nGfkqok6ZmN8KRu3
MzL8FP2SWFfUI5odo780Ls3WpX1rFu7m5Q5WhagtPUeEbu0Vh4e9oWtoDPRgLp0/GMvy102prKqN
3gCUeflBVCxfNzinAwFxF2b+RIqrIOrutGLQAZumi/RWgN8fXj2seT9DFdo1iJcPG1UU3/tJ+Wwc
35+Nfg9uT4khaU/y+ee4tv7HFApdwhbWfmm6kRmwUMUjTS9YurDjPQujroHfz0kURM3m+LoBNODa
yR0hzb3vnqds8dVOOrP4eV9LcYEzvafzCUwellAzDJTHRv8TR16MV+CGNlmAiXy+xTGQp4UgFLV6
Wk1j2geWDxTPooE2NWnahAPLM92lJ8hzx171wxJj6QfdVW92ZN+41Ypfu7OHQQQSUCXveHrHNTQr
AU7RphkUx3Il/ctpMHzK8eLCxqBTgQfzI4jEdGYFgdAbkSjsuQWNwhiSsr0zqgcIxedet7sfdvyK
FGLDq/E2pz4o1xr+AX90HPLmPt9yBM674HcKguctpWrrPR2aWd/gKYWJMpFqCJTIwoB0gF/a/X+6
fGx69G39vQfG1zWt2kgy7RVlYPNtxvXGm2n8EN5gvvgmDN0lu+k1k4PE4ktyeec0toZ71E+sfnQT
RUosti1gHdL3BNxVlQcP2Yhnc4ZHV/Ah0b3h6jKR4+I+g0FKaFtHnoaltd5hNNUEPsbX1fLNAMMp
Qn8BzuKmL3sU3dfjE4CSqR3cmtEvxegrZCdh0xd4TNGI9y/7v9vJThCvpx6mOYmKRAG9ddN+3xvm
o6c0i3TybiiJ4wVuSzUTbMV2S2Z7TWO/MBOUYfsjsdVCwE9Y2m0ZOwaPySTXYVf1lkZjXucI8vKe
Guzcb4zp4v7NGifQFwPFWzMwIlz9ZNFvHdwj/2zDwHYSPQAL2xxaNyV4A6F2ZicrxAR9Kn0hfzAd
WgTTOlEVhJu1QjhyNv6eXuUu4LjNFkCTnT1wCrA3yKGucm9PiWEO46e0IVWTel61WA4eNDltcVNN
hQ741Qsj7wk8PxXkuFpuCtugSfLPQ1RaSqUNWjiO0WzFv54unJS1mqRLuFDaKZmt3nMlQyXbvxtm
1LPeKaHZNl0bPIJap+nwsy2eQmpgKYrvZ2ofNPpvy9F9YfCpKhcEqd+Y1l+6QiFAWM4md5mDBl0t
ETljho7jBOcCaNSxdCWLVg1bFB9zpUGa2j/1JM/U0I/Up9/wZ8yh0ua6jqepKs8EXmgYkgbegWTJ
XudevZXew9MOKpI5UXbG+eiIWSM5lZ8ZKYGV3YnGmeLbTLyEPiiVWZNzHKeFlTOTuu6rykPdMMdq
mqLHyNmjAxcnTl3TdETJ3/twGocZaH2T1fZPJhh71qVGLh7H0zA8/hL9ZUcmnTrLPfPrcmYbpn3d
bOBrhHui0CBGhfAcqK0BlawvnzBQd8AKF6CYWck92ntOyklHJy7MjD+lRT0zoZ060DYLeii5ut7t
I4yCsveFBLeJ+6GTEesjQgov/0RmIOYqTYKI2XMiZGpuO+7sENkKfjl2JT/OPjzeQm5jNFdyGdxi
M3zQeOwAYEVnr94KppnUYQmh9o+r58gRCB8EJsTq9QaL5AHH0APC5T/DOxZ6wqdF0nqG4WoWARrM
axc4jrOV0+8aJlnX3Dpx4fGuR0LKTOK2LwT0fnsgfwi0ZlD0zF4voM9r5Pau1gjC4WJ5meflOBTo
pvOdx/a6uZmROcnt0u35zS4uNnaxs14JB8jAcXfwms7R6XS4ilF58/peyPpWfBVV5gVdwf9DTrPA
HP9q3ZkJawqUH8xAj7rckcMDfi78spZkkavSFe5Qky8tpVeAGgvfX8c0b01YwoFoCIPc4qImZWH/
FgSnpS6lt1GwYF2BgF1B8AUN1itwpddGkVoEt0nJAfBTLMKE/ozxP0ehne9JINqzOQuhg3mGpdfd
gPwMXbbKno3zsXH13euUJEzNsy7Vx1W0ECNIn1JG8vFbKMuOcnmqsPeIBS56cwjWzK+0sXAPxAiF
hiF5VZrArIoWQfSEp0j/lQ9LRUbeecVZ3DWf7lR3JUlzj0KuSJFEG3eisVqSnVTpz2KtK8UVPiF0
1llyUzSaJJaZmSIP8XzyRT1clnipC3lUhwsMPgDneIKbfowEgawvofND9vxodBhcdTuIQoZI2531
ifKleJHIGLC460hfpsFvnNIwW+n/oWx72uf0WM6iSnIQ4Ck1ugA90oppaPLbByr1krUGl1SGyr+J
JpB/dj4g7wG9NyPlVN1kRhzrh60RlP9zQO7XDqOPUpOBvr6YfNkMU5pCZlRF7pC/iT66dMEhmJjh
mFSGl3CkXAvxoTJlk4E4CCFhATpSskNqQ1K6OEhfwbjD7aszyqyi2mBPZ8Qb8GcBFbGJWZNHRCAh
ETnjFsSN1fvb5PbtkfsfYLuRreLUv3xqU1tv3S4l2EPoJxZKkM/Q79+hBLH0QpJTbtRGfzSTz9Iz
iMacsf6EI5axuySw6+XGR6aojAW8exw5iz0C4JK73RxD2m/dMvPgAnMzjXhthGPteRpwqxFAH6Cg
+hupX05QYYNRFB58A5+aAA3UmIgPaksZyoEOkQ3oa8AJBdyyWYBB8QbcT1jMFKrVTYoVq3J1jcCh
/lKZ+uM2tLiscPE+z0Zxmqd0Z+qRAlbo7L6ZED3rt8/13z8rqGZ9TCL89DnQea9dC3/o+FnYYdPv
DwUqEQQOAsudlLQtn5H/nWBYNh3NCLVsu1aQfDXjmlwr0pegz32BbxbBLmBntt8KTz7MtsNsG+Nt
aZI2NTYu9BD8npl7dfOLJ9vsEaiCtJGpm9YAjKpOD3py6e2eLGhUOb2SAumVnG58g/DDWqDTxW5a
NOPFZV586TU1WGpqOLEyUNo5iYIV10lMm2GRIe0N0VYVe5YHsBx3Ny9x48mhpeM6kKw87EvD0e8I
S+j2AX2NEfPBaMmGi2BS/0Itj8KA4q1L27KvYXCLl0i1BtBtVBtVQwXZU8xMBr+JX70c/W3lufVH
Rbxx44zAmesVKJiigOq2cG12C2q4gewBYtb4Y1eeSssdyQLA5rJ970d2UfWSqWp/9+yitHab625D
UzcefCjwvP3Y/bnH3H5uAqjYBmtpGVlqfCNit0CW2lp6RNxSCSgVX67uqhb9ck6lc+O6n+dIFpeB
ariYKFeFGXDKV2yrP82LUMEePTT2W/434lzQokFkFYQXxu8XJQM8hqDm8hhmypviY544UiE7SQmN
gBbfz4k5thTtQyEuxh6FjsvteX42wnmoQXcGf2g+qgbzOGVeGxbxzcsD/BDUWMyG3TvmvAowGWTQ
ZY2fiosDAmSvA2dUXPURNhCM0LVRB3WfrsfB77UBQzcrrKszKj35tIVZ4Tkmdcx2doMc1+dbsafE
ZSiEwaEYMM5Fp+lVQ/gHBEd8R1GK4CfI5l4wULU0oDelZIAoRpNw8AXA4HjDQs1IwL7ubzGetA3p
PpGLaK+akKD8sdjrVdOOBaaPSCFDgogSJMDu6ExoydaUMhOG2S5i9fgFpQkwxVpv4EuXTiQYIx0z
bWYDB63rAR/qPmwc2lcInm/C+GpVPj4DUEw5aQhmyGpcRd2kYQtY3mxgf13o5Yf+Ob1/mEvbqzN4
9PSkVdkIy009IyNE5waPA0HJVmRRZDhXwduTOjxDDGNAVJhherkpyN6T8v+5I3HkZ1dm0XzbFTDF
/zYualfNGAjJxRzGfiovo/llhpNsdNV0ezo+LgxL0CUOxIkO4n/GCUusWQYXxzpUGjOsN2XzMZ3H
/6VQjhElLWLP4+sqlytWwVzbzjggFRMFjaDGShDwgL2RGqL4mQrMaULsBMyXyfwNnpMNdfUkED3D
t1a/ysYT/DvMGKHgbXxf8xPfGl9Bn884NP+El4IJD/cJFLOuth5E/rgMDOKOlNxzyK12n2Wwymm1
e9iK/F2t8VZpnHnua46O8myjcHh6tdHlXWzIBQhpRhllpVDvHy75ikToXHdbh2QdDiMbSqPAELe5
y7Wtq3Z57JF+7Pic8cX30DLYu6ERT0HfgFL85qNrCbUoU/lCW1IuQ6WNZMTogD7mAc2CWQ7T/GCU
ZXhvPfIlnl+ZRx3xVgleAVAoW0eiyU8PpPoiZaR7kCFDWdtaaZAUfKNIMTeFBL7UYtSDQQWEonrX
Y88HplLsRkrN+nOW0ULCD4b3z5Rj2KsYGyPJjAvvjtkmE/LlM6QiCKRL9gLadjX+2MrNt405C7Px
leGHocu+sCPVSWPqI2q4J7ce1AmWe4cFU4RV2s+Okj8XEwZgT52g2b+SD1KFKwggIG2AuKfCicns
J6YDoRmQaYQwbM9ECkwIsMpuJxZWZiuu1FcxrXxAielmVZ9yZ1nhaSV8VHb/RHUCla+Juj7zpMEC
bGzBSMaMzEhiWvL2RzGx/t8JfmLE9QJTufxVSSHFAOVlq0k40SCnKxih6PCdLu6cGwbeQyJp1WND
QYZ4/c7Fxf2la0rdBbut+X114y1eMA1H0S7C96Sv/vxBTdKPHYNnyiLh4S7SzACUTli39ziavzIj
KKevrV9/ymOgEagw0nJbWfquFngFjzHg/5nUjLZgLGI6h4+t3vZ4bFVKRAiDNw9rI0gQC9YaoM7V
VWeQzclc73BKOoUp0Uw5cMgWnYe3K4KsGxAZJ5K0ItRjS+PJqqsLYSqcfh1ARBrGLQsFSRq2L46R
zjEXBHIHh1mmA6PolSoVBKzU5fAStz0ZcErYpl76VrNBkv/pkrkRixR/IfRBTGz5jr53YPWedfxH
RH+0UYRzLL+Ssgl0YJ8xLUpMGOvX+H7O45Yz/alpo3dXxOU/Pv5r09D1/me5zw6jmZQJO8OxOBg4
d/5ebt4YHfIZB/QRaKxQovF59hczIJ7Xc5KUXhznc3iGt7fEeKF3YotVMqRFKzX4mTeKVeDmU6o4
k/1apzuDEk8toseHi3mVtrUUMVNRUiX/TCLCc44Yx5+527RcFZQ+7szNaPNxBU9fbTN8N/21tVWL
TjDd/mpV2R1+rGveyRQ66yHtEmERKnGkloqFdeX5BclWvzurxwTTDEHfJ5kcNSd/aSirKtMtQUXn
Kl+C8MENIvRHj/deKUKUwNZ1dzQZxldevObCo7ur94LwhLz6nI2/2iP73mi1N4mgoFTTean3MWNv
jYgGapsM1NsVIEdOdwL5pwWlL2R/nE+/Bodiz4UWSKX0yn/nJZCHj5aDwEr4Snjfn7Efi/+O3+xn
zvqi/k7Xf0NKulBLuH93ehrPql1/g49waK/bLD0uCFvJmps+jEww3W+yzCw9EhBDgYMu0rPB8iAy
d7vREoQfgmU4sJixdSwPfsTqlT/BpIZoK73ei+OgP7Imv32BR5SQHuH9xBCYv6/p7jZt5lnhQo+8
DAsH/oKzAAnDquUpRts0hNzm8pmbOtqryMdMx7i9zKcVLQ0mAYSi+kZatlFKaISeuyw+0psnfNE1
67jIY6UYGuonZ9zyZLXcGUnzvSzcMmf6+Uzs5AQY8U61eX0cuBd7cmtNv5CpbRcHFHVkq1TXIyaJ
46JnW6+XMk8ZiqFmJsYzUt+ziMz0BjuJlVU6goXu+kmBjl8am/QXKiaqqdub48lDTID0gbUFbc0f
uRqX77OPtVQVK9EIwYkOglTfIKzn+NSasXhbzzupYGoRN2r7NdZyXrt+LpCAUQcD5Q1tDx6qBoGe
9K45UiD656Z9K00Jt8xv0Oq2rnhWGycMUya4gI9zx+zMpk1B6KS6N3zyXhcJY8TR7ILjLWT0mwie
n4y86T45zxPXr2maZ/bXpU5e+0OsicCZz5j2MQNNMcmNONbxCHeCVK/0Ow0tiT2XBSvMWw2Iiao2
Y1hJnQfgOSquhJUZFcjl9JHaqX1yjbi8dbzbiKXpjYhyy6kJWrTkhjZinW7jThed5D01hoIsfnU8
zXWrAyslmj0EsLcBtOIpiWVksei8SIxEFnbRENfVRIcl6HP3I+ph5p8Tc+wb8RNJQ5ONQjvyw4sd
oOsciTgjD6yN4Bsdh0dY04IglRfZ2Es6q2Yj8K5gZ1Lxy7noKs2zK7dlKOKBoCg2g/OwLfQRNDbq
OW2axapIkR0u+SEE69XgU1citWUk1j/b3+0JcYtSLjI0UzWZXZYUuP2K3sdNxQ70GPUqfJlVnrdk
zGgru8Q6vYiqDWd/oNzPpbX0K6PBsyrKJ6khf9V3ErRBX45ziDeZBRG4C+KAij3BX4xnjMSm/F4R
eIFPjofud9WkO6/NmzJqZFF+czFMvk2KasqIs1y/DQmvkMKhIBlWcBSX+hwSZ6mxKoqC1907L733
A4p/0C3nVImH42Yu/Ik7fODUWSMCAkou6iOtg5LNwwraa8N+AexnNFvrzTq0wmEuFJ0wufLAAxtb
MkD1yXT06nAleHczfNSf92GEjhTq3n6KlgVUYchdbwZGX13+9uzcGC7aP0c1494p/mz3SoqVuTBe
Mp86fsz4WlQKSjeFkQQp3z2wz5xtLqY+ZR3bVZbPGOazf3GDF9rDBXT0rJubnZ3B4fwIfaKukyFa
h0RSdzeXYzcGgHFZV2bdyzvzVbcrrt3v9O11wcnYYExapQirtCNEhXsP5cp+c+h7aQ3akf5AZlaF
AWL+ncH4b5X6pkuNB48g+jKHbI7L2llx3rnK/gvs6cT2xx6KHcMPm3M0/+n2bBxxy7+YzhIo0MUQ
XRujCJOKC+0xx0i8okfMHkf76oLlpl9in2HWclIJ1duqiHbsCssvHJHSDvrVObjAAdaZzuq45QA9
ckoFjgT7VjlFQj9li1k6XW/KrfsVtXT0eICCg07xTLKE0+u54cKBEuUsG+ZnnWDsf+a8m5tcNEEw
44j8Dq4d4yhteJdrHI/bAP1rJRUxHjMC0Am0LKEGg9BZnTfePClAlLDbtHCLJbfPFN6MvgQOzzsI
eoFUMWSREHTYtWtGfCCbmwDfEFl3ung6FYqsu95p02xAgdqBmAQsu8FJ0H2Sbqzygwl1xGWGjH1h
umySkAnrpXyvsKrTRHwkpzs6IDaJh6Bev/1eLfLmUyU7WKyMRi2yB9CAX6i3h7QB8nM9p7QaKafu
xOjjW4uf13RPskGAZj2sLweofZS+F+h63D6ZhS5Mky7yLTyY3kHCI3/Uh6tLjZCE5YhB9u70aw4F
WJ9l018iYmOsCpY6IHdXZvNvldHntc6ylk374yXPNs/615cI4KNYfTbakLszkks3IJJ3i/icYKqQ
Mquv5fYV8wQoVeCDe9N/d2AVjW2QWdHzLnr13cCqA55xfzPLI9/U5Re5u92GVV3dEhH815eUHd6R
39OMy3P8DXMe4kO5ZwjIRnzmtchBKlDVIygc6/X7gvRUYVKli7lCCUaGKDOoTOTy6cnGEy1UNSCK
taLE3DPK591DKmtzh06uZYww6xRhWXNFm0stNrlIr3GQfF7hVKoPnPEv8nVLJCwCOLTwD/0MOX3I
guDKREOrYHLMNQOPDgYS6r3qxJ2GM4QYvDzzQp4+w4LBilfOXRl2ugq5rq860eaK0YjEmVyQ7vgo
MxjfM5LPHVcB6ZQG+pwto9rkh4soFVrttE7kDm9k4Ygz9vrSg/qlAskculR7dDLy4kArZ1tP9Ydk
qG+VguLzMpNokkc7KxKaBm5exNlNgGGo4ACkBrIVdJS1YEinlUlxyHZl74NzeSrsn8QYIk88UW7w
JS5xUwsxJYyVUGT5aJPaLZrXGUjgPukvpmsOFQy31KEbU6JIl5mnRbgE5DyhSQTAGUf0VfmmuVIU
QnqT7u1n/V4j288MW2NVPBTTwzaY3iiuYihw3ZfL/mvVcchMizHJD7tiLKZWsQLjLEQuJjUlZaE1
43nHsJM8Y2GUw4YgKs9EoZP/bUCdq59GenZCupTZNHKHplzegHENexU/7ttVnLCHNx3E2TNnt1tq
AIk2KsSPpQYmdiQLYZH1PtfwhLQE3MMc0YXk9F68g5VnW86JYkIWIwSsKHOwvxOR+eW3oivR7aIt
qDpt/Ks+0okXy/F/Qpc+4ydWKotlDOQp6ZZqAehjCNYYEL9bU68oEA3EGBqa+iTnvTJ1y/VdzC5B
tlTtBbUm28IRBZRfZ0mcQ3bjMxIR2XAglcUezcUrK1WXS3JlNSWNzkQ+vWtltbzN2X5qyiaOGfQy
Gd7zBJMRF6M/SL5oXaheFUzn5hBxLdW1wqiVmEc4mtU7rWFenJUsMsGXEpkYwsjZk3ntqHlYbsx1
pmNBRaJvfHU8NYOXF96Iuq/46fU+E2N4k5zuLbpgaflVDDc8AzzslSlcqYQ8XtNPdxH0zoxxA1x9
9gnfWpBpmRX2pn4ewSYx/+vClA+8gtUKBPjWPhmIVARBu/aoxcrM1pn0g2N90AxbUUq1SecuwDVk
nNmgXsz3hZ1URK7JxRNuY0qWK86wjFOBW214n56JLUxuo8MkCtQEKkETDHpyUTShecg1fnqg9I5s
QRiUo/1cVcv1cPd4wyaOuem+fH13bgw1xVbbCJjKOqktzz/o/iyqlYZJOQ9MD+ha9CT7OWPYPi6o
e7emsuXECMtIQVuqGCO0HcC5SBKZr0pbAr3AkCGUasrbdeIhzHoJ50b8rF2TAQmXy1DvmPmc9+yc
fqcMnWi/2kLFtm1GKznnyp3xoNiC520o+Sbq++X7i3nNgBtfDpoqEb7v2RYVW9jGnhOxdb3vNBWB
EWunsS/0/I9dy/R4B9p5CXQ7qPOR4XJN7GSZmVlDxJupd15RA1A5/BMRyFqKKq15XIxy5HuePsDc
/5rqMnSv3w1HE7/d7rGvLSCmM19081xrLitystEomlBOXsm8O9F0mzJfivmqw4W0U99upqjr2PQ1
yAbuXUXBGwsMIIkcLLM/dPq0vTywxmk+RVeOAz5dR7TkgK8qqAcbR3z6hkQAl71Zm2Ej7taIon8L
BZfjcWLjdAde0LyO5hj4i3SKi3eGza0aqoQh2VoTWl6wRuH7Bep/FpINWP/lRkXO54PKag3pUu/W
Pb/PgKxvfjwOgFNt7OXo4sZux8q8/LxtZonIzq0pAGfTuXkAVQ1s1dvtSIzRK0ajoPqR/rV5IOhF
iTu/XQuqDlyebUQcCP1o9VFY819qdEnInSiINzUjuhFouQh/p45ZJSETmcuMYhvoaGCMo0k6RriC
FdsMZZPUg5KkwT7+w33dqjatbSTN1oDH5Px3sGf9Pbbaljhwx+ZJsuYjPwxFeL3zJZoMlJJ8bGxB
jNLZPh525MWZwRt4742QydkC6DY/gQ3EXPnaHgrAhgGlff6OpiZK2AuBDwSjLUNmG1VH5F2Bu8do
AFjmNO+7IEStSOzSvx0BKFjSyI1rfbVX2mD4mdezIdeMbUMEr5xrLqKwRYDjvTkn0nwdQ3a5EdeI
hYlp/kLjVIGmA0bfrAVtkHpfO6wAWGzeezW30XNY7bdQ53T+btJ4OEz4qmRVtO5mxhtOzkuM36/C
0BAyKuhBZskirMlgK5XvXio4MmxZU/4+yk8uQna1kvyAiGPgDYhip2FHY33Au7OePHjCyMbWPNjy
hvjXRFShd6hoRv6JisewZ1Od9iUiwk0c1blTQ5lyHR2Len5LT8frNDkLetqc+NULjFGbpVQD5oyc
4ksa53pbIaOI+81tSw/KtrDQLcYOIR+WdpC1RXkVAUEAKwEahjjjyhjcTaGiv7FECdH+9+FMtpwK
f3yrJJSBJ26wHhh2L6gk4yH0HKViX2WmsM4uw8EknY2kLvOgzpA81l2k3dLE5NfoqJrbnV+yKwXl
CMafd89IzDC0MLVw7aHM/UrN/Gm5D0KUADV2Cveiuq/Gsl9FcR4m9pDdKwry7oDcT8d9EJhdsBhI
W3UDqf6Ylc60lDDPxQIS/GZx45BK7cqPn7fcnNCFuySNfTVCX+6YJKSnx2b672gMmk2pNUYDo5j2
f4BrCIUv0incsR8er/1kYIeKnRrS7YRvrNc71bNzPmf0yr69hiT9pzbKigoUD8dnlilFWpLhLnM/
NOM1OfPq6iAF01Swbud+APoZA44CpqGn/pXJLhFWdyXtlaYOeufGpLtYLoAm3tONs0oXce/P7/DP
pJm8H3y1n7s30+8BwZhM+MPiyt/VnYDZuzCYTTsrPVfhiTvhQmddSwPqR3t9pW33lbQ0ubWG2cvu
ZrneK98KabTOhGVT9PXqqoSHdHDK0tu+FSwBxhsV+VGt/I7GS7NVMhpExg4MpaJ4o1dY7Qo9EC7X
QSpI2f3FJO9Jjgf/974DALa8sTZpgiisQ/CAYL0JuGD1EMB7M5t9qeV++37S3Y2n+eeHLBvWKiwF
Y6y/tfduk2tHfFw15YAsstf0Mk+X8T9RpiLaCJ57QzYM6MJBZYrABNLRuUmwWMHJkx1PGs3Rp8Yq
RrwBJaDuV8LgNg+BRnpv3pS+1ZCYZnShZDfm9d76A+o2E8PiGZw8NTU8Yh2uYAR+emVDVUTTHJEt
9IPuXrSmHKC1b3vBXpa5ZEUZ7oznjib1Cod+h02poH+Gw5TLqkFW4Cep945uhSHHu9C0uzHNGTxV
FCNwchRAKMTPIzFo1T+tpbC+xFwLL80ONE5hy1WrqnIn5i1iOs7FrW+n2cBCdEq5pkrRQs4B2Xxq
rJC1q/CYB2ImCNC9sFTy4QQeDGmVSnSirBsCPv2fv+6+EeJjNHMiT7GKJdZ8IVmawyc3a5URIP77
gGx73ZGFfejj+uegcXkSoadBen5GxdYKNK03CrOr6Kz8Cwq5ZhAyTLxdGwCSpNXK0LZAJLgQF33J
St9GKvw4JM9K2ML3N/fc3J+f+uNpZee2pIhvRqTB7MQT51Nl9vau9k15I23k0gL630o76a9EYo3I
eBPNgxtm6mwvIeeDC3HWX+bxPMGhCuBjnb3aW5o6fQLBkzt1FiyEqTsxkbwMigGLJYwOopQljcA1
gH8NvgEyXh94/EZXhZG25tO6a4M7cerYfZgYpdnuEQA2mMDPnchuNWyx6+m0oqL7lgiPan0NCT4m
LsIprZQyqtZf5K9zajxGUsgPyfH1YDz2U4cMydQuoVBsNZM1zUH1MrEPmXUGTUN22YX2iI7TdLna
1pUG/TP8ScwTwdnt0JJXdZgdY+8bkHtnuj8J2eLWfB4PgJKrS6OFB+5mE9BF6ELZ3ckgkamEwOTO
LAnyNelBrBohZ6Gn9aREPB1dMbfwi27t2M8M5YesQkRdR48vU1E7dmIPZgfb2+vBHab7J+7cqf50
iRPa/sP4MMts/RalOx+J2JXV9pY7mbqGNL8w58NTA5+LZ8B55qoftwyIvhzL/BprLMn3gW+3sB+w
a+Xe5k3uV5ELYgfSeY5AMCKjEGZiU+ogYX75JIk+heZ0hgXrD9TfsjwBL1D9n1qArniG2YdH95na
FlNSHqUjElMVu4HD1EtffONNCC8awRti0HFD87N61Rg+FPy2ezmncdIVgaYuZCIgZ1AqfJHaqNNj
+WVEe5OKQYVAjIU4QGIItAXuHxBtw4y1v8RA7EepxkyPt3yiO6I3OusLIuCrkC1jgrBqkud1vh+t
Yp00jJTC4qSyih2i0eDnAkNdq/2o64kvrxTlaymNXZF/Ink6XwtwTh2kz26CLXrlTJUBQRlbByUn
dMgTLSrfkFb404zmG2o750WuBqi2yJZhA3v4DXc6BKnn0UELaPvtgl2skK28GijUpu9fvXDRpGVf
9WAN+MdwRigno4SipotMxc+5nsErLAfsBYPkwaf8+Aw1sUmpTEjQO+15JNoq3yV7QYOQTHBvFIGI
dvZ9qnnUJk1V6wRIAu5T6YZ64+BC0hVDuo27r+oivdOA2lwatBKqMiWUhIphntOmE/aAoxbMnGpd
mBCoYw43T3Woq3EcHEGRCqKVIC5G59Zgl2UQKvdqran/y0IdebYghqOL1ytJ16CSQSayxsNXIDRX
CNpv07GaTmf5VE0OApA3bliUyOJoWaFFJlUA73Txfgdu5YTIIN2kHkBTMntFG4qzsSt5lKV6xrR4
Ii4cPPg0mx+Glr2SHIBiNfSd5Kk7iHYCQIEbnHBFVfxQJJKoFoH6E9zLZ59crC+naypDu7H5QQ3L
TAlRlVcy+HxI+OSOYRl5R5gDhJ3m8FEHIdPxLI8VN3+LT6RBrdmczN9MaSRDxPqnGOPUDrGqHY0w
ge0Ge3yv8Et7pyOuhvF5xBRuislEzNyxAPxaa64/Svfyfh/cUdaV4+/d4M9KOVDXIOiU9pf0aU1s
xpQPPHLZDQBzThNj2cPEczlGlxfXRIJK8gzCH7fDx0axMpt2jCkMJykq2atLClIeII9919cX5rOY
AEQ/ch3NwXqByNQbYIs0hEFZt8ggdoA+EnuMzeeSY2VFo4ojLDtvdQS/sdaZtbJN2hnhL3AlIX/T
tG66BZcuWrM4WgX+ptNSuPJZFyaPcRWl6Rc8s0uSO5XlEse9FEavMgKcGMSrJ3ztUXsqDqIAkS1v
ZMroQbqwOHmT3o/DuGGzbTA3Q+IQXs5IbH9jaMbF6vQrVweRnndfUOVHQneMjp+gIrx0tvTb4seW
bjwgUuwIQxUiOCas2cHodLRf47DWh58anOVD+/VPULwZKWZHuItpY2Nf4qWqVeFtLKnuL5YT5VLV
dXww+JkQxCHIyPq3utEqAhw2ZZ5RcHMeGjZGYUf/VhBbZSYcUVKkmtz6XL6XLP0oT2nFkBUjbWyy
GASGzUR9OkQzGn3JjeeuVNJQfBaM2biTsrZSS2oKP1yqBFuYV1ZjNdY+2AQJnP+rQei7JVJIEn+3
VArL2kIdXedqZPRGILWWbrh06OeMWVm4cUvpdtCne8SX+SdE3SxkijYPakZivs+FYSzUc7aCZIS1
w2ACIA+igrOGVCu+VaNLBpmlrNf31Wx7BTkc1bbycOqk0DNIIqDnx6MW+rilN+qZFhYziW7CtniC
K4eBaQXEUDLQY6o4406+o3pR7wsW/Vvwy+QBBrJ2+7HpYuszAHV+ST6SaYdBmEOUvVy0GzXoEcQX
dxOcGpIKlWqreTMWahTdzo5G6WUph2Sb0stWKH0X/9CaNxiK7umc7qoYKrLPPQH+lB5UAkr94CnD
q7d2BtidX2rK013jeRMpBGtvAKy78JsHUWNX9UJV+NxbKZhwD/hokdNRGtRdGuloZt1w/joq8gKl
nNtNWCYys3Y3Mb7GGHuELU2AUKL7SHDUz4mhVFWE7ckKru7jg7cPRthFSvJ1k0+gGdGOM8T9TynH
OHZZj3E2Ip/jojqEIdurYR9IIaT9+JrUj0TGy80AeO7cNmOzoOazmbi/mqcR7CPjBMgczAoJZ1ig
8QoMiPoutmDTDSaO/5nOX09B85mHCSh3KQw5I2ZD1A3mKzghpa+AGbPqPxWoZe3B4qk0ZkSKFm3k
giMRVgDoph7avx9Cy4DQg8AxhtqrXrtE0cg9V8tusc8O7AFlDMMdFcyFaTN27KK7SHAPtlTWQw+i
2msXjhplJ1NVYkMS9+lGyRsD6bAbiczWRvHrkoCYRgpA2I/NjJ22Usf2IweOxcpovD1iMkdYAbUV
VSvy3RJXk/EZejwoswh8zvAnYDyEEqq2nno8u5bjoRqaKbzproKBZApTcZOf7KAuG0X7VsvWK6Ea
kVOjlFzdDhMc+4Hfk0CgTkwwvYDSgTq0TvWy/gRGzOf08kdmjGCoHgtMxzB0ASDnAkRlIhwXMo6K
leHxgmoav+2FQy6Fa1PO2gg5vghI9TnrR4kJ1LkJeLRlfbThaR/4qTuWKu4v2AmAvu/xTTNtIkf/
n/Cunw3aO+LpO8fuSfHTuzD9nUbzSXHPUbqgoSj89V50Pua74RB0yRWDfemCGxg0IpmFGLPl9JTJ
6L/72/ZnUataTSp4+HnbIxmEyyUlPET5IzwKOG+2ZccxjfMY/JySz+pic9bT18hTCGeYYGiCftmn
CXRl0SKUzjpNbEZ+HIV9cD/emFcMjB+MLldWAMvdOR+Aqv4w3wgUIX0BrDgwyhBbUR+hA6D0fqUn
/yX8G5nl9MdR8hEVxVYd7Na6vxA6FsNpi1f8Ea4F8UkW3/cpLGttmNIhMoCuNGa67rpyrHgg85ZY
4Tk7Xfye957zc2BDXNtV2L38rklOG7v9I2FF2wmIhfHqXK4v/r8SNr8P1PL5lacON1/eJOGzYevG
20LmbrBIguq4wNIihVD2g8DigjR8skW2Tii+YEcWCouWYX9oNZzycXOty8ML/F9F8NXJe0pTdCGC
rqFNzLjs+fGHAP7UgWauaIjSCBkeQfwREej+dLa0b/zVEt+z+z8qnpj/eAbALHDQbosqKSSbaoUG
JWzXjld/Giu4f42Qx23kBZg/0yxAl9wgD4RGLIBmnSkcrc4aqbZSLcsbSb3hPVTYJd7H0Dndf3Mx
hDYHH4x1DY8hriQ5NIJTpFuawA8Y9w4x4mUhoOHJ5hdDB0vMQAUeB7JPtUw664FgOAWPpHA9xRm6
IrRdwBoeB9Y8HTNOZihyjTVLNYcvfV7gYlWuVOQ9t9uXMriaJhElK8w2Wpz25dZNmWt6Rb+gCacp
kuU92PxYQDxRCif+973yTZlacfuwymau/JBPmgmkbwqNvQoCpijIwu2FAuyPpbvXVoRd2R6nXlfI
vUBdybtkAITuXUnX90+4XvlR0bbxO321cxJ+oc9tuHzfAHBjg9glV1StTUpU0CeTU2rP6SWmUt+I
w/NGaAcuVnGz3dOOuQwUt7sTkVvl9YWAx9/wztx8BxbWOAEoBELoYj2nFMqVr9CkdDayDwu6cXAW
o+/QDDMCddF1/gjn/EpjVkvJxnFtNSpsej/NTJFgugWuhbqeBwQ1s4xAcBlaDaLwz571JnzjFeNF
HPDngXDJoTxeFJ6fIdAp0uNuY8Im9i7Wo3rg07trooJEqOLCy1Qjmav9hv+NVGatGVIBYHKRrgNn
5vBFpZa8aL/NyyCGZ2kUbtyP8aNhXjQNcqZtx3gZATH4OUsIS1ZjFPNcAXmLJP3550EwTwy1TTdC
BPJIyvaMIRHBWJWOfQZIk0gwTIIGM/Tbijg0cjGFAVwJYMihif5aM/Nj5TBeWJFo5FLUD4ocX/zv
uSpuXj05e0MJixU6PQUeQGNqn50HICYasU3NZ78qPoMZ3lrxC6nHDbmqdIM/Kw7rGCUGEWw8UtYt
6aI/hHj2MqZrvgjnLHdZXVQJB9mdf46qdi5UYBMq2CLkJT/uq8znmg74+rv9R+nzSd9p+ecAkrjm
58U74RSVm4zS7xiEzJS9FuEBHBUpjyGPbY57aHL4ccOKcd9KlsgsOn2dKiiCm/YdxU6uHTEWuI2h
Bg3SZUw9hmXAtaScYr6Fpl8Z1A7wLzsUqCDjtdWBP1huWXj1iC0yX89rDtsI8IMsVL+y/h69tRId
bHbCqywUnjt8M05TBsID3bhHTZpNtv4SsIojhD/TUD8IykjkmBJcKTvUl9zwRMT4GY5l3N72EeXq
vPLeG6WRAoJInyjCGAD2ggLAMEtYaQGVkaxCHUGaKfsTiHqw1barDpX1bNfg1zMD7weUkWKsF/fC
Q4du+MXimb7bnjWww1bDEbYJ5XfflGCAc33Tqj0ea4jD+cn+doNNa6JJlGVD7qHziMyRm/GC0Wyu
r3qb8WTeKtZ4wnnlXIV2eRzFDbMwkgoEj1tAd/gkqkgJp89GYm8rUmNkVjkaHhDs61DGxwBxWf6t
4k12wLGVYtgMYvtvwWkNxVXzL2PMhqR3D3sTAi75sfo9xC80N56RTHLa6ltqjKhR6fpQoA++RoGP
MUt7aBz8sAeOqEpEO+NHNWlwnLLvGwJMS2OQGd6/rqLIBtW+owxWCmP9w2/f2B9pJnfNQTjYO+/+
Smj4VwBwbnYnrp8HA/3/uoQJ0jwZri+LCBHOdLcY6TxPUQljpixvTKga+jyhhYQTVg4ibm233Hnr
hQe948Ie7iA6Jj9UYgypCNgIqnsIq4vLAICBGBuratX79PzOO4lW97/JnG4FN0Dq+EujdgGNs2uI
1JhrauqeGuCYQD4lC04bqU4MqyskduJBKoZAPjA/se44DEOSf7/M35brwsWt2FGwYD3chTgBoDux
TwSoF7lwMK4SRO9nmsfMPCkK1vEWleQLTzEP9eM3avs+VtEEV8EgGqMR++ltZQxQw0JuY853J4cy
Vw4f0b0l2k58cLtxSkc7M4HFkCTgRGJUYdrwgrnN8SU+Bzl3M87CgPflCalp0HiysesiAFpCL9hm
Yml4+ipHhO3zZEVDTjnIKtiEeE1jFrKPPi2/vTmGFOswMCzAyJQ5Yjznpd5CvcSruTR6Ky4IXZVt
9oEe/8cADrPr57HB/w5b08A7ZY7zldVbmoECj1J4RszEcldgYi71cOiU6ZtDm9y0A5PKuVJUr2pJ
Rw5Lr61ZQPkRL/o9kk0VTg775jDgCrEcVwVbudYJ0NMYeYkBY6KOUB4Tyy45ynfyNyLV1JHP5h4I
l8zzniomMk7XekEXpw0eGn3UywqKkqsa0a1tpoUDdn2ZFQvlQWU6+tyNumM3WvR38TA+LPknu3XT
ySVr+lIC7lm94FQNQwNNrpkjWtfKFb5n9+gA2BTeaXqscwndlsWzeHgHSk0lHQfP2luniosUAzXv
uszrixIqW4CYFhpHe8naXiOm1n++tJXOckqutdkhGMa0Do3baCs01wU1EOphvvu+gQpOCKv+UUXV
Pgct0HKmXwUNirlGKRUTapI3qFpZ1opXnCa7CRHAu1LlQ6AJvtgIIFtPqVF/aJWTn16zExDvnkJb
OtpRlP6Aq9glpv8hPE66XxVKXsiatliM1Vbv7Oc2BZ6RWOELnAqEsGdiMMNtusivEFmCtX7+vMB4
/IOPhzyKcka94PbmcP+BgkcuNWatiU7fNIIdTHO8CTFqMJh/1KpMh0V59pIWphi4bnAFWfFWwGfb
vbPoJZnVpvHcnRHEgBo8gRa7qPfTZGG9gt5+/Rhog/mPS9SOLYAvDmLuZ4qDjaYhOxafqcI24C0p
R/KIzfeLarInYFBSC+tmNRB+LA7kwMNF77DRYIqHDcog4vvlR6KJU6OVHV3/oFWDn87E4Vr4gEeD
UCkXFEMxjizLvHOb3hh8+AjEu0Qe83j3PdY5KUeJYH+yxHXoU7wnTIwNXZxCFzzqXAV9Akp3OxjY
7spihm3GRC1kcY2Nlu6Cb9cuvro3yxT2XIGggwSPqzNtG90xT9y8fOIyEfgPq49b9ZnGtJ51EYDd
83rack+Fio1q9tcJ8kTmhRdoXb6mg0rlmIT3mdxeL2SOFE2CK3ylcjbNJHFFDq/cnb/tXow/RUqp
uMoOlTUXlc6wa28KbB149uiEMEezgj/gTqEA3v2A5XxnGJHQukw3FO72eagj1qBbHC78F6GYz01P
+yVkEJkgJ3VlwZBdzo2WvD8/sao7mED2XiWaQdRW2G9iCY0i047YYIWZWLhBJbuaxQx3WjVNvy2r
e3qVLU5CCCXn1XFY+7TrWSS6waSgXb4zMeFDxJ27TX4S7YCkoa+6sDFjWt3E4ZkASsxhpVbGIUhG
kvFV1qkV4GFE/+1eZ1DgW7D2bXZgjfKCovhWtF7WC9NbrCpNwN6zJBgGdN8mXX5DNqUwyp/DT/BV
Dw18stkysWQGDr8V+KapHCV9xHbHnjHiIXcDGRJlXz7ZmVfeljqeQnlVpsNj969Rs0lGCl0DbnKW
mcX4IsY1OvHuF88G+Qv1eyqRQKRpAli8aMFImy/PjJ7oyJ7Teosy6V+5EJd45RmEeg8LuMUcYiAx
ELlzrKw+Jlwcr6/M2xvYTVpla6STxrFW1QlcOpyDjO0wfWksZA6Tkor9mBGuh31Y4VQQtGzRKkhR
cDC3eeYD8ZGxF2MpX26zfY2HJYlbwOxkrji34YefHqkedxRsAJFS93q9IMPFdfilrS+CDhRKhnIO
Z8+MlOapzYvJQU3PhRmios9LSIpV1kwF2Vd9n1ANhCtkgqgih3gVh0KuOYD0Oz/KCwJOaUZmuklm
uBEkLXlC9mSPdZ+Qc5T3oiBaqU5n/wwea9Qjq8BEpKDVIj2mFIsVHl7gJ9k0ixlOxDGF75N4UH+g
wJ5vQ1Oakbwbvh7URCDaVllrTXYfwLqgLriGYYo5BsBx+VSRk8iKDMjbMaF6tdbcRTEYlmuejI0j
vuxCJ8uRymTg/bQLGMgav2MEsPEFrCVL/D0dcVaPYz4o/hudrE3zqZYL3PEGnDX9trak1ZisvIvE
Q9W7vGiHl309nLDJANeVJFmEcd5Z9w1Zxsdu5TWTs6YWLowpNpaWUKrJy+37WHsV66Awlh/VCN79
nkD5H6U+jXoMRxW6y0wQCxolTPeTMD1eq+yIOYGcJprT38qkONUOqNB6pSvAUZoBUjoR7AI+l/2z
91j6LF9NKXHyfqjr4ESv6mDtoBKmhyb71XtbJmT94WMZcD4g8drY33dKYEPjWjCq8AnaSy8VSc20
x46xWvZc8pWQWktdJvz7FvFqp2BtQBmTnTINxguLuueo7mNPz7cxx+gDtN5NEqs/c/oxwkLYn0Sq
BheAqpOpUuMSVsG2NHlbgM6Qj5vc5wgWqHXGyEBzRpj9wMe7N1FU5XuHS9IfAMQz1i1tPpPhv+Kz
UoRQsw5+nR5EwLJoJv99wDumvKsz8asiMkTQUfbWothzhETp0tmlAp6AU/+tBTzAeMC3soItPuH8
ME1CNotBwum8ujCXMVPlprmKJ2It51VSfc3Nos7Q0P1sCrAftTMLeRAj7TkEnvBj6E8KvL7ac0hd
bWBU1kzKyrOJkW9RPehragG4QWKUoPX6b7cr9m+w3GI2ZF1YruJCA2D7/pJJKvmmP2iJh08S4h4l
YyHs/iv4jLC8CJfiVx+bWH4eLkj1aKIHrGAZ9w+NhMi3ZDS2F8FzI4K8haQRfnRZRP6dtHPh0Ag5
8u+0y9E4p0Zrjl50QiGzttC1LMuuiQc07TerK/GtwaopurPlZIYO9eiCWtyNhz4k0hDCXZ6nrahs
0ahat0Cl0yySgoTAjV+pzvaY+Cj3svX4FMaeo64ysmzp9wfblhg/EeqhhenqgKwTTx6Kk+QrnR/5
g8nOff5qxn/QifaGgXQjsTnkTUlwQMvl0oP53EO7tD1zlQay2QrfFiixqYXLUvG7b7LzWlLwwn3v
5fi3qo6WMD+yAYRTFzkd8FH0IbhI3BXTPWvehqEz54vOya9PbKRpsYsTGVUoMh0PttxqSLv/pEIY
v3RbcFPPIGZFg6c/9ZgYwhji98wVj0swj41FGQYGsPIyDrD7fv1Iu5YA79iPkA1ri0HOJ18/02tN
qaftqSz9dZ5gBbXyR2D5wrA4kcg5fDQPy969BE+1AaF49vbkpwv5i/lO5HCmG5r9PrEgLDmmMNs2
KZ2XXmcSa6lJEjrdVM4AOrvNR74RzDsFSI80Phm20EF2UBk0CUbDrGcl4vFh8obq5gS/CCuZtgvf
YTmlmkKo8KOT5vlSlEXf8/xcARUuz6kB+M2sxjwK1oLDZvtUiHe3NdqUdP6LOzaKjAMSMnL45k/W
KThixS1trUSwFWsb8X+Y+B8nQ4bxCpaDMLycdLmS0iHcMV/iHWboCq55vWIt5CEIAoK/LraoymYF
+LjWdrTCFPl50QsypKQr7rN7QDF+UHeDsZOAsbtARbECUIjV4VdCTgeTsZhPpAWAgNfOnFmw60jH
aBCNf1qdIdUS0EjN/ce5f498g1xEL92WI/LQADrDgqqXo+2M/K9nf94VnwfLBqs6bknJ5FCxYA0e
ZNnlRlhFBRycIV/ztXzfs83qGAm3gW0Lt3Ofd2VrS3zVZp83kkU4hZBdqI/rkOFy6VYLt4/CDKzr
+/XklcPUUNLI6MJeY+HZ2AsQba0VtoD+chL4CRffTyC6Z6Qfg/elHGz3/p6IlEnY2NaA5/qk3BBG
MJWtq407wBX88g6E2VHi7g5GMxRgQyaI4g69CqEqoixpgwK/iZp6rXPPfHhS0k3uIR0n5A++q3Zs
Zln6G/Tfdy+o5U2WtWcp6xiOFSHsYRIv5kDG5EpM0+cBpRX6BDKrQJYXY7jkuvpQhJwO9grBzw1q
c8dXEelpwCFIhLZO639amE8QNb1Lp2B3+X4X/5hRihTt9qwg5E7nMwCe7/voeEu3s0UL8uGZtSY5
ZJ584WNjuUebLMkvmYgfCwAC3tmzPjvn6sosYAyr2OPZAUKh5j4MjOSqSHgEa9lK39JygtI+kah4
knKRU9LkfYJVSNIK7RzevOlS5QIbRlVrwo/LoAUNe9etC42Ap3MgwjT7KFiqpbajG8esgCf+exOX
cf1oBJGs+cTp7gHQqurCIEGwgyp2FaCtMuHby+NXNNksCoxYIhQ4ipyrr10RHRjViqIe551z1wv1
ABJLSUeNeY4KWJtK9nk+K3iDGf8l/RXieM3zVVdFWfI46n47pTFB6GTUNpD5cxZmY42rkEDbhnuF
3b7prabY8pUTdQFsghQWXJoHhVxKrMGfKFt4B8CihQFFjbu2rMdRbokw3UZ1KpZQGjNlburaFYBe
YJhYOQ5pXtqnuWAtrKOfsSMir/PiuhAmrRcc1/9WhoUPnrFiSHXzlbVrMdNH6s/cg04TSMH13Ndy
DcpxCTn/t2qOmhklZPnanelyBhKI0D5d/YwSeFcHo+HolOTKv7s8nYKgy0H+r4OnsW1fsao8Fj+r
uZl3EcZUy66ujCjdnRyUvTICaoFYtxIJN7EA082ONqrFMgcsCftFVM1jZ2ETd+W61pkOwJ6bjigQ
0cLXF4f1/4g8nYmse29KpEWRmO+bEax6zsaLpwHJxLoaTYDZ8hB7kEWm+N+vyYPDmY3SyAU91tl8
K6acdpxUTKxA1X+AHIeb3qzep9EZpMd13hAkTzWEmHhk3UajyzOuAx42vc6Wwr/fVV6gJcto8RKQ
ryLPRP8tBwYzKq+y9FwftoQmCAbwqA8Kw+CJQSMoMO4vwK9aklp/HUuBfuhi5U8pOhDn0/EvPN0b
t5XwA2gfTmi61qCr2UxsSKuPuewBIvTIiFEmvzThHO/Vyf3UMMjAtdh65xbKArqZqRHNYswNC91s
N3w+XLir3RMDP5lW7qSRn8rx9TAaY4fT6IFJsLSWCfSV+oDuHJYx0/kPjx9AEFDjoslhMhGGyOc2
6g2udcj1ifykWdhBAF6a9RxGnmDmlKglIRwnasLmSkjWwIeP3kvk0ze1svTikz6Zfwb/DI53AaIE
vPfd3t45SqZ+8i1dNi+QcKxzDgOD5qUwlUui4sPFnPjs1C6RYzqs29vk8vWKlplVbAJTvSYK3//S
/otbI9umtJflBQFWkfBJSJfBoZQOT0+oAQeKg1UVVcPs1Y7/JrM41I7EgoCNI0UItBTvGWAcByRK
UKTF+Pi66t3HXkfwkb22Xjql4/4CcbafHL1uYZFn9OcqpAAxzNxUQxEF4TDlhOKETcedvk2++/pY
xPjnJQSCR4GZ27NHeDmzNpeqvPxRGlz4jhZbAvTqqg4bthddn4T028MlaaIgR7gjqzcSYp7R9l/S
r1e5TM2Gr2Kq8WBvt2STjH89QKfmGayCykuXfnTLHBBJttdCWqFNWaOYfBPeV0eOw1IP79q7x0GO
q05RPJ8wxyErCStCJbHMzQaC37SZKkBoBrV+Dtc5E4Fbt5H2MJok9F7iDW9v4qc+b13v41kejXjT
/mrwLUjkf18s2Z8vzcrqVMZ7DU5jDmhZhCW8ypx0i/tNbLLth5DHrDy3ezyBEW2iKkkUFFhbYuA+
0ocdOP3eh9/4ny0Oun9/WtpcQEmBAh6be6trcFYZB+AsvSC692sSor0E1ftj+33nn8SzPw/1N8rB
CHiw8fEC6BNCfCS/neiZlofLMm6GKwAAc+KWbo8btmh6VPpATmoA/kvuD1Ci0ZDttKqnGWBeHT2J
5LWz3HWxyVcyncR05VAGsps+WMGwsKwfWzJaaEQ2V40JNkvy89RQDq77FP8nZKJQiX1GKwfOMkQD
SFfpMFJjTOVftKYqs3VcndzOyqUO36i439pMbg+RtLx2V1AIFk5r4jBhTbKaUhXG0IrKC2eOsor/
Ea/FZBu7iR5wGMqe32iH7t0ubM1iOuKDcKri3lOnfYtMvNDKxOz8g1GskkpWQv5qJKKPesTDZ2U6
FRbyse9EiJK7qJ0bC24ChGblF9olLuSPKVlVYOdCeneJVKpVEi+Q+VcVgw4FF95NcjqlncZ2fnp0
equysa22Oiwh5X7Elv4Fd0A7CXyCtpYYoUSGCMn0Luc20pr5oBKabRj0IbfGeEMoBbRDVNRU85Zw
mcDjSRXT0032/9bzh3RMGW8XwAB0JObctTmucncEbe2XBi2otI2VBQEHc2Jux3sZJysISqUHssIu
JLVEA8HsjCKQaypt67tAlEe9FAqJ9H3aR+gxSmkaPwqJHWQF0kpWbM+Z/bgCbE4wJdY3MvkzmXC6
fpsvLP6ufYWnjT8d996B96nzApCOzGjM3kPgBo8DM3CDI9a/rfZZeAA9cLiFi05r73+E91oru2+L
5aQAnskdSFmGd5wXHlefRDWNkKgeOWtfJMSE16diqakRwzHkLjCcRc7EXHjyTej/xsSAwb9OvbEG
+4nFpuXU6kaO2Vv1r8UKpaYmbtY3xgqfvSvqcRTy49ASvsbZx/SBqqDoQZiy4aStpYYOGgEjvmcv
RwqQR2UuWPoUrElJ64MmYKzhnsZ+V5z4bNcizyesgJJcK3i2YRewzD3n8i+qWIJ7NWNbPDEc21u8
E3LN9n8WogDqlZH//T47Jd0Pr43uE3T3FjOBisDqmmreo7NCRd+o4HR17ZhRtmLYZq9j3bgPPGVd
zrO1f2aT86P4XhTO+YkhhJyNbrAfJzsuEkpPNSi4F7d4T0NT37q0HUNMh3qg3asKbA7ig5AfXCpU
nLtQGLMg00TiQraZfLal6tDEN9aTMlWZSA/Iwlo9qjraTHJGK5AQbsYc37hh/cm6tpKLhO6QP6DZ
XEoKMIHt5Ag9L/xW8HfGqvHwOfxXMjKqVstxucbLI2bkEKdd/+wDuOF/6XtksOx8tETMvmXxHHx2
7+PlwiZA/HJpHwJI/E/RudfgbRwwuWbePno7gl1jRKGsKbyD5mVQ2+gSlS+OHHaIjjUs92YLxFnH
D6rnsutKzL02QdXC6DcGW16i55j8/eAFWnn+JiqMCGSO7LkNW0z7urBchz50HPEXJyX0I9VKZ+Kd
pbgnVY2R1om3/hx5dToY5orH0/ou7ZN2sDNy5RUIKTvid01ZRVUWxh0EtBiKQMgXZMgPiil4xl2d
T2doMgVKKW7XJoc+rO++mdqErlNEpMqxs4S9wgJ2QpKqjClsycsrqDmIqo5+mrNTI/25x/EMfUjR
6GXy0WJhh0LBdpi+2n8iCgbdknGQPjk99BpWGw21ufq+xP2I0hVD8mcg7Q/Pcs94kdHYMp4+vPZ/
4Gr83BXZ5jHq0pzyAjxEgatr/tsrn97YX5XyLioaToMKHVzppMHI0O8fdl7fKeyE0r5zvEBnlWra
zwPy6HSw3Scg88sllJI7TIKDPK6H/y50fOoOcut2a4G3ilqKa5ndTITmM0PWZ6eWqJoyJejfzNr1
i1oBHSW4Mi7NRdMJCtfdBeuAoWoUTwGTQkmDAmL3/ycKqskWC9ktJbRbnQL24sC8NgOOuXuaPiit
QYpNwlJd6mW+db51D0/k3QReF+6dTcTjD/BpvgEJvhxQZgDeP7cpFG4AoMHm0ZD+RZN1EoZeiZdW
9nhNSwnWq0Cyt8OI5hgZcBZbRk9+h3vRIZD96dwc3fmF9DK/nMqEnTwuO+JtAcENcvzhqL1dO2De
RdIidrdEQIB8boCp/lJwiHaXDite/i5ussJSDafkTL8GOif8novc+drEL5+UESnHtaulFAbWv9So
eWQVuiZNeAC65gwhPlcrz7dh7CzSIVkOvGqE8DUX5DKzwtJOFIMHa8S/QQtBKaWQTVw+4o/5I4QA
Y8HSFhNh9lvOIba1eV9t7QDeDSE8LNd7XviERvzc22beVZaHVo2NMfR78qekaZ19Jrd0FkEcR4Bu
tkghh7js6Jfoip1OMKSbv6rH+uYEW4kevdJmmU4xH2e5YP9lUZBFYJmyEl7sSo1LMuN7pEAgJUbI
KhOFD6wVGa3nxYqVkMSF6rAz+O6gLFO4IKCgw03GkK1UxzZuuNn4QNS72uf+7d6XOaI527ZJ1pTU
iyasxr2xYYoh5P+g/nOQlUbSZhKeGOzuUl8X4cRterPkEzfpaZQYUP1EefOvTaEYBFonXb0YdHlL
8lLpyTK50/z3TQ+buvdVt45c00qmL1/swQXsCboZJgqYjXVxLl5ytAHR52KJbSr/fiVP0AY7wrSp
/cZcKLWbf2cCRqqQuTlPt5YMaBG3cvhp9wk9XvKHLnXTfwlW7iRnYLx4zTTMPF7SC4K+eKEQwW7+
y34Ix8uRSSxKzBNk94MD7XcVuqmVQY8t55Bnvx2dKxRnIpgsoaIFC2+Eg92b4147xT8e25bW1KZd
BCIa9DKN/lV8i1WCkS935QtlHr4q0O54gYbg1l+yDxw87iQZ9nmAq7TrIzZwIYpvJaHsAHezzW8T
BaA0PX3o6njv44ef9DVPevAM3FJ6+3p9+WiTJ8/Xz6IJfPhzM/M5jONujrunNRxOi3i+nbo5IpPx
jTUPzCEjCF7vS3ln7JnvAS4W1oJRFdbF6X6DLhdoUv4xtpXIV5IbYJGPSi9SZSo9oQeGWANaiu3W
nFeFiFZj4i5Nbb6wgUU5gMoGd6RblPz8aWzwQLh3HtY7gtvJe0efVfsZbKFK1f8tvQV+kcCknvXF
vin479nQfmSlUpaDEDhpog5E42vnX8MnYPGpuAaurdi0OYoRqIomauM+/hqS0FRfKkVJNvL9CARD
u1k/5+B8/vvBtAF46GKNrfiPOE1c69fmUT+IRi6t7J5N3kcBfgnf5T2miqDyjHebw1kzvi4ghJHu
FI6FYMgkldfuGJ+NKuS3vzZzJ32b8CC0r18yIdiy39HE9R8lQj73WwPU6guFww7440kEhpgw1z8s
jkwA40Jx+FoSfVERqEqLoNSWp/Y5/2wk319oJAT0ehbDW8wQsBAUpj+W1bHl3RZYNTJBKrK5K2yI
f/XkLtUv9gH+6HbYuuaaz3LbnoYLvSwxLXUQqSvqK+m7OveTfmazhclFxBQ9fvbPMaA1Jm07iNse
0zFw4sXhRNlE2ATLI5QjFkCAFTeU8kLCoOkAt5bc7wjXAudZWOhJmABZM7OOpcAci4kloiHCSsag
XmvpGk83lZM1pw58jMfEWTz+fPiO1zg3ePZ/9poopB64bsoKcuGs9E5vNfHpPouzYtsX7kzDbpDo
wlDKg65wfFapRAl1Dcyr8fecMyZ/hlIRaetfQUx8S+8MljUlwGdBXgU7oy/jsZwc4T0QMn7zRHSz
7ym/Wz6BOHfjx0DfrVcVxi/gdyFdtujw1cEHuIVeJsE9u68mcUG05Uh2lQhUJOm/lQmk01MULWmH
DuWwQqyAYe65XFgNrNe5Q81y4+Bx0/6dfsMxtma/R6VxHEoyEobx18OeMXuYboCZY0LFBTsn0ppo
/QDkESSmhbvtwc1dI0ouinFaG17jMGdwZhGL7iZcAEJjQRxu4wmfGoq5St6z478DVy2jiEH/hbid
OVuhLOQfSrL1aWVQJXj/RiUGuwrWgTqX15epCqLs0+WE+KuiAVZyuWEnC0vX8V7ImIQEbWVFtlgb
Cql0rsn/Off/DMssh6G2QkA44wYZ4J1BpdTTIjgzunZqoE/zt4xX8/VPMauwMBRbaoJ+AOZulFBj
sORV1C48ZhPRlWhFIvslJeXW8EXuQWzR5ZM9umFV3kAqoWUejQrWbXu40C+zHsQMMVgmQ0olYYxM
qGEwu1IBsJX7/eVhjLhq0Syf1PbIjW3nCmjL30hBUWh1L8RH2aUFQYjfJNvX+laiQHCVbfATbp+x
gyAtExuHEFmuOHiaDIJnMjMpCtoJnWph5E3CyJH3Eh6YVWUl1Yk0gZEj7j/Sb71f8rQZqts2Ne23
VduQILuqmRKFGhUSeXKg+Iusiy5akWvzt9//V88jukrco0/I5NeReBsh3mud8WJ0w6uCZOYqWpt+
TteRltjCqknse+3aJKnJ8cpq0QJstWpFR9+iseIHg1mH2liK5unrbKsznbCKadxZ8mDSoGueiKZx
PoNvthLjKCatHZw/6mJMfi10mRt9623k5ZHxR6OUVeaQXaI/ouPT1Nz0jVlzO+usET4JXDvJAleV
w6nc///w0H7D2UY7yVxxFGlyN2DvL7GiB+OzgtrmHX3jVNHa7CP8CkLu8NcpySsH/SXVQr65gSMB
m1IQCYVytsyUwZtbxLV4P4qlaKU7MtyRgMkFRCrvxmJbF+d3bWJn7BsUcIQc6SO86sY7y9JzW135
oeiQSBrt1FR47y9OH7++MCf2MWdvCx8itdswHGrAjlXXSEuJlajhgTvMxfrdRyG3CPkKupmjjvc5
7I5Cmjg3aXlz5NqxC8GmAQDFxemRhU6JRIfmxE4P9TKP/ZK39ABP2SFhJmuv0L8+4K5SfGc0djvL
Y7VEkSQU118hZNPuwwi4YOHOYPmplA1TrKpkbiMdHKyBF/O57KfnToQabJP4qBSzEpy2CHZhD9Gn
9JV4wTiaCVaxKrRBJnV7LgU+PlrEDfB7QujYPh/ABpoLoItRryIri5SU7bctLtC6KQTAJdiy/pnO
iVCsM+ISa2gbWrPxP83KplLXkzLUlf//ux10C/ssmJSid8mAsXSqvGp+lRFReisnZgKqH2ieUoUw
pPwvbSuZ4x0Ts3LdFQbhlFTBWmgKUiq7dzlORC4RkdT/7LP8/3PhR7SX3GcjI2t2D/VunHYZhCWy
qi+VmQ+IAZskK6RX7/Hekvo2k+7R7ky0UtZCvjdkff75mKCfZ6AL82A9EDFj747RVWYtxfrMra8X
MtPhFD7VrJYDXYfz7a91FI647gI3Ml6Yugjv0or9s0DJmJrqz0+ZKyxeirQ2H0u3A7eedAx8+xjR
9Abq+jwyEI0XaOlgzWc34tWNKm3dJ4M1SnIE/JA3x4EBz4vuf56zNsa4s8+NdWxKqUFO/li2YDsN
0G1qgfOijYvBBpP0NKp2d7nZWQzLwlQgzALC8y4Adsro9Dq8agVieQNIbhKKUss1mcRaFL/GVB5E
AJ2DjsGp9jkOPP1cGcWstOccQzqU16jaf+dom1g1Afsi5bhc6/FCAVs1a62vfwO/2gQlEkVb1VoM
MkxyNHaunxkiW+0yfKZGSl1FPqnXcZcM7xJV2aXu5ZMZWBT8mbRU3rTfy1SNE07Joxh3IJLg8oTE
Y/JlGHPCqK6yGHKQJUSma/QvL6HxILUUdsOT/F2ukkZFuTpXlJck2yt3C0WVN4Vpk/Xr1ENqOi0l
c3kc8DJ2cHe0A7JthUQVrirM7Ix3hPVX0dnezHAtFEnVM6U596dcmPWJiD8I8fWxtKvOHkFkJvFR
BDuMlyY52b7t67ztKteEwHfgU48/ve8m60Ld9npkTTEohqTVhqAW1FcXGu+o/ZxFq0wvd3pSvBBc
a9WXFPCYTL2Ic0fNo7YZyFF1uOMEtLJqEi0nxOOOOuHePmTlWPDtnJDigFt6Tqg5sBMbdY7i50q+
s/L33g0bAS/mj0ZukNhnZ9mBvhTKmEtm+sL09JwAyhU9ipBm3o0XF717hom2DgHww8gctDEHferL
LaE3uZmIkYtTyatGgAVDoobzFAxGCQTSRZPuv8PZUXUgYYiNiT+YPQ9NG9lWs6x5Y+4S+9c0jFfx
OPFHXcXE21zV5z3C59PoDaYGBWtZEedL5Vamf4H8dzDblGdwXxwBHO6xntcAmAbo2FvG0+W7nJE4
8B5gb02JXXiOge+xrAD7IH8/wBbYqWrIrJdLKryUDhabqybqQoMlgOtBy4BrgyqvoTCDJzRzTwy0
w/1X+kxNz0hGF+mP0Zih+plPNAAvZdYq9yycezAWqM32TrTc1zhhaSQsl5MsHwBOoteWekv9Q3hP
CrJhu3P4cclHLIEE2FOYVX+vyOhvutyjTZZDicY85T/dTG3Etux9LhHVwlLINdUnCRuiD8tXSLpO
ULBshyaR2BICL1kCQ15hSHZ6OIC5P45vHROejEsoTSCkPtreQvxrvocqZZ65XllzdFy8L672gUdg
LHNo43OVsnwlW5MFVfv6/GMyqXwSCCtqPuLJ2hxuFHPRDhiU9UM4zLOwdh1pS3A3fBAiC0O9w8j+
ukLW1uXGHft3FttwPW1GhVOUCrCaWPHxHGZnakWAEEfKdEdpQw1EuG72nk9FKmFpTpuGVa6qLGec
nJqXn2rgMVHWNM4yjbe/sbwW+1t81sqUy9z9yZFSvaTS93iufOYj9kP+RnRIE9NHh9ScI80FXtwk
koooHFp8Ajawos4bUBcAnN1PeUGlkXnBKX0nyi5hBIhQHVAsTxG9v+UC3e48RuxxY40KgEI55Qph
bciTzFg++ji2Ta9uynb6RKIWg3hxTCgBCM8tExmnCoO2cFSooRoRQtAkx+dcu+3QdOMCmVUkXFpp
YiSl18tsLc3xE+Z2DVuAtxSZRSUJdYY/oNAI83wseq5ZJv6cpFMdmndodFHbLEjkfiqqgkxZuSIn
0BQLMMd55VUSIc8PvQztAL73JEjcDN/F/JO2TPbX49wykCVG1XKpcIvL/a/I4H5IuWQIsksr0ama
IuluvkTh2ZEbM0crKXxHyM5cOA78UnMwk2abbNTfAgckOvAYsMz6V9wK6LCgHNBGA/Gj26V9laKS
pC8X+YfR8iLvCYOC6g7sD8ej5NCz5F3y27wIyiX6eeVMAfomtWF/Rm/n1EVtZ6ut33c6oRsuTPDN
InXS+nRiO6U1JsUIF1RDpMICnlFJzCks69f80u/MkpnlnUllV7Qa0kDiXD3P0JL12LvF1cXogwjj
bBcdgVFYiMVhjdIt5Xrzlw9s3HK5/Pvuh0UGY3B7zkMfyCgkYG06sWzyMNCFM7gmdR5tUizGs53j
4YdmdCXzuhqZ4YLNxt1rVpxHoYXgjZYv36O/MBcC3TkR1NwceJ2jq+kcr6f6kPuV1ij15BryXBOU
s6YkVZV/Q6/SVHqbLFK4l+8VLyv5lsjZ/giaDhNzFlhwOxOGBIn3Zm8aGieuM83hq1iknTgZJ2qk
e8UZ7Xr/6h+fBLbOOq9h48bW5l7hlhDnRAbBL8eDiboAQPmfXSa3cO9RBsZAAt2QViVnVu8bnSN6
jA645EoIqAi4SsLnfsPD8HDvfGfbNPtMpmXQbK5w4tQnhtYXD7I8h0vozJ+aXVDymUcH7MlznW0e
mMvPBT4boqsV+T9qdu0AbjTsKKt2vepo1eajcIWP4K7+3oFQHCNJ+lnePaASL0m+CLDi68eBMQVQ
fD1LnPHwm1vGTFMNHw7ssK6hncf6dpoqqHGcMqsEw7qPrVvoOrd5MRL3VDgwEJVsagpOjiFaXqIF
LU9r/0E3a6Ukw4s0uW/Qn/oHTLIJeGIB7vn96U4nHN5nWBUqoemVeYX9kAxrGHiL35RwDxcFBwHu
NR8GDCtwT+W77Y0M3APyE5dkJpzYYcEMiCkgTxnBHSDYnnXiKzHspPzv4rJmS0iGvG4BcEyWxoes
WEpZh/rcvTwEGYts6ENZI9av94R6I9lBa+OF/Pgb0r55e63Anpyu627HjfLq+VU2TF5mA9QMt0FJ
bSup7wUYQRzUQkKB6EKkruyRdt30Gw9u/hoa5pp2Nm8fc8sCOnGyPKImNG97Q62UTrdA4t4t+5Ac
v5www0iPDkWAUz99hHgQCR0GuMvelthL2YFhK/cRb6pi90DR2DNQdcWBZT1MX2UveYPxTXKd9Smy
5l7fS4dhcqwjcScoNxBAlnSifQwg8P169iyqowStzGq6+CbTdXkgaCpnzPH732T+A19PBp7uEt3J
ZRDBMddzU7fFUzxELizKm5JTKR9YLTLMknkPrd/AzQXPReLalyx//skXliIsOyPEhBBVCd9QVMov
lGAydY2yHg0U+piRTiDyZcJDf3M4wlzhc/Usz8v2D3JVeoTLkvIbh7zXYoEiZTtVh7BY6txFR010
6FcHcF+kF6ts2d1qDVUDJncMY0CTqovia4rHP+4RW/XcZBcgbANuaMp9TzGNbUQl2zq/mm53hrhc
MY8OZEMRsQzQvgt4EyZ0ExYGD/0Ai6Pp+ni+TxiG2Oa0jdzRbWIuYPNCDICdgWXzFhp7+Rk0OoI4
/RYw8+/SjsYB84ToPOf+AmTDLVMjI1jbw76s0vIRXDce7jI3Izb8oyEJ7Ll0KwPIy44nlmWwD8gV
WSSDfOyLolrNvEGU4uNF3FSVFrzVQyWKpvzFRCeS+reqpjmtoSSn6144r/6CtUvZLJ+PM5Y8Sfj9
NEFoi3eBq1kH/TqrcJWJki1pKlSJLjwRCBrXobYtfBpbDfZXQdZx6xShlTd9R+NdYICD7byeOJgY
qZR7RzmVgcvmJ8JVxFekWakeqOnv1cL3hfASa8lPTe+wv6dRtnfM1MTffKz6S3yqBYFNWDBDNiY+
lW6f8cMKnh7wvU7p0vCm57K4gKT+7vAn+1kq9/4PHKU0tKcmo29FJ4jvJStpmZZxSU118kvOq45w
XVBL2YnFWy/fhkk0wu7Dgv94AfNTJXSraojqPgAa106ntfS8GiAl/M1mCZffqpySJo8gYWSQJT6T
Qbs5iOQ+aPo7RgR3gbRlJRIg1QOvU6IyjHQ6R7Q68D0USM8SqBR37YOyB7NHJ5ZektoDASay7Ux9
eKtzQKcmSxQxr7dqMmCBlQcjEtluNDjuAWOITczH5RDATV0ckWv+beVp/r+Eb7aHuJsv0MsJP6F8
KtSSSC8t68mVlqAEqq7KGER9m93vpoyHLuMV3xzmLClfCEyen9qdhOTscE/ZE8n5oA1QDctZ/eX0
fXR9Nem6Bl5DtiSNpkrXWj9gT7bB+szY/iJc3lfgykOXYB54mwVcVcAS7MNBnmq7xxBa7FOiK1Mb
XvsSfRgkUkBW9XyvNlFB7FuEqSd4YjzvB7/i93x48sHGHpqtmh+Kemx59s0dpzr91acEOCpGIJad
rxmDdcHMlZRi87Mv9/zkKO3eMJAeLLETQqDK9v2ryA4PlKGghWjnkqYYmvpyt0IR6T2KYRQ5XPM6
G/vMSghb6Gwakvw9uSaZ6y8AbWRwsG/b9PuT9CIBrSDMIW4vnzjmfwh0zJHG9c21Uch4Z9pxLkgi
FfgJL4xSBteH17INniZBFxdOO2dVcsdB3M/yEGYlaxbN0AlKCIwKqeETedZhhU7PjxD4CBuAT8+L
JI+pVDUNAU7mUq4WN8tA0NrRTb8jDQYp7Vy8KSQx1BMbZjme/n/2hnpPL+saBvyA37uhpu46jt5J
OZf51IhNMihvwkNh7nzz8T2GW7dZQPr/N5DNsLf55HueFvBAFCMVpncwetTqKXEcaI7i+OimcCwo
LfVGDTa8SEZR0+W/KZ0OeKVbmRjRxQpiq6gZLUcuGeb+Q/pD+zt1gXSlp4wlNyMH81LRQoiQ3Wea
H6u3S0xFuo31WCdsBHl8o2CoBrBH87dJm5+nc7NmdoE69vYSSlupfRH+1pDZHELfco4ZI6NfRHxO
vW1fC05H0qOVK877j6ZjYMxH9nKEEEfBtCCGNHssWYc85SaDBioaM+RTue81XSaYxvINe3pCeULQ
vp0dgRPMP1R9/Lux56DBShpmkvDDtfit+QLdravipcpBHq4RaWlIr3V3ycSfsaJYKKGSteJPZzSV
L9525xgNV10yc92dGNRuYtkKTimEveDhaiBeAknI7kO1/4G5AacL5x8M9Bn7Qucso0mbULoPiaD0
JkMo/EKGstmsBeRnIDcm/X7pMGNXMPahcj8issmU9IELFrkoeFSsLAl53qHY7SXMyaPXgr49M9uI
/DY0YgEtljlWOhOxRfFweTt5wh3bUnmcwSLPj4WhqSS5crUBsSZewWzoSNkuXyKTW58PSLuh4LCs
g+8Ugw08IijG0PAwTKq3VcPRl3cXlmNJkni+4gLHNmhdkPkmPeOMFGXHieziBUNW9zR0CUk54Tbh
mW5Vnx8bTkDhnpXHxBfaZMjtzUdqT+KAuq5/b2KNT5UhVjTq3HNXlZSmln56TXGOqeOSbshFDNXZ
XxsYZMbWgZ11PEkv7cUQNMzpDQgnchLQxvlxkjq3pIP50RtXtwA+3bRE5t1Nvsi5sBQ4uyw41wW1
usQDqp7G8of52JySno7f1rbo2ctAhu6+1D97vDo0G1DVDw/fjEeebpJoE0nhphTf3/sA/+bLDrL5
iMI6BzLHlpwrQCpD2WQD8z5VaVHTmoFjsb6r151YJX3wxMdiKfON40bb0orE/ctxIWM21Wi40CaN
QGQjMbR+MKHIapbHpalm3C9YOcBLy+lMSOKtmIPYlmYSokbj5CCDeB5JM/2uAD2WmRsXl/c5GjrL
G7A/nfMqau1SMRlfI7Hl35fuqauM/G8iygk9GXddPxuhVlxOvjbW58uv6Kv9rQ7KWnI3sBSIGyOD
RgDXURzMvscIUJTy6wllezdXRMFbmKbFkGnlA74QdU+klYt4MsXzPQyOZ9peW+dKfhPkji9lQwzE
33gh6cpni8EyztBgv75GT/mX4xEBYJ5PXs7XMkVQlYtuBr5NHzSKPnrapkwme2rX57a0zRdhBk0Q
jOpbV5c8d89mB6jMQRClBOVB8RxI9knjj+YQKOWwwT748HFaFn/PuRlC1pTWWLdTIM4DzOoUJOXt
5eBvL++p/PilNlNWqTId9dsqRdPKvEH+dC1AreEj3glDI0o3HNagoDBBB49aFGCHEqtIJEwCYFXo
UXcHn+KS/8gUCrDJ/cdKmGzLDfMshmp0Oo7VLBrcBpRSTGeVAg2eet/Q3UzpoBYl1v6hKeVywLFU
cVa8DGxTRSmF5jX4tZ1SRsVjZ3o5eRL+7FndgTtvULatg9q+EGet5wlaNN3og85UK5111Mo4IfwR
xMWmHCXFp3R1ioI2b6sniHe7k5z8vQN4z5uzQrLFC13dC4bPFf39XHuLKVi1eiDmj+obl16VeGFg
ethgOCAuDda/V9sJ3sx0/pzybrndCF5DeK9YCSvLa7Lo9DJxsEEr9ZMp23c2Km6sTQ2OFQDMpLKL
Hynvf+w73aSpARmKZVn39/+7KgvOeRAHuzSNtnFbtxW4ZKkhtwLl2uRNRq7TjJxkbwWF3lOx0Dtl
VarInXgHPfSfBewutLTmjS+30KOVSU901efaA6ONn2Gu0EEUcVWsH6CDFFkYg5ycq1ACWTOtfle4
9Gb9kRBkDWZydx9SDK8ErdEplVQ1pjQ6ZYHL065grdfTBLX4RgPtL9ieVAzFrf1so5dzB8i5BgiD
L6uvR6ZUe8t78pqgTe+yk5NHxrPkYMQcBJibk0ns7UhWSi4qjR/aFSg6aOvBj/9RnHZJukPzgjk6
jU6zonOfkD2m4rmJ7GrcT9Th4TaYX0CGsWH2IMim600by/ulviD3OuXVROjVYq2+p2Bef+ytrzky
OMFJk/AAOGTIYNx3tPwhgrkq1T2R/Rz1U3FE1lEMQ2NUT/28MV2Eunhx2g/6VrqOmebHXnhfIogz
fLW73gQt/UAhGExXin5KITDgAH5L8AfvCNC3G38P9SyOX6g6ttL63PkbppRQSYVww+1ShWg63lzI
BdH4zrFG/8/V50vFK8wH8LP87IylDtWYIiK8v8KMlhLMB/a4T2qSyd6r/94LqkAmHOpaVxV3vF1O
Fee3arvJAcoVWaePNV4fP27fwOz+3D4XrCg1e+E0oeK7bnW5CcDaYzFEdLO4o5bXmiPVsejeXOKH
hG9yE53gjgnUIBRvQ+kSiBN0X3nVyT11zazz7cuY+L8/9s0ELGAKyJACwwNmSjLiksybPJk0jI+x
wz3vQdPoKkixCnW9wp/JwNiwfRC4ER/dFHk4VniMZ2aa4aRiaYkctAWeXSJecC9pkPBxNRZ7nBaX
Zv7Wxx0FUARoayuVa29jcyAnYlVZEWjitUhuHJDnrIc5i2dkUvCAqeiNSuNC5N5lgrn6ZjpSgCQR
y5JBoD9R6padEN+ZESJVtyO7xC4i0SfezIyNHYjnHELVv8PmiW4XXA3pgNo72+pYRLOMl9TFl4wF
A8FuFqd+8v/MxcK9s7C4w4NWv0hRhmNzeb8bCVIPmsbv1mU155d4EhtsdKxPGk9u82m2JKhFWIBX
BNG8+YgAio+iB7sAlle/IStHPfcc7isRKVrGC9GAiT13/y6mpN+OXmB19Ly8ONmabO+KhxsUvmjr
Lm/z5RGY+KjBIhFt4fWUh4UAEQdU5suMPFzbuiVy/xlXHAbyCiIea2Lgmq/XoFeucoFLIZLEmu7C
4kHuVVNuUJd4TtB1aWL9Rh4LXlSxUJYg/Dw8qasfyX9z6N7kj/AYK70fHuMl0pMl0gzBKioT8pxX
v6qPqhwTqwTo566a3mV2XUf0PWqMPqpRyPmfWr6kqbnGvmifUwUYZdcCTcwW3LtLTvs1NrMr0VsM
JKss2PRKHhitkPNECDTRDH4lOElWtxHHdZemupucSonW0dgSlh7Y1AVMB6kjYAWcX0ArS3AiGqG+
YofaHcVPeCe4NQsbr4zp6d4f4H4WRZY7Q3cRy696t4xuSkOXtzZa14Mjn5tP9+tCk1veM+hzlbaZ
tttzfQtFHKpg+FjkU4ETiRQLu+3+U1vwYbg2tCISnNm9ivl2oGs7LAQCVq+F5n4yd/pl0gm9ZpIH
W1nJe9OGA63GscGSkufWQvJg0wZ4zQGf5kX/+cMHr5dukI+zkZ2fSnhJ3eOyooTPfUgjzC+C2H29
29F4sV5FzqQBAEYQjOIlDcig5T42cV8cMkByWfZIhzWzhb9S0smtc/YbK/V+jQZVrKIBT1t3D4/n
TAZU6nhtNGmjPbxktUhla2Dq/XeOreChHQpZEmmf7J1L3Dv1GrWRukNarp7KLpCb/R63J9rCthCM
UEbIGLU1tfTy77LgG9oTi10nwDVbpdmOWv+zfO61ZFa3fAe0XAowo37u9+72W6G+fzpMAhUHvSHl
qpPPNo1Nrai/bqw6rUAa5levpICkXVxpKgFhmNm89sC5ZHxTq5034SY5PrDX4ZDhiqBy40ztgJr2
mkKZ3PhYzJX/CmnzlTu5/Lq/aQcrsen2h4xQucoI0zWOeuUoQejMIXcHolr/aOUZm5WZVnwNQL2/
mCTlQdTMUD3Qm8VX9YUkTQx7xrxtXFBNXKsBPRHTeMJVXHzmQGiqk+AaoCYtH0FevHhgyu4Mx3WS
iCzGKS1/PXIcxzjF5HdvKSsX1reIUaRmYrVY6PApaFaQsM5+ylnggkxwzyUDSLyTzB81R7DGN+eA
Ff4lU8OHM57RwdgR2BlYrwO7qsjCYazUjW5CPvae6yy6Z6LdgECw3Lwhkm0EwhVyLgR5zin/ee6q
uHvJeGovVBvjvLS7yZ5wVZ/u6N+d5aQoXmN5pF6wdDH1szLEfBDDQGjUVTrV49C18F23MaH+N2eF
GniccXhfkMEuduMVK0G3jttMclZ8XQ/exyWjh+qr5YCEhqKTeBMAEqFcubnokvimVk480GH8sjaB
e6Ri2pGHnPiBtDIcHYypStxXT8ASjJK9WsvUT9qcQvyxbWkvCMaGYFcd1KRUINoGepA4aRGsBM1T
aYolMPcsL0nn3zmRYAvSKj0nIoKrf9jAgcmZBtoJYvp85eWFNg9PXtq/KPG3EzmRgoAZzpm3Bqg/
PFwK6HEcSTjMWg2tJI00uLhWd+uVptDMcTUIA0BN88V2TlvM6fEn3wdWAzcioQksKv4l6pPvpnbO
N94NncaGEjLkUSWEO/AINgY3Cslf5qwEYiV4sQB8wPcVFvJZtEmJ4MIwscX1PfLMfbYu09XMdcwm
B8gip8J7vvyBfIU3hFT9APsWwiZAqYCXr+Y2eWjfYUWWJhFLohBqo+xQuohZ0fdB3+pbwzuUdoi0
bVhN70ZahQP8srnOjaHhNnvjhHFkI9brOHqDkrQ5OP+ZThRLCok8dQ8E1TVgC9AYNw3i5tK/V76g
11Cqi/UTGbM9xzt5MRyp3rWv4oRsmxq7KmRS35l6yZLGmIzGnz3IJ+iuJvM/yBkTJad8Xre+cGlE
Zxae/YBkxOOMBRm+cdDJm6vbV5DsiAavbSAwLAM75PsxzrTxXQ9If3dzaQDKEaxJjez9EBsy+fBi
mMUQB9/J/G4N4DZcSYhuNTpoBA3UO9+B98qRQrLTIKKGUu0S+oXwFCAIv4CTarjxXG4Stoe3Op9V
OOz1VULe8f369v+M7cA0Rk7ChRiWwq6D0BtQOR3f87pSGW3jwdmghUvWocct8LA7LsSohJuFt4uJ
NrRI4XtO9m+8hbjLgbZ+8PZtZncGkNqFBAeq2l3TYMJv6F5uV2Ek8Zmo/IDlZXq00G7PVGhbN77O
7czOce/nioccgelWz7j+AI/vMI0jhOWGMjpnDYlIN0S97obnLfqgnWyLkI9z3HfxBwIvX3uSSeJT
q85AQgsOhnV9DqWMhgXM4Y0jqJNMqrujzzCZmReGgzP1EsN7f1DB2fHCX32hGY0ONHKjuqg1xCD2
vzjhcwtJtodpJfNkJ+svCYyZ65jri2M48l09VOpcovCJcI9bNO2DmWtNbc+JZ1WPO9o90ZZbMYeJ
fGoEQEXs4JoRVN1ldNChbvkEIFKP75j+kQBJ7RL6fh8HAfEVWnQ2JurhVKDq1yt57bHbfN/aBksH
2bomtmTzTzyvN+fi1/iIdYX1qH9GtyBcgmqre5u0dHJRlg7BKMlOCAULbUMzIQgyfgZACI5OFye+
49ccb/QXOkXP2q3W5S62qBViwL8Sn3CjnPqgvYFhxRkzQE0iuFZ+ZjfNZCKBEcIqDL7yYTdHdh9/
tNezP1+xgFCPBpV6rfOy2xQGmsN4JBuNDjYMGopFN53huJ9WOTw5iGcs1Oqg7WRhtNwz1Ks/ekoN
hwaALwoOYI/3B5KIxTd4wMSiuBwNeD38LvO/2XYr4fMap+qMtnhgYBDwmpcZSetkviU4etRLmrYO
Eu9jWKXqnBaCA29zFxwNIUZpggdUg/wBtOTzOX/6zc1MCSWcAE+6K42OrLMO0GqjDS61YK7MAkS+
3HhkyeHRpzIM48iHVezkxFg3HONXamocmsj+2C59cKaYNtwmamQx3j027B3pwS7mrQRhoSJs3AMm
iOYfBYPWLDK05d4YtUcuHm6u2s17SMNkRXK9PmJr1zAx5/d46PSStmQrz+iozMRpNzJWCnM7kaky
TBOmxZx7wlAdL5j45ysvMDcpvgA7ugcPBQrhDi3BMc+p4Ymu9LBA6UbzZUVUYLSkwKtR8q+pt1W7
xnBtocUITB/h0gQocNRNm8ULBVJLKRfkGN84Xxo7XosqXFLrVW0kp6n8RNEyAbyVmWYfbzBrdc4J
6x9Echxy0XW8jF5WdoylR54QRT+pAvh18/Mv3cCer06LMqwf/dyfLddBVu1Jw3ur+TExIjrSa1or
G1li41fPDErCL+9aBf0Dnp/upXOf5njOzXuhn8mhNt0jVfxJnN+U3ZWmsiMdb5Anf7X8E1GcORLM
yl+Ej/65M4eFd9pleH6bObkNO970bjmfiCk2BU84CrseEh+a7Wf4Hyy31nyR5RKt33TkBiSvBlec
0V4V8i9OgW7capWxhJ4/ma2XaCEQFgyzksylKRmzXZshtqhFPLijUbHHQ4vFu4zOsCsjcaJXxpxS
epu3OI7RLQGdohioXcT/cP+zbmMKb3SpVUF1+vyWy9xa6997uGUd4jZMlRjEnKFUCFvFOt+/FKgO
nlXCZ2FCUHNZBKRlEhkn1VXGVE7+2ctf2Q9SWiIMBQf9qMN5cnrEaqpeyZ62NEiXGUufl9gO3i9y
QNxDFve+ZcIqrehWATehzrz/lnuH6o2/c11DcgxjUAHqxpuGWewE1zcg/KtUYr2wFiZ2rKsoAUSm
8D20jCV96g3QYOpiKogcvj11wbQ3UMTMEL5qWklKQEmFQRB4Wngig2DgS57+5QJeGdf/hqIXsGSe
c2W0Ubr6VQgLt9RaHkVWDNxcfNlYM9wY2TTNRwLv6pxIUYgbKtTFCFQXS+c37jUkNc9UP6Tg6DnG
zN3FB60ynMmsBhLghoPkd/N5muWciYuLJ1wqhs8WeOjEAEWoBWTEAqb4tXHO7vB2s06kM8lOd3ML
hGdARsh9cEYcYwNCn+j+0BQS7gD4bdD8WcKNT4oYGRjTtaA4xLHp/1TJQhj81CNcFTafi6BGWW9/
IFV+H8dMg0Jc74Gv2X/Zl0wWsaBTMeCTP49g/1B9RPaqj0FqEfDYV/s4z8I0F8xNA36JM1SR/JBI
xePF8FRAoLojXDDh1ZOly4Upes9C/wwkhm/270hFCq4PAO+sXH6rSry3smqhapDiKl5PwE4qI3zv
rR3vXf7YwJlIXNab0zxST95FY4L844AxUaZtYX5c+g8CAjZuyOPLuy0g5FpNhgVf93SGbhRIvKjp
zALLAlHZ6Zt4BqL7++U8MR5NATMqF51QMEY853nVkzgI/FGusDJ9CdYumaMPZahyg5FknVuFl9Ys
3q1Cn1VPTSbObPm7hnDBcDnN26h8wN970wQW9ZHJ3sNTnHKXb/XtABn/9AXvBX2AuJCH4RPjyAF/
BxJNXItT6+jjsuE7rwMCPrtH3IkCv2Evkh6xcqbMBkiw0kkO9Fj73Bm3d/91Rqpf7ssTev990Vkl
+c6W6VifxpoHsNHi8kssEV7HJiv2El5WTnqpko1lFRYBcWCTZUmEncxrFWUuL4zC6NByjmDgD5Rn
YpQr8ebhNzSo80BgxGfiasv35U2/U+NP864ctCCBqVi/72xNtrBdiXM4yopFoEMv8zJD0Y/FN5+P
EW+iDbaViSLM/3Wh5Pg933fquxIjVzkhAMLTkhK6fGjmRO/ug5teO396Jeg4IMRm5e0YlbqyS+ap
G+LuVo01offa5SvjCCa3emHVEUezajeqhv46ZOj0am9wf0UgyeST9d9VJwAFxSOFh9xWTk+dW2Si
5VJN+j3peep1/bH/AlE64jEZr15BBPDaUFcb2RXeVoZCBUB4G/CwGDqOAnvaiF1mczlYGgFa46WM
oLUtYlJMG4KCra0M3sVzLLBgd4nj83w1BUClLjSbBFAh3uxKYFlMPh2gwHRz3X45BX2M6ZwpFw0K
8JQ3iFs6rUXENPgsZ707GgoAYzqNggncN2CGVG9WvSPcn4XQx2+kNnB6jfRUgYsuUaO8VSh2S20S
KxIEnt8O9PZH151VNv4HVwrQ6ScgoXwnErQzFErsKqyvfHVI6jk/XoviEkeIC+z3ycfHV2wR7NA2
AHMOmC8o3q5d0IxyAfFqt/BlYkchsxX/D8xHPcNZYyleAAq9TJ4fMM3q/QmRGybMPaCkNtCe0qmo
aFEVOerBiJEu2Jwba14zv4ke+NaoauXcrenjkn1KCl5CeDLUgFdhyeT2/w0Xc7tKRb13C02Wv6KS
9JnOzmqQ2zvin0HnEHX8IvHqsRRuNFQKo/RL4/5Bvgk3aHs6D9duTBILak3cuXYk/Gm3vGMShnoH
jCibDbm14kblrz1Kx5PNMMMDSrSN4tqqaaXHpgxpqBd15joNRHqnsK4Phl0wv6qO6BJ0FKTuz2jT
DFfcK5WlsIQJLK05xIiJAen+9aO7FgcShYGaMatqhbiBJ8Ju789U8nGaznoLwBB2FXZpunHEbVw4
nUt/z+SiGBCLllIZ4qLw8DLsbAcDeaR3rmMT5XSCYjoG2PL7goPzmkyJLDmN0QIySRdNPQg8ERGu
QEPWHIzSf3bIrWaxRPPlwk/GegHfsYGkwESdLk7c3bT2EiteWKajOV9qSjTUbdnbhuOrf/gdLYlr
u0JrY2rSfN7kf2Pd3CCpf4qPasOYi5hAoaaaQpRjezYs+kuM2kB/iJl/Bq3N0qEpwPiS6/4o8a+J
uaKACl0gtBR3CyKmUMGfkHJbWkJ1Yuco9XLRRsVq1L0aMoiq7ID2ufe8iVr9y45wdJC2p8fA40n9
UwJf6aFRzMQpdm+WotUohnDcetiUVzBIT+ZiJsjn4L3GI69U3Cbbl/nKimqzHZUd7oPy4mPf8Pg3
mAU38Hq2q9eMcWuy4YOv+yZtUIOyoWgBp0WRtjhTaqgjM2/DuBul06ugKGrx/8PuDr7Hko8gZzsd
bKEez4pIkPPPOWy7GS2o4Sq9CpLS8TelblcNFaEQDBeDWb3CxoaTGAoFeYoNWwBXP5olW+F90KBB
e3dEEWo5S0KIvgnqmvwaW/dARyfmGNh296GzU0B5/yD5HCuF1KnREqlZR1ZwP07tcP4wpH731wPD
50HZCYHhxIqCprXXkGAQcLciPX1gtN3OTiSNXfubpHr/jqthTn+V6n47D4ptekvrdrBlbdmYmjkC
o9Hd7ww7Lu9jNlcQEQ4Mvv8EyVNxgeHJ48GREu2ZinBqgvFRdbLiic8b6JisqWzy4bnhUsG+hpkJ
pEK0gqGtoe9yVm0oWmax/hrfhhONGFYJw/ShtTiLtcoIYw14l33TkhQoavtB0LWdeeH0WPsZSUm/
kVC3Lojm7Od2mw1hl0J+r96KcqN0/k+7ICnX+rzsvyVrOCOQ9if3+aLtCzcoGHpg4+jEVoiboyi5
zAG3TCnjbwouKW2H8CpbgQHuuHuR9cHe2vvqPzyVxQwDK0mJBRtk2/pttajLANb51drqWPDQqljA
nitvsrpOyyVj3rI/MIH/q/oTaaAA3jqMxhoU8Vj806e0FNGx68grdgMzyFWNWujcvMKba0euCLE/
P/35R0vMfnMMlb4T//QvZ9lOguUx8BEOLrzek9Cdc1HWUl2Gm6Kgz4Thd2uyj6ns89ofCjOK/5kq
96uSMGxhLAdMpckTrUQ9TkKoVbEKxWkBHAdzpBTwFM/dCR+73mO83RQW8orPhipW3kAC+3SDolYQ
+od0JofT9smdzseVqmmyMH7DDR8OvQA46mjScYHhpzpqAxcAXunYXLu7km6aK4lYYRurz5lNt6El
BsIU7ex5QTmVJFakMN4zqgeUg/CV4PGktzzM7T6ZRhVqjHJo1OACr6P4dzIRVLd7GzXgB8F72XIp
0irpstnDDsl15HJlnC6Tts8uKVTznnRZpDyGGyEmPur/OY+Fh2ocKkEnErARcafowLHSn4yqiTga
kK6Bc4xlHrQSzhCDgHZPUWBw3VRX20hLgPeWih8TNjQQtk0KssbugnWVy0Vrkhm8Ng3t1lMzgqFA
XkXLvKLmtfwRakcA37aMdahsr5IPNlqPEzqiF+tILifZg72mZctPo/leRLxriYR+SXhKFuCB7JVl
iRadvbOsm1mKsClLwLZPmAPBWz5VLE+K/bXElq2AylcJFg3OpnEEKRyC+TCMh7DmqMk7Q7TI2h+P
1B8Q9UU+I7n0jFQYHZ7ZJxDZCGw0gnX7Ei68uRAub0q3Hb1Y5wmFLLVzXvmsgW6RRMattIvYRlaF
X+PHVw3lAY0dXOC3pqz5f+k8A0RZzUd7A2BhfOt37q2Rx05mxbQPn8mMRdpxYmLRr3Yl7hKUIJ+i
E6TqcmxX0xW8x9o5xnxW8Ii4YW6SpmyvJuQF9rFRKJh/G/U6O3RCsNgOdSb+bUtrIiIBp9+wyeZw
W4HmIaoqKwdzmX34WVp4mPbX5lIHmxen+pLLZzRcm1gv+MZtG51nQrCQ4002AWBXonXS/b5JX4Fi
t5usXeL20O+GoucmE3ExEo1sU2/+nMajYrsw29PWuP9uJ9mvRZdxgA2IKA3aSt7zcSXIuyXbVapA
y0I5xPcTLMkcPh5NlP+yePJxjJp8LC3Mr8shwShawv0AicJMLFXWJBAzAjq8jBs5QIUzzjLe7Gpn
4Jg0PDyTcZakiEWPRnKGwYKvz85YmHnq0vq1rmnRnR4I3MDlCr9G8cOvwOevznYK902KdKxnDF7C
sHwj3d9EdYK7ALgKZzm675AQx+e2NzepBjd+hDZ6MMJj+loibneJfNl4yfQYK23sSCaTlP5r7NjX
KQK6tfYFcBctJ13fZDbgrjrjlQ/gDUzrVz4CQjL8U0vyzDqnRZFRbuZ8JXguQJ/eXXG1mShxswDv
xzcRzpRWhZ5PX1IEIYmqPvCgwTpWHGuK4nhxseYlNYNTVbBq9jNFIV5I4t+2uKTk83MR5/zhTdsd
bLzdXP5DK+/7sWoWGqbBN4SM7lqgJSsRNcKrfIoRjw9pmMyScGfo6MH2uQ0E+kGowQsLTPRum1Uy
ysiGciBhJA48u8S7sMQqHH4hL3PzzO1XFltEBmoExPGUfvo3w26xLzbB/7bLeNVR6RGohhl+Y+dI
4+VFyTO8p+Q8iq6qQ8aD4PlFrYmeoALPs4GBhPinKF/IgPvXMZNu6r3PS5exKw97XjrX2ygr6rvs
Ws4PetWJzvUevFK/JFszbK8z8pWtfwlMuO1ZVZNvWX3LO2QBwJmD1NansLMsUex+NvKyD0C5jbBV
VtxKAF9ZMk0wpcadVTK4LOqgoL+2b8TZvQmrIQ9hN2zasYRoD2uZPLEytaR+iWqUVUGiLzNi9aUt
JXxPzS1BiaZ9UZAjZypynzzXf3BVNWGJEPL6pX9qtI/jBlHhCWMeA0gCHk+P/p6T31qHff/e4F+q
XJW+HmyEI6P+30lhRRRElX+lyHox0Q10y7wPdpNn4e15BZZWK/qn8me60j++reb5/+TG9CKxREpA
9rsm5o01CKx04rUQjryqxDzr1KnM+VEEeoq+pZug9Nm07VNl4jEoybq1Hp+IwqdPMydik06jhAni
3zuCxICA58vR44Rgt7vBi0cCKudT6L1wjZOAGOOKHK9LhelPt1owVCuztMRgMyQJ6eIiwSgATinA
wB5QYJtZY5jEbftVlRm2E7syga+nex9NO49rgEDhryyEPVzQKYWhYmk232XBuRrcjG1wM7Pb2Eg6
MADcVodyDPMQP7hxkkHg9rsoImhXhe51HuAFX/0TfextegDmtDH84sV1BRb6Cb8cOiwIgTtGt8wN
9654tb7ZZ0Sd/3hW4/B4QGLeP6z0TkiOBaqREq58w3r4MKz5bZxDXPUX87DmR3atI/Q/Y7Kmdnw8
kmUhvKQBxnaJDNsmfdc4f7lH4hjupHOs48Pi5rxzEdPdQQtq5/m27K4vyf0Z8G9v2hQOTG9big2Q
oFM+/m26dLgslI7QX2lI1a4yrDq3ZMNZp4xrtvnTKYWKQgqz6P85UtwOIsBzbHtaYicTJXBRlEle
sSr+pmKfPwStCahVnFwdb/Np+wPSBszkXdJ2NQAelaO+vF8oV7in1wLfN77QKohgoyxBJriTTuBF
paLovorGp+pwGdCaxBPEmS0QQYwHd8HTHnH5PlAZR/faK2jMt8UEjrJhz0H2WChkUYNzZDkG6k08
uBL0Emk/LE5VL8AbmSDW/Ug0OqNYbWTCK2ZRAuZxZ/URtinwCtwAdaoKW+TqZ7rvHu8oxlUvZWd7
B44xSMxeuisIEepzAdyKYhlYVLtCiTtQHDlvPWrCipWcilN33WRdljR4TvUp/q0f8chzCmcog/te
/St2UyG4C6ZE9ajPSrcVc+Z8K3QFVNZz2j5y/UV3rq6J1/9eqMoquqpy3+E4FGwUbNYSLx7JIvIa
25oENF7vucHRp1levinuDs+JlKNZ9PCEofIPIuBgeHkOPQg9U9+R/JKsTKyoKlRhEo2edsRMuLnn
cR3/wPdkFnFNl8iX10S4vpuGkKW2RHrjwPoqlmreKZX73MlZhLum8/Y+kVjxtPB29yCN0lmd/hYC
29rU+W2y90eorl9L/y97VWd7mKUevwFyQ/0kugR4eanM/MTQnPOU79TDv/J6lZbaY6rHk1XKZgNl
1KJZytKtqMcmH3dVD5CkOIGWHHQC7Ktqy5jE+lnqXAdlpLNBtlf3hGbLtX6n9pZAZzykPU24V3Th
0Ynuy20fIV7wfG1al6eZXdAgs2thiawzpAB4BHXZBlVydmiB35XNJ6GAJGYCkZC1XdCXscjslp9U
JAnfUdfl16WgfWPh+E0aBS4Kc4tmsJhIhB//MgKtiEn1yX1UwNAwsiU7E8HfnAmhclFcFbpWx/vg
A5p9psBZsrky5FpI6YE4fS3eOjqaM7V1IT9Gxt+iK6aprDEsDdfl7ZqfDTPeU2bvcqUmKnvSw4hH
FQtjJWCrJDcEsVxgzST3rp2FP2BPCraWoI9ycF9e4QanhjHUmsf/YTl4rRnq42xJixEOWXpbTuvj
ON2ihjbPCL9LV0nZaJnjQddUKUEwhVpByb0AP37FpbeN//J4AGB+9zT7yE7wiiDuM+TnTYqruZun
gn2OfILI/9s7EptezSpWrYOM+aOdpuAgwCnIdGcQ2PbfpOrF/D0jxmbh43LC+QGRNr/3OV+qmppr
pb8yZKcrq5NuoQwf4J44+FSloXF2wv7lUBivWja6hD4qeT4eAsilNxdUCin3/IXc5fBjG41jXSh2
uEKnqdHEdeRdp/9Uhz+x7vvLdHyNhY2/GXi/4996sh6orm8oKMNoFXZMPFq78vvbAboxgsh6OtVj
uxuIXhDWXWcbkMmDyebAJP1UFj3RnG2Og7sU8EcQLel4G8qpS1XtCH9AznzdzGAN5LqdRrhBN+iW
5jE2Vf9WoQN9pQRls4CHQzroHwRjK56vHHhRHyUGfZt+7EonmZACeUQvD3mqUbKDvw0WZEGpUlpd
yHu3XKr1VhxppSsfXTo81TYFajIcBFI9n9UNQqOLogpXsOolWWd2Qf1fKx17ItUQ4wOoWkcq879A
wNWLvmmsTnl2N3Ct+AGe1Y97S8XVFbmkNKcm/JmnJ/QXUzCz0VZwcEmUfJtYPNAQ5XHBK9UluMz/
Gfbq+raA3YGgciodb8874WzjbZTftfidNpDH8JRE4dqrp9z5KpIBnTiXH3429lM3cVdCmRsefSK6
ZNx1Bqzlyh+A8zriHa++khK0Q/j0ZXg88v2ItbLE04zvbCh4XjhvLTmXUs0FNZJdPSs0CpS6O/Lp
oPFxTrNw+zxIy5eojJOgtl/Kb8m9dh6dc6+aPDponrV2pGR8S2iwiYCzUp8OXK8dAZSZhqaA2+UY
Mun2gLp6zxmVaN43NBbRJXM2qxEEzAVUI8NYL0PVg+sXSLxTJUIT3jEda9Yls7PMYaRyZK2Gmmjq
e2poThVWhBoEGw+/67/dAoogyKIZQg37LwP5i0jvA/Yo0CRdQ9u2Qk+DRiqM10B01sF2id3u98Fp
QMdua2VOssK4xnBKyoU6yEUNIGdP7I5SBSn2Gp1q/+fOiQIiVsyKZEJ/Vq5/l2UJG0bZNPcrx6QO
ZyLROVnZQ8JLgHxZAbPgTu8T+dsbYlgMWcOGwlzhi0CHW0uBjGw2DwgMMSvCNpMLCw9SOZvOfBCa
lJnmGJ22SVRI/jS8+fAqkEg8fnIvWlXCnmjzFrXhYQ+4r7BqXhNE3L2AHxKFy7uJBaQGkPZnqyik
SPOwpEESIgKEpjVD2ql+KTrirjWMUO00gpJz4Y9vSKBuo+3w0iWWsoktTLh7nn6s0eeZLKPm3Pgy
6MTrWSr3ztxwSPDPnsibAwZpR9w94n43SMKSnCLwQns53qdedGeyGR6OrtXhL9Lp3XXtALiMa6gw
RWKpE0MwepzX3OeIf1jtXMYDocui4eZ4ez6Fl9hilnlHXCbWRxFeVSOARIdF6AT2xModVVHjhT5P
50bv6RBQFycGabQlY2PVD8oZDFzlxoSM7YqeSGFUB7ZrRl9/Stto49XuA6YTsblCZrSD6aG49ndJ
5vyL0C7szp00xj4OnU2+3tJrIFos65BsZJIoSIgTdHRhPUd3DZcLYxa8c3sK6IytXdow6JmsbiyF
9pgmUIVnJs7ZHChc3DjgjiwFbQjPoRaaFURti75Xqatdgy3goXVNJX/v5EZoELXqRHHnUN0VIzQe
j5MGMvVLcAmOXIIERYybjHTGt7fYq9Jnkok04c6YeoIRgR9HOlW1gNXd+GUjZoSFcm2mynclV5Oj
CcmNJevsBvkya+kxRJ6r2fOTA482o2KI8QL9ao5w6ydcJ3zDwknIB0MKcvqupKRTUOGLt4+fK3//
yzs5ig6kp+XSUe9Gb0+vv0rnZQe85/AFKJPSaEsvbpiRb5Lsw9Djct6BV2MxiYO8C4N6cbWMPV6O
0zSvjfe+c5tOcV8r72oFCwAxQPo2/U2tNhN1ZtYFVbGWA5nY46HFaeYosYBYcDVXOcXU6ydFculv
vqylYlRoleRqHchsLYBCZyriYmqyTeP6kjuYB6Naka8SpbthpHe0qntmkMOC45yBO3JIGKYNcu6z
v8o8V07L3gl1oY7iJ7gL1y3zg3109rJWijFsHykFRcASWg26kxnmY6mKqTsuYHRXwE2VBKeW32wd
4kxlKtIXp7Uc1mnTwaq5pxZHY5Bml9g54UHiFqlyDH0Mn90L1PDEGuFiG0bWGpx+fOOKZhahJ8wE
j9F9T4DdHgWsuY4xfneFx7/6ZlItTX2f36zOfwv4zefVwbnz0EzZcQrbz2BVtpngoIncVSQ3fVlH
g5iEqRlCzOIY/rkOyMvh7V8EHVx7LVF3CJgaJcI6FnL+AdlJXUGMH1VSms7oDONMgW4M1Fw9N0hQ
s/CcWyl+jS2f7tUzijxeded9xDJDoXM4nZ9sYJpoa45WOFuEEAhe0Lf6zXS5+3/26fNLWSrep3xp
Oaleep+jDo8X3w8ikq7Mw8bdxq/A4FvYKIAmVcT0VUkz1J9FcY/7/gqTaLYSHFef70pcVj3Wa8d5
FNlB6uJL3ATts2Kc6DdiMbDSR6XTIZXLa88JKg4FpVSn6s7HDbsG6u4rzdR3LkFfvM4462K7eZqS
UKKlJqr48zpcoBbtggTTEUWkwkEPEZYebYjxVyDDyGl5XtT6r3ou9Un/+x6n4dF4cEZN06MKHEnN
Ta1tNHac0BtGRvrZMlve44A8DgRmPl1TKwTlamz0wWgQ1bgvGMOLPV5181uyAh9R9wpeq/gcIe/F
ijC2+kBdOXNO+ljj2Kdhga7ki4Hepxh2JGAv7oiZYK66yG5aOI9CvIzB2Ztp1Ss/CcBI1gl2EvgS
xiFtNmD3+KrIRh53OXj2TjwNQc6s3HQuqCdBXxU+MJ6D8dbcqOVxVc8gj5qGdecJPMR8E6HP7AJX
Clv1d+DiTJpqgEcNVnoNk0jMDG6FQLmqBgUuSsoPEFiClSVpzAQRNL13cNcNcJMTq3yjRKdvyvjr
e7oRgEiPFCe4UrcB6lO/qIxZpNfPW1RWSEei93al7146R//dfy3dcDgmtknqn0zC8yk3Z7T/w5Eg
zvrjLp/s33Cpug3kD/NssfXo1870i+eKrSjYlKhi8/P7SJd6MEszFD8oiM9jFU8nmu8gKRSot0E6
vRkMV/gtnG5kgForJtSzag7TLq3jz2zYxZ2sEQI0sYq/133Buwm4jOoECsnQCIkBC4V0G6re4A5A
AyAD8DW5c9Y2v/2k9gJB/gKa/bxKTkZW6AZsF6A8+Ov/5yWXUmEz0OL/8j6U0K5LLMClGQt/937G
yD7NXYd6dHJs/Fb+Ng0rPNLIAyejbHvvHsfKcVCXEcxf7k31uGDNQlal79IGYLS8VJCDfk48KBM6
j1RA069gbVBSMp7mOUVOv1Dt/srNxauAL4KbFzpD4v48vItQ9jg5dO0UmC8E4wOMEna5XPBDucgX
zuA9HdoKXAcLVn8mWf7bz9CG5F57TmsqFRtzuA0tRzaIs1+8BbsFWYJxz2DIqIZzH27V4sH17wxG
417y8OdfMAbfb4epxJsZi7V9XY2hAygNN1/Nx0Cghd9GUB7X7ZyMBJ8XQN0tRFH7GvcZMkI1wZEV
q5TkbQA+h9FA9EkraaTQna3s+wMGjuNNR14+vecVbU0alZZIB+yYxCkUqvSya1eyPCRxYeOFpZwX
+8/83sqWIObnPN07iVn2hNLzvxX4yZ+Kg6MBg64RTzEsP5Rxcp3dvwHAS7D8K2mn+PHAYK1NHKea
gzA0AwK5029zX7jD59gxnD45VlhgITbMESc2UUknJOnSU0Lj6a+j1uaWcZzAIn9wjfzgCJUwIkYI
ISz35P/AwHx2hESvuksNNCLf/H9UApFYGHomSe2JygQFXmnQaFXsedQegfGafCWepP7HOGNf09cN
0MapinOKsa0fGfot+jc5XM7t1waqrnQExki7n3CwOPcCYMybiQqKsnjI5s49POj9L2cjle8QwGDg
86N/H6NKrLw2lFCDn/QN95R1ErFgybaK0BvgzmWASNnitozOw1Jf5m+oMuwB4TXGIGGGI6I1A/51
LFj9MLKHSjqdqlpCcxur0fvfBkVmnqhlRqSe3QKeRI9FSyQtQiZhl+l5iDz7eCZS10qsdQ6O7usl
+hc3CvlM1FvCZ3m6U8kNR1ohQZrLQ9RaJzrViWGMVUD+mA/mJpacO/dApp+xERojTuNgkUTrrGBP
hlNYGEK3+9G2n6yOQNsHhNy1zvkEf5JcF3lJIMkZHSlvBT/C6z7pZ3Qi6LWdk1DDzL7/LiLUVgWL
be2j9n5E7p4D98QzPomxazjjpGRZ1q8yslp/6mdo3ldk9K54yvnFSZb8RMRA6OX46pzU1LzRqRdk
atCOlDoKFHv7RCwNGvv7QXHFfFyVNoG/+mSshrH5sBs+pDrhZondt7cjTfPHfzGiarbobAVLtAcj
al2ysxTfyVgo7WyRvwAN0NOB64uwaqGUZpdVHLocUeQTxD4UJZZ1AGeInupg4InBbXcAuFrwY9y+
OXHt7RacX1aPldQGtPicDa2ePHexGiicuuHA8iwNqrNQonKpSnclSavUdXeGasNPjvZK+a5vHSOo
oIIRb8xwfLLhoaGn05gJBzB5yokgJ10cl8zzOKPWs7NSt3o/sN1ytAqKqV2vBhR/l1WImb4jQuj7
lKI1x2FI/zQVjSi5CDHxrahkuNTzIMepo+hB/lJQf8d8KlVlYMO7Aq7FzwzHSghe8YUguuQliitx
fuKynrqpPHQmUK8Tfh09qI8bBQHAtBY9occivaT2THuOiBTkpMRjOsGgXx/4m1klawRxUbeAMOXp
IqhMyFPIV21VbO7JIhVgq7uabQ4JbzwkPnIyrmsoeCqrDe8P8B5NZCdLlSuyUmXUc20LhsbV4OIF
XiWrAIfHaEHWJi5C1xaTDzXBEdIpBbTC3F9NomJA3B7cw2QUpGYFhNlaez6xPwV2zKI0+/Cxa1rU
Xl5IW9NqrMoNPJT1oF34XtR4jtroG9cbbiMPSztAdeIBhdfhSu4wginKcFkkmTKRAJ4ZF2Sawgv+
DTu5owzRAd7/Me+QruBu87Wd64uQAaCNc9WCHYfwp7QPBMCiEBB2S6CIBBhZijJN9g+09pL1uWAa
RrWsnUfEssLbIhcSfYaxhSY4PACCkIXTC6dsKUy4LE+uU3tiCuy+qqy5uUZ2VPVSu0X489uqQYLD
HbGyzr41E9CXDx1AN4Gp059txaNk0zS6haJeaKOdU4KOWPQCa5kPStWJB/5LbcGCgm/meVXq5cOi
OlPJuKrfZpYnjMl8Ks1DsqTnckAycBAVMkzrNE8pvIQhv7RIf54cFZzgjQv7qEs89ghGZwrbiJAI
w8jyKehKOx4doLurbfZZnFQe5Rsf48+fG9RpktuRR9/1yvqrOMU/t6BJZBK5OP9zN2fksxHve7VH
3YncUAmk0RwKGqASX+uIq6vtRdu1gmwwQTDHFIrN4IKrqoGM1juyQ2+I3IeOjPzryjRojeVsk1Pl
1dkYQu8dyI4JMPV7Jm8mSOMCCV6IHb70A6fKtNNTsMFgjoIE3CG776MfsUUdcsxKpucmZGhaqG3R
3o8BmuuKkShfW90THsfEl3YpUHOemz5CRgnithfyOaGFTddrO1nJS6tDN0tVUpCmIVARurzAbLR3
qx/vEu78IWk2lM1D1VKX2cu5XkgjG3AD1z3r0uXqQRNFO7mW9YYXmFnpI2X5ZXRkwPbcIhFLoG3m
2WMfgThPmdtcsbrKnsYflNMpRvVcrJ/h2VtDezd9lQjkne+maVrG+OYM/giEmADRwwlgGJfE3q/M
GQOtFJJSZNZRA8Y96bNIdIWr+JPm6O4dWZ+SmMiqytTKs9iFBFgkOuI6JHWojsfFcqNrOjTPzPam
iqKL+GHNvrClEndaNTI4agiJlJeWydyJkjgirooFAc/z0jh8+wACMGhRV9kM9mYRHivbQhUnP4jV
VTsRdrMuYXeyoy8CAClM/zLbQlDk/nzYQx75qQCplia3HgZNWnoGKTBFpcqYdGnGsi2ZTljb2/go
Sef00D2yDWgbXlaebknEIGZp6chnSL6+pGli+/iDboJro9zgfMEV8pf5WINjT4Z/21/dAFO3Iwu1
d7AGcVw5eIddPTTXe7cCZqcH/3a0XUZsgO8NbAPvZT4nTzSLzedWN3FyhOhJdotB8oGrVJHaeD7C
pHaRY1uYUkvqLJya9aW+XAc8odN/O9vl6fYKJqwVgLFUqMJlFZouBCnwqbh33yh5/nCKJ30ZKIfo
rPZij6e95aZsM0YKL2eEMDn4+j6b+ejibWBmyheTWTIz3twNJ+rOzO2M/sKoc9kGIQ2Cru3+FI6+
j0ThT2nSEqONJlp8IcMyYckpgciAYtrz80DQebgtjnTJi4+paJB+/kZQ4Vt2oD0/s4DVRAFULZiL
qdCqnigdI/Oey0RuEXjfX9v5QFWK6w2fFCLo9zVnEMDrbfkfgFuPtOo4H/evahVEpL+D1Mwr4cX/
koZ1u9folFtjF5KyJMvitpG5SkeQxQ2lbcQzKu2L1j0pw2Kp+acPIblx+Xwz2r7hco1LXSVd18j2
H2TDXKbhoT9WJ+QY4ie1Olcwneit2SfJPFrdOZ4H4PLMbFU1p3IfiTE11Dg84QsxXeLNrH8a0JOB
6bh2a22vrJUgYuzjRpqpeINWDWOo5hfERZIsLEZlqvqDu0xIsv+Fv19i3fHjgiMUqX9tuE8zVbLH
k3z7BLATGuiwr71y4emTfLMbxZADpNyfY/FsO/Nlb2EsGYzXVTp6yT4Us3JQw0paPtIswCS96mq4
/nZPiTcseU/dQc6bKVtlEpAQoCjFU41Gye4GkfATJ3e57X6WvxUDEcoeKCFiA35UVyAK3MFBe+Zj
tHMBeqofplpbuNS+7vrFqHo+X+bHmCxRWjTnMz763PU+NjbkfrgjVlInDMK8hETLza53nJTqZySg
A288WW1I2VVwYkZQGT43Du7Nxz0EJ5i/rFjT3Ewf1NVBaGoxr8voyAqpcTc0YM+uUcrVq50gkIXY
x1b+H3+4ZNw3AzmL+pHdwzdx9FFPQCAS9gmcPCoj2FMHoaUw8TaZoMtJHgsBVs9B4U6na/mTv9Hk
8vxsIvG1v+mSVJh+8qF5fDCSaJbstvvNLds20TsW0RmbOKDkVwgnDvzZ+XhXpb7A0py71d4VTBw0
IybpGJPLB78JgFMNHistGkanPwCSY7JQGWVXuFICDl+FCK3nDX9GbQwXgHl7C7/UEhZG7qiAWzWz
4SzqOTaeANtzF2u5xBKbpIEqSaV7chlO539MLHVusLbM5gvYL2vZ8nhIUNYMsSR0vYgEKTr3KDPy
SNONjiA6gGq5m6CLThRHhut6cdjxf8CIweJYiofgPP0VYx29PmXabJa3Sg0xaHxw7yqIlTyVNa/5
tWyVTD4SjBMzT0PgxuCKTJkGv9Lhiq5xwJ5SB5rBD8kt1NHWBPaMSfqK1wenzLOVXRlJVtU/8otW
9664d9SflhS6fJa4CoIlt4CEpqKbIjWuJquRnyc+6T8GXMHSqfdDNfShc+pB0UG3zEd0GmtRy8qr
+Z08G2Ke2ZTex+GjfYtqzulsR0Vj3Km3uTCOfyg+ChuBJC8mU6yMdA7ts6lkfzkPOhU2hMxyeKgV
DP0CiYHRynuxgh3uuIGwXO+tl2Pva+6PmR4YuEfolxu3j3yybDA/JQMKqhn4fmTY5RVEPx4X7fL4
7lwktE3eQ0g3VlHMZiQxF46A2vMdABVbupz1+adlEV/lwbqgnV2UriAixK+v68Fw1A1Slf9XbXnS
oEYPbUA5ERQb8M2fCtAPLlGrbaW0t6dKP5/bkh26XDQoEb2ulOZGN9V/BsgWUmZZ3VsbA1rllTSL
F8jPJO50P9PlQfB+ZQymbE27NFPNE/ZhcyM4tvBx5uUkn+wLacEhOXhLA1Xupi5HAzErRyLnIdT4
XhIiZHCr/ShyJxQDTsGKYj779ggcnnlAeLLvnIHRgr1r7t17tVTeXRnJr0oU2mQ5dgxrOFDxdt4m
WAonh7YaRBxGwbSILF8fN3DIHegNOaIFhItCOQ9Yxd310D86TDoyWEsRSflt1Q2j1lUmajrBF4Ho
zP9f0aVfOlW1sy6WTKNhXPjrpOEf4NN7ZGc/yJXPLqMMhSyXL0R/rcEuWUJ7y3xnM/2r0ZcHapwY
GxuJo9/Lge7vJWHqNXT47fZn8Vzjg+oOzLVdulvvHi+ixLPAvL7OcAmTqgu8pQOaEcySoNdBZkvv
mq5M7a1nqhLq/7bTJWEsy5qhhZUHD8GZKL/2rUY/8EQjrxsrq2rza/PlTEbnGkk67smTd58weF09
ItNszMPc6CgPfGCTj3GBvAnKiIpDAV+1IUjg5y7JuoGGA6kC1GmORVTavFUXUiC3Uo0/6z+CqRD5
d6G/cGgsJ2kWtJUKKCw/rvJKzALAe4CMHlnS3AVW6bmDGFir7h/OJCh54w4Vl6BFZiZzmTeOK2YW
FJk4tcFnZOEEi6L0FN2TUY1FMGvs9En9w/faRtPpepQWG+T/vWPmRQMdPnjCQBAoZJ5/lgnLk0BM
KIsxnkcyGSJBFECLrl2hAO4sC9YbWS7H8nl36awbrMTzLRk7kDacqfAJhE4vbhdoEIOpwNIMrFU8
xyjHBfIX05litDMDk/5Fi+3oVWbYjmhdB6a6y5NlgxIMOPGFFUsf6f24QTBucrw6bDsjoCrqhSrE
zScb9nPohzALTvVMVcwvkNIWwi0qxkX6yUCdyJVwcHy6o4ZcIa9v7weOv/VfdZrSQzWPpjzuHhRR
/YVtQqA2qoLPi9wrVRy7rw2OfDhGhHFkLd+zAmGW7o/3DaiiiKItcfoOb1N8rIf6VLmMgn2ZD1pW
KWoEVGaNFCYz6l0DyIHR1aynIHPdzMIqT6GsdMAkLC4MWsLaOHhxaWPO4rWQPW3s3Ytm2Nbg3HUF
gMj0vhdXkm2YKzqUoTDshGbs2JyPX6Ce8/RCJWZC3ZVpm6ZGJJsQ7YzMbgEldieQ7uzrz2x+YZTP
XR+ROz/Cshqvby+eG4mixwQ0FliHrMLwidzNtW1IXbqi5IN4xuQF3ihvfGGudMu2fVAhcq3iHmDe
rXIDmAbUeE7RfS3UMWodYAuvJhwFGnL/u+9MHf58vw++JID8NkuvP01Ufqr5rHEXBT4X4jlyV6rS
LGuSLpWBOIt6o8fwyjosgBq3s6Q1/WK6krGgibfKjdlpBwHsfVDGGqiM1vWyWXNb7587ueDSExhg
c8wYRSEPXo3FduO5I+vsSwKGSEL7CLdT0Z6o6FJ3JYbkv4ScznTrMxl9BgvzB82eqy1f7hVJJ8vM
mZ6H2KwkWFU8jbxMo3kQMaDsYo2NajPOTahKERIPDJgrO2mQIaW9LbzSPosfkqi0dVYJ0CLvi0Ut
aov8yv3dpzmz9ZJS3HIFOk6xAF5FRL8JiI6dtdWLWN8BY0cfkKZh2Brh63vG2YOxhIM3tQpqQ6yj
VSddmPrFTI0t+nalc3pKWX5ljY3oVxdH9kNPgQPE0k7f9bqMhJ/vZviyOF18QgbLTsmR6MrSomDl
THC2AIjkrsSKknlevsw495U6CLUPXFhVFXbXTz/QZFhli3/yKRQHmnr0hj8OReOM0kWk09lrfs77
k/b2aCAZjEulhE/wLTm55YO3dd5AfkM54biaU8ubem0dg0Q9R3XOzQ+x61meO46bb8cjJvtGNhc6
mgyHTtfITuQ/l/bZ6w4N+CRvDknvgkaR7iEmeLLJvd+Ehs+J7+XcNMm4SoP8p2mJI6f7rBjhQTjK
n359f9dInfWisWUX5GpXlsGfccaKdlLVNQeuO9VedFTGZ9zowmKnanVXUvvmvEZSQMYkd74lrVVR
0DedWkLRByesVPJyD/gJFxSF8sXx1MjERk1pMOpSdkj88g809jukkDvzEF9rpH+hz7kSPeNy/INz
U/7jCdfCE7tYVVYvqEAWWsyVnZ/qgGrrf4AY3zKYX1ivlJkN1QUfnPrfjLJwIQ/nO5wsIQ1s5/K0
yKQhyzsCy5WhEDBorIKwfJTTj/9S/MIJMuPfRTw3uhUz9RpWsE5cZ/8wFwscs1D2/BURRGA2r27H
lo5JzmF0/dPlFxHRWAsAjmHo/YPIp2Wu9nGrH5b1GgM/xLtCNq/tuzw2xIjhbbjdUvoDWRzFFCJ2
Ue6oewGSkc30RTQSaxeXqdpbqrN1UUzxkaEkRvdss4zC0V8NydhTyN8XosdZEsgrVRGLvfWScJVa
PYzPpu+crKrmU8P9Kyb1aqCNY8iBvbsTZiqn+NWdIYkpu7VcleNrWt7Jzvc7H+aI21Mqa9I4AwDX
zdZscWkjGzNHCi9vFYtO9moLqy1w3G//oKbke49DWHrmELzUEj5QgBEtirTThXCRULPOUVWUPKLD
nnyGO5BQ8M2LPIhnKGEJEf+p+rKJjOmFbWp8BzA1O1Sohn0DYYSiXKi/CYyJ8O9K7hK8gXU+Y5Rb
Uay/RsaDFnep5p4p/YXqqB8x0Q8T9qSChBMuwKSYpvLX8pA6VEtAjERhACQm8mGdds7fq8ZownFm
JDISvW6Hif8eZYRObYugOdp8HxekJMjQ+lLqgHbOuoI5u6s9XjpCrNO8460dtaBLYRSVWhimnU+O
1QO5rpKqoyMn9qk4Vd1ciNZhTwyyq+wekyUDlFpnO25j2nlnhx6JRdvxcg9cqErsGX9EjbPX12AH
TSeet/sQX4ebi40cIJymRfn7TkFMEnVurG9uZj7dmRM1vm0tQ6cYyTEltuSYHkDmAI2ejhK8K9Ap
2tC9YLKWrPUJlivZmTiBQs0ziELfN8W+pDLp28sgHj8Maa5f4mDTMSK1hEgb0blpiOKpGjXPXmJM
JjbkqG22mCcyQPd4V68G9W+n/WXvrYcceOUSAYZFqX/YyYvIUOxLY9WEynA8m71+Hbv8oFCUK4E8
HsokeSrYcef9C9hdpTiW7VXDnkC8MzNaVwYw/b77U2aICrkxjfEDuYR6ZlpRKxN03t9HqMbaVdTI
fkptjl3Bp9mP5ES6F4wpFPhASCHECh8DOMJBGRYT+oraCEbgEeF8RK0LRwdCTQa/2n2q5irRxJcx
esqzlFkHtADSRiN62BgvS2a8WvQAxoP+GqywEo+cNBgwEvr0gEwyu0NTFHx4ZNO8KoXsSNlC/NU8
ua1bXpGh7oJf88ALXdVTeJekmpzhBna7gnsHL8CW+LrU5Sl1oymu8uawWaeyvC0SrhQ7UKvM0qng
l2ibE+7BO1oCoWB2pC/EFru7h4IFc+daLfFNKuaLc9FRSNI20t7yMtRh4c/n88uC+xIpXXbL3ZWF
JliKyypXoWapIJd+lO0UvoGPSfeEG4l8qhQevp1fz3Ot1Tq0ri2z4mFdsKfNPtdrJpEn+X42HZF5
eti44+P4Q9fklHI8v1bz9A3q5KS6TLq7+XU8pLQP/myWSAvoawMoXM8gxpnVkAwE4eT96jA8KLw2
jDcLm1QB3Zt6lQsPSh1nkqsSoUYGdvIPh748+eghx7eOgyYOLRact0MVYFT5LfuHAcJdRLEtvv9y
DqSFY4rezhFBwdM5KQi5sF/mAx/mE/8PSAtmJe5/EqHYF7MrH13uEQqrq44fhMiQdd5Tij/T/uVZ
o5UdmW8tPmV/mLLhnz4mfl2uYf+fFltvcDKWiHOf+97j3+8FthqQu6KmWra6ZzRI36GiKOscBO3A
t38nsveOCSM6n3VKxFtlpZWWzWMy1J0tRIbe0eALzhUpaDmFoXAdVD9UL/QJRfdKJz2Q84q2hGlh
ohfkWhZvJEpvudHSvjCC2ZOV2l1SFJUv/F9KtcvzqHdzRTzHEECU2NaaoyCcRsiFGUrqunmom27w
WCWzkwDybDMdqgTPc5O21NCFQcZBMGiifZGjFq2fAb28ivOZA8u2KTsNoiQikMMClsFbloDG+lY5
o7NNdVFGe8FUk8klXdjg89XSUxh+NoqXAE78TcUom7BYciBmgZEZFPYjDkEnNUxd7anBOhr2ei+m
FuW3UasQSEPUMSow4MojP3/3T6GFfsgWeG65kITr6lJcF181upr2CHc2b3aCaCqOgnFbF44R9y0v
Crr/ZipFL2jUh39lo6wRd3GRTdVdb5OHwT5sryJq7d9V4N0ndQ1YvfIqJQzY7aFKjP9lDWkkJakP
Cev5coNbIiCd7mhHn1u3E/2nnVdBBCIvPusWdaJxjyn5E5HtuOirWudRJ4yGWRi6Dl2y2dS9Tj+y
Nou7f6IsO+gKiIH9akN0RRYZeu16VMZ1MQza+WpFSxC4ZOFkhu+ZQtGKV7HN/QzoesIsyOfaAySH
ca/Zwax4/H/R1a7OHwqdQTmLCkuBGsv0mVX4Y2YYilm+G3Y/MrnGCyML0XWKH6hIm0uiZr9uBcxR
NDWRid2FeBid8fgLLNOUWFSEQF/vPA7MdBUm6FmdmibT1mKW5a0LdwnnsJH/83rj8eR7N5rWtqp5
kyYc9zco7kMrx51cwKnc8+N1zGEp3BmNfc8qvjWeQ0KY6RvBsL2Vv409ews7VGt3E5KxDLgd1CI6
vRmLhZCkruruuRrwrhxCnMXqmobrepmNbJ/IcMgZ7P4l0VAxc0Wpg70ENmXaBf6XLI4ljHnwSuet
5XQJsGBrb6AeOrCKU8Ihl08p6HeGbOyKtTQrhHG06DKvCPDhqPLZqLvh8DvWdpdzTauY5NN53bT2
zTXxYmpV76exPbbDpGyA66aK5uwpmlsaHXqFE+q8kGiW+FxK5iaLtn4Eo+xT6/dotaFN2SM9XZLW
TDNLnbotbz1xIODyGJtxB2BPSPen3eYBcvRr0P3WKRAiENhurSC2SV4nhIQKZXCnsGLWOexVWCst
YNIM2lPApARor5l/a/MBxprG0Ww/iwkhgTX3GQtkj0vVPKpShQRTaFSJtzMWtMYCQ7hZ+rLz7TcL
PJkPPIgc6TBWzJaWJMXFs4qGNUgDDywXiNd0chRkvEk1eZrLLvDRqL+hk2wbGUEwtNKcH3xpTIKM
8t73DQo4TQMRRQfKWv3PbqqhPSIkrQeOwU2edA1NNS0n2CcPjb+J/J7UQw4Qiysf/cWEW2Ow4rNR
xiwV/rgGasdxiYcZ16J6grllNnv2zJYS55083WwnDl9Jq6YNQMI9RsbMz5hqKYYQZKlJx9LXMHWB
3jbtOYz1nHHDucykHHmVMoEnkjaNyqZkoIt3Gn8Ixu8a54gFaiIjfHx3uSAh6T+eaTfXh8+XJXPN
hubU/gZHuJ8PW0B5OdXqyfkMh28GwL4CdUZfyNTTyV8Av8VYUAmESFohoamVWP1lDI69f0fY8fZc
ARqRGiDpOEZeABfuJ2AGKcJxQ4kdcJeIKljJPnyuMwo8kGunII51zekwb/Kl5T27XdT+My+xQx4x
+JBVDJm/h3TsZsCeDF48rTdvCzPg95L8cnD+jR4vzvGz8YB+mVcQt0Orvxgm3q4X4KTKvJKluEGy
+L69DvNL2OkvFqtP3LgmNdajHV/laBf73JhZffRrJE8isg7eupc/aPJNzQvlrGeM5KI/f1BaRiRb
0NfQiA/uvPMzfFAcOzROLhLPvrP9GNypYNdeUHJAmtCLlpjQ0wLUe5zQTlQ12gPi39ernep/U4BL
D/HVpiy+7hrCBMiLKI8PgJdctBkwcBm/04+c6ICtx19B20Lf7CBzUAz9FtT60x0YAw2zI9c+Xloc
l15MJMMOHyB4JG30hrd9Y4JpoJdA3KhJJKfvgwGpdlt6YkXhWfY18ydyLhyN/OI7ayqdZ02k9Rs6
paHye2cgzywZnuXb1u1VDYaozl4N6mg2cEKuQQp9zLMqZ1+NIg+sx9gmra5fuuKsi5uOOmdglh0u
jxR33wBLHYWHMztxTbUTqp07/cOsWxs2J5oL1+QVq3MTdRX8xEp77ZQ4d0xuIwiMom9/thlCfYJV
oax0kypvplAURTqz1adsuIcMpQKT+xyauyB6heFkRbabG8lKe+mc3ab1EphCVn14gaORuf1EdpGa
p10urY7T4EAUgxvhLMoxxnsTdOz8pKqyVu/pe3ytdvfW471cAmCge3PdQivJgiyI8DdsViewntNk
ge/oDxv4I8se/qixHiFlZH+ot0KhObTRW+P7zUOWNTvF0m87fhUEP3aGwZkrbMr3eF61gBlC5+BM
FUsmWOG8cFZ7biLCKzEDA6ZaHEiWRq3Y5g6M5HvBhC1srmvfXLSIEJn3frXOEWz5EWuw6EjIbek0
ceJYigCBsNl5bDuCD5YfTcr9DEgPlqa1UKat8+/YKhxCkJzA+rizQiE3+V2s4EBl7eIRYlcb7g/w
eQODc7ntTVW4i1DzNdBOdK57V+qNk27Th2BncZZE+SuCMRzjdpqc97vP6o5zWSD3+kBgcCEkX0iw
0BkdRyuk9muc0jUtFmoe18YpFWprTbJ0A4ghZGVzVafcyrJaL4qYf31X3LiAfDfcLbcTVIuY5vMv
zvIe+uvVoSHdLL4S2FqYfNHfvhFaofKrBMwPu0G7F8Au9/w8HzXSpFs/X/6T4t15ovYGwLjWa1I8
6yP30MsbroAqlQH2sbRfSt4NImbmLK8L2FdYAX1KIZFVDX1l7iPvZOJY60TtWHUr3AAK26BNhoMR
jSohA8dpQHnwSY5VHk1mmqi4d7bL/FrA0AR9ZAT6d3YMr2TJ+CWij02/IwOMJELofbDxSpkQUHkf
oCyTXLSCoHL5iYhkHOh6bW/vKrZVttXrqfnzbUND66CTe4fhMMbAHNbJCBolUUFEZ2RjH0xLxLPl
iWhpcTzZwRMNE9k3cAZqDTrjnuLak53JifVJlGDK/nuQPVJGdFi4dwfB3ZhOEAFmzcM5ApeOo380
M3W1mSZx2BwjE7vNmG0RAN4Ku/JLTgVw6t/q88p/yZtsEHcQLQU1frMHU27tto1Z0oEaMMGwRzSj
XF9FRz6dj1gJQxgFyYaf/oDzMZBkla+Djq1TWh54KxsUsA+5a9yOKMhkGxjHa9YTl8rL7+CCQoHD
2JNKUwKp7cxkI2Weir0Hc49dNusT8o67o2ePa8lBpu6f4xn7j0IWXvUVGLKZriE6jcnjqJVUob/g
uij/3dzee3R6Nmj8Csz8V8NgvnGsf/4fY6Qf3/13XYKQ5zVfORa/3JflYxTtUvpXnMI04+LKym2z
i6GqfKXJKn6Oh0rcH+5BFx2uPMSrczogBCTfD4H6zs1HnFco2E40wvZlshh3ONMpIqQ+dSmm93Co
84MUZBTllxJBGyTAgzEe5/3nX2gOr2o0NumkYa/JOuRWKe6n9LReyjijQDJQtspe0gcfDrjGiPLR
SggOGJlSguyIh45pzZ661frCw/Uqh3bXzdgYExkpp+zN0XPAIHpu0YkxWCNX5VvoIAE8NejxfQkp
n5mb7ETkhvu2heUViqJyTtioe5YKcWRtqENub0SGM5anzG+s5UtNE/QzG2uIwMI5p+jlKR43IiQK
YsuNwJfiUQgmRn1oh7E0cBRuivY72kh8K9d+06/Fu/8cpz2fcsyfFEK+FKh05j4iJgleCWAc2lK2
iD/56rIsSUYPL0QZoTuNXdjhQIf+bqt2MwMIVI1WcLsa9P2DOOOdsx+uiYClu43TGBlioF1q5AJZ
SJkfpyPzKaH1+ifDtnYsBYyA4LXypa+LZ+F9nJ1PceOSnxByeQFhHTprRHsWWtfNXfQT1218pNTQ
qhxf02REaiTv4asXC0T+ODf5HS7HPwpg2ssslMhUok4YsbR9uFvB5z2jKePMXt8paw7Jv8BNx+/p
vQ0K+kSApBjHA4NNefwf3YlJ8sJ5ELbc96kt4ErnlIXY+pgXImYa7OL9b5mbprf4DKUxUI0dXGyi
U6l1COnjbCLLef+67bsaMMQOTBo5yMDi41iaAgx4faPHcNMkI46tLyHui8V3ntu2o57m5xbspN9+
OQFigOaSf5wx6UkU3bF2e4O86KmU7wT7PYTT4Lr1+OoDvWuaYZ3K7d2800gsUuR3jERyNziwlA4a
Bpqe4RWMifmh+EOFEHhv9+eCkPcxcYvxSk/rgT6j67k0YVDYiUKeciXPYOPNaORQq8eP4P3ueNBl
9HfKgDEsHFUvH5RYEBCUYhbQKkQUr45N2ybNQD0/wCwnWFQqR6XfPkvtg4b93Tjey7jtqzRVIEvh
ZlRj1doqPRfufcwQfv33nqZnfF/mXBvVRG3SK3wIJIKgxBqxG7YBz0ma7+4RCr1YvHiZwukPmS6H
QwyNH374dCjNJcOh90cyRDlNu8eqfVhFjQRLp4SgXjSaoHYY2b6Cf0eRNt2/OVByS8d4b/GcDVAM
fHFIyvx2P3t3geS/Z5fFAbiNIz92hvmI6L3IZQ/QbOxM18w7VWwMppsM3si9YNuMCXLhpwk82WjJ
G0pMpg6PBspEbL3JCU+I3UFqJs2PZSscXqZh4WzcBhscv/nWWMCIWsyJJWIGpgRmO2axSx1lzU2M
Or8BSO6i2I5n8zmRjrKGdak9Mp8ApJ+ij4GdXnHjiaBZUTNZR9c+uZGd8sV9OUkUM4mrZtQtfa0l
HWn/ZN3Geq0ZVjfjycc79NHo6cyHGsy6COWqWANrfmPU6SWdPplDJ0XhOUwIkqRncV/lJsQR4dDf
0M2Q5nB0IiqHYoO7IFqpKeUX+tZY1AhuwJTgpGmYrkP7AU2y5zrgvJXfld3OoVWy+9/ZAzni0vPy
GU1uXVH6fc2lFFhj+sdPzhP/E7O+3V8RGoHqfcNGD+x6IqjmA1E9Atquh/2Bvv/nbhkuQqrJuDfs
ImNwvITYYJWfeS6nsBdQxXTFIvaJ1dDESyLiy7j8lBKxO5SYtFN0DqpIP2ovCugbkXYYqmelcxuc
ReepOKNzJoBmnXTWwBAHNobaTgUpcug0KnAe6nJqXIdn9e/Cepzy/u4xgIvqApq3a/WguDnDaRH1
M/CYjXaOQUZOS5nJ732XXt6ouKCeeK6v2NdljQIbDcgEHeDa1KjgqK7AruQvFwsKcynYy8HATxDm
F8RTE8CjGK30vLfUFcGAWagecfKFrQcYfpslE1/hqZbamxx4K5e+tUFtk9qhiKjZVkllLda+2WiK
4uVmgturyxpUdzYxNP/Y4OPftjUn73SsRb3OBDIS/D6a8LV7WtbkLF53k7DV42QWdjJy3VlwK4/9
xxD78Mr5kqyRwl45bvY9P5gs2ZJ4ebtOg07B/LBphOeRuyBK1ZYnlArl3HUjPsHifaHCR7JIjGze
c3RYFWGfQnA2kae9h4FABsK8/w7t8jiyockeWWzkMg38Lw1DaW73ajTpJzWKwGKdUJ424Uss3fUW
b/mWOURcD7hOz8+pE0UJ/32+EXvXZLwJik6R6q8A8Lrchuaznlz5FE3Vadq9XRFlR43t1oxZZ6hd
VqBkCTtcxxj9DEQJm1vjB+G39poV2r4wkF4woyQlKfUWxjiaHIptXSGXyoDvnidqfDmOQDj6hmo8
pPL7kgVVaE7cXh++l1geF1mycrZ+vkqZ+cHnkZ9fhAJDh5M5feqFlJ7q+dHWrc61JrZM51ZVWlf8
gRaB8UHJAAe94TCjTtpN+0+NXHnhORGEYMpxylUjx5OnMWxb8PTmULftNA77lNdzq0Bndsz/BzXH
WQ5lj20xVjTY2x/xqAqegxHiDYXPNZFf+VjGRa8JYXWm20xWs65h5I3k70kn2EHfFmCvewKvkNg9
IhxVG4AY8d660MWBnFJ8DGzZ0fENrtsy2NmU+jQ+4GRMimIh9ObCYzjlOogTaal5DgE8rqtUN5/F
f9GEZFbArFuWJwcAhx6TrEDaUpBLmrWwbF/uEp8+b2EQ4zlX63lrgXRansn6V5IVUAQDoy6i2810
DkMJt1GcK3jVrma/fHwEnVCPuuGLNI/0OC4DbLqW/wP/aOZUTjS2ZxLx649+wCpUYxWSrc1MIENX
G6qkbpxOi6ygD92UyOXLVuUp55LgVR/JEEfNqh3iCOxe9IRlVQHXvpAOO8fmAvsOgMz5pZ3+DjjK
Xsd/zRZV92h4fEgAl+AejaDuAFO9mHmPhWiuBHS/y8Ax7LE17uChDNZk9154jqg1pA8dTz/o29Eb
ZLo/bDWxiMBDOIQgN7hQqiKVcsOT28C4LyZL+L60BY7qeqonrNPW/XyFMdF8QBCZtEbcIldJkMSe
AdTAJnuE3maC0VaPzLcRoX3z05VcbhOFT3iN/bqHpWwMxnrvFuniRYLjAstshcNgNBz+3GCvH7u/
4TPHnFac14/5bUtjbwp8YwbaetoZR7ICzTNaBixJXug08iPI6n4vykapyg3CYCD1AQM7mT4ZlBtV
b6g81wS065ty6MNuH7DoyWATdIlTo17yBk+dHPZW8PL6cQQSvrfh+AYvRy9qvqWrk5zQCN0ysQTn
mTqynW6HDaNb0tJiEc7NF2UEmoP7XrloT6Oou27iGEBZ2Bw6HTiGu/vAZ9my6ltfgz9VkzqHA+gM
4BJsrqNy4VDgjwjCVDXn8AfjLGshDO6tSYxPFpfDo+YD0n9Gwez6kH1s+hU3OxQlanyMz5zCBA6q
fKDqgFHh4iQA3NHRFngbGlp+r5W2EQm0QWVbU3wDtO7SmGRQWcE20ClgEhad65Cxcx9N+5JEm2VT
CNhZQ3IEaZ1VJTTr/dGGnsh1giRNwheYPcGGQlxojyGLTYg5rS4L4QuOk5HWzScf26P0n3cbfUGw
urcDkcq7JzYSRZaxkeq1KNrutvI3VfGaFmy1zMAd4PohT/zpedr848eY5d5UTJKl6W53GkM38x3U
pENuonXBf3KNiuNN4qE0JDztDouLPfgc3XCd5YwU5mBaqFexUXranM/SSauVBgqMIiTia1S3Vv2F
Dq+RMexoCsWrpERi73sLEnkbVKA3BY4RjgFyXsp7eUlW4OACOs24XqlQpFnPHRHH7aZ1T3Ld9JP3
ck2qUwyOs9773KrvDnbmArrLi4EhY/3KhkWf0s/RFPS7jFsnj3kJ0qJjRSvoudcb6XkgjyvwR2+i
prsMxnAl25BjTcKNs33KRwrGT6yZa4RymFqpL0t7EI1hBaFwNH/xwlp4GzQyKFp+o0g7AXZDX+2J
ftl1nR+/ArFGHajsPSi/sbDQi2BnyCw74+dXnSwwXr8yPAlF+w6izupSnTtTnspEZb/65XdnYneo
yKA3K5D+mb0U5ylKgvJlscX1kipv/jVZKLnuC/hsxBZhD8Pyen6/j4lzM5DbtEXzE2tpHQ6wNgIY
kFbrqvfsegp04D3unBvumTdxaL0mhVRhk7tQ9arfY6r6oah+IFmf7RKCXd5dX1M1LlLZ4T6Y33CL
Emhs0iRFWXVSgpxrWC9lb64kNhTzvIADJ7kE4/Hjr5Mk18cEkkwfQqNmK5he2hYC88mGTHvJFFER
ah54okVP4bqwlj5dyDfIGGJEmFvw5IFkt5a5UpsNuZItMxZ4o5nId/jNRbyKwhaRagCwYEwn9KNu
mZqKUb4LFCqj2Iillmqy5jXF+2CJCmfevrkj9z2uSECp8oNRafWwNnptUQyTLHWdv1cNuQoIiikw
R1L9KzXu86dYcSkhmkRxVTvPMGObg3djI4khkBA1P/ZWQ/PYbkh7/d036DjVY/SHcDoffX4f+O1D
MAdzsvfXUklJDkZLbjmg5W4tRMIOso/tGHbSSYBAVz7UeqX5uiXZk5SxBLDGGGkwubYIHwwgxGHY
MOPEHBQs4gUeo5HNFrhyhhNhtSXk2WxNymkZAEAq9OZFLYwqmvxZzPLQ3WfYFXEl+R0FgXmM3BnB
Gyd8bAdOYi4iq8ky1rvQlUjbvPj/8MwllJlw8rcTtSt0NJW+co/JCp/PCFQuJdIA6dZbdlSVZzZT
rcj02ZZqWchqQ5mzy5cVSy9APq6OJOvquRl9BWTa/uhOuS1lVSB+7i1N4cQKA+Vt8QH7hkDH/AE4
aWhRjI2Yku/DHn2mzHfpOa08wvJ1gaeczUUOstrjo6VjMVzwTYyrO9yPZ0KzE4IZNJ4kFzmYgnaH
1a7FVgCB7raURjYgRRhafXrmAXb5JVj5uPYRfMPlhbzWNCh0vS9R1PrC3jElW8kfwLi/rv5Cb+27
lz2ixkg9eXdVtu+gE8exvSf0x5Z7H+BFFJsmck3iTyhUvOMD7dnOLHMvwJwgpFp0llYTMF7HKh4G
d53aTV2OqJagXEV2I1oWtwbnPh3wAlzADbIgdHRB9phKOXVIoOACsfsaky2Pu9Eer5HPqc7GvXGY
EWCT7/UK/sTLACsJYaYfyQdCC+E7wJCRh1+mXbf2WIXnELdRmwtDhgVK4CvGPNzRHriFR9045M5f
y3HxyQJGQHEzWMIfsP9Y3FfDvdF69B/lHyZJ7LSIMa68Px5ow/1hYxOxmzzUDkzx3jx+D7zXnFaf
ArG1CKQJ77LBM7t89AYNJ/o3gkIqWx9G/dBv+aWJChRxb4buSTl81Di8TfEDy0NwfWcTquUf8oN2
oN3wWv0Sh4WvupNkDNeq6jO7nsDwW/jWd8JMm16L4jmoXeFsM0HDIZ9deeyUtp9eEabeAy0xBnPa
9VxVQIMA4YxVEzheg7UcnZD5YMeRP3j8Sej7OG19RENlcW5O7kJko18URNFR25T1jW7iGw/2U50d
OAJD3TtvQM5ahFtl9EiEmHrq81ZxqVVP9YHM+kKk7JKGAt8sxVM7UAygS1igt8YmKpi7DKeZ0qvG
Cq+J5WVHy8kUn9kvHMXnJJk6nvHuNYz9iIDU62oqm+fjgs07pmqo4qSGzlpKPUZeDQmn+63ItpjQ
JDJeZP7WstYSuwaDpWgEdVzZWAB3vpSMU5tRlnXA8SH73xJoOcxvGRfxfp4SordlPfUBPtgIv0Fm
8OzeCprXJrJaI8DPxObCu9umidizabWUs14SiQYGL7ENQJABGp16lEEuITdelZcvPHAKmAoxZdMT
mhm+HCs//2OmlyUBTPzSuIo/b5tXWkNjcR4zinRds1978a+TQQR1IhWCdhoD7sy/APcRUo3/Pp6v
q9Aoa8mQwEF2vFDjNnQ/r6+To4W7exI2zw0n/nnMt0ukuQ2tBbJRd1VTA7HrYcx7rYU6NBTFWyyd
nyDyR2SiQOp2Zu699CECk3d11QghOCQaSRa+7w5jTrs805laJEJ4IKhxc+DI0gHnQ9Ue3HaGebZH
Gaz1laxLSmhptV6F912G8na/NdcDspt35+v1qUmeOa55uVTxKtl6xUDKFrGig4d+UyTcL6HjUF4D
T7sO/5czC6h/GgbQyoC8M9ccKi1nwG0GhEvIhSCumfBQU5LLBxVhx8WC20BhoYOGSMFmzRKVEkZ9
c3ZEF4uLmQnkcS+doC7xHUX6gAVMSOaOw+xDEaBJSoZNmxkV419VYG8scZjxFmZtnz+x5iQvmOEY
U1ThBpcx2bVVCCpxYtAu7/ulDmiHGFw2vAkxV1swrTvXBq38B1NlpNgmWx5OPRi5nrQZosnoxsrK
K7KbpSB2eM6Gf8R1tmLdMBPFujjAHUFlGxYzhJqRazjlQ1wTlmYKTJhSVhew3WiNYRS0L95JAS6R
FKrygY/A2x/6z8tqx6B5ayn+T/r1oQedhmDycw32kT5uSd9m8w9Xnb68bffwVqIegiFJ4mTuSjST
CzWF3HlqRpJLMBn2Mk7igJcljtk1XjKq+TrG7kT6TYBt9chDepoiBVArv0tazQnSfmtlDVmbkrI/
VWmGyjzKrxN3lIZnBAjTG3qKz2lbFqW3pKMlJw1D312pGlNJyUgZIncINdXRplgieI9pl3KXTEnm
jVMNiwrPyL3sHimlGf+QyaxMaetvNeWhX6rWjC5Xz7fDRyvLxSDu3m4VEadvkZn+8sADPopU9Npk
QMmXlnpRujJvgnN93s5FfqjEGhUj+mpPUI3kOPpGiP89Msj4xvkdTsEmf2l2oWUBNFnnPv9s+9wO
nLNEbeDuX2YTux3Y4UyGFQAK0Toqhk4zwauRuC1WrJqaA+SfL0EJd6F0Iu1c2+7Ez49mbOT5iTjh
j1WpdYFdq3r/DEfn1O9n4I92TC52p6+yxMrNF7xS7n7EdM6MzFTVxbkyoaZv4FQZLfSnlPuq+lSh
lR40tlQhL4sbedXcwvH1UMDWJ0CH4TfPZGkqDdlLHXWl3kUTfqFqUPUpMWbMuRp75Exwe0Jz2H2m
Ti8cGyiEN9IFQc13nSX+toBZXPrNnIKRK1EUlhlcAk8W+IUQRX2tZJscEcoO4+i8OHD3KvxKsmH/
pH3BODdefy9GGD2p364bcVkfOrdq1Oq6Xs64PMHGutqQkUdzo1G0ZQNeXxp0CZV19sSm3njgR0ln
mf9ZDNzPnA0CpOXf06LBP2AXjmB3+v9/bEHft8mT6aWZdeercShANyq+TVnsR9vqGCycnlx+56rq
OD1zqrgUZjDAfSXONCEhOmP+TPQJ7xKEmjmrwQ3QWOHM378bN4U2OxYR2I1M0IeZYdk+zH61sR+5
yOxepR1JvujLwgiu29KTz+63rX49qeptEUxkexMYQeq+zXqdATUc/cFq2ptYjqDvK/liA2BnfDDc
snfewZZ0tdMpI/yzMwyxjOgg9Qpc1A7yDoXw70mCoKvcH3kGjbOSEUNXRSJbCnx08YPJi5dMeuru
btPDqwHor7Y3dt/stRo7TNr4S+SwiLDeS+4Z0UN3xbgkFBNkSCajgYPxKS069iEs9zx6fOliZY8s
xRZ0UktvqzrtgNff/fKjU3jxLyEP4de0donxwwNGuMGLq2wmn6EczdlPRuY7SNrA5xtmmcMBB7n/
zKbe45NADQ7Wr2h0SmfgcVmjfFVc2AjibhwtC0NEElQs45tcDpM8hf7Te9suD0P0oZ9nMGwYx8cJ
YwU4w/QPvQl7mLiixy4BRn0afLbHN3gDrdtcFN15MC7kMAeZ5orNq+0R+DGg1PEQVcc4P/JI/M/d
3HoF9lMGXiCmjfSZ1aC0+A99GbSuAZZRV9F/RxrIHA99LuIDCHFgMz/b6OviLBPu6/6LYvv+OKzB
qU2pxkLp087W/7vAislQzftbAC5Zo2ksK0YANXX6CQbULktIUqJQhKnIjndM9oMVZ2PtzRwkQGw/
Cne1YIVdX7cxGJPZadlCjF/ONsP/jqsCe+cdTGhaUIAgNftO89gcZMMyX86W4R3K4qZRjQ44Cs7W
DJzX1N6BcRJu4LZcYsaBf2JYriRBIQCNcz8sT/Mzf5Zf0uxNBePndOpCvG4DLFFVXmb44xOBikLs
HtELjcuRTPS0KuwfWyCOv0/ym4X8Lau/nGlJ93G6ClcnV60DrZzwzijUt62ty6OI0tUJYKPm+VOs
2iYtfmOd4wbQpjYq3PXiUGjxLtT88mXykKxtuq2DhIzJAqEVd8yri9UYRsm7zzsHFmGaut1d7AI0
eVRbloFOg2vblfxvALhmQDvomtyzXeprbimZASmAPxMXkxRQcDHgg8lvGnz4GadeN8gxhaa4zFR+
pM0633kOmiRx9wtnrZdVr89qE7nHU+v8zUaT6ZnCSFK/5Tw2Y5+42/C7uzhwJ0jfc+j6HYlnXhGr
b6SBHZEnswZ5B7rwlfCwZ43rheyDFOwiBF2ZYn7bxb83JZEbiXJhF1rmc7wAw3guarJ2KF0YjrXK
G5q8n/lSbZcQu4Rn8CAHdVkbz3AGLDL4qNya57A9A/6I72gU0aUGAqXlSMiXsVcBwStY6NzWz4JW
VauPvao3lExWWL3UjJzQnA/BH47JWtHDRUIoXsnzVOnjYXWzWlEbB/qOUPelmKCyuY9CMnKDGrJc
KVm+hJUEm9epq3ISQ1Goqo55I2+SHnN3too+Ydye3uhO5DrUEjVG2D7W+vbRyD/s61/QM6ixpFTr
XVMiXyhHq3dxdcCbWxeHd3I1LY8Gapw9jbqBn026C006qLsMxvml/NEdrHfWExy/7J6FmTlL3Qxz
wjkZ90NrmKZ0aQ9pB76JREHzVVOWw3bBY+tdOSP82jt6u3I3PEcq/abkaXqjNTKLkU1RQDZb/VFs
D1ddACN6AOLSx8oz/XHZqIYJQUixcRmd+rpy9UFswEg2C3Yr/CamWwLXiDXI3BbLSy3c84eBAw8/
h8kDy8EEnyFg1G2AjSW4NDh3cyH8Mc1ayRhyRmtzMR7VGu6J4Og0qRk2z0V37Qk0pd3wuClHhQnQ
vOV/RX/H65rTNLJP/QfjFh3Ys6hfYBbPZj8oXverjrfxzBp+S21B0N5g4CjM8aKUv3tfh7cTysXQ
n4gyo6CnlS546BGD3u+mktkoWy2Pb0cWwhCGh4VGjsdg0xyUJsQaBuILpUvOdxsZcWqT9rdvRyJl
OYQy0bqQ+ykT/KEux9IGD/GNPniuIxNmbnPUh4fKl9CCetqNV8arT8giqQLArnaVD1DA/qgtvIus
mijaEssedSfMXTF94FrT6ao2pHJmqtaoH8h8J7b0wD2SR4o9EfvV4i/bcwQm6I2Ihc14fi6VEkQz
/0T4YnDwPxYfwSjbUlt0zty0U+EyHPWgRp12f8p2uh29t6y0kZQNX7ApO3JlSFfs4zFD45sLk0u6
/U/Vu86WXbg64vaByIul5+QeoPL8paEovQy0QWgjGFgJZ2fwcn4cxN5I0lLHnBVI1XnJmM/v5bK7
BZJtalLN6/LhSfTvciBCXhDV5pui1f3uh1SJM7TLm8sjnQE8okkHqu21Xyr2ZGnhO32OZa4HVu5o
6s1vN7vzLwGPHhEMFDscsHF2LCeVYpDJiOKDt+Y0nhjnh0tjN9FVGguepF+biEigdTSVSoUhqMA3
Wojfnx27y9LEL8LPcSoD/ZLyGBoq7Zk/7tlKC2uO83skdb7L46uEp7jcBG5Jjxzh+JftAiTwbExD
cRueFkXbwZnWqp1dFF9wbdr93wdJrlZBBpXqaYbX5Fj8yIt+i6OfVZPpqxe7hbrZhAxbGXfOgEZ1
0tUIeoVNtJzFgAI41HRPNS+vxMuKgFPExy5dk9mEFeRU/LxikBjG1npPvkTbY2Yz2ZXJCNJOLy7q
ubtljwGVtZ7VcyvamgjCxdUiTCNrxAT6jpTevSMSZ/akU2z7H3vhE9lW6xj5tZQ03n1RfRXq67zk
cjosPWu9Ip06L4bpFsYx3ash3q8BxmdItosrWkaBctmTqe848QMD3MJE9MyrJUKuTV6Qn1x6rqbY
WVcYYYptHgfvHRG0s5VDW0mV/+NzwhWQhgUREeyIWMEqXnnXVzchcGK5i9PtzHTUiPjqpuITDKRY
0JDj/bskKu2hBowbY5eOWy7gryxAWZdEILAkfu8wLHz5XMFW7DKh9DKvW/lllYcznwuVoS4hWKfR
XNxW1rcysM8kbSECOqucBFvVANJgLps3KBX4EVohDr1esOszmVOnOYQq6uY5sixelsamZ2DMUhwz
Chpj5ngIIT+QlwD2isr0yF0iOOodWYbL1NAu5AvR7izbyODW2XLFBWrMBk4SZkiD4JPszQPfyHIw
WmI0Qq4dADlljfqEx0bYduYzS2wJYUFlbF8CH/cJJR4PF5JTr9Q+M5PwYfmsTiYUtxhtaWo5Ugij
DWrD258Qr9kEFS5HDr738Ecb6W9oJJfSkr70dpw0fkJuO4wv7sISWspQtKZCrx0BHl6xpXgN4GCB
cn3ylJ3pCAVpostc3l0YR9dDjGYHQpOtUYGgfs3xSrzN0pqpo9hYAHyEc2kU5R3sOhyeh95JCAq8
0V/pwHnrs4MzVC7GptHznH63gBc0n5wE9/Gi12Km1ZaojZilFmBF2+akpuH0KQiIIx7gsQu41JTf
5ZmZGOBHdMWF1MCdNnFRgNkMwQVziaL/u1py71cNzoeeBLPWE1iv5kijY96j3OfBvpgtW309IjCS
O49HdvPHMT+t4+4SUWxHHgZaO/DVDeLY3cssH4a7/9CNeatcqqNEfMcFf8QQdSl3+7DzYluFVOJA
fup+KCFDciW7lMBw7/G3GvtxlcGilAX62R8bK6D/3ZFpbYKl75Px4QycPfF2JMhMqPV8+98GNnrt
8Ovlb04PYdVvj5ZzOGInoIkMmQvWsJznO+uckk03KDKSurDziFOxlXHQt/UViq4OmIAhzpY5TCy4
/3SMWp0T3GIj+NPaXqy4jLBX7CKAG9UK3I9vKIyURzTC9AuQn0Tmkw9/FSnWSzZw/8AGFlBOfeVg
Czh1zva3qi+EGkFD9BKTp8Xvrmu/UIlbzaWmxZWEXB7Zj+kxWjbofeQJjACeuTznLP5sFcZbDYSO
BxGJXMD069TREeHb8hk1KkFAaa36YV3qTBztmLrfHDG3tdqhUow3Krvghb7JdQ6+6UrCTFXkaGO/
APflhXtdpniXy7UrAGH8cmOC2o7rYBP3L8xWxROIIYo1iZMLeaGkUE4A0oPMkwOTXiKcFXRejc2h
QK2qsLVIXVVemcW2eD/ygXICEQuULPptg7rPyybd92IYO7gqO+7pkcpJLEw+gQBFtHcnpe/JjHOD
ht94Db6f4cd52LrNqPY3Mr61hn3q2AMcu0tsH4kFKzB57Sso+ZrRS7gL1UMbmpgMG1eyETnjoFvU
lyDRLDj23EQxQg3Ug6HD7UjBLp+RW9G6WJRWQmfR7MvlemR4eGnPSqRzlS290PCXY4JBFkyFDvcv
HskL4jXe3k+QvhRUssGYJLmfjFDuXPswVDmGPXfB3ikIqw/C9c+Cr2QgH1Vo0Ca6KrI2DwdFV7U9
iYyRRCs7TwIL1N1QgVTGs6xYheGpiVm36MN76mlmrS0hV+EqkpHYV0uFBcfNZgKdV3HEv29Uk2hH
Y19qK7tiN3fddG7BlBTqhfXtg4eNOAkLfxEnSaHfMimF2cyRe6F7HRmjG1T0mAn4c5HgqkJLf7lJ
zO7C83ngE79ZSeY8IE4/3UG1Oyrn2gEvtMbe5ihdbA8HBZ/Ge2A5ooIrhatH4JznH1HjViTpcs2M
dhGGYcmzX4+7TEcXRw2YLUUO+0K733CGEj4c4EwAzECspE4wLGbdBI21p1iqRG6rPCpOPqtQZ0oi
WcaMsNsf2qhbB9gUP0mLI7CyjoL0RB9NgTZvrmfwJIkGRBZ6vO5tToEsSpNKBIgEBqTTMsaPr9nE
XS7In0vTeJgfEhxGddrqIW6AV/lqgyvCu604cbw93nwhyGju+EUdTbJW2pa4r64VeLBGPBuGv5VV
1FM67uUg1iL5K3FtWxFD6V8AcVJi+4Yu6hPtdFaabrDFQpAIbgpaEcamyu7LiKUUSITAc9hGX1cg
1GiRIWoCh2rFrxcAAXSaXplw4gRpZ25G8/L3xlVMRDD9XND3Dz/8MwSEBS9MRcTTMWxdNp1i10gD
IPDbw+Fbt3cE3LBKGRPXcyotXEfYJhQI4WpYhd7CmjxcG1qDjy43/8RSOPHOWpYYPKKktHQV/GvU
JrKXEICHPiMmxVwg8TPJP2C+Br0xO7C5i1kjedjVT01fX+sNL0sHtA+/5t6yi3yiguTX/SUNKTnP
sHzVeuJGt9HQScaAkUgybCS+0XgeAKrcedPcJzcGOFV8qJoMu7/Uj8ZrAEyDRWtX/4u/AZg/zwvJ
42R5hZ2EQCuwpx8M0SPQKl9QY/AN5GGH8hyF07zAkm5KGUMwbWvXqeDt4boffC+gHiFYw20qac+M
5i2LXUe797u2YDVx2QswsU9xJYaoah2NgByA/2d0K/Am8jKicZ6fMDF2J6+A/6j69TPiNk1dI/8Y
E31nsgrjmfbB0EXlFELTjwleAVjNqCjYqALHAbATmqNmqf1Mez5rAEnZdA2IUhZouuwCq9JwooJc
PliwmMLuq8SJ+bkXzWLkcaHtsN6scTnmMliTveEqF12oGnR/UzU5IQbSx+5B/hwmvAcVa8hCzqE6
IgJkOwNQLBSnbdovoONjNhQrI6p0icfrI462DuNaiv0oQ5lE+Y3Dwpo2iM8yyDhoQD4by2EOUu3J
95jrxL1Jk8es7YSb/nq0D2KVtRTjSAQ52ROsyH858R5jDL8hX3o8fyP+yNSncYRLJtOf2eBGVPUO
p0iqwoGImpdmhv0z4WeQUuWbfShdtUJWHlnZMmZcRPFO5cpMxNqDtrnfbY/Ozx91TqHMEHQM4LjD
oOYquk/qYpraLPocpLWuQYlL9baZ/rBS9N16yW+hs4WqRcdwX1gFKgaVb35oVXxRCGr++sCERnAy
mIgiZZ5pWZbpcon97RbvKI+gr4iG6CXFx6eFkY3dhOPJ+McaBL7JRLX8kEDgvl0tWYLpBtYP+AQj
ZYJoY4PMkNZD7EqNv5zqvh3PmYVrFqskTIIM2w0uKslwndRguQXXxtNWFWTxo/gYyS3kyHVcf4r9
NSVDkoOMLdjqxVy8jQelOnFxetDkaOqdQs5XEIqB0rIc2Pg06tyqwmDf+cHWtm6HYmBZJUrnx4nF
NB9LZjLtIZJ4ft2I2m2nu/S9WOAKsuRFlgeillxPbgpWKHjgc+Ilt2VxstsK/ndwzv0x1s3yH5CR
Q/apPGoon9V+gNw8yGwlN4/jn/HxtwVrOkx0772BkBImhYMAInqnydgdfv336Lqi5mvfLNwxTPJJ
W7qBEUctNow7Ob6bg5tw9mAeBch+nCz8O7Ks9iQR1ndD4tzrWuHBEGp/UZYZNihtFd/e4FegSxxq
Q97nQa2gf7eTmcet1Xmpal6/CZSUNhTQ1FNgGn6yaHUvDOKjGLIy4sZNoyG59/DdmjidGPfIJ2Oy
0GfBlf2eUxS/WYlhchYDTt8+enBu2t9GCGMKKj6nuL7d8tG6zpqcUE/izzEiMZoKNGFg4gJDRsyQ
7diWokptAw2mxjpx3yd5mDIMOvHuqNCFtbTkVsYIrVJjGE1mlBGDaAYkeWrHd5d59oMBDMXSV2GP
B0adtpobHLjOzkarwdSadxTzmhh0cs2qbC+gsveo4aYKcvTQ4t1LIgWFGAX6cLiumf53na1y3mP6
Tz4iAwlm7c/nPPK0+DrSboiMwt1NN/C6C6+5k3mqO/DdjLE4gFRcu7eC6qo85SKBqQBDDooWnBuY
YIKj1xUIe2+oamiHv9+KAnK08bB3a+gr6br2m5E2DtuXDoDRrQk1I/7MpWQ+Tvcba00JwZt71DtQ
/Jn7OhjEfj3kwoOC25iuV5YUO1aVixids9XcJWsSdp2/HLZwT55UPjXM6kCEmKz85W6IogRdq5AH
bALzQd0T5tB3dn7sh2UVLpZWUPnyZXi8HjpLF+1pfitzg/98AcwB63f0IzGdYbDjakVxt02onlP7
5WNkdDhxxONzygYbIjRZpHSF4kEv5P3PrdpaC6R+/9p4EmSXwKf7Ec8V7kUGR5z3gxJqV8ADrABT
SSvCu64XPk6uBDuwS2W6S9+26EmtSBVUGTsIF57695THjUJHSYyx/SLQvAnd8AYAbDge0zijQ8cV
P5dVoydNVy14SpL3WdXi+GtkyoRPW851rgjuKzt8ndCrHLj2gZtsqe1KY5cNq03i9qRBcogrzZnr
eyPLUlGRLqkEtFhyBTxy4ObgIOx8E0Ic1Gs7pbkzPZ2/x/Q+/kKTi9un7yI4FXntEvRRR6HMKCOR
feDAu5WbCjHkNDQGaPfjduoQp480bRfvDtHeGiont5asnEsrxQ21isaiuCXKNPbzpQB7aAPrHrT6
ssBOaX7D/L1ZECc8URa20xBcJNQF1Qwxiwp8cDzlTFYQnIyhv7FFMpr+yD+NvdRI/qLgAQQKD7w8
HNtBTKX292AkBYSOYdTkMjc7G1lFSHFluWCpSB2C3X1Atja3nrC9AiJDDNzF+/B0gcZYIiPV4ZvO
Gxp23x4evuuwgKNA7O+p0VuN3dw6RKOCbVCJ4I+cmK02fC2xrIbbW2GJq3B0/FYdBwSQl3OskdM1
dRlYVJ18mGaI8ookekV3uQs35GP5xha4ofoz4NtRYnfl/Cd8vE7smoxlCB3NhDpI9ZLwJW68+lIe
5k+D5dRu/1VMyYQbIy8auPsuWGRg2a3ku/SpaVLvjk9aUVwXXAhFBRIjy3SZdrLbqifO+ooKYEiF
YwvxpFp99yh4j807xTwW/5vSotrcY2st3xtk3/SakWO75HERKqWpJqK24rP20Xc2ZyNpWT0fwHLY
tS+A14ixs2ZjpHkpWC5vXVtFGmydYvphrfikZwSKrjGV3gbWJR2hGoWCmFPXx5BLnUMCtp0WNnS5
J8YFggHeN0KkqnmuF2YxSl85W1Tl6MznsMSWS/ZrPBlvCnjSOB557M1ccq69nlFkncfMbv4XLAcH
ZQOL7B3s4ZMUpaxwAoNPATZ8h1F++Egxzyc5P1wgNpo2WTBX+Q1+qBNom+CMgfXp2uJjr5iun4qI
D1bt7lAkrVazw98WPF+uYfQZBlL7OwPSZrzb3/0U3dlAc5VK5hDsmHOr/FMHSzBKRHMK2IYsBcTA
lqQx9LpGo45AYo9j5fox3btS37xRGysrEAmalmMejpXxvJUkbowdDSdPriGWKMp33Re1F4jzwL5c
TXOyo/E4svZ44DSrmr/BtluSpkTAJndtld+FGqD9CtReDCdVc5E3fPa7yuGW31kD95L3QCriAWFf
CurKsGuYfzt8NHImY6xB42dfS8S4wpw2Tb9CwH9A59COgktxhir1XmC2ivzDlTlvjunBVRqeXZJZ
iXbz4ubOvuE4wVouOEYfvvPIEIu4E9XoEhpFOVs0M98Z/VMCR1a6Tenh0UZOiKWo1sTpRTjbtL85
clZVbaxuj5n4y2lliv0SknriRQ+T4QFtAqZgxXX8BCD7kd4hULDWmFOFVMPn60onIVSin7Uzt5Hl
trAKtx/py/UgdSslwT4FrwWfV+r3bstMAcSwAv85B/rILHF+yuaXaHu0vtKBFVsTV+iuMcZ30fc9
+V4RJiAqbF9hkG4KXh/jT7+NIhLhTLZxMENTbUZzRE4tktTmxYHN5aap+wXrKfloa4NJBca7Iyj3
PFGiiypSvYb1/SuLO6EqS0+liEsSrU3Znjc1y/I+cCuNslXwO/+mQ/T00GA7MiYaaMHsYaRf6eRD
E+tQr/YgcMsV6ZR2TtwqqQ5h+adrNyVbvc4afd4sWfcccL4+rnVm24ZuPGqr6BvPl5SI7rtDTD1+
6q8KxkCLp1Y+QT6c3IDfeegUcNQm/2fV88AXGn1+7+zGoUu3ziHwyUoghnWWHlk7bE4As11eLJHH
qFWr8xfy9SVRfP9nuBXGNmZxmr8HH5dAjZlUIUNFShtGukqlEBaipvr+FDyOG7gGtEbpGFxQVIIZ
h08MSw6Pn87l/Wtjmpz1HCcF9hB4t4F8OXGQixH2M7qSE9+M0+m0uIlnN1Xzb9DPgAaDPCL43xRJ
y5kbih2uoWtPAWH71eTqbqbERcKWRIFFtzXKz44QUnRhLiKtYZkXbzWcqSIZSdK/6Fmv1/gl1TW2
8rTE1wqyQoFQITzrBVfTo9B4HEklFMaP5JDhWjL/IiWrFgmZJ1qfO4GK4QixP7Y2/e70BZOGH5Bj
JXjxanPU2sc63zCy+a6u362N0qgm4kYACB8RMLkkQ7T4PWKH9C/yZW4I6W7oxIB/7jHHYZ1GwKOg
fPt0UHwkRPTw1/GLfwFYmaxBi91oZJ8V6N96UmeXihXbs8C2vOLh7SqKUiUiajjlj9koEYkL5Xd6
Dcl6AZl9qL4WbjiwR78N2gOgiCjbnA1jZpyoq8w8+6xgI8spnvj+VoyEnjzjutdkZ6Tx0djNEDKv
uZci2x/1ZUjeWTQ7zQ0Xq6XNEfJdjPQEMR2YL9fibzNuPKTws3+FHcBnf/tr7cU0FG7M286r2ZWx
qDwu+fww4U1tui/lr9kZo98CPTgH8n/a0Q0OcD9rVhb6qBfsJFJdGo7KqaY2kVatQPKc8pMvCf7/
0Sn+1Gczz4f26NySascKQfU5mJIgAxJLqShhkAmyDq3HGNEGTGMriWnWER8MUyzeF7i2X88cEkwo
SGQ1XHTi90wbL2/B6M8dm7sQ60Qe3lJE4I0rI/kFm6OYQv1ihcGtd2p7tXQElXW9PUNmOs20jD/E
SuXBKoByh1nv+bxWTiYRiKjOMUikEVaPpV9OJ1PCltr+dhNLQMyxd0tI+ekJ1DfmGT/uDpmROD36
tIuK1oB7Z7o2z75ygMHM+uK4AXZ15J0Fe2npUfU3zXfX6MKEfAMbNWuScxElO+vkWDktg/0mnWy4
o3F5KzCerQK0t1tfM8eCc9MU9pc7NatkyeJ1eBpJlqLkuBY2hHx7KQIX9PkEz1I31FEDq3501cl4
EnVMPBideBuU5vN+77+/aJUlcYGzL+4DVJNL613KoDu8SpwNBurvib5upvHEnqootTjhi6JdRNzR
pDR9yA0B0poMUaeBR8lLurqdR6ra2+k4W3OBZ2/0b104xUF3L2Za45lzvUKxHp0QLRgs7KoV3cGM
tQPEnB7ssAVL5iwAVGWHUQk5qDDYJoyXWASIZVL5UcTABYrINr1gBx7gwPbgtR/SayVeTyB9N6KX
CxReOaHpRxYX1oU4Xj3ld7sFFPFkBWnt+0q72Pu6H60IOVB5bGnDc0Ojpm+xS0Knzo0gCnJTclB8
+beVFxmvxLLOgnc5GeBp1ESJ+XQV9oFVcbvbL7KQJQgoPEIxEtpA8MQEQFFz+lEHylccnuujTo4T
pJK0F1z/dY9GNhFJ1GnGzJLwNkG3ffDzEWH3Q0qnySiwaRh9p+qBjfsswpMUzK4LwuRhOw7uaWa1
GQ1DTskym/QNt2izm2yuseOB5hl7Olwme1Qwtwk4j7A8KSSzfwuNj7/n2PdA7DeUDieL1qCTBbJ+
uTD6A/uEtVUU+l3ow9EShnHUg0nWBOS0n80psBoqOzVzL1JWrDrYSmmqyvesNiBW638PrOsNd1bJ
IKM9wQqPKM+sJzQ04DR2oUmiL5vJKxK8kEqJ0eiWa0wHxHC8Tp3WpnSXv0IkFhBXsqJY+lAf6WVd
aqfFZo1uz4eydAj7t7hdlOauEx6jmD8KG8uT8w/fJShqJK1YGhmBUET5QPglWjmpD5OSlmfQdBLi
thlvB+S6wwhwaTzPzdyYWbJIgjC6kJpOJjRSbWx9RL3j0CH923caeEVHIjX3rFuNHd/jM0Bl7Dn4
jxngaBVVu9t7Ej9SsEmAO0YZ4x9Uq/SDQc2ndVgnU43fZPM03tpSza2vIiijKDDO5rhq7O1J5Q18
cAdnxhI+GtbDtoudm+PnPtJ6WToV7wW31ED6ctK3v3hBJaBBe7B+pHsumKkSfTvfIZybJDg13ryL
vkJflePEEeyO38FL0HRvD/qw3/AyP+D1Aa5fSWA+NKMgdKpuWttc2Lbtcotkq09/JsgtYHv9bBPp
PNw6EO4NLKrzEKq2Em1Qwq+JWgh0mD20Z846TqhS/nnAKk69j5eV7M29/BSZXWfCJe084Ozxm/Lq
8naStnVhDFHK9ovWND3x02hq+0m1+LRqDBFjFCuf64HkxJ96WsNCRJ0E2ZQEIrkrZsrxKBSerUPO
y+1DDfJ63ON6ZXMQ8JeXffH5J1zjkdQByUwPSCw8srnPb4isdcz9PBo3fEmHfZkVehb9eVT1UHXf
hEXkfNOWnuWXjIxQMUVWGblXBvV0xXgzxVc1KLVtPja4f3AuxQIriKDq3vgYYw05DjnJzgER/j20
gkhkGKIHLYSKedJH26ZdodJBcHRVCsW+Gm4ke/onPNIfgx3Hl7VYKtmvn5iApbLbPLZ+Vf6fSDtE
f51ufa9Sr1oueK96fZC/eyntrKJIgfQt82GMCI4kDyqrzNrQBCSx5j6wu4LtintoWXsx2bUTRNTF
hy5KMn8eOe6N4fziP7v5em+ZNkGBu50rYhmnwbb8eiwX98sRa98JdgWNsPu/TcbvhKVDNb+o73Dr
2g+ZNtq8eVb8dj6QF5VBzFaPu/QWkFedhVNE3bZgnbW5VV0Dt9bdI8xQu3sebPQeCAhNdmkVor7x
xP4qvH8xHyb7B/QUMS9kSb1gSXeM3A/2XtEyHjpsPkEqr4D+GdlvydyEp4njVsQSj51ihqIW1trf
79L9t/FuKOIeLLMPyTQiaVetVMaMDsf4dgxNGi+GwMwrjNwU8N25O6jP38DYguVjwAq8ELC5Lbkj
rE6jHk5ujt30+CPfXUPyIpL9X9K7mjHkfPduGTBQD5OKvLnVsQ8Ktx2VcHYC3LBXogjn6QyZkWeN
OLjrxZN427SSa7Wemij3auup5kDB/ia1Xx19zV22wu9k3AsvBJiCdqJSl1lM6KNEY0ZWLijD1vuZ
Av/D5QnOG33xyoSgdWD/+pltsFUPO04pO82w6XcAAN+HYRuExLu1Bn12lyTAFu6hsnN2ShQgZc3L
lidqzwV6/BQN3L2QD6rMZvqAjMnYubdIeX+oIHziiqVm+yQEH/2ZAvvCJOI1WNfduDS41fSA4siI
6FXRDf8GEGuRfR8JzC7YYcjuEd2u5pYSyAM6r6ww+uRxvSnVc+zkIpSWtydJukELuVpbj6+elwc7
si9ImG0KJCVURSrANmO11CmHmLNjnZjh+z1cRFaMuFhn+yYgGLyynNArR8lMd63Q67VRMPmUS79S
E0oAAJ762TU20fc1n+XsThMFG1lpT0JPmIlaVG3IXMiWaokCW1vjCDmLIgj3FzhfinPIzFJTSxaA
CsBqdO5atuxvFwW3wxRSsdwJNXRTZtQWiePXD5RAh1FHhuLa19O3YgedcXjUHKqIX36KE8zHRgUV
xq7hEC6ljVvJWgDM9t44bIdWzGty33KSoadcJ/0SumGpHOKjm49OBGcMFOPJNpgZSPCzeb5QjBu1
7aiwKoOO2E3RfAVuIf0hg1T+OvDty0FgcGIxz4JLckCe5Ni5MtAh7b+4Yf6WWt1pZ0BVSO79HRLG
XXDFm1E5yA+DHByjpL8maWmePyZoI8oIgQQVEQelNYEGiorIdSDpCI7kdD0ZgWQMjeDvTg4ejzOE
8plv59mjUira8xY1sv39eWepHzKkKHUKmIplMtppZAroo6xmLAoi5rDvgFWvVM1SsVG6ngyBEEgA
EMlqYktF8Kw3H8gCMp5ZprvszPzP0enURMIwTQIcbKXmxi80M0/iqEbjU6rrzLuMVrXuS1TneGnb
46xhYuATB9yyn1hCoITczHZCLqlYpkdGSjIOf1bSvsdg1AuSCiqiuAn6T/b0dohYQ3J7Zxx4H/S0
YvGeqMDzAzWrJNBf9HyZOG9zc9atzVfEhf59jj9x+HLqt2mlSNrVzCmUiYxSAJ5hblouKOectOlN
KBI+TpO09xYDPyGXPZsmLoxcGOZi4DkAIL3Rjf0eB3zXc4iOEQEP75hnF25Dsx3y9NqT356Pwkv4
VcX19Alov12VZ8pQA8heVWKoJX8wMbLbyFztRKM6/w4z4C4PfM+froe7umyWaxUCk5nvSOHafsxX
4w9lGu6y59TVy0A0up88b8xr66WGBOX5N4Lppl7+xeYXpQXqADdRPfKc4OUvM9BcvA+B3nUl1Prh
4tTHzkQQg4JdixGetQTDcIqk8hJnF/B3rhrbJLoWqppPIk+1nV6E1n1x7voaj7duGeVR084RFIkD
RCQnSOQ8HzHldATJamVkZEikHNvI1kyNp8Fr8ycuqoQt+w0R3jEH2LRAFaGtvyh4gtuSc007dDQf
MwPX/NU9dFeHdjfFYwXSjkTtSocIWsv9TDgRVjWZyDhaZwEcWNHKdmyRupsOiIZ3GFIHvw5QXdqB
y5KKiWUFJNn/U8tb61SeQka9BKem5WVV/A6mI3UZa5tQmRJrv7R3oA7N/qwSeEkPOaGVO5tF2bTa
BQHGS0sc5ajzn2v6mv3sxePBlUmh7HRCcZm1Y2JzIwCe++TbxmRbKLeLW4fjQZoGB91LKs5pV9cg
sBRXspCsm4uP7M+yrnECyAp6Nsly4qp7WTM6vN0uwsYSMommjQBlYSBeNRMmaI27RU2XWPoOaBmN
/vUiLhyNXEH9YASqfr0+5VYU5uPKqevN6ILxdcBpDlElcyfYDPpDOfI0lL7w3SNL79F+izlQxOlU
TUKKP3ud2tS+MDXoo022r5ovzXo480Ds7ZGjUM5M/hsLLteSLoy4acbyAkLZ8Vi/JcF3A7lOM0dA
wCkOzduRVSrOoaRasKS2gWXwcDRomt7CW/ZrLh0jK7+NnMCqw0/Oa9nNWm24gtbvUDG/1uRRsl/B
gCFE+vqjddMCZdFMGp084kMIGOCV6qUwpSGIn01ZvgeOgKZdcnwGfemRc6jfYQiQrJLtOO1x8Ae0
rTBwhfK5CcmTA9+XkDW2zEcbFyA6wduZ0R4QV2TgiI90hvfDrmkbtriQFqFeFAlVSLV5OAtAYSmu
RAG0DEPGKJl51dRkY0dkiQXKzMuq2iusKaWjcx4rFr7riInaS4z5rR0p38ILJzZOMcGiEr74sf0a
BvQHoWGaEwI6ajyMb8ABdysxtFckWiGRovrcnC0kq3aB3Kczdt2Mxxsl5LWz/ZjC/9zjdAglRTMv
CtOPaPbkjFo4JFMdwQOIC9oyumQjGNEMEHs+dKduRBAxgE8CNDBPtZc3VYptga47lZ1BigBqTIgr
ivPWYVxzBRSIxM0E7FuKQ7KFT22IaX6vEt0hu6C5SlMRUlBamboEl9KGohZIwo0inKCE33wToYgw
ossloAjkw//BWRFbRjV8aWkHe3QPuqCpTgVsJu4XVnF6b94FgPx1MtyixT19C5vbxGUEd2gweEto
ZZbJ0Yuz9mB/YHoDlPPA0tH4JBoBQqaOnv/bFUYXUSglyAc7cCNOow+wRIE48m9Sp6u5ttcWC9de
gIRYxx8gaGYfpnqq9pQcq4C53ux2dTzhW8EyA82NW+EIoA5eeOzUJvI++TJDXgD0l7vwzGXTkgkP
weN0k0VeqWyhRM4aN0c/JTwi2wk4kM6/L61ANKk2G7AJmC+P9zWDptHiHNTo7zvc3QsIQlBi+/Ra
fH3KbLR3J6lZSiaLY4e5Vy1Sgc9AA/rhu9leSh6XRepbRj3FtcPqEjUd7m8vBlbO2NTklFkdUeB7
sYgNxMt2WUm99WFSyftzT4CBHPq9fCIwVx5AtFMcWAO2VRsv2+BeSnTwIJVgG2/mAqrvkRSurauJ
VEDJBWoTiz/SIFyUUN0RRFFEsy9lzR/5xxy9se6FknfeeBjRLkiILbjafqIJPtDugETNZ3FGo8AC
dnyWeOEFJ76rmpa8qDErTznpKp5BiU7MyQZf5kVow+pQP1uKaIu0A4AgyhefTxiBSEe8OB2ShWhx
Qr2mLXBJKD6y2H7tCV4z1oIDVKRgFotVtVbGRp969n//ChEI3frfN5AKgXfDGhyRfAo860oBJpIU
fRZCOTr2G9bdSXn5JkD+QjEV/8icXZt5g/Aaknwd+5nXCpEJJdMO70r/dP7kbiQ3BYqC+UXY3bWW
ZLfYet6tDCnjyk3OhHAxM5/1VqmBfNhjT/OeXlEupHWJKPyzEbjVU3S73Fxf4wUzPSoPu2ByUPNF
PSxvvlHnuo3p2BD/gp1N3llxumkEZLw1PoYKrG3fLLc3x7wSBD40YL8ViGpNQCJO2pr3Q6fs0WeO
IxQ4aX9dhLQCGqxiiUW5a1+x3ZFnrYSU/hVNdlhTgoFKeoEAjlEgFv7F0UNU2ByihKqETS6piNhY
NHrQYAsvXLSWD+XNWST3PQjsouQLUvl7SUtx3p+h1qLtu2oAfS6H6XIfGpvGLfk/Tx5bATxEOO0j
Q2cgx0snpMNfWa9Z4O8dp5mwD4uTxSCKPFMEKcBiU7o8tHYhrQyFF3JJAu+4GA1ob3BJTMu2VjHX
JQFQ5OBTOIRz+hr4kN1vq6+xSPFs9X1NqBK3/aqERBvKSIms69/xqP6R1Y+Lvvnzf0Qevcl5I5FV
hfdTz9USOYyHZjqvuDh6G2z9uvUQPXEflYtnFJvpIverUwcYW2zSJY6MUgMpcE792fMn5e5tPxVl
NqYwTnm/0Ti8OQSTIgUaRsHhdgfVoKY6eJRLWcX4O329ro5zlyTaiPhY2yqMZpvK8eik88qr1XBG
TmrT+IujV7PRTp9bftq4g+/4eTzUy+/WgLuLFrvIu8cOZhzsgEpDAw17Fa75oHhQCJaoKHMgGULF
0ZsBggFPkS8wJGk4fYIVKU0QJh1EClMVfKks7YN4ljqYI3aFwWbSPjVRw+hDEL+5JcMllYpJpaNI
+5ovql5RQ4nvs7aso+olH5fL+T0t6fYQiI0+TiogbYThEBDWAq3PJLMbS/AJAUEp38WUdsiszkG7
8cerEE4s2CxiVtTORw29TOVaN+Kp23I86F6lhbBlbRwtqXJ2mC+gZ8TaynuJO4hv2pQ4R6TzPRm+
7N1p3aGZbJ8fKqceEGWTamTV+hkK05d4wjSlMZcvJdUdZ2NftTLFytUDF6JF+/mKjaDZdi8ZUolm
cuNhsoq7QnEy6W36NsCYEZKb53IiDZkYGvstjha+vWMrujPRynog15rc7OvrExq0jV9c421eDUeI
f9yOPVOTUgDL4Rm+DvCBhIBOYGanH0OomBONakQ5GFLZVpJS34U7ir7sgW5oXpIq/1PC3wBseXHf
UsZUDLgI+I84iRVmigf5NA7Lhbm3dmdNZyTDQdUiD6j0ZdyhMVgtDhE7ntlsDdeZsR8vOEkcUW4W
cRIPsJihen9TKq15WAYVRDwiNGirq76Q0BvHgBi4NQ3Q1QxCJBwmfyAezf8j0/vpLzIhZwKwfmAa
ZfCREx/8NzzTRWFegAyoWF6fsimWNACaVsZPFrXVwiT3nR0C8O6DOnwsTWFIEgT2SCZnVpTOAM+9
bfu5yhrv8g3G1XiVt4ar6Qk9Ow0EHtP+Mx0MKuPpJMqlfx4atU5tJZ+aJEd0jTmBmdSUnZz5IxFg
MRNWcV8+i9x9PAJy5U12RmmtEJNSsKW7tsTvSg7kYJRQ42Rxmdb1fqG75T05UTpBwHoQPbtvC3pa
Csf6r6in0KYmjptAZV4njjp4uKcg57ghUBErh0qmukrj3ZSM2M3xPhUU6FCuJO589WhPHayoptEf
EGyn5fRqoYLzATdnrDvOs5N4O+e6xtyyAUkWtK19f6ioZoV9QUGDNxJLJW1x6srZtwGqJmDER4xt
dU7A0q2dk6qMzC/UsESBRDz6+clUcV+P/E31vMki/kXUYtKigrgfxao5BoPSbCEgEoLQWd6q8YKx
u5J/sAvtz0EANOqPA1J3cY20JxgLUkutnvnpPDF/Kciib1xFsT6UHeL2tZS2kX5CJ4IcfIG6Vxt8
GJxG4OHaH5BIuF6OP8MdybntImoWqEyAPrcj5iuiUUOgGOS1BhUCe95bcJehk6ktQXCwGGBh/tOz
q9HPLFn7Wf2a6hz5bGB1gIHX1zv4Ig0IRFtGvAdz3PuYXT1bRg6duNHYxpk3ACofh876lJWy0K8E
R4XOvVnWJmFIiN46hnVJi6PExAVSry2QQutJOMHHhpTx8Tgsytmdmx49AhGlgcWb5p9boy5XDIPh
B0DjGGuIc9+XbhTrJi2O7cro3WZ/rrxP1DSPYsRJ9DPQaENdVZL7V9Rd1y/w0B7rS4bXjHRhzPFD
XiVrUY63zB4lBVgXug0HkMaqwcf9vSky353qZlZKN4gsupW2GgeA3CRt+uqeIfnsMlCqddUi6JUW
aicxgLsmSDSqdnvkIyE4Y95Z+H6fJUeoq+mCfnm4U3SSLrlHhc2G2ciHLh/qVlvz8bcID5RwaoEQ
IYcEL0zwB4OpluSfYWePbY4IWe8vCAsJI1inCUPiYK/3LWezjxa7Dyqf2ZrijEc7vZLYXyj9DcT8
5ztS8f1dNIaKtEac7+QpYKNth6m+5CiRAu6al7x7vY0u3QOCeCV+V/xksu5XyF5fid/FTNiFkhtQ
0w8qX/hgNKCREfOLgBXgVabwxHCBllxYhTHKtnF9QBwCuJRjDRUeETtMmKz/DZT3AOfumM/Ewxu0
qiDSTfTqfKLcaLZxO8EysiGSV7AvJkMwM6hxgoaMQFBoNV/mydSvCGvX6/BviufGwBn+K3g6CdFB
JiqHi+k4LZOXH03UpATLyJSAXXNG5H9u0cGdhFxAYnzfDKjYv1BZRZixFp3V3RokRBP3PLhYAf/v
PaJQICRbCAA2+vDnwMSm4r1fXsrmbKILQD/RpJsyFCWao0PSd1MTyuAc6+CrXtmvrk8wY556ptzI
LG6wbAR/pPko/m9omT1JPcihSCol060KAI5102P9i3fkwh7dW/PKt38t+o/zjmNWzx3fFHHOkjUU
GPmIGmWW9s2rHOUeHUGnSgjr+5RmvtO89ujPcyKihkyc49HB4LrH4n8TV967jY2rA8BwDbsC7H5E
vUfuk9bYWM0SqMl6m2HVYKO0Iv7yqU9/Ri631DY+q0BJ419pWxFqJPOvGFRlqMbra02zh3uHhpNo
wPMPwivUujmkFbel6GY2AgkplwV74XkqL53cZ8L7j/a27Z8iYu/tHFi53PVqVQnXCfDxF6bRAlQj
Gk3Sl6ZOsc1tTSfJPzp0S+2Zq/s2OnVVuYoCjzBWxp3RDy4+D0KXCDea7wLTzQ2sJ0TziHw4YJg2
ZKmpao3Btxg+pRaySIlUmK0oRz1ssbdZdq0gcp8M/MEnq1fsAmCKNvseEOROKdJJ6Gpq0b2KbPLb
IDvkK/XHvxh/5DiiL2H67/zyzv5M2TAyLzLO86lYvQtApDIjw0MDTQxrtWaiIBThabfKOb1vmGbl
JcvXTaaJkL3YHVZwOSDtzU33XUWhcjGIxeZijrcc+0sRZ1dbYJRP5sDY2eh0i2wa8N0g90mdn7l2
V5OuVD3xeFWQw1v4ZZhI3sgs9qlq5UeqRbcuN8x+tL7grGFBUI1lUDLlaC5ZbqVmWrTG949TkRg6
JBIVOfEn9kWfnNimLx6DoKLQGwZb5SUd5foORi7tKd/BYNdTkB6AY5RpyHWsS3TXZtcRbiAYkcwZ
QA2hgDqCXUnffH7OaaLTdZwSRit+i5kTD319W1KNzzayOKyx7CdHxfiYhPElgaoyb1joUOUIp1zO
/KTOJ2Z4Uy4/CiDM+vQcwa23awXthF8pmQEH7OEqd8dueUBWXkIvw4V/91YbMfUAMwFwFv2CZ5oA
esjU0cX4GMkzP7J8NvNTAFUpbEUNd3ImeUV8uSMRzO+DL7wxuaxad+S19x3RiLCfeWcM0LQJMt4K
JrRjpagOOkDaTmexOBSouJDJCeFtIrFs5HvgSm/zbIrbfdubt5Tu3yq3Xz9w9rhEpfyGNwK7epBP
8sBZSrg8rwi35DF+zl2dI90Q+NDhkwbcXEnnDK6LGWG4vxdeDkDGWPkGB3Ce+8TRGeYBYXoHCIDM
cxfjH69uRw+/MHJEZ49mmlIZbkm3yWIX/ds0s8RLsHYTtTgI0lvV+HNIjfsM6euR6dvm2tsqmflc
VgAgiHGcLZyXdeKDGoTVorLcL5uJIQMXZ9/ZePIpuylLccI8wJFSElPenCxvtv7T7PRdnIKC85u9
9MVYkWiyKCHvG4OgesgQNsV8kKVDif6WAe8GFRJQPaRtJ+e4yxUmZm56XvjdB/mOF8jLJ7UXEAXX
BYKFvYbxurfcD8bGkneqyJQFTJTI8kJimlKWp+pGNTp2ykGwzEd2SUGMDwP/h1Vn+/xcH/8/w3VO
iu/fohZXNm8iWgSYjfuZ1jgM+CRP8EgNXeEGLWgi8U/gOTWLj4TwkVKEIoBJAIyUyMyjaPLYTl1t
3xYSyMJVBmFrbO0mHAmS2Qk80EFh54Q9yJ9fFWqOMJot1ArlCKTl4aGJmdPuVjIekpaBCCwsUF6Q
YOhDTg2A0ImnG+UWA7Ar00K7VowkJAhvqBk1Wt3YkaWhnPRjgjyK35iPBeYSc48zbLVoqqZqZrWo
RHj+6538ifnyOGrI51XNUUccr8pRt1BwaRK7QiljwmTTBkPAvgxh/Igpn+XdeZasdP3bXfGhHOs+
8nn7/ixd1DKips9vVc+hLLxp5TZJ8aRVnG5q19CKHy7zg6apbO/0VlteMyLyg2Q31fuP1v2/+XcI
xwxWeY+t9tAHWdVlt53L5bhfsHptPtc2JeY12xiwW2usZNgoVt+yAf4Shipvn0aCE+xwe957f4ZC
ZtqvexlcaG+7EMaSWvl4+Rz8b0EdzY4xkkns/cRpm89BqQjTO5AjWbelkVBxfUp4ved3feq4k5VV
StILBTHAEOxEdWN897gDX0A10jFvd0V1zvbdAKp4RkgPOt9lEv/Ok0yzTvvwR3wkfg9SN+QFy64e
+a1aqJQQ/qzC7ByZ4D9WZNyxNe0wK5JE5poVKu76UVdFzUiyMbFN5fGVO7EbPnSLc8StU0pBCRtb
7YnW/dpKQx9Vnrsxfe4wMYss+Ud4BM39Knvwh2MuQn26ugrsFLZqYXT5wrkH53EhnLXPR7vmhZrk
Lnw5yZ/HpPidd2et41UePsKT5kr3QwfnmKilE5EkERzJ4jj6rq+O9a951YVQZzRQJWqlDRwtW6Je
DDWUhU08jI8HHFdww/9NEpVopMVBmrQunZGK0cxHROtdtBJlZViOGBuJOWDSjZ6qcOQWsrdAqqq5
YAm3y/PtcSY4xPmg5QQ7p3Bs2tVQmcA5fARNDvPhKjxyz90S8MkeZK2qPkApvfl6Yvjx/TiE4H5V
URyq8SQAhrecFmjofdAJ8/c/4ALzZa1v2RhKRffg4+35ejQQ7fGXtDFbI2I86o+iBtyxiepATfeM
7V+JhIDOGi8S2NxEPq1sHbT774mzyedqZrowGBQZD7Gkn9NRCI4WUx0hfGJFO9RUrZSrGH3vzqnw
m4sM2ULiIaaYAqWKkJ1FoseE49yC4eCCNIOg5+fXMIfQ0JXnKuh4OMZQDZ8zeUZIE45vCKDsZDEg
qVSkvWYcumuUrleBusF/8vObyLD6nujn208qC+XnjU/ctKPuefdLqWRk3PPMZWuplUXiDmuzgDCz
Bh/rCH3MR6HYiwHJK2VBsfaRBt8MUERndxX2vwuwfBFQZgZikeyvaB9sGKqjQ84ECHwgmMFoc/lO
cnW0rKKrjKJrn2dtbA1aPq4D/g0ePZsmnilGjgZMA3aMPulETktGO4pFMu9dXcCJeC0cb0X8d4Iy
+0wQaT1kSGFYiKgQndBPjLSApEBxVWsblyrukqH8jbE7WR40Z/mJVEyjbcVo0WwS4ldSN0SCxOh0
KTHUbmWjH22FKbyg3YldaVtWfpurfR2dXt6BfkgqmTqQyFXlDUBdpBYBxqD+LylCzI5KTdmcM0ST
9mZ6fb7URsmUvJCRkiEEbh3ZruDBF9AOp2tChYOM94bAdiWuoqJ5tzybjt8vlFak0noZ1gAy69+B
/FLctJ/xXZh4ZkQ6wzPISB7fMrh6zhvIAdPCz9JxBKok8v7GM3JUsbmQSDc51yt+5YBqpqPEEtqS
4WRM7cfzu20N6wpSk+YmalgB+viunGZHOHCK+gKQMxRrE1k1+hfhJlFyslOqZquu5CSl4KJgzVtF
KKlvt2mO63ZjHIPS+lX9g4f+DrQuruXHTnNLy/RMXHIZ1xoW55U3Ht3ZIOEaV4y+fP4o7BdgKeqV
ll0RJDk9/ZAjET+WJzrnPEvv0vn2SeE0ZZYiL6/ntCpnx6MwNgZIDd8AdCUiqTcKXCLaTjgvA3hv
2mkEQFdOfxkVV5Oq9jZvstnDC7fFlUonat2Ut8JoLqD02y0zqYMuS3K3tcoHG/vEFP4MXpGLh0a+
L39mP8Y//aZ1vZLc/S2zfrgTo+8haYpJmLDdSfOBqjcFEONXpAanvU9NOTVK0UM0nkef9KlnbzNb
avnNCGkO5RPmGkmK7WM7UK5ngoYzLo+/gD/SogxuEmBpYT45xJQA4woz1Za4QUht1Cm49qmeGXnZ
KSPN1F7RSryteCJs4Hcu0aD5MXuCrhhPL9Yo17dIFBTFSCkzbUsgEj07gWeql18KDiI7gz7Jm51V
PNYKg0id7fy82L4H9NWBexHboDk3rtHU5D1FjZ1Hz1QYhuFRn8HunCjUE+dTeRSFKimS4Zjs2nEt
v6GI2f1XMFgoGILfcXnCSYYG6KXoYE5B2S1Ew83135v6W5mTBWQhU49Vzg9WlDkkagUQwQs9axSl
4O8B5eX78boZ7mzA16zA7sgV+xRiuBn37wm01+PsrRaCABfAUCrOP9+4d7GsoF5xBsE/qYv0nPji
MusCm+H/72542v4l+iRTUQPxnJUW6HHi0Klv43C5Ur+MOn1uei7Umd0RDKgtsnsFFRGWoFPd9mOk
3OTyRmVJI4ci3yXCr4K0EVSHkozM6hRNf0I7FOIP9Ot+kslKvy0Plxt8wdNVZthJ2qlgf2CtJ/YY
YC8KKSv3/0jworg4XP5BC+dVSyxYqr/E/AN6sLNmOv3xcYZ+yRgtyz9aOAqEknXoaJKEETNtc7q8
6CQG+nxhBXhoRzrwPYuh66+m6jD0j0pGRupgQrGy/AKUhcVy5qFy6WSLmy41qNEc/HVwSg438B41
A9h4gWgbOrWE7aj47P60BAF9AaZy14IBJnhU9HjNMx6GyqNWYpjOnV5lYG41AqcQ6YQ5H+3XJvot
ohR083Bz3BYkqar/ynuAu99ODRMyD6+qM0g6hj9ScnLBR5vkqKXQ6MRTXh/2D7sVyKG+uVc4jzRV
AwKuiZsgRNdSexgvaYCHFdoIIH+X084tCcNd8V6nPtFdwqOyBprneBYXPjBskzJYKvHLb8tPkwcO
gNjsZTltE3mTS9bPhXqW9N8wDrTkeiyvBsgJRDhrkSYkuarS/YRynKs8jyqVqrCJIE13oMSxoWeH
yBZ50rYjfFtW2Fkq/xtYm+J2BJA56iU7FpAnGQyrda3+7b1gEhkHYUH99F/V8iCo6MExr7R0ZhuN
TFW5nhuIm2xgaxjvaaIkK3qb+J4xBccpSBh97eHF0amgoVtPWvKBOGvfxDkvekm2jK22tmVPyEqu
fttxQUmLpfbBbt8Rqgp6cG7c5dgpcEKoQ33k0VMNE3FDVEX5UbIw0WIT1wNVdMoRlEjj0f+GlWRR
H9E34GVtk0gqMCJAKpHAADKAu3QBeA134b5187qzviwM5f/GwiXDTnXSNzqyUvrPSgSJpZUQQ8BH
HMDzaO/X0oWpjiVvab3IBE0gQMqsqDHVUX0AfBpTTTNduhhTt1OwAR+BXWiqXYLulwktmHk1yzW+
VdpWqOcHgVDLEdXOdBVIhnC/+uiiCapuCvthTGj+q5+OhCYL3zkR9n9BukHejgZDCzYYnd8FCCSY
wbjozRa8lFbfJ503p5zs3wmFyXDVgrIA3CWYLN6enBEQ1UeyqIcIUpEPmpABND/imz0sCYUatYYt
M7Zvm16K8MbfyUdgU9Mgl2OirqwGdoCU5feyu+aE9NU68Ms+l6EIaFfX4UpaP18hPD4Rx/UFlaOb
mD+Er8enCKlBCC4rK83LTJ+/6VwgRI4L7d+h7olqLR/IPaZPltdxMbiMICzW8KJKJKw6hJbMnmmL
Am1E7zKvjTQSlNu8Eby4H4cgrHFtQk9nbObIRgJLDUxMsyggICAoyBCz2VCNSrD+XvW3EGFGZbm1
ALhEX8G8HPho9lk+37G84RVLfzAyawD+ztmDwjVNTp+LtD0U7ZxOIS7TS+FQ4PXh06qEGfVN9JAz
y61hJrwwhoi15Oojmi84mbyPo2sYRM+cz17OJ/xS59utw4l8kcUwOK6EI6VT6Cz3x0SeNW1uTT8G
2jxXdpdmBuiZ9cZmWn0HZ8zYEA974PYduSq3PdZazHilglO+g+XwWxR8+3gcN/56QjVZIPhdlU6c
i3WkTeiIaKGTu4ZUVzM8pp00i68Z2Wsr8Q9VBFw3m330HVYl5XdWV7a/JejAkKD1lU3ANHOsQMa2
VmbVCVlp52lnnon5bCfuzzx2e5Wxe114hWsJZZIkvz/hNthIgaan/pV567dXaKhxY8H9qa+1ghB/
qFsDJuAfZxf2s3dt+5lV714AdqbfRu9MCYe+tsqM9SJJxQ4iEAhWBT1Lp3afdzgxyq2OmIUfGIvC
ujArSgs5T0KNirP417eJDuRhBDJ/CeFHDhbXm4z+60bBwNePvKx6wrCaDDsNmtEJ7GOlbY/FWwVw
wLhD9dUVoiQBzCJgC5p/YmVTAanH2H3DNVo+Wdbwg2ttd2HZsoKCq+JlxPQLoz9/ZfAzxxV6bvnh
w7XJNkTSL0rXBXAW+LMNpuvGAyDbH1zy25sfg1NmuNcrdQj1hGmBYLfvHN6CF1GhdpZ44VVXeiTm
gvWe2S9J04e88j2e3ACVaFky6jajPMKTaO5bdP7Usp5mqE+qDCI2cOUkgCUyXXybin+i6nc8blz1
bBegqTJaD3HS7hG7NiO/pt0zA/4mrm3NKgfFlYgARNPrXTdvWjrpC8n6P3Wzq3YrpvMJEM4VTUcn
tvs8qLtqWV15PbSSPirJcdkyGiEpsQZf4waLGGSMhNDSw1csuI5RWDMimPEKfRZL1fokTHLul03G
+FYbTj8kTBQYnkuf4Id2hYfxefuyGEsLaLwVCe6aF34F9Gy1HYEki66fpAzgv0XtBkmtTyerPMpI
G0ejggAmvcGXnIktines4E3xuD7pExfmXpOhKTuwuMTC6+Oi/LtlPA4cRwWEcSewxMKH9tmTM71X
QcqFI0Bl6Yz00MjvZh7RYB4sAcb6EDrcZ+h9HBQ2VLUWKePyn18l5PHzOdZy4q1Wg+/0BUtVSTkB
eDIZUuTY3yXdJY16tHA75B+ZV7Ldz6FeYsQf2Urzm3m65L22sxrW28tjxbXYLwrqW/NVXKt3T8re
PlVRTGfBvnoy9+lfK0KFAYpzVhG1JFpX+oP27dhLy+J3V21gCFNxienw07Z5CeMyH0T3nhnlQtYE
z1vo3Otxs5i0BPqKcmVlssjuamWXbC0zw5Ib2xvCJ+SFa3Y74QoEkXfe2fuy5uA2Jx+QdT2YQe3x
6w1J/I9mFU3jYaEnDPI4jMIBjwhI8MCYJ75NQe0H3wgU3kdg4vI6J8Xu5wqeYd4alk+cjVpQ7Hp0
vQSw5gztISQsnsottLyWViUOeqPwiqDHiA3FcrZrJw3kUWSva+8HfX4xuXw4AgcO0RGaXj6QqMu1
xDzJrECOkTCscH+uAWZ6cUYch9kcRg1c2n49IhLz1hxoxqQGBWDhh2216uiZPBHWEaPRgdV1nXao
fD21Z37hGp4gXro9td4kPz6paqMWw659KmbTNCFN9BH5pNzcOx0EAClBBELr9ZqRdss2VP8KucZH
Z+OSmpWKevYn2bEBJu1NhOMMJLmeQbu6NQ2wuuh4hUYQro8EV4HVPzXkOXBYRyFs/wZGppTwamrf
t2YXqZn1ar3Cya0gDOEFPnckWP/MR0cdISvap9BaepH6yknyzeQ/+vd7qnlvlWfX+dwBdFjRFP4/
B4sug3k1U/DAQAqYeK+PIU8OJZNsmRGE+scQ6hVcfoaeJtaVUk038OSWlmjAJsA9wQkmz5mdNHQ1
ayaXACfugP2hxCpNXuuBKuS93qAyPviH1Ox0HNWNYWE/TFQ5r9OmTi0SmZRNeYN2QIXo9uwZ97Kh
mchbibyUOkB0o5Rtke/YrUU8L/MV0ByPohe8MOl/IzADruzyqmeXMxGQfLH4DfSNQv0s9E7ktCtY
nBgWtKUe2+6GYrfvvDcjyD/iElKcmq/SjpaACHDWFSuBknfy2+KRF3pAaUR3zyGE36MSnEA+gqok
by7ZLYBbgg9/ECVSNftl4aavQo9Gh0RPJ66nDPkddt9qsU/wkbzwV3OiKI7JTSO2Sk7KUJDQPhxg
PkEO7X8ZdVuLF36boA2LG1+ir5stn6HK5xVgYRSDocdic+OCISNee+LbIewcaDMDr5FphXcnabWG
I/xngBxL7oFg4xzK4soTdYyzfoHWPmEojyyZCncw0bH0dR+/r81yuE2sSGnKBpQCtk74v3tW19aa
W/MkFluodakG2Q8Ur6lw7r5MKTTL29B40yRueTvpYlZfmmMrrw8if31pD/LPQ7wGAUQdhLS1Irhi
++dLn1JzVG7LVAzM1ONJmMCTm73rwrBF1AEic4l6aNnh4Ues0wkFtI8AXmjJoH5v4VcvnjPWeuhr
kS3PlqyV9Cgx4gIRLpBPCaysxnQgjFZhQUfqG3PWkiKWuuY5grfmYC6wCvP2/8LiOxE39MrGxWQn
PWQvOCmKCM9x/kjj+z5uHfBeCP8ps4drI1kgKTnTe077kx2Lx9Znyvw4cIajLSkw6+O+XSqC8n7Z
nj4SDJDDj6949V7xUeTVARFA+ZXU+LayAmtz8SOTniktVgAPuDJHnkZqZbT9R5mvn0gpoIpLLx73
5uuirjDIQm/irThpsu8XCK0tla+3i0vFoaiYF0EGrkz+l2T6QAqmqHGomHBOQ7YwqfSkWv2nOaSJ
iMEMi+tdOLg+FppWMLlRBvubm4U1Tf2jN+weVHQ7XN9d8Vdd48oufl/+TjSbR7DYh5p8X5saFW4G
vyAddUZmLZYPliTLnsSVIJ8ZPMBli8u3/QMnh2s2spnzrOYoy1yYRzKV4LBCg8yajL+Xqrf1dywU
F6ksJvPYpg8DChBJwH6gojIxHTzgU58LfsqEzVJd9aeP4hERdm3beXhZZSgwdjHs+X+U7lIfLKo1
rl9HJnxgZosLme542JQ2ZCQreLQf5C9rlZJ69oKLA4uKoT+Z47tWSYKDgKt5Xelq0Yoze1cDtUl4
DYEbPD0kAl9Z0iDnIQP2ZGjWQJ5nkNiKJeR/F9qTUlff7fBxM612sJkFQc3m29p/nDuHkfN798KZ
5IwPyHEB/dht3j+R/pZEs0OprhROLD3n3hb1fVkrK5uMhyAKD3xNACqRmgYdPyvEfWfYm2rW1CsG
jIIYW7gfd483L2SNpuigfGzkfPq02PlP7KocYbsNdU+pNZ6qTceVCfhyWmQXPUvrjbZitxl158py
tFyyJdjBJl9m1bTmDH0M3iaf6F7gd6CoIUOHkpwGQUmHiLj20jzCKNefxsLKAEYND+N84SHU2gE3
nrLe9E09JjWeiKLgef6wI6HZPW3+6IW9SIurBnlGyuIEtSD8Z+XWMW0UtwHo8q0+0wo2x47wa18J
JY2HTEKVYc0Tza1oJjAX+1EMmowPWWcyUsVY6FqZDLnZ/vbpyn9HSLXnnILGKyeSonxtfWbAbDq/
uba6P+eJ9Fws3mFRlYXtJzvbwh8EgerTZ4aQM0N7AGrIZ+UT+CuHy9JCEU8f6dDcLROjP1z6RJGe
ElKofBIFLZgSul276asFJ9GGZR9P5TmwXUYnffx4Ldeb8n34zCX2l4WH7ty0rvlHltofSm91nvZ6
8C1hiAm+CD5VDIIdL2B+mFhL56YKPAZ1UeSef6R/WUMg/a3hgMQUE7DWHYQobKFqLxAzxgJpwIz9
OMVAkyC1VQQNZegRN3OCGARVBRNk/fahKxYJVfnB/q5JYlaOEVt9pnPAvbbRb1tFbuvfW9Pub5J+
W+n4cLJhFllBeX5prynnOBUqpUS3Ce45K2FjtZn7ngvn29g4azCifSIy1RDemzKBq0ztsI51NSwx
dYZE7sNwkUJJM8J0uoGDZneZ0LgCrI8qYb0JD50f28HhdfS+7A9wQNn+apqhLtOQSqKEtVsSCmyD
N4qZB+HSaKMcx3l9h+8yPvMrOoZAeYbR/1svZhAMmYm735W4OJ1WhX2B6uvP1T9XBRgl87Jmnva+
K+HvkYiqQegPVZGyH4afzwtAh/0lWKQFHilXpxZX3S2zTcI0aCgrggbJw+8ntCudnl14GKXtEsEl
XBtogPgJpZQYt3MjbRCzioMXjdy/bz+HfzDKrDmRc3/UkzSv3OL59V9lo1hRMMtpHw1AxoNU/tSJ
LyK4vmBMV/o871PqQGLDlDg6k3U5XoitI1OJezPiA9D1+utxCcgItF9mVLMoklbGG7nYTd2Y5nti
g9Kzjuf9F5hrf25mFIIz+B6M1u4eCtyij+miySeEfhHMkzj99lRN5KxRzhZb1sycjqH5uLfPaW3A
BY9TN15tMyRitNScxHnYVP0LF9rgNpTnXTCjzhTYv6882wfwNzAVislwdvopPa7QyH7IoxfJAOfm
rmz4XYsyexodXBubjXCNm6QrFxOlvjQ1QvhxZPRV6gaJT+o7nPNRpC32KV9/fa+skDWHZDhz0uMG
ECzaEfEuZCHpIlcR2aZnN9FWZO9fbi/hf72d0BLLfQVB9XjyTZ4vd3p0I6DKJdSIXtXzpfDhldIs
/E8WePnk2jU+EITq++87rAzzvN+D1sLNDJO+IIbhopGliWTEy/iDousoGiVK08ZgC5rvI8O02dke
fdo+56SDI89jcep5cHZCdFTqc5p2Vk9WNtE4bICuwSrPySVrouScqGvXKqiV+Taf35KglZeQNwFg
up4Ab5U6rmkgcFwn2Zk3J4Aj18lzUQvwxcOx/Yy9wbwQiCaeI97b/lYiCxXoy9QQctLwH+itQchG
Yrw8c7QtHWpafbhO6Ru1cc7uwgObAZziNocoI5kINPz6g5O+fZEQMh/4uw9XrijQqvDv81+v3B6c
zZPh3wun5BDfgdlJlufMEXbwPXksdDMPNHx3IPGgip3iSopDe3GDxIcLPTuYdZ3M1SWBIT2WVZpg
MSfWIKT/mR1Z1WbH7PebcUmb0ZTMBuWtLdd+f77BOcs9eJQia92PLXoFBXSckYhjKp+lAe4OdgX9
/97EjVkspi0chps8UW+lnS4kc3e93DfEcBLTo5Gz9aB4oHS/JG5LfBOqIDDiFkqIAqTIK2zBx9P8
gJbjFnBIKVwjtM5q/k4fuzKFNyqEz2AEP/auMBuFXdOWTx1bfiDlLo++jBKxmW+nBYY46MamID+h
Nszjni3Sa4HxDn+jUdoyI7O8cIJKUviMQI3xjypVXIC0R35E90xr+lNxYPzqb9KFMfXT4Yq7XiDH
ihDdOFhT8YQkoexxU2hs6tLETvUsmqsu07QZ0KqwHXENnsYUhUfsW/kgS99tzl2qKTFrMED5pXe/
wDkJ40NSXGaxJAeljCPdaCVgV9pNCov5Q8D1gjr82EMMfp//jEv6Ghtk60AD1PXmZN23drtyujAU
BIvC0BsGJpk9lfi/IagkWLszmePT+iuipfrdRsDG89I1uVxyKVKnD/d99MP+cn9Mv7lrylrOoMut
4CoHcF823sLkFZrN7MHVWw+HGXB5XOlIQthZqL+MReq9YSHKWXMjQsdeu4qMpTtakXWml6j0vp7d
E8ftNnGQBLPUtOYEMd9U8xdNvPL5rmpCgusYtmet2PFOIWZ+BF1xmYV8xQCnnO+5b/sQxJid+uS2
11TeforUl605s3zdR8RZIWHStfczyOy37TP6HFK9ejsxhtVgh22czb/BNvWlajRvSm0vHnTmQ2hQ
RCu3I9tfeYH+SgQotM9rve2PQUzlUbtqMQmjllpleG+BgImyr4NiECoY6dFODuihPWyaJEOC/x3W
ysP4hjp+ekrDYg8SDB2dJ7Nfxl5sDDX8jd2hCXm3sd/eG3VP4b+w0NMyvHfkUI3wH5B/26/ggzHw
SLPZw3aHGhiLeIdFAVkFHl7ClN0/+/KOYKI331OllPsy05oU4h+aXpp+1i3Zq8SX459azuc12Ro9
62lMu+6kAiiX4UyzC70UTeMQdZmtnAhKynse4qQmHhZ/rrPkPKuXJcBx61Qq8mBxEwvomGkVHksm
8IQirmN81c4qYhc4o3u0eqb6ZlBPWEbLkLSaf8xI00Zbd/bRCyI9cFcwN6V0cQwzW3BhsimeqUMS
ErpZuyYwNjWsiSguqA7eKtufzL5ibAmPUan3huJpzKn4zEn4qgblnpGtU4F5jF0yO4TCIY0pHceM
cljB9jCwuWcIpbSbYcAYtD/0R56RWeTn9w2qeLecMTiJzioLMXvaB7pP7t7Rql308BIfx8xkQK8d
qG8t+PT6AlPyp52hBMKo0mn5ItDuMAsImbQTGosX5JQNUXCjR62MTLzjU0QLcqB4dCTIKUnmw/4n
t+IvzWG1UTOeZewdvtV6JALwvGCS0aRw3HSYEZYG/zwRnM0K6dFrTM5nENid3v6iMwUD43X1PmXU
+g0dvjWnxcTMS+4hA4+M9jZR1onOw2fLMf9ecN+l34Q8rtZI0zjfR8jyYVqUvw2XxErVgtsqfJ57
Kh5uUI51sbzuVgLyop6L9I9DQWJxaBnq7SK0g3+/SjlkQJ+1ZWKTqtChaqhZ6TSKsqvb/uSkHTsm
IKC3XFDPI5dfiypK3rp/a1uR0Q8YiCd5LHo5z1gf8DwTG9f7hzYSSsWFH5MZRjXA9weVpmEf+Mjw
C2+Fz3Sx0lz7aPWxqBjEfRnBn9idRspa6LC4puMmve7GymT9CashOio0CgGsPRZIJccFoAPFieB0
TuZdE0DCSwTN25FXt18PJHYHRWxe/B1TiaFv7La41NVGP45VHhKtt26/gThhrZTca4sKpyUuHocG
N5AkZRotWaWW3Fenyw6WEhAcAKy4cKa+10uRgOGbohNsbI0hYBmSas5XAa7sb31aEIWEjUefUAwy
mefps4ddy6kqkjqp++vqBhaEKF8fzz70D6k+jT2NvtqGHtgllGb6OqpErfIvO2NVVIkWiYO5My7V
CgaZgByN+0S28Uxj4JrgTbh7w5eGV9QPUJ4iLl5OM4a+u0zJR8ydfHg6PLWBUxBSQQNxwpj3WLt5
scxMfIKeQDZz/J6hQKKzucBOhtY4E3wAIVo1s80QHplw4wP0R/KmoRbfHxmHBfavFXw5zvKCGwkJ
lRFTnUouoSqsWZGLkUAFxNyTfOE1fZb3Hf01H0R+KSRKNFEoP6+VyWLY5/0b4LAMyB1pRxBL3ScN
uCkwrzmW2UlCUgfJlr4cpVeWdUIZnGI7ASxZf6jbPHjodnU3vaxTOw7aNH64a3cw+X0qFlY+enef
0hb9dRZfzCkID6R1hMAd9JLsB4DE3ob0bIh4DdQ4CYzL97HdSfzyt2qthIK4cn0hAyAdBJuNae5a
aDerY6q+QHTBUIWGPeTSIdcHfM0vcqgQfxPrgejgkqL7z8FN7gfKBKwWYRbsJeLfosTeqDyu4rhz
5w3w1oC7IKxOtKmnwH/wUrEWvYqPQze/3M0bIhhVFnNtwPE8FRembzmD0ykzL1qT7Yk3NvtwyYbc
QlvBI0WP1wy/9SbOaZhyIQ8yqRg/cY5qiOvEFCQw8aMkbOptIsGLJH38n7REQc2pSIeuoXOsXaj9
I/UMdhMj1nZ9ZXOzn4vx17DePrQ80oKlcbkamEI2pLu/KpEQjs+cFT1jAmJ1vr70p0JyPUh3i3i8
bksXlcY2sSUt1AMGxlKBd0NjLEUOFEtbkKVbDhD1P3folSegT/FRqFpKg2GCTle6dEJtriNSwUGr
+avvPcBTceYFDcxa/WVD3O9cqdv99OCJKyWuq5O3nHJCzKzdKOJhNUjcm4LgBBxzfX5c3vfeoC9w
97wKvErgy7Ru7mTjaHZOg/LPSNnnIyQzbg0LVCL96DCCTSvFL02c01L/bYVdEnA8ObQADqmQGN3m
QuLp9Ct5JQYXAATEsNKNYMsujOumHWc9Fkj7YacF+2DzDiug+WnWPLfb1lRlYh6OnYwhfrH7J/XB
mwnCXHrf+ZEoXPwvyqHcwAf5Ru7bJxfZ42cZ0lfrNhfsfNYmgDVMq4MazeDhDGAOtj9j4MCAajBh
UEsghDV3jrfuIeupH3FtB69qbCyZBdJ6lyo2ycT96Hu9s5Aq6zmppLQSN7DmZP63enFW6VvnnJY5
cy2nSPvVcmfsf+yHCH9ldPC2SOfTftvoAXIhnG4HNxcuxa2OQ2fJ0ZHolkTWXZeFoHR9anR3x1Jq
FQP8vvXUjEVNH8XaErwv+hAYbo+LJVHXCLOSwuNry7QKrKBVG4aMWLBjMJkfu796tZ1SYGY1ZWbc
tPG3jMhf5xXOF1zoAgg2P/t8Gns5UhXYsL8m+zjvrQdOEjQpLZQChHLI2mJzTwfNKkC3l+C/nzRZ
8M+V1Zfr46ihqcaSc9hMVXKuE9518Cy2MR+kcHiqwm0zggavLkW3knYKieGGSr3ccCzN4BoHGPDM
vW9Cu7uTwff3R0Jt9Z82x9wM0rlOm9ZKVZ9a7gvf2hahme3DCnOUenmSMCKt0u6SkaXY17C6Witz
dhsDj2A6CByzpd37KDXmOhZAZ9X4xijch0zqlYaFRKyTr20z2Mh15NOZAJARHp6t4TM5hVyQ8UTr
DmCAyiGai+w0DrhnRLmkm1WonUiHRIpA3fkNfj/qcxYCbdR0UA3P9h+kUULeyAX5IRIVVjfi5RsS
1pySEGkr0WygKy957OH25v1aUW6FooT3oMzYFZwMECJX7BG5O1lW7kEXKD7tI+zzEBWsZZN0CcSg
d7jYR+rn+gt5WO4Ilgwgf3tDMJV108e9cbRZoCDBXIC+HIy8SpvWMwKlzC5mtmthFO2vVNWYNM72
p8Jde1mjmPurTiCcOCpdUq1WxijC7Jwkmi551XmwA89RBXn5K587BqCZJ1QYi8YOOVCjFuqIuHom
AeoIb3HZsAEj9my6cDLRvBUvj8/bWAOU6V28FmKrnuw81RwdeC7zxh9FVyjFJpMojdpNdOZh4BP4
89Vax3HzatIDB5QK/+L4RXHQFxqHi+HcjoXD+EJm4O7DD07UyNAtj295TPUhaAkI/r6j2yqPEqn2
PsIJQ+xCRZduxP+Kz5C3oOUOP+2I5fxVnPfxHcomlA34RGobS2reT0vgYd5yR9f5N5rxjyAf9bWB
rQvFlMZY3OR6nxEepkh0YNxB27+3QV3i73KSVOLiVaWBbdDK9aWq1LdTit9LFYFu9yyXB1VgYR1t
E+B2c6gt3PPY7j7vtzisBXmHZvWwbLhRA8us48JyQ7Q4GYHNUKfPRtGd/mEQyrSg8eePCkfkrUG/
zFTVcONffF7JPebhru1fDpwsERAPbk5Bd0f+x88OLXxTxvnEKqBU87n9jwctnct3SXwkXmDJ7hNE
ibvczgNletKDmOjHFZ849Qmyp6iaj39otbY9fZqMoa+4mn4seuXHd1TW37GHloGAPCydVEl1vLQy
okvVXUfU+nKlATPSELlz4Ou0FzfgxdKmuVwzWyRJ/9/WwQZ0TQtLv1snAaXJLyobJ3xQ2qXoUsbc
q3UHSGB/0+BWLJxyYQLTzvlxIK0qNHfGdmWyzjRNOoBDa5NoSFaDqXa0Sv7H/dJeHyfctCkLwi5F
JVTKhJIb6NlcSLi5B0Rtm5jSfWjWSufadIJlf43wvDq63h50S7oj98sbEg/K4CsXPpF7VvAr24Cz
4YvP+V/6T3KiGzJOemwsYj2PiiPEA7WNkjdBu3Xfxw/YsOn0VGnQ+yvtNcvtujsEQFkT78bIDMto
6wknQxVz26An4i7QcY8PRco04y/SEHXqPsdZ8hkv6Z1PqrU15CuId5QB5K5xl7ne9QMhE3+N0X4Y
nksFNHdZfkqNF1/n5XppS3aeEy7+5vUbkA2OTUBvRRqCsCBpq0NlkuvW8TuRdbGOoWZ25Mi3USI4
n6meuEk5rz4n4g2v3gsfZnTje4Jp0E95MQKdM4DWEkc97/oAbI+X1OT05A3iJIfQfM13NIfu29HW
A8cKfkTm1EMwPvYzaA4Ao/E3fGcHxFVyBC20+NhZlcSNwc0cmGf4VuXeuccqz4Dkuazt9jxDw6zp
MdArv70g8QNC21Oghbv7t7n5OCk4/cKTn8BqIi+WPgoo476Aestcdv7LAexHyJXS4QlHbt8X86w4
RQYMgUT51DsyssJgZXOvfG70MCBFdbyT023bm1CqhPZ07udDMAmlhyrTtA7OTO43fvcY527tn0/C
m8QEIqU+5lVzc0ZrjfdLBWcRLcGHmCvZMiyX8qXNou+T8Pk1X6n9Xgd2lAlFxw3QBEMMwJNysrjZ
sJ5M8sCOAL7p4c3y5WafStzNGty5nf6G21C0T8n0Mzd1t5sd6XL8GF8l6+KXEFqB212geG9wvM8F
zsOv/Hqrs6YWXBtbw7T0snqhf2K31J87lR297sT6w/JAndYtWz4/cflsPpKyRvKtK9B5eOClx6Iq
gIg4GRX1/kyM78Cyw2rWJDkBPGwPwkEWtBQebDoouLobEr2n1C/hXqtELq0GOqWc9A2uLUTU1Xbh
v5rtMYAS2LdHtB0jdGJTfOfBkFrhwrWKAtZ4HNHojB6LNTPY1LnCU0HFmq0odfwAJJvVayZTvXxr
+UY2O8AZ9LUnK3sFiOyssHyDxxhzTjIv0o8fdyfprF4wKyKiLBeIftJbD8elo9Q32e+D3ErvqPFM
v5d4ZCG+4eV3yOI0Qr4HSVTeBTSUnjK7EeBLo0TPGcSuuH3K/CwpPprrFs113jV0rwsDGYvzJa2W
A99EKnAG93vsS3P4b4FkkOLGf92xzrRiYXPGX5tVUzqmyjmdI7dLwmEnt4FE3BmY3FjEpFbhorKY
oIeS7np8so4zKixvda5PqyuQrRyucEHoTZRRpS3tr6W4qUks5F5Xc+pshi02unAdvM0uGTJXYOGJ
XY6MiBRofip0eZU9KYXZ4KDCwK0dGV1hSgafLix3OLePleucDCSt6WVhxuFiqb31A46Z0s0Gdl9A
C/JQN5gH6fJajSugreEMZ5Dh0V5KFhjPFcOll573iJY0m2q89+mI6TtFEl+lR+6aOXSqtyBO799V
bZ54bbRNLXy0Q2Wy1qsiSEfgSiRGGMk237vI7MOL9iM0hSyAy0qAK4PI20Mg6A20oLJESv71po0V
BR93sFcIi0htGCdEEz4O2RSTaNDxU0m4Pi+4oHsObDs6wqNm5JdJUzOUcRurwoRDKoRvDxcvdJxZ
CP1+FLPg8YuJLRzR3VWAwZeD1+F02wrZbOwu+Tz6U9AAgr4HL0oqbiMA91Th3GZiLESHKyCpD8cy
y8JfILZm6OtXQYc/tXnpNhFL7SRnzM7Apckzni+emCGtFDkoTQ1PMpw1ddnN8I8suEN5ExP0WQ1R
l1B+rLH23EcWQCzbKbWHR2YCM8o7VIsfqyUQ613gpR4lpXut+7MpdOfO3tvafBiX93RWSdsgY3nJ
cNOwE/e/0wpR4c7VYQyr9HCuI0nbrX95awFjnm34Wes1Bpn5RbDFGFfAZQv17pF+UtnLUn8pf/wI
lwPJv9OtoKJIj4C6oCLZFiTByS7BHt1MuHhdd+fZgZuC22XG+THrkdLfRgtRO0V7yxl3yeOT1753
iH0+P2Uze8+73Pq0IQ+rYOLOZJO2eACXKPhFtCATGKz66pNpiNv/k8cKNBDVMDfxnbgU4Sb1efwf
lwqyps+pYNQMXEVdQzaWZ5KpieQ7F9tKmHyCZAHbMXr1qtCncVL5n4noPKDlkdeFgfr2Da2gWrTR
5jqUHaf38AV3x7VCWqBCoraJPwqk6t/W+pjGcwlvqKBLhVZrK9SE2FSPpYVNqZyRtqY8Q2JjMoV+
S2FVejxmOuipZnGrwmdQrZ0OadRWQiRm7Um99R7hQQdPztJn4rgc3ZonZdkMZPc9bD0FlVBESYgQ
2c9HAQXkydMGnfDqSQdAENV+bsMJ2dtaB/Q/dznVNcWnlBe3X5T+MF/tvEcAiPnx7G9ICLhpThhF
RyqvyJ89VUQFKUG3IhBaofEdiAtF4hgD6uhH8GxwMoWBSbTwWmtgeLMRfZIVL18s2S6fTUS7ZMNo
p5kUc2iGfxKyT4Q7S7B6E0lAAA1wcZQ29PBOx46F6kFBQvyAK4CPmt6VuRBxKX7PGnyEekZNbzgz
In52qxiNkYDX7jzgKoupqmpHMqWDcjUQlN1VWwkKiaW5SN6eQGd1CJ5SMKvkmwG47qzuVhFvhaP0
WYWnpje0qskVaaSRlA1rixUF5ROzj+HO8XQHnfnaceeYGDQut00tdaBAsb3YC4GlhKTUSCiZGUq7
x8bAPXmg2Z2tbK5Iwfn02oPnX4hIQkUHUToDSWcQ+4pxv15XTwLd6pnoJGOcsOJi/QSq0K7EciEv
BhrJgz983dJ5maU3YnAtfyK0gyGzqU8nrf0Q9wc3pr2hWRKlaQvXz6PAXcKHah/rgdbdn5VBH0tZ
JhsP274S+HFdHCoDxb0ETxxDCsuCCUwDgu3BvCXAST3BCLJNn+E4Z+suPNRx1H62u2WmmytBjEBd
MriTfoId7YdZijkrvJng9bBBjiSGk4+i9LgmQ7Ynu69a9059msUfJgwK1tbQuKRPjmVynIiC9qyc
Qeo9myzepod2WOJA590U4FZauj0nVpaDrYoJJNnj0zyY1evGgrzWGF9anOZtVuB4HZons7PGyvBa
NBmTCYjT8b0hVYKWWvekr+5e66KerOqT8H8uxlPVMX5/Jiy8vR6OH4P48DSkk4/8usOk6K8rLY/C
4U+0rWutedlVBsNSUcjd9b+Jlgi0ecNfrIG3xWzruhdQ0riRzaUiysmppVLQGTzJ7y6e0LLJu5mg
aTJ+/0Ctn7xQ7Aq/Q4vuXmcNXwDxWUeuWT0fNGvk+Jk5XiHZNKzyWkgN4qHQ4jccxVpLPx55HKp8
wMS7EGUwmkMOkagpYI96r7Ep2bpEIVG6qpIMR241EaZ9StUbvHNVrnq1Dx3YEN1uQlwsGvDykiTB
ymv8hUbe1DFCoPOo1DC+7vAqTW162t6Bwb1oKwUrGa5/NXMJolGhjSKb+43EH+Xa1SIlBBvc3w03
WKcmVMaamo8QLJCFKJp9f75t/BA+vpJYuQo1SNGepOLiQ2iEG8CNPwQUSftHY6jroy14L+XE5who
ArERyGMs3ETcxbbADVffZrz85tUQagzxe/CcJO45JRuIj+XNIfNE1IaHRz+ZfR00fKG3ZKa9EcBC
2KVEmgWktZyaE68OPgS0TA6Tua3ctgKT7t14v97jgao/NhIsZwkbIB/eeVpMIkLo10fz9whKsN+i
cr38HLVOrJGVyKKSSF+EDCDkaMNPKvBOFHlfdUfzhEF4K4UA78aJXqWAQdHITvsjaRwF+g8zWpvU
o+rSisY8AIpWf3iZPz9Uu+n+mx/22E3EFi6ts6K9pCbdSlMIbbQ+vurSnNBwOF5twzdx9m7fHfr7
Xyqzo9lnZxG3bbsNQHOKMpZrkOgRWifr8Rd2Es78vnHWNTXOfXmguoaAaBgS2m4EDg3HDDoKfFug
Jd/sYHLn5nkRNPHxnAeqH80ep78VvZdaBZTp3F2+n/L18+J0pRySfj67dEj/ZA3wJFCUmMgThWy7
IRL98Nh6BdvY7jr75IaIbZbW5Zfc4hakcC6Rt7w1KWJgHkf/InoEFO1pz1OLDwNRgaQttqD5ZsC0
b/KM1SfxOW8hnFQRh7s6B3N7KPpEqWOzc33lh4RJmNx9SGc6QezlE6ENGQ9A4rn38pRs7HT8rVXy
DLfKLTRr9IluBqENR6O8X2886O9YTXDYphF2DzMj7l9o3o706Syy7NIzV4nHNdmUgPysSHVq1Yii
ox/PhtonwyQSoksg868o71a/djGgxl7XhNu1Zq5/TfejMBJmLh/k+8S9Cj7dzCthrlOM4zk3EcWS
gaJ87uvhFsX6Z2EgBS2p2WCPzjOkQ+MkJ3wxEouzgux3wI0XRulKoTkVulhIY1prTJmVSyJg0ANp
SCHvy43k2bpFRI47OSxNFOynvO/gmN+08lqRImycyaKfazYY/r+0Ea2/iCKYZPTJNP4MF2uic4FQ
uPk168J+CUEYzAR7YObshM0DRZKJPcoeURuNDqDRcL4Jd1blPos95WfZwG1Q0J5eOvZuJvh0m0oN
XN2uhbE4pdB9Sfn0MGoMGlHueBSXwqw7deLCQyo0kGJuzuH8qO51zzhYr6IZ/hXaGOVnOB3HVfTk
tcAu8U3AEHL+iYkeqIKFzNltAQfyEo+RuRbTST43QGMUwRAazm1lTQKz41e8+HgnYFjdruty7BWv
qU3heeeSALcY5IhEl5j3jSVCEB/0CgCgUnSxfo97iqzhFLAUgLX6JQwDn7tX8QHEWhEOLX3aPKe2
arl1iscGIYxBOBtIjtkPHIyawckwA8O2orS96VKXEsCnlbYLuBPYW4kqKKDcQo8Y12boFLlIUCUJ
NT+5rI8ErLRAU6Kvvcd6yH4tJkxAxJYTF+qtsDiRkhs3Hpjc3v8lCbi/KXI7IUmTEB9Xn+tJgV8T
oCPpSStrQtXSdd2S/ADLga/L5m0E/lEeYYY6kc6fDTbvnbItIrvba4o/4/50kkrE7tyBYxifJ9CW
PcRA9EuGA9IzPTLOXlL7+uYSTLOQ3qqHSC5VFWOe/yoOSZvsQXNuEmYQ6ZxpnYf3ok6XAkKWTWjq
wDhVdF8WdtgWYxKzpPLlRd/3+StP4oSpPWTZsfYuNf3pKU+cOwjJMP3oixWqRgKW4Hz2HfnGLMtI
qn+6Rt86lKxy985TODwc66jhdF0C4zbCbAg+gJPbOQYwqcs/2wBVXfPAgJkY9RyBH0NGjyPHQ5jf
h4L71dKh5boC022aImrBbJq590MCrOrOdp0Ohz40kuufWSPPHNsgpkRlNailfnftUhaE2qKYqO0p
3l8boLU841tdTJkJaq4212c/crk6SxmEa0bzycbsb5BrQqti3yLAlXiM0UI/2IudM9UwE9FEnY36
vRduOLsRuVaZNnNW8iPsSpe763OLyua3Kw+VJ7MQR1KyxbXFcZye4qbUojPj1ypWskCw1hDVmOPy
noCY7RbMrczBobOSKFpR3osaJ3BpRcGyC1jiu54xfUtdiFg20m4QYcb7y5bdQpdagbuaiHwL9j5E
9Z9N8wCnTgZeh4WV+IkKY+eWv/PhaiWOfguBi0XFn0CZC/Zx9tbgYnnLZ5lMSQGmjoaxTeND4vLH
Qr9X0HohjNqtVYKjIQOgPmZeb51WsgsiDJM1plqqMn81EctIOp0bxHGYnYrpBX+bMSBkLGTc8NBt
A1OgFYbSuRdIIXqM2GSA6Q5Wjrk5EI7dPFdi3CK6wmlQEXxT/mM+FZNZIFM8GOnmHyE5/Wz8Ajvy
+9eFGCafg4k3fFjcOljxshgdx990ftrQGG0gs4/zaZXnhVEX41sDC5xeeK+DsHmfS7fMWRngjQfQ
DVBAv9EtgPZWdEVQuraJEv7Lm5Ii9VHLj1tHKmslNCs1hvzrKfZVSh44dEJJmgqCAf6jDwXaMWxm
bjQyW+vtpmpzIMkmN8xKXkUN2ewmIMLsoHskSU8ALMS7vpiIYXimVKTfTrQjLXwTAwLvX4WLg+gz
890C2MLTAH9FAZxK+kjnMb6uCEn+cRFUN5q148w/JQwTXoIudPrYceYUW6QjaK0RNhB99Uga8NdX
37XGa6rQY8zzH6JHQPkE2ScFpFrZcWC1y7grkI4JJxY6nAuFWxENG4Q94ZO/YWlZT3TwdLishe6/
b128oOkwwsEeYWjhQa47dcsFWByky2+U8zAaUrB0lUdWdZZMCNoZJN4VOyHevHcBQEKF1U/KNTyB
2uOBWVpGP08Mykrveq2hd1UxO88Krq3ioDbGt/A1v1kAOKfDJtRyeA9JNn+c5B3RZ64ZqE49NefY
9GNfms51N/ey8IjsScYVy8hSUEzdpoApxvZNBg7Tr+oIShTINdrwN3c1O9OzL21emAGXW06BLCK6
YV6T63Oyaq08oJC5yTNj+tFNWa+L3Mtu8z2x/5PcL4ruD448wFxgXvF4C6yqTY08vU8f8GA2c2Ov
1ehbbkm2qzP0CqVoYyEEkT1/M0/rlwkmiMB0KDDgdlhsg3SnL897vyrrZiPm+As0cX2x9NZvLDma
t7IafXerEwLlZko8v17F0g8Pxat335XHXGhCca5NNSDR1Ry3cVW4PHCsiy2ESXMOvgmUQqkvtMJw
VBr+yPh95sXkwwyVfX+eAiukKTEEWtQVyEupArMYq35PtE1/+FgSQvg6UKyqx9kfC8b9WnGhk5aj
tZx4WeD1IGlEMZEROv5brXjtpgJNo0qo9KQ33KTRSkS/KDPSfGBqgpnJiX5JFriOmA3JJfRR0K7v
49IkN+ChlqxByreAyejiUhxZU2jGJsIEe0JErIt9tZtw115RKpFiod5+2EO/S/VMgilo3QblwRa7
Wu8O/QkxuwiDpORZGSWNqLQ8ymU9fy1rouF/Dq4JFA+dbBSpAszsNzU2tbD8hMA8uZdJwhxGju0y
E3bh/Uuqj3Zei2cNAb3wi/P8mq66hSPzt5jZGGlo3UnToguujHXuCB2k8LqrsELHx8LuGGU2GkFo
Sq4uTlzSAumHOdqlJoLTTYpjb4uOwGdrqngmvk2QfWPsItGDHAAAbcUhNjKyCYWqohY95CHehSH7
2oHpXfRoOgBTIGSzETNm9uPnWHYVqk8QmyszsH7C0BjmXUIFU1sDIyGA8Q4dMGWDtzB1dNG6bA3E
pJGGcLHp6EOPHqTHsiqA/ZPc1/s4FgWsV6irFWw0EQ1oNE62NUy4vL6aPt/A3W6TUUDlN4ZjF74n
XVu+1hpPLwCQLfTFXZoTkpwcIr4xPpm4ILA3gkEBD5g1TYMtm9zS/gEMo080taNvnEybvRVW1UVL
vE5WFDrROo7ZCZOVoXSwCM0i7tTuWqIM0lS84hUTrOhnaTFdF2Zk4KqNjbpRNxf7iTfJB/Csj42N
4N4aZXV3zEyQcq6vfrh3Qzi/JkJSbGNlCs88RsuRa8CwpvrMggiCI9ievcHhHRIPXZgPelnedXjp
+nBf5VhqtxCDQj6B8OPLqpEfg23Fpti9e06QCTuVM6TI2Z0Dxdbiv0/6GFEgRoZzCaTb+lD+Ne+p
T9VoMYTXx7KS0JXLLa/cjsg3OkNldSgC7irNMbAcpzW+oPeM3t/zbJCBNfI8LOs4rrYCUN3yyO5s
5XKHVRmYh3bqTu0TAAAT2ZGstWHuqJZes/HXTm+6hgJRGlpDpmpVAXmFC+XnVq84Zqx7K/XcYyaM
I1fkzv3HZq5R8x3rcE+HmjPYUiazqg/BaEpU676A/oDBNCfhoyvM697f7ubpbhlolSCI2ARQsFsj
tk7jpVIQRZGsR4tudxEMw2WgiDseOAVed+VP9a0MsohabumP4mOrbTKJlCC8aq94kNrc2TMW+tyy
xi+sSX+M/K+WzDBcPH5KpUQ97Z/8/c9tfKX9c3gJz8GgbyRYvby8PMg4jNt8hjrdVHSi8PGcgl0h
mcDXzderBq+pW5ns/9evBtO9wkFXnQ4iYLplA6iA9TWXvHjq3XHNCRl178+3wfgnhUapV4CvSk1Y
x6V6Jb6YpyVzIg4d3WiRF1RSutTwuKsQBJB0dAAnkJRqOeorK6mNiPdw9BzoGz+1ThL84Kxc3AyQ
zG8UtzONjHTBCIqG7jOatjdaiw6r8BNz+DdWGLVHdKcO/wYzBERmEpiJPuOLImpKSKgFOWaojHXt
zdD4Au+Fh01uwS36oZEbYi4LDi3sJTUEcKWQpRZ357UVykc5/oW6VRELh/SRzpe3eVB7qvfpa/Bm
+6amxtuJ/YWanpds7DAlQM3H0fkcgiqdWII+URPcEtO3IuA2aMfuIvUYag0mMlDSXGaM0D7LAMkK
yIrP7tVUvxnUtzpvhF2i5iSwgIHRVCmjzTgZnN7GcpoO62uwaNqMe6FNOP7vgIWQ8P2k2isQ4EOi
T7xxYsMsXMEGFfJkbApxEPPK8DNQ89jTUoX+2CT9QBfRDN5iG0j5NR6Z8pqMdGaYgmktsrT/bqT4
iC9vaFeBmZAXgv61Il/Kod6Ml4SA9Q39SfBbz+LPfBDQvvk2pD2Bz9MiqzBq8uSjEXDOC2y6gnB6
B7TRSZfqFbKekRdNQaP3BIVaqMP+BbdIWslQRGRfXTYTVrloHtx3bW6IsCQlsCQ8ZabVcfy075C8
PwbBC+w7F7DsbWkGz0Ejtu0J7W/JFWX+VNqP5abU2T2+NN0La6luenteafYl4X21BLN1vTbyrJS4
KALBWKGmquQdEsIT3K8K5p3hw1+OpJ8koK/0VkgikG2EhgZYILNJZxRGAgnAJmShil9oSrXCVDUh
9ww7zrkseiNtTUldUqENgxPZPXErP2L7grDN8DogkInJiqOSv/FsDiZXol1IiSJ+92mjyfZSEK00
6dH4ALPBoruvhUdAvwHQ6GvD9JIpvq38cJ4sYkzIg4yWE9YS7+9Akw6/V2uYluZQrsEuoJS31+5E
mX8Hkm3W7YQT5eh9tIvVJbVp8noHtJlHqiWNcL38Ty3Yzwqiy3YfidgHF43KANdrcse/IAyfr9eg
9I4mCGCe04mw/mX8Fobr4F1Nd64BveJFDuAUmY1olESaK18KHcrv70s0e8shnfAaYi5WKA3Jy6NU
14tt7MmE6sx1kgec6J2D0ThwrwLLm93HbgslMCaRMnyBYqHXP9m7qfycjE5thd8fNBzTSx9oOI58
tXXzN59BHSeF35dRU/B3J++5RHFPFGgUPTWW+4xx+IbH5srNQZ6ql9xjuDRq1zn9y89JjziB3JoK
yF0l/T4KWIJyReM4CNhWm/qRXtzXG9tt3iSvNoZg1JJBIT0vxE509Pvpd0+PKrrXTLQIEaT3O/OL
XQP3nV0C7+UOZ3lho9Q4M4qB7gFES4gOrHK4DfCqlQheA0nyKlwLDERxdd/rgArKHbs3iMEYQLpN
A6RiA2iejbfmf//fy9tAYOOF9axB4X/3zaGn5EYx9jMFsulmq0h5DIjV6kssKr594aS78D53ez4U
aICQ9TfjUS7fCBbu+svDrbQt52XC8/6DtT1p9INxcVT6s3FWm8la4f9eiz9qizWATNY/IC8DNhzI
LMULYbVHgUTZ2VAm9TcSPtDbj5HWzKZX2fhTWKuNG3Jp2Y9oHKg2Ww5fTRubHwO7Ruev8rT481ln
BSmLn981clRpFwt6Q/S6ATJqvteNCBl6ADN9CBXhazMUssrm/iKXEb3KaMFsN+1Om7nwV18WKPxW
rZA+xVfb/fj3h4elFEUWaugb9tHq6uqekw5lEbMwF8dxx7WkZvmZGXXvjFvEfwj2+GEX/nGb5+fL
K9/9qP6FoNeXRkKpluzxTmGw9MaWQNlfwBzj/0MVs8EwvmFfbzuC7WazLr/cjkNdlc/5mw9edOIy
aqqv0CUreqNftir9wDd7jX82qGstYX9W6ram2HLG4D5J2EaxNzdewHO6Pjze3B5XqFsRK2nraOHP
dY4aE/OMnvAuOQQL8DpFs6Lh5WtB6kbNb49kai2jH13oci4gCjc9jcUzBNNEg6AdBqpXnjtWZcar
/AZW8o74wnyfHMQWiDGi8w/q6iEeN5xvsg1meXCtZEQtQuPgCFJENrGBPC7IlpFF+esrmVqmeyzN
pEASDdBiI0IRkSUxG8+anE7zT1eOOOTGyiFJFy1NGLHLJMXsWzRKHR+ONuuYrX5pubhDDYonpL3E
dVR0eJOCBj3qocqKwIowMrY6v6ixQhlbKSW4yq1REG+fU1S80asOVj1vYLYjSpCeSZrwZM5lBTtG
A5joIqxEg47i9MzwnpOjRp/ewavoYj9Z5gcsnI/F5n2cLkHS/dnwdxJIdFKrH3KkD4vBsK1e58Fq
YF67bH780UhNj/2Wu+Jz/49xlqwC+zKOrQP4Pv0aQ3gs0AypY5s1bK1p8glubTnq2aLy57BqLIkq
rxoDf7j1BV/ZJAiPs5p0lc28ILMxrvmDFRDxU4q2HJRhVK5ZTUY5Ec6RLD4sCl7m9vwsfAGodKnh
34gWafA8DvUJqo5/mmUyqUB7zMNGHV39RmS+hL05dmtc8SQVCn0qp+m2Gkx2QhwtQ7t/q+O2xnyo
sCvs04fmU+yc73SePM93fAYD182JotZq3i/SVnqRczsuPn5lQbweTASRFNc/TDOqba9Ryzay2cX5
qZ9+NSzEJxy+1D8WwrMfBs3x3PvfM6PoEaThszkZgPVD9yRUBH7bjSoQLEJwVc6S+z54V715NL20
qjP2IaUpPO4leAUfajeg/tnp71sOMXJEbQd7TwYO8vfqGNFtS39TjcIsdxDySUePQqpzAnq7J9bA
NuJMMkXGsgUEzJGdIhDqBGd8BcWuocm0NccS9XK2NXBomF/YwQr01KWoKuWNwuxr2XO92EzHyo+n
md1XKh7t0KE9LFhFWFrWqv76wwgzDVlAKnJoncPCCA7AyEIyhyUB+TNk/SQfuDc46lMPot9X4Uc+
k7tx/K3vzCKzxXQuacjdJs5lfhSlfNSor6WqwVS+F77ZX+xGBTNFwn0CCyW4Qy+gvpn0zY1st2oA
sQQAIeolu/36xjLodKb2dn8RnzRZ6AqGVWVIDZ5hMUZFGwLMIwwDvLQK5sYaZTBCiIZNJeP8jMw8
rMENayQ0WtjpkeSmqP8VWuE+YbFWIbYw7NpNDWHitYTlmQn/E2qEDPViF5J7NLA/xVI8w/L8qCUI
oQYvPpXmg0cCZHi2Hh1Z2YXXhJ8rnj200HDM8ePz8o11vmRkDt6KP2xbJe07ywJZeGM+nf9D7heK
APq3c9rQzng6ZMRzvaPjkfMoTomtHxuBMNEy/7Ak149Eooef2CGbo2di/lNrxoO57hvnVEj15CVV
Occ+KGK6wJU9OMa7nN3uSQCBTsJi3vvaFYl8nQdnIBcmdIrTSWSs3XIlzR6M2tNvaSpm4fd4XfvL
oj88AV9b/Ht7nZiCXXaJL7NNd0TH+irD5bXmnylzsatPdJvFlQJ4cot/HQxYcDRMV825ulZi3FEX
OPm+yQ5bk1bmEsW2adohw39QhsX17x5bV7fLapt8EGsaTlwpH1QvUN4kzAKGOfSHO+5/spGmUMIm
1A9PpWCj3tbzNAp5Kuqk+GfREzld0oTcG6PJnLZlbBY1YaXSUZquHtqwyjSlBDANTiYW3QwoxhjZ
36bDAvYc3tY+UzAq9NDumXvicWAYgN5FWVJfNF4Op72nND5pk1Ca2/3i7M1niwlQUat2pj3TyprF
tf84CGUEQhfzLqVid4lJxLyT+MeIRy8f681AOnrmhkKxKDV84dRaovq20tyEOEltxvLyYgTIh6rY
jJIxhjTjXgJyl5qIiGSpbdwwB418aMd7vS0rZLFy8xJtIcmSxaabvhTXmBv84HIRdjtpbb64mIkG
EjybsRzadGQNbjbbNnPr30Wy98efNjAw9mvdBg9GGQE+upgfOE82kyLhISfV3XZqloq/Tjou9z62
fytRpYQ6vmFLXuJKaqfJf3XvzP2mLYhROK50rWRLrj+i3v4NePDOpJoE4y1YezVcDtx81EmtSxiO
OWBjKjEPYHMzvjCbyZ3wgIEa0P1aOE+wmQ0rItdnyqZ8wVesm1xa/6SM0zcfOi7w9T+ORYaroA9s
mVw+1h0oRBprZgeQNJsx4t0O9dQtfCInjHLc84EnISA8NIB3iUvmpEBRy3D99mgvr1FG0KWfNeDl
wA97G/JHYX69kKhCy3gTjFzehmtaYD1KW/NB7QR94JQ+8n4g5juTCMy8EK1iF1wT4jkLOxzEaLm6
Cfv0fOwbMKIKfYmYCvcKBXi24q5gNKNdLLPcRJHlOrCGF8VWt+Jvi9miiOMoE1+xVifRQopZgrEs
MCsCduN/jgkbcq+uj45cxx0Za2cHM3jsIF4uYK9JWjPfioVdShHoXhGyVZWgswA/6yv3/ELRK2iX
tf7ehJt3em0BfYHlO2AvFgmHAg9OXzgXQVrPQgG6KBum0JUaNll7n/kK2Tw+gRjOPjwktw+XLK6v
bF81+gXMXJNasl7Oku3f/u+CD4Ei8pJEdqUF8gAcov2lhLTv5sjaszTmC41uDjUJmObKsFMs/fAM
LEYcjFy+/Z0CEnvXp3Mbt2MbP9VgvFlsAjmdj22EDYSEGJ80CDaAPGRcSikl1O6tBkdR1jayq5XF
NxjzO10uvCTjK3OEK6eErSa5e3en3LQ2/0OLCG/OpUIouwibHDjRIbHMEF1+eNC/qD3QLP++CU9X
azzSCYWA8mYdsiw//WSvW9mmmXxHnUo9A+teN4OMIcFK1JltdAtHBY2paU/S60rmGp8z77knBOMd
JGpdbp4adcExWXWNYPQSRFe1+tSG8mami3zOaXiAEbQsr3tq0qC0QD6NxOV7fyje1vmMqGaF89iE
ZZ66rEVejCX0W68qICllsLBIuWiu72iGKKe9MMZ2C1NHNsosjl5i/22HdKnR461SW42ZAscV8AOG
JrRp22+zzynWaz5wgEOBp9+iRAkw0NDdO7VKpHC0PPvbahPctzKoPGe0aUStwK2s+AEGRZySaO/s
s/2Jvz9ty0ARIn5HzRK7H+1eWfFugYGTIVw1ChEvHGyBmgfK3WVGCLcpezIASUom/bDZxzrIeXcG
Flo2d2hko69lWhGWduvQU4UWdBXKpUowuKPmXwSkGHGfSfNj+mQRlP7sUNOByqoSE2zX9Tx2kTYn
0Y2OfBidQdO83HJokf70SEsi4pUF2jq/PURnH+6Ct3Dn30+dHgmIlOgMFhOdaI7BF8LlqLd1GMco
sa39ZoVdJySOS58qX+iF/MnZi+fD/Pb11d35iENgIXRNEYJRlka1GXDfkOdbBF+eKXR/34mYvwfr
moq08NtT5wIVMx+5Pb+PykvfzVPXMEdd4ULJTibjzd+bN5eNEk0UcbNJyKFl6SdNGxSQRpV+qmL7
sfXnjymGzWUcQyJDDziU1iwgIEsIDj5cuxLXOaA5L+FOMkdrneAtmgCYWbNwgyLOlaf9GbsqOhKP
fXD9Tr6kNmC3Vgr3iQQYQmBTc/AcAZH9ihyJH7YSMwhysfuqt0FiWdhd6UM8pcX/u4wHBJSDWHp/
bv3NuUSn2cpE4m55gztUhfir3ehV2PSqR84qSo5qKqruj1OjCGHa4wXLdTkXsHFuXUY/OAwnwg4c
eF0qBTSIEp2wxQuhXfSkcGZi/2A0Lb8fDfCuNC6ajTISOBc/9oMXOueJ7g74BbUddVAIUEP+MF0+
gTIiaDEbTav1IIJLpFEbIvDKPRQZc71ku17ZvX3MBeLcTTcg5Hf9IPJAJdWtjtrF0y14Bd+pB8Sd
gRzMUUn0HnmQZvt7oIIzcvFh4519oY55CzXcxDNKvF9PYRBL4C8c6m/npPWlpt6TGK/MwGPEB/qb
H8u8uK8fkMBHRs2ph9E77qFXH3IAU9k6b9+tAGRd7wQsbUWRVVbwRSjKnIPYw2V0Ag2Xo7KpSai9
M1svYuAvUqr/tIfvQe90SXG0iplkVXuqm3cJCd7V3qip3TGPHNyZWCe+DfJdYZy2jyRsfkTtuLxK
oVl065jlToVDXOWhedv3/A7s2s1xdEf7AC3cFy3E64dIKMlGf/uaYts0M5cijWfI5UWLnMe5r8KJ
TQPtX75vpY5vLmOpkm3k3AVXSksmRE6PKPoMSdOuZodsD9bRCaJtyAjnquVRTlZBY8AV1ZFZ1FjS
erlrpn8oHZ6ErTHHojBD4fFgJg1F959AdJgzD9hF5WYMGtcllKicbmXp+ZXn2l68I3xoKBLBi+Fe
zWfXbgN2D/oD6qU6WWRKjHg0xqvRDRaZZdNbmWaDGpNv9cgw1i94fi/ubZgWtaS/XG2K2fezsUyq
41RTcRh9XmxdyxGm+D36ZmfDqE18FDhzzU3lL6CdjcheNvtDcm+VLpxVM5P7ep0HmzTBF6SfiEop
uo5K5ack+Y/Gj5/Y7tgFk7UlkwaZsUKiAlP3fLSonqQUu6jXwYHwHweFxEUjoexPt59r6Wzmvm70
6mjbwk6ZMrtZKYezdvj/YO1xEGSgS9Eu4PUQsYlKu1aUFC/SMJoewGRvsh95KmTbw0mY0Y9Bviov
IN8azzlPR/r1fe77xSskwqqzFCHnalCXsJoefoAYiJCha2hGNTewYwG9ol0e9ZiAny1cVIHYla25
6ES5/j6DZqJG/pjYM9r+qtiorYe0c0+s6P+PykNG5+Z9qM775j1mcqVXTljyUzz7lOpsFCCtWTmQ
JFI7MOjYCg+qhBuRGsEhsVLA8eE3NPChqqfMW6yWf0Sbn7HQ/e4IjyxfTd4pHNwAor30yWtg54Cw
hYVxsDRpf3/r5Byj+ez1wR2Gf5FMPDAln8zpvZUJ7Jr9a7y5DV0py5lMw8c4AzpqG4YJVu1K173C
KNoS558/69eR5amLDfGRXzFaGqf/AfKJQJkKOM04vi5IuhexjBYOK9l32VrsoBatPXAPPEbewAgH
jAEy9wz+PvEk7BLvxqZXyuyq70x+CJvd5FuhieA37oVYD2HFM746HRrpg0CIoxK6S/X05fYwvc0c
h71jjh7NWisIEm7TcvP96kS/fep7n/oTTBfhHB4NLOKLq1kC9ZY9rduh8tMROxPcCcY6d0fRXBC+
8xu2+LpJk5632eyOumC5rNzy8RdwwpzQOdk44FyQWR/Dk++pGNeyyDzGw2wpHompTwneieUhsnrv
PcjhUDQe7wERXozulxPgeMtg476JelEDdadyLUAGbNSUI4pv+aC+tTG491BMjdcLm159fcR7LVbq
qR0+ywm7l7NfWnGm+MBEJNVfoe7pImNTg033olOIOKTw8qRMmIEQQF2sU12lZGwM2b7yKLuM9nRe
tRw4YBq1zJbgpFPLcZWPJbnaOSUmVTip8wLivlbz4CYyru6qa2wpH+stxeyb6phe6VlASYzNpWk5
I9jUPO8gp8ecFgJ+Qv4oX+FRLniKXAxLx66KOdM9K8+n6pnNhtLQPWEdQMGuTUGiohsMe/4g8cJG
yE8w0Le/Wl+yh5ulOAKtsbz1HNzO7uqbcwoPvuOpPHCvchAUhsjKdHAgdlkGIJLeYy5LHGYY1NJw
zst5lX75V43OKqcjV2zATJXE58EjTie7lJOVK2G/LzNzDF0jOaoXauCcnO2Xd9vvGmChWM72m6P4
yQRD87CLJkzd4bqUKB/dMzPHsKexdWLsJITjT9nCTJEms14nrVChHzipQt4JEKWTTrx7IvSpXZSv
bZZRHmwdxuSQlKsS/OyIGyghHW7KfKcs6AhVWZHeWvYHkFBgYFGjtdVvUmZKxO62QyQ3+G9NnuVc
DtQgxMegBV/knivme9Uc0glsUTwwUWRHf8iXcpdzB/RrQMuzJ3wKaMPpIrCfCUBTiG0DAv0jJWHk
W30oaoyPUXGzgXru5DwdSVl/v3NVztR1zBAxDVh/oAps2WVe3YW3FUyANk94O31D9UsDHsSKLQ1F
ONFG9PA/A6npHYTePqeXP0q2kSgj86HbkWaNNNEBl4HuvtwCsyGKajSM1zW8m1g6O9fvzuS3IoTx
JpPlBacv56zzr3CzEzVEx2pl8w6FSlwnlUoqaion7tAb+B7uyYifKUylXmtHIrPwVgohxqNcTsTR
4fDQUdT5JLY1QYMX2v0aUvGPj20dir3vcRe6ZNUd1tW+j+1Yg7sfkQlFWyrsgJU3fz4tDDTUMhLR
kOYmsl8Hj32zZFH4TIWdBd/l+7pB2xh7QWhtrbOyZKFiSbaO3dmaksUpDcw8ZNa2/fRbXIKdujhc
CY0WYcl46XO4UJta1etVVMeJ6vK4k/T8GxVE+57AoyKOrMSEuAGmiRAYedR1IDNuXhzxTnjSdWRa
CFbkFNxL1Gqk9l2FocARKIk9D8ztKmfHZ0dPB36pnGZRn25hKMvHdJby1MsNOpKzc+6YXjSHOrxJ
+v8y8Rp6qgp0YWyeDuv1NPe1MeJx6iwWWg+Py+3kFNYMnSiC7EO42lVLnmD0IAsAzPNoRJ/ESMfB
uRiHITMWkEo+R/IU46klqFkOQnWXuyx14LU+fAH0d/bcBLRDjTqiZgTOq4MXgqGqPlJ6QKUwmmBI
bLy6ifu1BdK/6UzE4jxXncjIeiVMePqE0YDGoUS6vaO0WrG3z9bK+hoOnijN1Zx96cWl5wTPerf9
9GqWxQuBf9s1vTJ+2yOIT2tB44jR8zBYRjBrjQWulNG4Ec0g/CgfUMxGOaAvpwr0itlipY7q2SRM
v77jwk5HN/Mp2wH8MvEX4hD0fJDI5/MYICpJGYV+VrQotLVLz5K2qRCoLcucchl2F+A5uZYKmy25
2lAlVW2+zB6NTYo0zsfQWL9VaMRxdvyVJBZRQXMi+OSGPQVeNO0ozot52OyVfgnijlxgIaPIIJGJ
HqoZ+kdtrlodS73bqPtPL4lUTXK+tr471yok2CbufPRUwEY7M8jkPLxGFFXjl/gbHidI/8YKaulJ
w6kd9w8QEx6x/Xe29Kt4A6zRGY/vk+M5R5wDSRBRBUkrvPLEYqjW6+DsjlLNWFBJtgLGokzM/ByL
kkGpq+xiwq64DoaGDfJTr58wPOS3matO2hHWTvAfjA4hYuYDM7YtnaWt146KJMGuT90Izl9nEXqw
Hyuw+q7kH+6uv53LirgqiwVornUj6judFAxlc3DEwJEfMXoAE1QCBPZ0eMbVd0uG6moXLVqsk8CF
WRo8pZCp+kbFFVt+6zas1CAo+Q7FROBIePWFUeRZeHSz7ZgO4mdSXRpsjn+q7raDWpm50Pa5CgQj
E1kqZQ7s/zEhXv8khrdvqeEUY2qT+abFq/LaR+8uYH1GDWUU4moJUtQEgNwxnqjZw2z9y2+jWOh0
RSLQa2bd3NIdOYqe+LNdZD0bOvwoUJOXKXxsQOruDHHVJN7SN1M0/1Xs/w+gBxudUyim0MLt9epp
tlAdni1hS23Y94jkNmjKZ1w1fxw9u6yBt6do3NZLD/3b3opnd/dQVg9E8Ui9IerslSWPNEIlkCGa
YPQKIeteqxqkp6eFcvMHG+pqTyEX6r0CYSekwFtzCHXySjkYnr+SXJi35TyAU77AiSbsO57JxTPb
NqLqB1DKPpEPQB7l/cvC2ECcwnO35zGoHzbFDI7agEAnehBgh5q/iixt3H3BW13a8xBfRdZz8zuf
pTyKBVx+M5l9XeoCmToIz0MFwOuoaTW+ZACxbfD59MplKkhkEE923qeWLeuTN2j+vxa1TjFRQdKM
zDzW40awQPRovn+O7lh3fLQnBFDTWizJVHbeXfl9IHIeG1YllmSqJsb0WM7flDGAfZp/2RuBJauh
NHRvdIutpuhbH0Fphk3G4CWZWzMPb97KOBOiWiDtj460FfZKyggRsErZG5ruH7+9ATMuzP/BZJhG
SHt7EPJQnBhWuM7J3rJNUR7kqCZlyYU53I20Zbv7kgc74bFZxrq7WDhGZb5wokMgrLpA+oOHmCR7
ifqm/4Plf+8Rcne+DkYWLEHOsTGj63NkHclPXWxT76lBDYcIDMHIYf+8AnEsDgdAD0akfiYx5nxs
GS4LzbIy7I565xCDdBvNfVVTJgidvuN4tdyGjBPa1Xxc3qwgDeT63oojvSulg7hioX8AeYQmX+p7
qjOFjW2vJhgakYJAXI2cjxql4J+xdBimdSlm2g06oEY7qUtNx002vT5rTaG+Gqh463Fe9ei9jbvV
Lac704Mrs4TAo8Az+ZUKuvKhRRV+ZOp513gmoFz3th5FqA+nQRs0n0LI7OivCY1oMSvob8+vdrMd
7CUElOp43sGswD/ajYf3ol8zsmE2lx47VFCOSbrEhGrQugsH5R9Z2HSrJCHsaqPrnd01dsUuxwsl
/CKSvSap4HjTJEfFtq4tblAXR5P1BtFFozBN5ON16qmR5e8GMEwz3vt2rfHofGrFCIs5fKJviOeX
adZaWbW2J1Nj1uYY8lHqgwjfOQH3CZKPxD3+A6DKuBhhoViqisj8/R7EjxzVwlPpJlSXSab5pUNH
Px4gjAdTnAxFLj2fMVo0IXAEOtJ2xVgnKYqf0IZz5FTZ8/57YjQaCD8qm2pwKq5MRscz+Ll+jmqY
SpgDPuv4MXaGw1T88CsSJhf90retzMIwu+u2I47pS8ATeoo61EGmpm+yzXjE3bhOoKT3TjzVuGxO
VUCbqf8O42h+c/yjCQhrqX5qPkY9HchTNa3DSYBe81z+SebUopfZm0y9Tcy3OBXXxj7HZ8I4G7+j
8RnF+UsSMhGCHX6k+sv1xiUGOTvQi+oWuc50m3APBvMbNX+VQgIFtKHxJYwZPunaq8Lq05gd6y6B
UppF3EgVQdCKA2YpFaC5Nxsu5R4o9B9H7RV0LrnZDRiiGlNYaO7WHKaKXQ+ydmxOb5nIrAsAtsFZ
7kmKyemhuJoaZO1hb4M6S7ZDwPwVKFwvv1nkhvHN9btm1x2mrZPYKjGdLXdPl5VN/pIbH79Odq5t
c+UjxM1/P6Y4w1uaSo1dT9OH7xm0Ko5SjOKP7JASe97j7TkAaHxdFWv0pfifRzUuNGcQgqR9uInW
U7+YyzoKqaqE9N34O90xw4LzQsFgimAIBcTXOXIMAGbfy7Jq3UrfNw5OIRpp8N5eOthss2qWSZ4Z
kTgnXx41Ww8tJc54MbNeJcu5Ob6u7JIQLyj603vLogzSe9em/SbZcomstxe+Ey1BUuCVHLjuVhFl
dKJKgVbWQPcK7SbyE1tbyipKuRIY34Zp+IjSKpSxGxQ4yXEZ9IahGY99LDoV7yTwkoutCsFYAo9T
GcJmTOew8mTRMiKAaR22WVqpyZMzsmozgVekHCszJ3hzzTbyRCvNGMrRD7xzkdwzZGQh/azfTtb/
XIoLvDSVbVij9nOcb0DmmquSIirwWR3qK6ODMPIfrK8gPQCKyzqKCV0lEFLyJBOXhbO8TbbV1fpX
oE0SO7OEhdp0v6T0NRbJ30KeYjriml+uhgbhAw4zGLG8hOXZPALnlgnlyAdUjJ0D1nIkAc+o1yCE
BILDebPvZ+pw+HdUsvNXGUspHhqf7u8Pq0RcehKYfJDD3C5QOLep1CDSbPw3CJyjmpcgHiAcAGGf
jC/aKNhgF8OQtGTKZqHaSuJduVhOxql4nbEHZxOD5AsguFiT0eKz44/+hJu/1PTRzCGFZHtxEK/O
Y6LGbrr7UVo80GbLJ8JFFV5Co6PR15PcsAoMdD5/ymLoIyE+fnM4674KE9RQImtpLX6z9X6BqW9y
OH0MAlyj0xOei3VodGaIBUVASOfHof5WzST/ofg84NYOtLhZ/2NE3TDBkx5+O7RisddUFar+NnIv
RoHIbj+dGxnlLY34SJlljlHvfzOUGUif1wJ4RDlUyTyaMMSeakN/nrX2DntKCgoMYUqWCM/c8r4C
8iht4MN04HgfY/ugsItntankZbRjTQjBvwRgBFxhxH+pRv2SFfEberzY81v7PS9LjabIhQnGd4ew
a5URQvPPL7p5r/6VJCgfiprdDhxjf3ucae+KyYHxI4M0owKL73E4pxw705EbmqLeQK0CCfY4jH9P
N01bXNxl8/7HPP1AIyqq9Btwz+lDCaTj5ufh6TaxS9LXuiKoYncarckoRCnAqNl4/iAhjUbaT04/
WR/jhWKvbGt7fXsrROgWMZq99FrKWyPQUtdhW3q84LibUnGgqhwprN+ysvrE4CeekyAc7tchBqZx
I9eUcSO4DIvLdrvSW0ttJcyXOCk8yr/eyE71kw3uIXkwePXxsf5ntIEGdAMOVULpDkn04CAteDTQ
NOf7FFfC9kXQ0sDIFTZ73XHJOmmNvDPquoFQJ6pBkrXpJPM9S7UMzvH4AxZ7InJWZoj2D83fxIEx
1eJiy4qB0ldGi3y44dW5tfU+GiIZu+1bEtP+43/acXigtNxMxAJWZuylaP4RZKizKuEdG9BJ4aLx
xneSoHDShQWEcJTIdLgrkGw0HoJkk12AAkJsktKIF9AS9uYMek3uT8Q7XGMkNLU7x75rprKJwocw
Z1viYq2Gw1799iBaoGpL76nrbvn7M664zV14hlz4hrUS9SrFUpwwgfaT5gUoe54BJTU61obKNMTy
NQ1Mh7My/qQmdY9vHoTIprgJqLYhMbrAX+vaasxWS3fsDltYsi9oON/X9jXY2ZNzXFBUpXBYxWvx
TlYr6ur8a1pabXYHOVM4sqGpz/jAIn/Pz1WhXn/IEUwgcRQFOEDw/4Eh7PWlXVMNfW5AqKYWxGU8
xg9siahXcUy+YkahkYr7tpi38sRTQn7vPntrR7AJZVEm3rVFlvs7Di/kvDv5RuwUeqna5ZPyJg+N
QavCeBym9AC7Z80aZJ0YGuz2ymcQ45WNHPEBDorQwTCZBff7DisekXW8pGmP6nMWaWH2kadChdhk
mNXVWIPV1YF6CYMZPGATJMJfilkKreYUjUskFGVzhTU2V+L5uThx0kzPCqPRbBUvkziM/MNrpYsg
HiMq8x48enr0sXu1J3vgrWdSPWzj56TXMnnQjEkfZ7sj986YFjwvCm0VU2BeXhA4Tap5XsMN3m/i
8BWvOnwf/cd9zK81CnZRoZIUB3vFvT7ORXnUt5A2KsnytNDsuQSppCj8ozqBdnbsJakj4cZ8jEeR
RQFzdnACCwn7tpe8Y2UUhTyQQrGl1Vrf8UL/em2s43yLe+UqmDRTPka9eMFb8/KwEN2Und4YkQsJ
zZM8eDd+eXTkxTBT3LIBkaInC0GqrUTl8X0s7D36b7I1Tuh5khZK3w+lF8f5tC0Tt2kOMuBU40VW
cgbqBoL1/W0yd8onffs5r+Lf79qerJErBJXMRyUXQoGn6zQfvSSvmUr4/vvMpfxXzqVpRoM1LSrK
ICjkCsoNXV9pi5bZHLG7mmxrxwG8ZySPcM63MuLcfaPZ+5uqdvha5iXWcrh6lCfP/GB4TLWh0R4h
U1w5XGCXSXgFLfOWLXJdOmrv93oYBjQpdbQRPVPqZaMJli8kDEMKSapZCn8c5x9nJqHQ2RH2l4jq
Z7OL70ueOmi/1XnZ3rrIzx2CQSclvpijZogO2ZG85SHKE8R78cWIMLvwym517p+UeL2vouTC6l1E
/y+pZC+SjIIbc89gLkkNGxpajWqnRGGiEOoklmNnfMk8ziVT1wP3MbX4FzALaINMPYLIbDBOk2v4
mk1RauaZ716IY2C22ts1Ej0e0xuy1eXLBYFVp1whgjCodxm4o70yb36SgzXYu4lPAfyc9MkWmfoQ
9flUY54LMA/wkgcGs//JBjg1mmKKe5dDEaG/F+GrW0IMng9cDd0xsJLjbSPlb7Zole+O5CZ0HqHY
nDlBTmGIsyqhyZL/86rLEVG1X/Pj2eHq62iZ6ni5Xl0OrmoY6i8Qwmjt9GaV2PfSMm3sPjLpy7LG
B7V/xnBecBqsYNmorfC9kl5PGgaJuvVHrjShyjJmv6icP4dARgfQFqvTWUX0FuiHfGx1zAcOtGU8
eE2Hhmn7xvWRTxiYykhHkJRFwsu3qrswyOg3lnq4q1koskPGWn9isb7FgIckBozpitVlb0/gWcGV
Kc+t55FtzzGD8b6tOQ8uvwi/YNmy9LcFNfjc0JPZPjlYo1zsWvUk9nC9I3fFAW3rDZBTjFqnSjPk
Nb6V+SN8LBfXBC6XGzNslnsjmKrncBvFBdf8duVynrmjGC5Hql4H2iWSnIxw5S9s7vGKaEePB8NC
GaSkXc7YwDzz+lx2gY1E3wKweC7KKqbQ5l1pMLe1Dt4e3KsYFFTjJi91OnVrDc70T3FVIpA4LzZE
BAEOosOiOOC/BjrlHviJkTZSW/u6oyWvkt9anW1YtTN2NLSyooLOTTveHp2d1tJf2a4Y9gPwL/nC
9cFhB4mxQJw5MfNAQmtKRJo1A6tnAutFYawDLm3y3CgVPSfqEZagYy7L6laog0YyclqbFXd6huFL
xQUaQZsujflr8Zqmygwr+lpHHc5yj0SOwtWVb/61qs6VH+RsNdI7apOatOiiSeEwPTCmEJlXmcxt
20eGZuE9baHt23Y9/2OrSUWsZqycC7nkMAkPLWygMp9l6BXudVpKm9P1PI2YrIm4zu+lpwa0tEls
6MworVw7eMDq5O0NsTRdcjWEpI/t+rOAIs1kFac/VjlDuwuJH9Hj3BV5iwCYrVQJZrUbBmcWoYMY
/b9GDdhwKcEGr5oxjKS1jllj5AGQj40PRyoURWRHN+QnC7jRdVw3PU3sMfcY85iY/evGucgDyemF
A/M3hdUoopMfD4HEM7lo1qkmDktoUxj0b+RndGes2ut5sqrYwsNC8zsOL+ZiORroriydlSFSCFDN
NaxX9UPA20WnqbsUYXbwDPdky35KqxoZWGZ2A8NIJBAl1o9e+K7KeYL3MyU2gvaA6ISqis9NxsaD
xqdaOteZ3N7yV0HTdByPGtTrvhPqgFTIf8V1Zph+jTVXqYsA2udWshMljSHJtZC8qNEdFKe1rmyc
oQzHn/WnZ8PZe4f7uSTeH7/bh0n5O9GARA1yNscR/2x0MmoGMdjLJ/0wwk2S0av5HJn1N89kORK1
SmiYHWKxA/evRYU1YUmaMOvut+chs9IsrwWXkjbLJ5vDw0iQA/94+l/EGCOP2L8EASOXvBHQ7aQT
y7F/PMdxntqrEg9UcJzmkqYpT62xhM1OhDN4E19cv1KK39cZnBr31qezrzUvLs8IlFO4VCVpv3yH
9pQh+D22sqXnfKFDg/8UH6kWz/AIr1Mj0VAJLr5PzkW6QKM5JQ0wHHrpUakL5zhLp99slulzkwUc
rppeoGjPYFew0jdqP+QAmrdm5aq5d4CbxghJ1AofBMdSBy05U1hyg8LoN3gWEM8s8qAE8wooqaf2
iRiu4IwKrKVhiyEogi8ZDiuMzEbBkVNcS05uOWG0e5SEJ0ZkdHSgcLa5c+q2cAYTmEE7xG8Iu2Ir
iXsEEgs4JSQGADOPO8yIP/6JwIq2z/wgIVp2gpdeOr0aXZHOi2/BMbcsXmmlSX4Q1kRSzx6eMQmn
bRRK2YVmwNNGObIDul+ftGbL4NlnTkkcAp5PBbp9U9Y3NDf3MITGzb/yDxQhH57n5e/HB5gT2b6M
dLsVRKTHkoNDMZXWLzDJrETt34wpCHtKtuIeJ/hTAxxxR08ggbmtV86ovyWGMFtr9V9kipUu8qjT
CyGMCrCR9bmC2loy/JxwyZHiWp4wwEV4EWsZODaC7SvzahAeEzcqIvmkqjQ/7krPx+qLfPzpx3kT
Api7OFufGQv98S36ifwKm9L/saTcKjAPXYbpzrVnf+pHU5ufD6SBWH6DikgOd1utKUZN8Kg58n4k
CLtBWW+nolSVeVWRxznmLxvGwjCFm1bRTWxjFCmnWHAWSVKMN1g3ICsamTsmD/rf+I8M4mW53+iQ
UUaCy/TqqVL90KFfE2YL+0uICn97Wn26dfU+Z5+arLODhJvz0bEmGxmTWcZT/m7gx3p1vz4XRIT0
VnRK3u8tBqupk7+p2NQ8Klaiii5YgKwAW8nWQlH60oW1pS4X1q5I/UKcZk7pk6gGYrktEbO7T6qF
hGwI8NhTt2GZPZYHc62WXFwIxIVVhebYSmUk7/fs2E8vDdsJqVxb3aEMotkJFjU81cMzYRUPGEz9
A0KCX3F9tTzPeuvwznTgIWq5ICIIEpTzuGiQiMoTJkUmLjcxakHKoHFwa/EXcu/+Bc4ijXk80k4C
BNd+JQkl+ZBfNOXQDZybOyu825moP+vUqiKTJ8zZaJVvVRXBBEiRC255Qlemj2M0PJy59HN5WH/H
oztFpYt3FGjWrVY22VX4xL7vvLtPBl3U4fOqUQK8BldFWzecKijUP8OCVjqf/ID4WIcPyGQENCfQ
8plSIjtTXbR6pdUzM5s+TgMAAEuiYjbQltHd+uy/uWbMSzYXQQMZI82ss08jpm5fRYoCC5sRQS3o
7GcvyG4+kL5RyglyNGJXUcxbRPD84GVVirv0AvaEB4rqiHUYl9/WUYo7odkx3G7HqtKuiW2pXDNm
4DGuES8lbsH/dkk3W+KwcHxfF4dRi4Xj13DLOsKzVze+m9YTiU6d9rB+f49v9lLmy45kY61PoAI3
wlfSPYbiOB3vCvyc3kDHNO6Ipzl9dPexlgaRwS89Addbbyo1kQe9Qis+ISM3AEu3tuRnuhxffQYq
5KCcx4INq0ZTNfyIDXzp6ATdNxuas1J+sGnR3CRPxxtMc5zYfdtG+8mpJvFJM6OdtidgG7WvZCNj
GRudgl6HKC5AisL7YPz64/8WnmTq0d2R+ZGyGufF+hmzgw/tltfoeqABiuhvAXtMD+oYB3o8Yleq
1rFU5fff8ss7Dtjkljrfu8SGfcPIAoxiYRQWyZetR3ypHUFsAANI+4+zVonxzeubngH+LbfOHT5o
XFCcb8ti0wNxwhJutW67dsztwNxp1hx+3pFr6l30vDXGvYUqCpkxmq3O35U/5lyoNE9RKhuTKLG1
5gQM95VLApGgb9aRXaME4FrPdhPBMBBWtXksgPu8H3AhoSJIFQMGYQxpSknvsEXDAneCvxYZXe7V
05RJvinqw1nhHO5NH/PMTXdCnzB2w8aSwG0ExATc8d6EVHcvSX+n36PtSbCmvkObJqo7Vmg7Ds/O
u79EblZ/ZJkwwgNEWMnqnARKG3fb6D89xfXZOQXr58XTOOzyHvQh8WuW5JOxewURtkM+CzvBCe3p
Aq6OLPO2fYpDWT4k5QoTy7HXluuIXFSNS+jb0nizhef53uqxnT8G56itz0zJmk73MWjUfD8YLzjk
vUoyGEGHODLkQ3SGZiErd3QoIIaTZbLeN5w7Xe5T3MpZLLmReVAUrk92UsDPDcilcN8YXPG1dKvy
/C5x9kDYyCqLzIti07sxjY/n6QtDu87m8HDj4yRu1YAuEI9v0Y8dWOZiO/idtK+GPmVDbBsK8pqA
+B+7yL5SYxK1BP8XEszya08ifJmVsclOkzL+271/tvoK7QvuxvcbwDJDfYhOg1R4RbT3yaxNJmX/
WA06BDvaEbdh2965V6+bINPgFWJ0tBkC7YCdwTMhFT7uuds7PQJPo+IK9WV+clzwvkDzp5TaNxw4
YE3Ys3OL65ddnL1uH053yYCOtw1xXOxgLT3GMSbKpVK43b9ubLE9eVS9zb1Qe+/W+El1oXiK0S06
CvrIlJOhMOdXRtisp1y7aBPNbkjYR8b4KGydMuiM/UEYE6tMMSlCaY9xM+5VGZD7plPyjuE+1I65
42/MuNqgo4aCCScSJq+4YZi8Czv1ETV+2or6PhroQLeSwysViHwqaK7dEamourB7o+fXm7qv0AiL
67sRDunYw1m1fH4NrDV6ju7vgTQiEskzLVGIdA+7QfmkKeO3vPj4YfTuNGaYKH9ybS+kwG5GReqh
FAGgFkEIHbL2jyrKy1Bg3ZSr4/b9EPtVmrEot/xCws3WMlnvjzWFpRrFIz5u0xBUYlbcofbvdWZh
DCT9wfBgHNPSVnXY/lPfapD1yv1NOyfll6RTFbt9DiIF79v7PTiwhs9Q4f0nsGqOgWThJ3AG1YGm
khx/X2VoI3aBRnGZYScxTup3cr/bfcORnA0h75jenKCqSCH/CXl1XDZWZpMCeYEa+2n+e4bxWUH+
nNDV7FxhIAMxpQtcYXN9VUSw7/TGsZPYSqqujwigVpVj0iJ+hjp4NS25Hivn8yBJJhNtKFHzuvWN
U13KQe7+TTrhaiAhjDnO4OHbL0o8hSWDo8U00VYaGHMeTE7cn5oaIezZqKZUr/sOLnblzqrb+rRg
P8h6GxbaO4yvOXO/e/p98opV6Nivh5Sdenhbo1Ct9hUihTY1gfNGX+yMD+jf/dA8ZYWMr2r6zVHN
7NhQAYWrZkaEh+1Qs7ARiMAxsTfO+wlagg7Mc3wY6ZANN/NXnRqk7GyXog3nTRytvpF/ILGR9PSC
reA0djFd6CpKXQ5Wj65Oy8rKED6BSaeRplfscQsogC5n282W8drYrttE+e7Bqg9MekovMrxRgGYD
VHphFVJinJgJ+GCVK1wMsuprBYBgIY5+GgfFGniwfvOT5nm0wTNR+1rejJNH/RPS/JA5kv3rWviV
loBihy8bYAc8GvKNicfMLQ4cXS2D4WoEmn5rmC1sMJkn2Tchp1ldWsNJi90kgJnGlz6ZV7nTNUMt
abWG5uqmH2lF2/zYso9k8Zt9JQmbvgZ70puoXH18UN1hNgmFdinr4fEEob/LLlsnQPV+ymziOnC5
cnmUTR42D0A4H3nGPNGEyX5XqUEzgCF0DkcO8dApfLHUHv1vE8bXYsPmlCBhSUbxcWhZiBW87pNj
k0vR9QRx0slT4tlG3UszsrXiEnz2VBSlOAblojHWaPq35Mnz+OYfgICVVbUfs5rnpPX4FjQnX3u6
zzD+68Fr44uR6cfW3QuYXHDlUFErzTimwWj5joYmylL1j5UpaByBOC4LSemwYak5fRT5+b7+Y2Qz
qR4RF3GhN93gtu3qJgd2nQIYQ9eatJBoOgiAF4V8Yx9A4L5RsYuBVlOH2J8CVNbRoRu5J6AB2ZHw
YaAHIL3UwDGp8c1jNRlB3oAZG2uPoRU2LfLwFWyDcftXvbQEYcCyV5VNJzRD26TdsZUrtnEEOkqk
XT5JIyE0+2HWibHqoq5uw4vzTdNEWBU3aW4DaZL1dP/Py92aYAzItNYZ05Z/USpxh/RPU2QTrc4U
vzSc6axscAdQJHotp2bm1298xfBSltFIrvZ4/uOn0JYmu2/7UOciwYbzimsbtrVKJtwmvJs4e2lh
qy492+l7lIXZwP6j+FpsrghBT/jkbDJRWHAB2Qw6dDU6irMlQiW05XJMr4tKD5TkDPhsv0BRev35
syiI9uL1X2rgjSrDJATPG0cNdygGpUHgWM/ahKPwjb70mxxIXOz6pS+GlfSGWLPRr+tldlNy/O+z
ei1xddy0UAvpnYB39ZK44s6c3IhS5mr75vTIgP5zLDbjjc7R6uy/9rXb/dxc0fGUq1jbBb1U5Iz5
cwGxIv7CTNv5K+f9yDJYikL4aFVqh2NRmFtLw1xNbWrewk+SoD33BFMgF5eh1OTT02KnPj1T0bMg
ZQoBo+ww7bBwIrKKyxN2gN3aRSZYyEejlc2f586+PRTI4EBy3e26A6cSVZqWFML6E3HkfP48pDa8
bZzOZWrT27os2TH1EoblHpnxStrGCEf9alANJx7jZyw5vIpwWW3I+vni8+j7YftLh2aQrbxkc0bp
cmPSN/a/aDvGYtYVQlZjEHStiM27icTKW8u34tM8rXCj+gDDKZG/jng1IRFVDH8WT5u5RvBDlrv/
Ay0vN5vpQyLeKjnH2+7MYqZUfRK20dxAComlNXCU+HEQfjeaTTM8As6NH+qspJrcV7/c8mVojuzU
iIdFJRW9QOpjCvQqKFySl/gR+xBthS26DeqoUmrxn13+f7acdaAkxCEVtjtzX99xfFHhJ598ZRV9
s6JqkWqTM6F9f46Jg9+MU33txaDwbbj+QKXEyKeR7ASWmmNzn3RBRMl7bNLPkDHS0qn7uaKJ0yqy
m+MMCbOD9ZWQjAYNd8N4A5+cQROkcvd32uI4kDHY4cnODc6FKP1hTRbyBdApb9kFyVuIMIThVR4L
mV7OPQNelAEM86IaJi/b19dRWY6pu2F/eIQF3O4312aFCsYhktXdZh/g7IbyGgV+/TjF5BMDF0Hn
I20oS6VJgs4oQqBxRptGRvIu/7XArOqQFFceSb5mWIkyu02qtpZcXulw/O5G9Nsp1mEYfCSfFqtS
xYX5QLXsdtRHTYFK5W9X9FbICPiVK646OjSPpH5SnaCIAZQR+Z5YLB2Ek7xOhJr+5EdB1w/+GB8k
3+6FN7cbLMz6di3/6p5oE+qQ+J+3mZnnigq+5HIKJzW10YkQ2fevH174CbwQ/jZ+KEpDI6L/2dxQ
ZDpY1qAGn1O3xStJKwjpSOA4RevObJPmJTLvU9VApXKBuU491S9MCCd93jtivuPNVWRFH6z/L5JH
XsgfmuN2FPxjhcknG9zwS+YYWZ+0fZRJrdC9ludk6GJdBBNUPx2YXcg+8SVWKJWLtnE3tT0eobU4
zHJKeQgAskZR1aROSHmQ/t8onottoxaLGISZrd6wxaPLTRo4VXDUbR2z6g4wSbDfvnuuqJZHf/lD
8Iy88wZTsMQ4PVkkcHyQOx/Pyc3prZpYKcI+znl0kv8+RTRoHQ18eRLLB5fdGyJFP+DPSPboMd0x
dnjykplim9dnqOuiZgP4Nj6Q++dmwctNgEDJQxyQaoCRLdkCL/Taqtwhq0Fxo7zGMrl1+W68MkX1
Yo6B5NHQYSKr+OMp9HxOVwWsvW79qMqCruuybQoT9LrSkr1vNYFBosIPUoUga20PdGP2/VDz4oYw
NKbNaykkimP0wvoBFeJWO/Whti/yngpYlMPXXLnPHzDzVVVNS9aAhPUmyXHgUpP5u9HuuA2g+t+O
jwQtSjrCNvCzVU93MPiCy2rxdH8oiRIQJkJWLR6HCIEb3Ig2SSoUWdwY2TPNvAhn4akHWhmRPshM
XbdCfpBnjVuql/lqfdfKIluUXi7a2rOFXV+OxBNPRrMeRIpOTLx4Ih4vcjIvItLUOYEz/PONzf3q
MiCqK8H0+Q+MWGhbXILmU72lpQdjyivZEQyM8N7IkcifJAyt6Hh7S0hwvpb2emdAz5o8lwJjHE8G
lEH8FcpPuRitpOhMghGmshBjOd0ZN8mTJvWq2WfdZBsm/gu4aUBJmnM9KKJopyAbyDmfLpjW/4SH
ITXAdDLTeFEgfTvC8w1lef24CrdX50o8scAn1EXFzE5Xan10cFcxiTMStOfqeUdFLWyhiy+OR+V3
4ZAna32f6q2MC7JSyxlyJCcyzu04ygHW2XHxrfplZoivM10scaEfu/dFHpBaKmumqDpTVhcAwWAj
xdFeCk7rvgsI69IMlVsxkngVrpJQCg6i5w7IkfLheJpdpCYOlEjKx6KbvOpPgRhEfGf/A7DVRea6
eAo6OfcXaQoGABAgi70LoD+5M6KpE/6uvDJ/BexbfKD6nbYk56+T7AOkPcKiSS7O9vRLqJIe3Ozn
RkkNYPEdbUky+DbAovoU8DviCAbnNNczxz3aKhLvE8Kr5HHPILOLSuBHyjYbwaSaY76qdSn/AuYC
pKMGPgrMpqj/N3nhRcAXwCx9OQcy+ZWtldBpKA8ILfvUyaJD7scLnCLuTPkR0uIAp72yqUALjir4
+oNrw+X6pRsYYeosJyAuIIcXzUV7smCBo3H+Bv2TJfJq/fTPGOdFzhAjAlg2V7vyBy8SeaXa4Iun
m6ywM+vpiNs7swM8P5gNFfgRUQbL8oYnJis/AvRBlHdyexOD02kGo84MpJPLUVNrbkont43gWriw
/q4cFStfqaA827QDjyLSd6wfrPq5g0qkORngKgtnv7i1MLL82jgfYXsiJGBkMPwkd57idG4B/WNZ
R1EUQ6JouBd+Xq+LTYiNbpT3p1S2GyzICtpOQeF7JgyooB2DEwdF0uWrgBXINUO3FBomQUWLK0y/
Zutz0y85QbGutq7RBUcREVb40Nzf+EJYlJSWj6UdUuUdvhhOAn5QfmENilSlmAbtE1KyEsw9c8CF
V/OTycMpphFFDxjgueYo047hNZAtyFdFyds7fV38qrBBUsFi8OYcs7dHwQxEeqSf0S4MDY+tWZrb
fOS7RoLdFv7/1uiJROvw4rW+LC2ff6gRmVmZsBUrwHWTGONMsXGUjMG4oXWc19wVx0u2hAXeNiE9
gmSaXW/TqeCvq9fsn9amD9pXxIguK8hzVG8aHa+60taOLB0gp4PXwZvyxnuR1OeQ8NbKfgZEFbt3
TqMYrQdp67pfbXz5BqQ1wWWXMqg2LgjFemNAlgHyqqAMGdRro1CTZ5CXGIJggZUxszwfGmqbvDHp
KuMFPAcUrthjCsVLYR9pFlLiDZuamtzI4/ENTXHEc3SLUcSaXO80434VN+py5Gs40prTPq9HWmVG
kXQpQzkuIz5mm3drOVmwEkL9GswLqXQOfCL+/Dqie4LxivmMQiaddA2FvbUZOrV/w7LQLMOHnWO5
jK3VsrQtrfihu2f38b8wK9inEKCzfChPoO9spNBQr3GBxoCvl8KaSxB+lwcN2caGkjGTbElZrugX
pfAJ2lm2ltQcgzge7VLBw09DJfw5HPidB3G4B1XjQOpcogbjFG3skOTv4cB+z5fUmwjo8FnVG9yF
TYiUqIBG6cZs4f3WtyTv2EX2UYbowyw2V953fvETpyCsbXcqhD5Eyu/1S8rIWuyXEsCK3Ef9vDzq
OggfCMDKiZhzPtsSgNEtmHqm6bMf5A6yzcorayQLEyaVbQOo5mans2SqjAD5qNT2rhrnwjWuFp3J
Hc3LOOyyKhPPXN8cf3WrdFB+cbEXLvqXJpRI8sAcCZiuCy7eOBjy08OUnESGquIdCdSfSm+hjLf4
lkBtKb2onVDqSErGuTrV7hoU/G5KH5pRAI7fV6XUDByRzTBOACA0SqfasXiO1WKYQR3Gdu+wgENB
VktIwLuhRtF7WOn13eUfvvzuIGRhCQP/KU7mr+ft9JN57OHDyQB3LsMTyzgX3E2NR3W3LfQA2a2i
VY+HeWJe6DvcHwV4O9nA/rQ1szeRUHd5WBZAnjdXf37btMgb2vjQ8hth0G82KCNCPxZKn3Ie4gfy
tmmmpOrSLW+fOBMJ6gjiDtxVeH6VZS47aPmpU4Cd3iuq7mxoNqQH9UJqGipwjrJqUiy0XJ932tbJ
rUJbFDKm8SGglD/lIB7vZqL5zFy4pBiH14+l3YIOLvoG2IijYFxWruwwbR7h45AJdmAmVOcbSZPL
w+SV0c3zhcALdY5eH02pkUVoOvRWlCqoZ6kmPAxvnaY2CnkRMRXlZx9WCQT/yWb01SeWrgBP0JNa
rvGKr48v5OtcJ5zkLSz71yKarVHimh/Nn6qMtGxlN+D+/LoLNzJcddyLuwkZwA6DOec5CNUffgPG
xYis6Hud4WtGKQ8DyLhoDEcf2CqMa4n9X9wyBfeF4elhnS0TDBYCn4N2zQxV2kAbqGFm9SZx5omh
orIMkL8dc2/aGNObXoKZ8E5pnq4HPGnRR09BNJLfTFoILf9Z4N7fH1lsRnDixyR14R+vwEmrcM9D
JiS9OMEW92LAw7e0/L+Ohz2fAco+qftyZ0wZdvB0F9DNVFhdr7ULfb4/EUhAQzL1ukplL5wLl/jq
busDxI8LwHm+58JE3VNO1tbXPOqWZwmSlb4J6aQ8Z2hHmriob2/MXq1PDIpByrNasOsKxj5m9vj7
C8REEZ8KASvkT1gZj9wD/SGFHICVhAm2/n9DAcWs+xkY5VPxIVgFUWAOtDINWSZ+hYLgRJ0dxi2y
XWU1VoWZ1uCddMrBXWbrr46vpgx/7m1Dm3qIPUvhbwTscbqGU7EuB1u8p/xlVBC7bG1TF7SRmcIs
YqRWPBOeCL/+HEaLmFIYYiY6+wl0iq+cY488BAWqxgApK0DEtHJWZ7rJg7IgP6xP5aXBnkYpf/DK
qiR108kyceV8rdySiPoMp4gGV6jIgg64jYj1kIuQv6Su2/nQQ2Ez9M5pc2fvHPgLnZL/WvOA2rsq
eZlqGaRy05C/W8Q6XYw1VxWoPTPA2wnDGZMSxk+qs5gy80ATWkDXeeykeZw7ZZzX0bn35lFeRJHH
p0LG7dWJvj4TIqBopPpCVYgl9YsHJUPnc1iMd74z60U4stJbf92pVokRZJrlSfsIRm1ncHA60yyK
N5zybaoimSd296N8udEBEBK0NNTTGW6NgZEd08rYgi+nb+yhQMxu2m229CPgS/ogpBKYOzpNyDZp
SVUjnDGFgJLxgAKIwOQNoG4B2P6SC1fAZhPQHwzSu+6SqS0FxyACLnaDA2mFccMdH5fkzk0oLrOP
LsktFtWLq/+1sB6bhvhuC0NPwkLlHA9iwqmi125qNrz1eAuJVWiAMki51kjWUgq02aU6Vg7bHfAm
TboOrSG3wCe0ZFhboeUC8pGwySVJFzwhVXQnsQmQ2EdscuU1e3oJn1fXtI5jKL3gx6h9sW6fbAMD
X6tmvoH+Z64uoIoUVrhmzbG+ye14cJB+yfCghBmZ6vqmKOB9PPxE8d3wlpoK1Piw/AAdtsYso0KS
0QmPWlHNSgWSAu+3g+C+EnpqXro6IZ7q6M6GoxMtLlE9KVI2H8DiddmQBikxeARYuI0GFu89CBb3
6sajhLUqEfnWPX7QclEUgHtL1lBKGmmdqLsp7/3Wh26Tw2uxKx8qUb6l7mAkGcVbGhWTBHXlOjQD
CCYF4mkA85ha0eQQaOs2Vv3gWu06MdXgCKSiGejEoZvm3qhRs2H1LDT9N9v719j6icG/Oja8QoMP
DwTEp0SgXeW+pwsPgA2ftukXNRKKCS0pcbgbd6X9be3QK/1r+n3QsdUxkLWNJV8dSpVKewT5U7Zx
lRKsBjw+X16ytkb5JXl/+HVIWwrMAvb5qtmvdmOaPb9qJGkYXmL4AdCXBvtHaESpuH1vK4KeRQLO
4J8HOBE5tjB97L1YEOm5IvqW2+b6w7gv90B61jWe+MZPHlIBcQGGX6REBAocVV4cxrClMPZkB3RS
2eLlD8h21zenVAeecx15xRFYdjJ+8k+PreSvjDV6qpR7C7ZHCcya9+O6plbOc5f1MOJ1Y4Uczrfh
d0x7CwWF25bmsFy1pcOfMMNhJnRdV7p6O3ASEMelrIZ2N+62RHi4JQJUv8zmhLeRoWlV4M555dia
QeSROA/SExbYbWOGVPLHc/QPJDGcU6nhiBJloftBkGK5Fuj+AKRqt71WM/kCaaLu5w4+JyNyyJlT
9MNCNLVKq7VzM1BJzhXJ9OxGogITI1ChB6VxWgCXY26xwme0zNa8OQaRteXjm37qEdZ4SrwiQdjc
tvdclJXPeEuXex90zTRg9apXOeyMCKD+NSPNcvPk0Cjwr1/Cj/CeD4Xit0slQ/1nh1y53GIYUoeT
Qyuzwv87hPiq46cRmNS59Dp8foqIc/6pXGkaa2OYyWeSyl9Qhw5AQQhBHclGJMjjHOCmo60+lYNH
R3RnsCBlvftDJUT0JzVWJSmC8gnGwXbvIMl5vWFLvmqi2zCYDtRbxTXmV9l2dCbOJyLvBYF28Ptr
ArK4TmzjkvGni9kl3VsLAubDUyE1jLwVEBGvGKn4BK2ri0ir0iQra0GWVMXiyJWykD0jCTWI7fHs
FjfusOrF5yCtSWa7ALZ9LFzLpusf+rKGYvJFsaXOJkyTxsGd2jRY4gMoBUSppdXJ7KgaAYFR4thL
mw3tUxN1sJv3DpslstIjv24gWt9iJmO/wmVjnqr7RZVMuxKrkEF+yTa35DNOWuD0V3ZViyk6uedH
IXjcxkvIbyOxW2jkSK2uzSfErPnkNrL77nmwBCp4JWjWluKadTTQ4OrVKjAHAnG7U/P1as3n5G+D
vBLBWPVhdg66Jg1WYQmBgrhH1EaKFfLpjyK+MaQnWx3MtCp4yfpXb8GBP1nTUWk369/gfz4ciWjP
9aUHFdyico4Wpj/2EYHaHBxKFy+qTh6+XhqV2h9fV1dDIi0Xv0mjoIJVKQar1YR6co47+Qo/huvS
X2mvpZxZiMf8jb/5DRWmtgNEsXfPt+tX1DTNW5H6xSgG2gD8lbuzoIXz7lZ5OZSZFarl3yIpDx/M
5QO+2399kFrd1aVL2N+CQI3Qn36mnxBdgKgSTG8Yl6Y9/0Zg2bW06LgFAALEp2+7kOnPiZWMZKNv
q+wO/4CkaSffN2IY8GLeSm6SKniRCpfQqWu/ho2pBMvjUIInhmyr05aa5k7m7ibY4JmlREDpBz24
/ZinYmQQvfgpIYj+OzZm/2HGUt8knJ2E8SauFPLv+kDMypSTtXpzvsqB6cvfmRHb3GRbWdRcrKmE
0FDCq9Xl+MZyDZSzkaQvhJZFrI7KFvS0mnk1neMeBXgDunQ4GEITCqLQXpHNvfLF5VxeVs8rPhUt
6JlpS2KdTKXqUD1Srm8FMBe1l0Bnbcyjy1CgxoDWGdjZvk6ImStO8FJa48kA6ZpupEApZbcmuNOJ
Ba/uJrJ88ZYqoJ1/tbpVllOGaxnlJ2SLI8bCrTceU+OdHcVsiHOj1tU+rzTlNVEqcX4IJsabhNzE
ni1ekMT4B/bMO9ZP/THe7U/sGfEuq8JtE+LPpdSoVJvg7eGL3B9JDAjYMf715ucdePfb7/63AWYX
CnDswUf87/2uGRZVHqCMqNOhNpiWDTbcpFfI1yAuT25encrjc+2Y5mb4WxTaJcYuN7wdsIOCT2Cz
dZI9/dSNzUa+sM8x0w1D1CI1LIvihBnCzRv7k9yVLPNiDKyBcG75v+fcQ6hmWkVxwz4VOHtl3Pkh
KlqnK0G+WuA6ycEfjDPQxEiR4KQcl8KVutN486PuZ5qMAAJsCU/Bg4S8COTGKt5wbnHDRiPP9nSf
5n2v44xfjV+7W1RqyYgYX6kLUHzL0LDSgt3qkEnBkkzZOqTmO6mJruQov5Of7wzfEvnD1wzZrYIp
X+rlDQ47Kg6tHm37I2N2WSw3Ih5Eftn0HAwDkkvpNSAiWDkuisQqADqzX6ldeLg0DqEVdMempTFi
eK+ZS91hPM6WrCTE0FLKqZ30EtQo85a1AcLXX0AKzT16MnE1HtxGZrQueo03GB80kmhtAhLoNws6
Camf2Uuptrq9XDgv/fujTpehxx+q0MmK1GBajSQ/J60k8lbr1O4t3nyKZBUus2ZTFW1JPE/bt3Cq
jR8wdUs6w7Vq7E4/PYenWelY6Wc3W4xJBXNY5+HSfBTzIUTXqYHRF0tUgwSbnbBsUvmr3szrRFZs
STj44Ke2dF1suSH8t63NhhxYfZB/y+MrJIHf0lzX5BNbkEgzVWMuM0CiVeQ0eGUlY+dlA5IuVg+r
h4BbrG5Yt8MeKATYo5TbuaO+11GV25+uyYYcYljbpSQIlz8Thtc6dnQ2IJ7ZfeVGshlFP5wrP8bi
/k+chgiXsWaJM0xk0nyMY19c4RtW3NcSBtRCQygprySbEdvTlIDs/CfGApLEe+6EY6ndTM0x9Kl4
U94S9mKxscS7TbNn3ySi1U8ILFzkf4SK08j/yaQtc893+rGN/zgvuKiQiL/csXW2gfkEJURc7XNZ
uTW5J7UTpn+1e1K4HRCV2TNGQ2AbeUo0vsJmnWmc5TKZLablXX1/Zse5Jx1V0h2P7w7WM2fVsCTd
nd6bimFHuF2G4NF+/62ceFcWgfYLFrA3VUH9bTGpVowSktDFUxknX7xoXTR/jkEAUAMtqaCFTuRV
KdpQ/0kGpEH+XLHF52y+XVd5VvIaIdEUKFoRvyN1OPaCfReSoFs1YO+zd3T6kPfbZItA2TNMY2cX
sfmOyIOm/4bmT1KwhY7ZqI9a84oGafEkQ7Hn1gqgTkdhjTi7vK2/aMr/qKFPvXRq6dFgw5kC5DLb
LvIWLIgmdz85Bsa834AVXPRDBf0tgOYV/LdRuwwau/g5+QyUK4o9lSnwL3rMORW8J/JTX6EaAFXB
O6ZaAxoN7Y4eY/QGlU3zwZZNATuq764W+VB/4q2TRdb0CoO86gLJcqAaVZ1yWwenQ3VPrhtLdwOf
v9/dN7E8DVuc2MfZJnyzUdgHAoYNBMGoMNbEm4PVUlX0BYDjWlSYOUKPgz8LFvVJzSDNSdjV1foX
hYD9XAPaOcezW5g3OVLVZDFsxdRuz+2Knfjxuvyy4fdDm6wsJnUDGGGJLQnuI8Nkr9z65oZMSH+z
vkVqY3IBq1HY0bFY32BNzE9VZNufgiXQRl/StGlS3m3sG0ApjUdoPUv3/KUKMVXHlTGW4ZANZVzp
9cef7pg97Krk0aIHdON5vrlDxb4AJ/adaEi2Ys+2Ty2Qie8SYIIYjB+RrT+Cwp09QDMLzK5a/W50
k7G9jjuwwb6pUtvnmimlfodPhKtqdjBqX32CI12bVESwtUR1oCctZo8BHcY5NlTGJYLQX58Xc3lV
vfuVASSwHXj+HXqUYPCDTtflIL8ugeqUlG+Le7EhVb0R5khAZw66YImkb9jyX5nCThRPAZ3nSySZ
pWcddkdbR8kqKabdNGH3q2SNXOCn81wmft170c62clRfpumj7UGDuIRUXfyGxa41ejrL3801u2Mm
83A73TutG8hwOiiSCocqQ6KMgvoX86TmfS52T065AVHOd5p3isRHff6WZP2xzUht1McvpAyeE9+v
FtXAYdlIsIH7DMu8SBMTUyIyQpdLZ0CaB3vSIrTvTlWMkFaWTvy/Bn6U/KnSIhKENDU6rxzsWCkR
mBa81q1G7mRl94lb4KlpwowW8JbCrx2HlYQWEf1CY4Q57at6ekPI1U+ZIzgof1cTeFcO8iwZ4XSe
S3ZbJGVCNtTK9ZFd3593LzV1twAR2Cn84SaM+Jqd8aDXbJ+wfM3iCaQ6ePi5D6GGWhHnK/HAG4mq
43n+sVbFIOCCG2q7WYXoklyYazNKDQtv11zTfCGaKWmKu5zdBD5sA+FYuf/qWI7Zsl0tnKi0Ahgy
zc5pKuh0qhZy4y6evGYNQoQy2gv56+I6Lp6ZbnNHapPm3llqgo/cJkqC5ReEswqITaPSZSd2r9kW
7KHXM/3KnONDye5UvLEgf+qDP3AEt/k/GtpgFfkXs9SDayFmt6ndNmdk2ViBCNliSW8vpNtPC4xp
ihy5RL+e9/Wm68GTpqLXK0fBKeWgrThaDrsBDPek4TeanFPCBgE0ARhKsuE/aO5vjC6m85bpw704
Kv5OWHm0jKlJb8LiWs82IjsYTRkTrOva1R1CcL01xLKQ6D2r1m71AdzfurOuoX6FXjHXb5ghLyrZ
un+aB4PcE0c/Y26qzSKvZwVBx5fQN+gHgzv/Hv7e1XxZg4uyoqheWQSUfcyKtZovrbEfO/rsJ/nq
REt4ZeBSf7JGfQWxZB6lirKwnIjeGuh6fm9kKozmcQRG5dNQ0EwSNcgN/F6ZoRQufAoNfagbW2iv
iUpZhFP9xJa1bVFKXMrwESd86yS4Qnp0P+YXoBPvLkFFWacsV/p9Jz/WabrbzGW8nb4NCeUPBt2v
hmANWsSFuAfXHhJgy/8A9s6Q8FtB2yv4pqM0uQELEvvIFPx4n4AkkkkmC5kVNJNI/JD7T149wl54
YWGDn9VAeC+LNVursnO0lwZMy89pb8wj4Fgrc23toEO+zWmBqaKqVEcc/lbYOi55SYrh19wtzfYk
FwBFsOIUx8uFe7YHmMxTogNYzzYNqvN0h9ZTxQV1rVJ5rJKZWgxAecS9lJJxPL2BdbUJwjuP/dMt
v4+vF7sBwc4GPWlIgDCfOXNA+BF7cOxVYX7kfYYJx4xpHQhHrkfuzyvMeHaHjbxx3RVc/1y5ZHaL
5OmZWgaugGB+JfwHZdMbGTq72Pt9hEWtagIMK3LKG1tt+pf3i7qBqq9ZAUJIM7WAkdVWC6PxU7UI
T6QdvyWfk1fNOHy0ldJ5Bvlev4vwBs8PqO7dbUg7kWao4cznffedSt69/w/4YyZvEtf46kucH2GS
J9kHZWK5CiCsZ0f12WgPkMxpdjcXzzUV+l5lRKTljsnmO20fAe+jHQ0KSVg48VpyMnF/QgkTR/Px
OVdq3yH85Lq7qm22glQ4MdyMIBP/zn7PJmsd90kHJspav+ufrdw6kT/yBsiD8VM4wtDRMVCG18Sb
RUw10Ne0gHW9KqBO0VBl1CGi6GCD12EMxQtLTsMIRcBbmLZvfYCboM6JBifEWTIYFx1/GErftpgG
CqiF7AKFjD417Rco5snO98Oajs5Yx7DcPFMygLRxqMosIpEgneTigKROo86URR9VtzfpDUtDZ3Op
ROBJ5HPTXDfl2ZDkOylz6tAJWYz6F4zAulAaToG28v35C11pFvOORO8CAU6KttV5PixhU0TYF8uX
XBSMdNyXwQvMQkDI4nD8qTJ4y2q0wC2zbTFCY0dEoteYsCBDpwd3bM8FQBWCrVH6pbEYpV0c5Cf2
SYw/ISdM442nbuFKXwgtm4BqDzQBkdlcl/IgZKnsGefRyXH7qfWPnyPHNJ25tkUuL1k9JWNUarEf
y3177N0eg0R/BnhHa7JVxpRPq2wRCuhmdxep1pteVkKgiFxjtsF48xG8EohsEQMklm4Xf36Aw5pd
yG0WaKnjPVlE5DZmVuC55n14raFF9bQGl7/cNXYfzS/bGTlul9fMdCwi+Q2KFurmdGiGlgylI47X
ygtzYnqkeANujxlMqpd4MJOvdCLgSkfAJ1NCocYd1fRG0FhaaVv6sVcRAX2hy5S+Yn6Sw0elX4bH
vIGjoTn8t73HJvh7FnvbfviphN5lWnZdJppl8jWX6fi0tkBABHLKwepLQHLhKP6tZ2yBnYMcgOpW
pqzcyftANXOclP0pHjzJXuAtozkNvkzF6Gwt19S5nYglrCTvOyWFsWImUBbmPOK7O6UK+/6bcjAu
Oq2omkcNFrTCZ8MNaYJkYNcVa9pHLDXYV0nUv0axkfevnJjAIICXLG22T07Cf/O5c3tyerpyU3xR
7JDrDkSdOkOS80uAHkyskVj55IgDvPMi+Lsf2lXTlRIlD7yBtoixcg46XPxp8bDithNyYFeWMKn7
GUQe89jGBq3qPe222/j5DEwRH+Z7KkwwXDYRmLnPncHtsjmV1065MKAY/mAX6w1TMvFrQFRl8hce
TB0dbcfscbHOBuGAiIhnK2GZVqcctySCs40g4i9KVest3RlOL6z71/eFq9tFKJBgELYumeIcjGMI
OJ4NKnpOxTS1RNO7T21UXoiKhZcO+Qd1zHeaEMp0ko+A9SMJ37bigIirlrQRa/ugpLSOoLrWk31T
QC4jzo/nM2gKXTFf36cQ9xrJyQi0bQHIp6aLfyA6aGht+9+VL8ufbrPLZ/nSiKPGSr1qUmXSwYYl
EwriRPQDc93t5yi/gn2ilry98uR+7D6W3gvFmxXfWwOnXUdleOPtQp3FDpj/bA8xqOMyk2b/WL7N
aZuKCOFP4lApt+N/2bvv3eY+lGqt0FwUhaN6YRF1UtTec9pBoGYVtB+5xcDJYr3N/eWNkejvpNu3
34evtzrhdTNR2LnXPR/gcV4R8jfOCZ4cqy2Rv4J79TgkuYl08tt4eOsAI2KMFKWdGFB7afcGGUuK
iZNHxaI4wKO+QbzWc+5wAC0MgXsF6hDnKdHH05GpUynpU82xFpbPqi+ZlVLdgk2huqLR/KsZ+AtX
urVE/4Nne7O6lopt3zWrgRhKurQDUtu+0GHJku1QiDDyDKv5I3cCDrdZ4BY3XsgupFV5+qtZMCjw
59khw6GW4Te7qXTNO+yR6PZHVxkZWjnJYoXibzM6/ARen4soSlf63+MDqjG4fggPr5UdJwzwbuEr
s8/djPTrqpWqvxXbxK8bmwc2CSe7LtD3RUvQ3c/iGCAw0qciNWvOSN+pOno9vf8nSPUX9CmPyNE9
YcbBDy8UwyR77Y783YY2zLRhzuvsaqXGbBT5rDT/wnNazA6UK+o1U2I4jwMLDAVXPwjvArDr/IxI
S7MZ52UGd3gGPnIf88oNnvs22PxbdtEH9p9zaGe5NqGl9Onpjby4n6v5hgxKmcY0mFKiBTQS+0al
P/BOJZEBEWYUB4iOIVeHnAbA+Cn0XNR9NJefAGmeWDUo0+XClEpBWJO4LV0kjJV1snXon1Zd20be
LRJhrln82NhrwZBgiDo83O1fAxtuj/EpOc/v4pesoBmOITvHKDD3Sk0kHll8kQVOagT7EDrFX9UA
troAyYGJWJxX7mjfQ8D/4tySPhx5x1FhILxah99Gnm3Yx6pu7U7TB6/fvJyTzaU/FUB26Hsjslb4
CBCZI8mPTvmSJGbdrUkhp6eYVonPTB9pK6nUrfgoFB6dSq3HKusu09VtwCADhPznmkGb3pQG4o1+
d55RdP9AVEeTCR1qHEk1rwzEHFp07yb5XmsbwZZt0q8v26GLSMW9Ns6duSVFEJKkFTmJz7SzGAYl
lU/HBmYGaD0Xf5KYV8fxL/ugvVhVImVF8ypOWVEaiR75XyZ4L5yUQ9XloAKvZ9XscD2WzmfqZ3BC
PHVPsRmWGPzv5L/wkBoeAbbcp2+/ce+9jJLj3kVUczKSG59TDEG2J/YcHq5OrQk5n7sCXo45Wwll
v+68eDF61fYyPo/uwsuOS+tIz4ro5fC6GJSEtDM8s7vq+4l4iS6VWSLEOQrIa/dhCWSKdsbA5ywy
R7GI9WXyDY6jQQVNlaOO3dGsgqYJeVKyA5u1/VacsbD8TJoyi6NhBDJZJb8JcewosxH7PVFcRdVs
SwUdob2OE4DOrrgmZHkR7WVYfZD/gHHwzZ60MYh6RYwKsUmdHwPpuqN9nLOXQjnA7b2h5dJsKsPp
ij7mYUTxVN42z9iBXjB9ShOTyOqrfIBqGV7BMqlKr3H+RBlQQL1Bpl1AtS9ADpYOqcICCAwuTxfX
pi1Hj29PwgOTA/Eq7xUbDuoqzY88mRzW1hN8Fa448dU30St5TG1FX9V4ahvimCucGKBCZH+SWqrh
6Aq/huE55KIb5k1JT1s8Rnweo7OEZp6ylP82mr1Ph7GDJCfmQtjgbQDbZ28wiAXE3NlkQ30rJlQU
gSg3I9qqW+U6eBuw1VfTlHssiJSRc2BE82N1J+s/hLJWZ2GHcIcIvxFyIkcYn2+v1RLPEY2ALgLQ
1oY+lRGRindJWQQkHjIFCtb51cKfHUks7FdIw+ygLCERRYhVq8d4QyNPchB4Y3d+lQb11FsuvxiU
v9GV+nwjxH/00sghbLsxpqhgRQHt56p4fMjr/dzzN45fc1HXwnfKwcqrvpFgrUNljkaplTiJCBMX
e5Cf7MUssj/B2M31EqJwOr81zghKz6u2XnkHxtP+bWbBqwTNELB8OR2Gd9ltiCKJHtQb5S9wCz6s
73GNx3f8W3VTf/s0MwhBmsU/yTMs739BTxc3u7AkARqqieszCzV8hho4IbjatmDQlFirOM6sr6k1
EUUCJNRmzg/OojUXK97rDmdlcjuaHikEri2MTHwM3H5TDFr4oPdONxw85s7E+ZXtqxNO4IDgXods
3T0sfprYWxZ0I6R+91LVig3/9c7rPrHKPqanTkiHHwaWactBqhWIP1U8Itg+tC1kTZXsQ9F5vWcC
jz1/bfzpfbmpL3WOkPSEbRqZs7HvxQl5nY+wkCpMZnYjHl0SfGnagsHRd0pDRKmuMK4HZg98Ro9I
8ukbKQlTVzPipxh5EYvRkE+Uh+CJBF8Kuk14G2i47QFCL2E+87qKRfqbTn0L2LLtkDC8ugLZpIUy
9JQ4qdVLyyVIG6rZLInLo38kL10uR9mfOnPRYBvW+NLgzfUyxPFWOPVoFexsNnkwm48E00dUD1kH
h6AKf7dCGjZFrTgfEY9xeqhXA/EXNls+UdTqBtAoSsJl3IXp//nCSyk3mRbpWa2F+uPcwIwA8RQg
xL8Bru5dzYVix+r9ZjkiadT3lt+KN78RvB4nseFXDP65H0OSmF3miHDaWM9E4r84Tuzx2orM+aX8
YV4NmbBgKEmmLvtd1qaVhaUsJaewVOKl3v5xSyTVF69XUEv2+S7o0K8a2JFSvRl6AschQwqh7089
sSKfSUUeNGdBVwcxYhRY5XNE3FWmzCe7tQfYq7vk/n8RcscX+XhkkQ/lJl5UIne2Jdcnvpv5vlkT
7Wsn/hmEitrlSPWyJzR/AdyXOKLDiQV0JgsVuipmO7bZh7HmcVsHImKVZdAGjkjqYVXzg8igR66K
VKh70oM4xZTY6MMFjNsEHLffCwSCkq7ToDKWbKljJrkL3Do4Pm7IyLkFFHHyLpoTz620GLqbQuli
ZwMYtpcBsv1JDIBzlmdJNwUKkFcVavIggAGXlekF56iqlMnOInCwUoG+4kJPfOezn4EaDYHE9W4X
vWotfMJ01omjagKwEoym0iW1LniILteNf8NSR2BzxRc9VNIhtxFjmX3BDg3DA4PTsAz90yonaO4o
+phZuPzStOPlVhLwe4mhNGOmcdsMJH7/QzWEk4h0FV9YFeV7It3LDVbgcI+0h/+A/epkrSAeoTtp
qEDTNOyLksbXyuEv/npqrXPx7mq+3EgwD/AqsYGa4YaHDcZxdmIecNSWKyayx+c/L9hHeg0elpbp
9PeRjZivAE7sZiBy6YLkh3UJ6coqmtLz2alprE5pT53Qxe0Gtu74b0byrrvglDwuHSC23h5noZrU
gMzeI0HPYzY6wWaLDH+I+cTHRxGIVqXbirBVQY/TkCvPKDjU+kh4HHmmfOVnrfdLs27SVtT1pUDd
dVz19yYns605YYug1S1OxMXlqGHpPj29zZoVHzvsYTlyqV6akCxWfI/XxO1HtbruSUIs7TuBnFYB
du820YKO4RlYksJzQastsf4d1T/nTRqon6cwLKXD2tnBsZ3Wm8jAWxha/6aZrfsgr0upB7mOxpjj
/aHEBXPNYU4CbgnFcryadM7fZlxdfSgnfjJbwRV3JLIdljBooSFlOfFOHM+Res5XOrILf9bsp2on
ZkWByYMfxze190oCPlTSoFnMlJpl6jzcxf8LcUMczJ9ythHMSL4Wx0Sm4ge3QADdF5xRxhE6vHKi
Ox0AcRzluS8M8mxaWfhKAJ+6XAIxYLVJ+q2+wwie2JX8ujro9k0Bz3a0KmgAhHgwZ+x0TmTtWGOn
qNvFOClLhc4f5zQ5+brY6bgEk+m1B/0S44s2As8CnPkfQH+YroCfKQi6mLbblB/sbiLSQIsF6nlq
Z2aQNIPbQOhtTMyiL186k2JKkU4luenkaabxPXBMc+AoSsOVZ9PTsHvsCWae1xYrjh0dStYUhj1G
nyMyXVZxt/oUcSwimZaChPOMCgmNiEua0atE+SzcYYir1WHYJCKlKoa+ysftnDr3ptupTBs8OOdJ
beK97Ofcda6hHCKOM+8hoFMw2Wh1LwDjnUKVemYhYXkin8gVHPvJTm2MC7JKNfvLDVL6WY+lIaVg
2jI55Ufg3agKWcyVL7Z9SV3q1r9+LulQmgogypKkGkqFGecYUp7JsQEj0WK/G2fLWdB0dZVVvK9l
R4sxb7+dLD8QGYX1TJ0ZLa28IRuV6ZCo8Ilk5kkpCttqC4qpURQeNU8GBHiR+YQM7K5OPqZKW+TW
S1MiJw3IH2hYg5DpUt/t0SXYJc6NgvYWQDlCMUzwo1rEsmImggADd8UDgVnPE7/IEmVz3aDq5OV/
o63/gPPIMiEc7u0gCCj5UUqgAe/NWXS8fcG/u6e4Sxa7n4uEd7Pizgh5hiY02S7jj/oGqah3y2qE
N+95p3NvZjw4dEiExdgKzVgi3DGSNRu7WFCIva02kNML9MzZ6v615eXb5WgVW4pzOTijaqQPCjCA
Zh7Ur3zmkwQoX8Lh2IUl64rEoHZacuuzDdZflUGYaaM3tIDeCbSxcnQo039uxQZZKtc7XKfRelLe
n/yovnoQdpBqWQv5kzU/6pU6Mk4EUUk9ptvzE7TT/qBATJBUMww3Lvq3gl8c5SpwO8teN/swI2c8
ei3M0LfxPWDTgg/OonMM+ragvsjPZjWYpYDqO/AAFkpYPIxOtiLt9MWrUqgvPBAODuPLTr/TDygW
Yr5moOHjrCalM23XuHhVtF/MTce6m2Mqrw5bUqe+Zsv5am5Gp++sPpeVTLwBiuXK4GRaHNLhUCNC
NscAMyoMZpabHQBk0PdUIvVmfuBVvDyfRtC9Ppp5ddYGmANQp9ThDm51j1c8fZt8K3fLw45CRBge
ki4ATkPKMQGiR0iOhcSHw3Aj0Kl+S22ZSUV7charL7Kd+i56t3T0fciuaDC9lM3NXNo7Am8LPuBY
ALVPP4b19vFaxiaTwiLFfKKoWUoVWw/88sZWJiRg+tIliBele+LTUhgTORJpnKTAviFp5kA90xTk
9dF7qZmcTMen0GOIpmNqyW+iGyEQCDJI9NC7uU2BIQNmxZ3CMWYkT53tuaUw5JO1Q8qTBipoOWKP
R/gWBeYSWHY4kmNUT5YbSzIJIM0EFO4tx9fnrMlCuJlCcJ/RG8lhLUVlCbheTJF9Xvu2trdWBrdh
79pgs/lERy1y43rUR44XbDxf7zENYL3qHggKqXGNC/qYfs2PTycq9wwwNIQahPqCSwXjpLQa09XO
I6z0Vq6sjWxqZlJktWeTUq4c2LRQVGVOlJEXLJJyUX2JwEtacpD2AuHX/e+vaDP3QpAj2sEZyN9P
yyy0enBXtmVsLKRNlS6AJy6Vz9XsQipvG8x8U+wbqYY8rSJp/8Bx4+ZHrYvGII+Rz2Rt/bpGcBSk
Rln2ux8i79BO36oRzQO/fO6nrtp+ixCxbnxu+jV+qI2eYHmohyD2yXqKvZ6ZpCkuxN+IeT2nU/2H
bOeSHWmbUTrmOPlgYHzg/Gy8OA5Zqfe/gofesa3VFF+DLNupsyAWNOb3Q7nElTDQ33c7dOuK/fMI
TDieL6oDOxu10ZKS8Q8l30zX01PNoGt7JBGeQmVPE19it0VKY3qAdVZ64aqUT2QWW4jbszF0hzdt
dVsP8aIQOFwO2yYdyOiXVfmPjHxGyMEznuu5pdC8YMktWhkVdp/Nii4ETv+7QFwXPwxAv4YlB+6D
FsZ+Q8CC7+AZLaXhSxsDaI0HJxmdQ3Q9eI5WZSmSgX/H4Dvyz5kgz+9ds9UeVCaEBvn0KjM6yg2I
3z5cJyMdaStKMDg/UViDZqkebY8qdpDb57QOyyYniMR7VTtTx5UYVFNHrikdhv3e7mcZnfyzziTZ
A1D+xgsptZQrFY7pkX+aC68Fjp7gpXvmhIbwTGcE6Ekjg2gbCnyedva0frEuT2omHW1EChdtUIK9
ddy9ncDJydIg16BDU/dP0CsaHCjPe8XPEK8y03EyVciJlzVcvVrM2fVp/iwnM4ibZJhhQBM4UvkE
GymT/8KqpepODOrSpTbUhEQGPEHINNRKnyA884aV8s0XVnHgwowjtApRg3RQmDgq9Z2WvOt4fqX8
NqbLOt5n/BhDE4x4546HDktwQzPXgD0ydGnr6kbi+0VZE7fRaVALLQQw39B3MwfiClrA50E432MO
42i3F2+yjQsmeLsKDiprsJiWL2QUO/4WTlUc6OBGk6Zbsa/9E2eREqvSo1JJX6ObGpcnjVO/5GTv
r3ZNOhe1HCuqVguCqZE3VsSUDONJoruxOPDKu+SEGwJoRy2vzIPA27Tp0paZva+d3XCMzCPGX0aa
FGSX1D8AouwQkTJSGorI2Fp2tz8Fus2E9i00ej4j5p0MbtrUCd4pBhd26IsPioMfXnYQHRAuii2I
Z9KGyXbqgNnC//yjyURUAChQYdgLRJEAVKodvFHk2f3cEdcFKPOZPSCApcA0GC+YSx6WsVHs5bj4
6UAIemXkCXt1TXr5Yoi3BMDTQxkCYH+gTXxnh5bbw+qkkeeDd+AWzEuAX2mtIcLW5CWmUlV7gTlv
szx4Fsf/vJTdP+LtSiCJ6JB8bO7doQUn9hgNrVOmyw4ORFp549Txm3ovl6GNsVdc0zWAFG+uWS0/
YTzvHcOQubg980IaMkICpnL6ojap6uHpxOgKjfn0eHVhxKliEkbuf90xgutDlHhqgtcHXZxnf0zy
UE9solIG1dfSFcEhctTK82Z7rueL3BvobuBfx2RmqfqQwbK0YIvEi8e2Z+YdVgiH+64n5PGZyVTi
EpJzhSoBLFM6FP98CSSpL7t472TeZAjb2Ab967mbJX1CFi7yi0z3Thfa/yhLm2j7bvyL7teK6Jpi
2pOsy2LsmPtO04EVlUj8Hz2r23mTjTbEW37d0FXrDizOfOzWnWzw7tgQsyCUpCFyJkNH/SwBS/ir
SRq4y0zt4PeUu5kOSmTRLpauTRZjNruIPazdKd91a4UO+Wn74KPpfUJhWCS7QB/C1KYOCs/y8hMy
HALbSFrO6w/yx+CM7IiY3c6BobJDzj8aCDsmmZzVjAtRYJ6r0acv/iLACXvD7tk32M9snLBXzBHN
z/o8Kq5ZYCDY50Bc2NxR20AZdE8/k0wjiJB2cCdO3wp3+b2hRP6jB1hHzp359LBObL4phvHWx958
8LwyRNQSt5aDTdDytgTZW9P7F3QwpiSZyD0iOWLQePTj+nV89ynDFJOHBg76mzNVQRTF8o3tTqxA
ZUGVHqEmsKi6vrQ2Yz2DnmS0qQQFOcpwPHJy64hNgDCoEafORtkZ+VJxj1Buc09hxfoKwRctGR+1
iRpNoc0DEYjkNu8fdzxGeajWy9huE7G48OjHTcCTuNXHbyk5jB3WfF93SPjgCcPsVU0peaUoIV8X
iLQEP7pLQ2sJntCH6xJDTZkCR88TaevXPwmRfC9MYp3BH6w/qASilbnVhbDrVdxA322P9Ufqp8kB
PCtAsAftorwgusIAJoiFbt0NPJfRlg8lrbufOCoGlQft3F6HTPzQegFSLZZ4OT643CfQqUkdrcCc
PT40lGWDfjRjEoTdXa1iMZPYI1O8yTOserE+jxuG4SvsBYETnWdNBaUlq3st5diAdTffQ4qviKeY
MU/h4TkdS+eeNP5f51l/UjytIu1xMqhlRLgQ2Vb2dlDShgvZHNaJR7Yf77jY8Qk36lmzpvLfY3CK
uZfFPKTWXmGi2uPRmE1uK8G55n9VNtkLw5NCuG0dNfPyv8Fgzi1U6iOV4D+q7vHJvWOf+yiVi615
lv/wscQc8GxOKl40wI7Yp/DWcK3PlNltUqk9CXZgPbO2Sq7XhAtPMsKkKtpPTvaMuJiJLDMawQZM
Nh44Rv65mtVDvtkW4+3EIjEhB7yiudJBVatbS0Zcj3443ph75yUt7GaH1HFH+7VHMNE8dlqhfOwi
9h4Za2uYJNtE/RWgEgzrVy4ZLI5kzZeFsX6PdPtLaQj4LW2ElQM4nn/NBWuFrDx1DwyGccTb1mux
AXU46oEHSvNVAMv6MUg0F227eS51toWTUMh3fKwRZJA5zcZMnCgOToPBeF7V8rHyxFkz1oFTvdWj
pJ6FFkmjsRmUeDvrpLoSsOHysBphuoWV+8PFRLQhp3YYwjg85WETonNyYZo5j67qEfw5UhoEByyt
j2WISHP+DgGp8CfkS4t26Y7jwq6BhpUy51yramlpqbTwO+NkNUalNhiZq4jmTJnMRD97/RLF9v3R
4Shdc2sZX9Ef3+oh80DVnCNkLcZHeeSR5UgJA2bmk1lvtkwmMiIM5DUFLJQv2p5cfP3KtjM8gz95
EvKhQNm9iAI+5cRmgwIZo6ennrpw8gW54yR2IV0wdbgBdKYSwUWeAzXhm2iFyqeUUteaNgmrdWLm
rnngojzwIXB5J0h6XsieSLfwckVddD4S+GnpCl19k4i4fJUeGDOenoxkgzjcG4zaP+VALnFh882d
OxdoZzvQgODCGRZ5dAnaOeol+cpiZNmLMSqE0sOiLyIrFt9CACN+H1kdLKyWwfLyw4b4t7xe3u3G
Uhy2c0pNoVnaeUaJ09PPiBFRZguouAz7iGORMTCGzoI2Tw5sdqyNENl9+aUHPgDs6WXS1Yfmn09j
pYJtiPHfRF21itKxgewB7ILwgcZ13DsHtN0K/SXmscbDy5rJKI7A2EThgMa4jB4W8xU6vLgCQ8eI
/v4xc/RJi+BcZtp3JJnlsuRHP15Rpc9duCINNDO28bT5XSVxxrEJ1Eq7f3p4r7XlqwaKNNQNnuhh
nrRo7mgvGx95oQLcWchQXyfF5As3Odk/OUaoCAbOkdQEtZSVqVeq6IHsTp9v/IIk8+od0RzGrqoV
iFvHvlnRal0apk1WEz+uhbu4XnNsxT2qfWtwN/MtbbKZ2ZeU8KTSVbT6KpWcM9csFKh5AXFnxDpx
MfPzVNpSvv+1quWDVGmjIa3+Q8Z2IfSwgS5KDG3y+ZxVtXHI6Gvr4d/BlVbHB+Dxxc+IUgthxCmL
NMQvuXv6Q1rYTu2p4v14dGxAdMjC9djaTjNjGImEw9WNqgXkVwskkImIHp0ze95xGI1yMo+YVFgd
N3uUSgAPZBRahwM7IXjnaKHbMy4ftFF/EaXb2zbtp34+Wh1gWvq9Ppxnppjsqp3CXxPsz2P6OdTL
iUKF5jmoWFoUsl4Bki/CMM2k0HNc8AHCYePHiv0zQc/0Ol5LlSlC0o6z8yECDG/iBLnJlIVcdk/e
YYFzkxzP7fIhOeGcWtZTFSp3S+ZeYAL5xHDdkZXCc0ghtmRZ9GlO3DupXBeNNwMIHeTbSfV8HeXX
AjbqW22npPweeLTnWyw3nUSFzHP2GROlyCoroal3zY3g5FIcZQddOI5rGUaX3vp3zKzAMjotTWBn
m9H+Yt1i8speC3quVPy4fQ8UyDjDPHSRA2ZL+mdZ4j8zsZ3sFCnryPpscNa/P32QWi3jezgLkX7y
pJHjdaBOdmsgJTJlqOrfBh+ZZL+Tpu3DhTI4wkmSPo5GhbrkH9ceF6NDuJ8gy9ptTMeusVlRY8re
8UhR3oKxeCMOS27DXVHkyVoKM9Gyo8m5g7rp/xH4P8ap9/gGP1vpSOCFAS5YrLNTj8fPuKIh1iDK
YGUEmbFJUBY7ujeWKT9aEur3LkttjUmhNDSZy+gTaKCvRS/CBAPWr9PuYIro3LwvZAc2iKsvZLOT
1xUaEdku7hYTkCuqfs1tD6Swor1AqqJowYiM3LFNuLN1WYmAnXffclafIQovBBR1YFM9YINyUFYw
BD9R5VxZTfRX7yX+/1MGhT1qkGXjvhzq741v7tqD7a/z01t8gNWw6Nf9pcir8J2eYGhyq55/5cwT
A1da4pO1vQfe7YrxBAMaUGezHsDZ2RRlHk06HDIb4D1Yab4jh07E6LCMRvOWoJZsqvBahNzXu44i
Xma6Wk125uZeVQh8qbzqnxBNBZpcDwrQQih1l+sM2H9J3XQW988mVXN3C8XwSwVLvbkt3HovXbVq
kPLfBDxtQ5a2Yxfoq6RS7LW1V3K+FwZGSQGrBhXKILoV1sTGbXV7h2pk20p9bgJ3iBzvNtAGeusW
UdYHB6l0Ih4yHhyuZMGVZWENhPgy4P1hbptZk3AeVo0JAoPFubfRcNY5PFakdN4wRvymlgIjkAWg
cRLIXYPbQztweZqomtCXBWrWhGfAyfDMOqKAXlW4Ne3OAHkG18EuvQv2BjyytQWKkKYP8ua0CLlL
NFK4HDMIzEzX49r4/YKbbzuM5SLgeu8pZxHXVs5vmfEuUPaNyQ6Wr6DOdSJIBgMAozvgUxIztUoF
570vuV5mgXWKf71bv/eIazvjZbt+PDDS4wuRrD6p37W4XsCqgPGbpIackwgf8kSpUoIIzEcnteRw
TCjqpWYkJ4isZZKkWnVtZOlmDZURHqhGJ2BPc+sBfYpyA5/lVGXBj3wESwEEVY80t/DRMS/XCAKT
qYXzgu09hwLo3zQjR/sbiQfTOOOSkcOdPg8KqHLxu7GH7RKBuUenYoIznx6Wb7IdYHNg0ZXmiUr9
QhSig1NV6lRlmnoevgNE+Bfn1HwgM1jXIm/SeD0Jfl5DesROBvtVzzeiwwb6pHhiZ9MhAlzxlasE
EjaJJ17qUNp+WZQc+ILmfemcnO/FgRK1hubN0iLqEsHHGugUGqKXP6DmDDSCrlAQxGNTAyM1ijmc
/rcwAw7AjHTv37ZqPXGUP1J2Ye+So8U89GQn/zyFR6+vPTlJ4twZ56caUZTD4D3hMCrgTk1R1U3B
/YV3dNMxjmGemirsSXxv02nGmiGbJQkhH1XMm9Gi9LiGvC4SRJw8nzXI/UnzhTYP4eFqnprbrI0A
smei32AuTDjY4oc2N96Cv6sxCVZGKklBfLN9SDivodqq2T2l2tBocr4GUaCSrJrilYsSiuaw0NWi
WAVuoVJ7Ip3B/Utawr6bKea93AVpT4eejwayuBV62NZNQTHJ+qe+WfTCfjhdmSJS1oAozoevQ4Wg
Wimmvxaj7fqhfiPJl6j1zMoSozpev9EuY6WiUVliTLUGaopWQNutyytQWeDGc0DTBcDvnB4z0dSs
eK1MWF6Ti8Z5gubFvSkQnaHsU29cnr7BpeEa458WmpPRRnrncXCbhSy4qpPkfeNzl2M1VnpUloHk
tCieOwBDjfa3AHTR9bLB6eaKkCRqdgqqQ8SX1EcL0kqs2MaeZh1Idp+0YsEirVSGgCH8+PxgrVRx
yHhMkYVYv6ps3ewmHc6IWD7PrQvAfDJ4UGfSdJCd/8fdN6vAFKWT5PSEF4SKDjR04fhsbgXtkpDH
KjTMvR0lNjFRdSWNFp9axdcBZwQtHbfeCkzJZuGlW4PDstpl/5R6k8PnoUT5hCrpVIF4+MvuKl57
LrRb41ndsST57zhDSm1UhAACZMFosjwbTVIgaxWbq56MIJ0zUh/kzSc7JxX1hDUfQLBK6eTVxQIK
YLTyr8doVELG+/sIvcllQLxGHcIfH0HnYndMlP+GfiDaLoWIKnWUTb5owjki5BQeEdHGBBVHKoIL
WqYM0uEhOpyVudx7AsXf9ANDgm663/5WJ0My+AwhWh+4bT4/qlOtKeSDl0B7JkNgzPP13amu2bHm
MEHzXbuXZIbfs9xDbm08829Xe7CDIj+cgbfsnO0qLH15TaKXN+PX04KjlmOCR4zTonfFbcvaMSEu
NnftmRWNx/EI3DqeQ0dRC1KGvMVfzwsShtwTPax4JZ72p3cUruKsyXG2yBb4Ihw4Fcl22AqqMNL1
Pe3Xchll4l0sSbgIWiFSWslzo0OZNmMNAE6jKp0T+4osmEJ4jIHvj4dW2oQZfYGBZ+j2FsVW1yjJ
AcUVD9fbzt+2GLm3hGFZ6EcTXMniPM2DxJyODuxGUGqFNM7gw8rcVDD+AD+datgxXsY/xsiU6XTt
Bnfqmy39FHWZGolPCqZc+nQumtHCV7Ot7ViRNZB3X4xQ+GlBRZfThxeInLiPv1I/6Tx5ozIp2vU/
v943R1yRgWm42XsIVbk1IE4MIPzrFAcNzTDgaIFuShNNCOCpFZ7M4RlGjDIa8QPicJLiRnPJxyUA
96jdMIapeKP823kf745oEMdIhuNioNRuxWSyjb47A5rsSn8YyjBoUSsw8w5pvRRf3jCGBWbN92+r
9lVFPtS/JwCN2ddYIGqwWi1pDw8lYOYN9PaOAF7ZcO3EjKT4EE6oU+DzM2vcJUJtyMS1m8SaC+1D
bpWOG+LFJgo8vFwDV03OBiocqw/pSy8aY3d6+NdPBCWXZ/uBJI4nrqKWOlNcLNmOSh1cyypM78aM
EjUiPEjjbnbojg8CWX9v4/5+TfJxk/LqxatdNdgMicmp64Zjw9mfCY66LeM+sYIz7JM5z3mpGvJc
ZRYTPByQ1WQx9b0kidDleBEP59xz4ot5zbeoFT5NPO0XZvDZTuTbF2/ZPfRkPIYnYlvStKRPWlZt
BE0/+UUDJXuO7yjRvxkmjaqAhQCoBv3OtWalvND2DfcmzLDpKBkdgTT7wIti5NHUIC9xksqGXvt5
uAUhF73tRRaHkhCGD2Ml3fHAIQJk/b9rg0YU0d8SvuVKM5QgV7rJ5sWLGfpiyAKljxcRi6P9nuED
9tK/KEaXNZaBxu8KEvy2LqpuHw9OkbYWYKljPqDCEXw6hRqFAm/syIKWOSRDG4AmYxpthPOxvGIK
LsYYzdW5DCpX+AISEDD/UBzKPgbcqD0kQpFMB0ppMxuOaq1F9KcJlGxIXIiGBt8dfLnYAdD3TO5b
5DxL8uW3Afwh2YCqlzwSGrS9eCJ+xuhSalLOIRZGDnovNnu2LH9GcSt7HigIO98pH5zxeYhEIY6Y
NPFQ4blfyqYmG93xPL5n6AnGnRT83dBJzV580hnQrS51+e3ZlFXu2IwmUz6qqENMM7zOk35E1Cd6
kb2BOT7acZ7wkdhrp0Qb105ZmDAnKdOICM7kVwa0zPdqVVJJxkai7CrohgzsogU31Sh/x03i2OrZ
7KYNr8TBejMP6ZWPgy4qRaIhxI3Cr8BwP7eD/sQnIuXzjH4ruxBjfNuQokNcM3JSWLvPfk+lYePF
KsWN968LzhB6Woh4lpWwJfVJ6uH77fJUVgUGW1uLHgKq/6VlCZfmlRfG0Iqpw9zPZnh9BjoMLQH9
7RnCrLPvV31uQ2TpKmgE0bMIAB50sQTvZAv1QtXlcMLspEIfqGQy4AIAOo6rO7IqSGEDIHYv5Hak
uikNS4grfmcn/pYQhz1nHbMiXHlW9qHMh+iz3n9BcEGCqtyW1vwLjEnQ73cZ/miaNVX5jLACcAum
ynbqpxAq4BsZMwMNW5Gf/t8qwpT64C/1o8mZavj7waJODYl6llusLiqfKX/tzc8lgOcpFGig0nBe
3RDb+3e1YTOeU09xxDe1Xx+ZORxh3MLClzaSrTDH7UfFj+w1YCTdVtMv61uscBacFRrrfhbt9PfX
QNhT6ps1QGGVbnzn6teDbWaMo5ySlIzf2j3J6iQSp5t4phn1eJpRYFnnS4dgbCH9feZ4+YoNV/ND
nnDK6fYOwIcUnRByP7XjetjlNTl6zpmo2hvMbZRyCm/dmvCpp5qGQ6OttBa/ODmpIkUoobsttI23
QYS1gjlYB4JLrKt8O9KK4js3T39IaDfJB7njqZu+YmZ034rYWCbID5eMLHyOFlrfNOEO1n0mjf2w
1qeW6OpZAcuIpvEX1+8yOoLTcdLUDLt9EUB4yL94+wX0Y6XFhFmN4APZXNp81oQroihU3pcMKNX2
YYWSCGRgAltPwW0tORMwv8mx07N3r/Z/NrgPdqbclAJyYUQ2CYZgbH7DSUxsawNfVIwEbQ746+sH
bvXiSrxKkHwNGrA5sRof/YMylDblZmlE57XmIYa1YZ8KLK3zqyZVvRxG+sQkz+2UYwPJ5XH9nQEC
3m5iYtm9ipl/7ULybjoRCfllqY17BwgFQlt6qrgUBkwfLWOckMQ1GPPrHc4HpMmq1GMpaSa+oyOG
m6vucYmbtTAuKx+sYqHgce0gbeAayRtRuFMuWk68NlyZeGrPIVIuFCaweJZ8MBT64q/bODOajPf1
C8hbZfZgWd7ahb3GUu0r4ghghDnb9B+j9/2lgSGFQT95C9W1Skdo9x8cxCZFYQCn2nmBH3hs5brU
MJCtfQZEBu5H2ZjmoHb8ygQeCw0Pkz9m4fFtd7PuYa4jpdwkgMXSK5aITLZkpOSht4FSNnuR0zDH
s5Nr7AUe/E/O3Nhg/kFgW2laV63Qi+TB8k/NKIQXYYsW7OVRbRNBJ1exHF8Q3CJyxoVu8FwGHDMz
Rs9t3ubj7pRsoB+TQPMBPl2AFrGelGYDIe6oeSxTr3DmTQ9OR5JhhHR7pZLBJJm1vkWQf2TqSRgh
vZXn2Th9Fh4W9zAtBGEEQ5/95pmrsCVGIw2VoBGHKKO1F3Q2YmSv8ls2VCLHQzM05uTBYJU0ROqe
xKnpyU17Tw6xO98N4UebcdU00rHC2pZnILC1GR60Ys40lMEGStRxs8JSJdZ885QfXw+SsUPyE39n
KHGGEgwQEyGWuDz3UBdmSGPuyYcZdwM8Pg+SqPHVc5TCpInL4syqrHdHomS6uzKwhNxRB9lXWuyi
EviowT74fl8AD87OAFz/xjlNJa5UdJDtO8y5BaQ9DBEMIv/dGcc1GQfD0bB2cy4ZcVv2AwNWdbLc
PJ3kTQfhVOsWmZ02aNezJWBSm9Lo2vTE5G+7H5+gsPZjmFTFOEHMh4GFiljefpf6GdFGOL5l/PTt
8wA9la6mOLEswELdmoghRMxT9KkdwfjqCntwAeRH8vBNMBpCD28OyizSRTgxL/rcfm2jG4nY7hKO
sH7bgk06zRng1H7uDnYm/KFSe9AjlmjqzwCyCk5kRu9xd6yrJcI5cnDOrb2l0uw7k1qk0DqsKN6x
VHgob74vxFgZk5f2H0YmDYbst/olmRhCDYPewdV8ZUkLM6PdTgZxCQjY3U3v0jSX3tr9g7R3H8kb
gUjVogAzXlQrh6ELIyxj0Smfa8hD9W8F+qT7z625wRGaHBfgHGn3Cmfu5qO4JGLfnWcUkPsI7f78
1tldcEI0dHpSs7cfwFEBYMvfwwYzUDatELtT7zFY3lKjGnbD5VV5wdwWKYRN8YYf37ctQtidJTDc
SyC0ugS0skVkZiVFLyXwVVhACqJUKoxWTE6AjnyZFkz9YcIbzELFeytr9nQiSuCqW2cHbT0B2gX+
P/YdhtPctYTKqKY5d4LB0+ck5JOuTbliYKtCoWXjj5SegmmmQWMd1+lteqbiEw/7vlY03908ylXD
ymLKr03jvAejU7NMFIfZGPQAHNmcxEL+8KDE7TPpoyVFez3nZUexFRlR07XEnj/Jd8x4k27imIIl
7x9LoUR20yCK0upmlZrxeGV826AJ5o+mY32ZCTZAMT3HddYdZ0M4mxnHqCAwkShZVdBqEfRLde3X
Jei3fygEopmx20/XXBQiSELYWCGO7wzJic4NInL/aJeCBQnOnMIyVdsZzvrV0h4LXQOzdYfAK+0L
gbJKmxwkuI6Td1YUaPw3ahdjrpyYznUPPJL5Zp0irGob02PsETl6zdo45r7NxeDBdvkIm3x0aqlI
LcLU44imPM3mfIjBzLiWuNesJrqUfgOPpOhPJ2hzReopy8YTHkrhZBOw7mEc+IVQet4+5kMcGZf8
nVtUcfM3zUkzCMp5mGj8b7nn6z0A9jwV3XgjmqjntbGGjfx0Z0c8448wJ9yqYY+LgRyNy0FDeBfE
fq7mCKagqZok9NnUbd5Li7my3kI1b2qzxKC7FPwqUQKb9ALXW3QZxve1MpWjr4oF3zMtvxMNAEBk
gX3PMJKp0MC4Ha4CipSmuiUycR997Bm+Yzj54yGtT4rEa/cLVrmHQz/+U/Uwyd0azMdoOfTjIXLb
cp3t0UUQjfU8M8GRvI/EWLDT8Xp+czOL8HPk/u6XzcDdV5K3cILx9SNprfuYmQQU/9BtSY1CPjQn
zwdYJiNW3H7QUcQWNDrjD5ytDj+UYcNpkLW1rqMLWNSxppAnqycB+z4kZ7Yn/s0ZBkyFIhbfv40a
k/4aGhRzL2LAx0VdTyQnDnIWuMCBZdWALLlfkOJlULOFdqutTJJ8vc7dtKMtA27o4jrKJbwWjywf
e5Hw3vVvirV+GIdfhwzwEJNdftN+QjIK4z8Bz+33hwahBp6+FqZwXrcAPM1sq50oC1fgnhEfh0VT
RWR4sozLNGoJ/IVoT0vPepa8eeHY+Z46t2jTpq0peDDEYDrOrO+o/I1ke4fGAkQdXoU9wOsHjVyv
aMBX03+sYf66IuA6+3XSx2vc7Te/zPQezXK2yWSPjBIPuRUzhFTcnYhBJ469o6EV0Mm+rFEzOSvp
YUe5NXWjwva0B6kGC15YbWZXbotPvgJ0P2J7pqc4nz3Cy1IKRkLRFwHPnGC2KbUjfYz6vhz6mvlm
W7EmHCCofiZnqn9TvNb6k9yPc9oV4GB02JMjKG6VFR6moBxG6vAnzJ1N/PqbJyJmi9WU+rpx++h2
X7gcSugtfaaOvtyyrw7QwHXA/Eb0zSGySVXiUMM+rywfu/SmTp2OxlggWKKeMunMshta7+bEqHr7
yBybEGCAe3jEt8kQ6/9L2eU8rJ0ETYBZky9FN4MDpCCPkiPZ1ttM5hiGJykz1yOULufjKznmt6w3
Nm7Hr3pvDaR5Lq3kRAuAGwGE9+Te3IE3Cdv9BuxOxglrLgxvaBz/136WcVoMihAx4QNjEGCCAMm/
jceVWzNmJhK0/MW5jl148lWCPNA36nY80z44BqCBWR8lsbJ/FNGqlGSgr414PzuR08rKEjKmK79j
kMpnwqDBtWjF1QoqKYKKPG7KHYIdM7NXS5D8TwyZ+OmcfDOXDLUuJYHu6DGX9GamL6V1eYZu1TsC
5zl2DXj6qFRbpDacx77n3DTkY8SoyAwOeSP9d5fdQfYc54/Segz+V1LWkZOZWbE1iTJrIy65HvmO
gtSIP8izIDrHA4xPXyNYwG2zyqSKDI/eU/Xj7DdvanzL1FpwOb5ap0icAPkJY1gnATEgvh5DO+zG
SQx7nV07/hSoixpcFTrWu+oVWi8qH0svbo2U2VgK/GtFmA/SqyOR+fMVQadHHds4VgSMm7/Irds0
vK9uao2EniIfJN0x+0KBh4Io+N+1HJCRvmLqYPj2SV2zxZzrrLWXEBLkuEI56u4p9QxT6o0eERcm
RULmH6qXGSYvDgEUQJOlVraWjjmZP7l9J3Zi+/akbA1Gvm53e+j/1UA7p4pb7gV49L4Paadfb7Wb
KGn7wPaRQ+v/Ke3YIRfiKr5VkJR5F5NRhzQkKe8dBnzHNGfEhrngLYpVOP5MQmUQyMyNI7pUPOwz
eBapE+u1fiT8TTRGKZ6TzofUw8p0PhNnHJGx4j63ESWS2dSaazgNcVG1wvqkG/j1O3fy6mWAz/em
3vILKvapHZh9WPGaTrPKKHlkPjtspt/Rx5JONPC8yqG8m/TgJvfIBH7aVQZwFYEm3/6K4eoTs32c
Qe8KqihF3pN2F6sZVOcT0ECZP3p8x1jo9ZAHzb65pnxs2/HID+Qu8LjXl1HIi7h2rGATu2b5Js3w
LMrEnscNz1STFTAvRdSK+WyBjF4BS+nFFwMSG6SNp1cB5tjELkz1MiyPpoQMjTVDhLBHIj0Zzbr8
s5EOOiIdB5oAFSxWQLiQ5Kc45o63aFqiG29+zp7sAfg7kLO+gAG9rpWVw0fVfLFD7JSsxox4jOPZ
+LEqk4CxwHBuA4EFniun4Jfvx+dObiIUbwxbyEef48O4y19R4ZY8IBmW290HUQgNMMlODPfeZFCP
cPp0RQOmihtF0Dm1krnO2GfqtzYkUyB90xWkCO6MJHeHYHsppIIgFSyX2jn7U4OiUZ7DujAUxV8X
Vy7aZGGSEV2ydOrb3cvCfeV+/l/PCHysFpUqsCBDJe4LVjw0UvMt7+9eVsPi+t/+UqAjsMErmhde
HXUFaAyWbP9OVFav2KeOVjsfkBkcmjOE+UkuQ8mbW91MeRfXaeogO0EwE0dY7AxE2wrj7QGE4vlj
x5b89UJUcOCKHg9ApQMVUV1Xm0bALkv4ZH+ji5BlBojGrLzgILL+wBP/64JBoWhdut2dKXBEolwS
nuUC4GTiss7e+ypTKb3AbtrDmT+FyksvR3WOK1jiM7FS6i8lLt+Htm8/NoA+LAeoH8Gdj5NWo44a
oTJ0BCx3wX98qLdlUkLQBIZWZca1Y4U09ewo4pJ8Zxrn99+ZqJwgVIqeUaWJlPRsJ4jnOdg20nwA
QbenKlxKWyuxjzlphplJ2bMpJ9jX9Z+FEIEQ7R6UnL4MSFnbV5TMII4dQXnnBit7l/Lw+5WxYGqe
M6mQm+BZ+ZWRXMLMtNweasM4G0wQnmBLW1FXttJZob06Rozh9G+Ojb8gHwKxdjVLwBzB8A4e1VFy
ohwXn2vB7hdckBu7p9YdudFZuDLO7Sn1E2rLr2aPuavvvHWgy8Oq5BHRcJ9Xr26+fZaK4aLzqLmh
vKPoalX5uezSKKlmXnR2tzk4LqaLmGw98N576oWpMF+VjJOe3YdzCyjTC4vBdCxXMGxYOsEF/45f
j/tuUnWldA0ukC88XYBKbLXTnetl8C5Q3QChXM5rd5R1aJb6HCjvT12wg3x73f1WlThN5Jvj5hXY
9z7EPF6rEWOBFZ2ub0DTnGY7WB0S74BFGYOBgnVzCgl/FqNAJf96ByNltfdLMyvLWOl9nunnWtB1
knmiHoLhBT+ixFns1QLD/J+w8CI3Ct1ZN+1BE5lixImxFlN5tMwMNjxqEHEcPL2fMcQdI94C5wp0
thFPYYlQqKM9JrO5wW1/DBFc0v2W4ihiu3R0AHGByjxMEMw5KeFOdR3SzUgLD+QSuvIdTwAOWsI2
ogn0i2JCBun3smUq5Exwc3gXAvNE5yGVHX62dqyrX4KN540f5Gz+1hNVpxH3D7Nz+zGdK9G2DlS4
uPdaUf7MVFxPrlO0fvMozuX+/71dmtfQm8/A9w40pk05on/AzGaY+ChQdNAIVfPMyhIq+IbgVfZu
u1gIUoK/5IhgMouO05fP+GielOVASdHxj7lyQWjUS+qIat7hGkwuXWf8MQKzA99fq3jTD4vHVzPh
pamS/AK67u67TvOs8r7ygEE5i15JE2ZhH5p5ImjvDsassEJjm884ldtQjvbRI5gOdXqzvrjsszqX
OgoBIu48oDFIUe71KfxU3lir+rGQl4PZSSHnLK1FJPcNGgMIwM0W8SxbgxRuvg8VkZN46L/SvwAx
ddTFV5F0Kddg9bcpPJjGbaXHEmjJ1Ca/gqtyelrRtvzQ8xWvjHSnhFPLkNYu8izRuZjCGe4tqlNP
bl/AR/a1Xj5l37kpmP/pjjXTSUjjn4MJQ2sCsXDc7I3CbNiwazBTxvUOT4xuMcLs5hUSjQ9AAsYL
CBtaeHUUPDMXlq6Z8CZSMaXY1WirNJVnI/nch4i2qDFpBbdXBxQsjLgQhXJlZEmh+PHMlTHj6tbL
JWgy77gYJ11N3F1J0WNHzm6nyzAbe9KvykMzY+yYxPQ20Dd6nSAnDPL9DDm0ku5UVrNB/qavSf6p
rIexqrBD3ARwOYf4eedTHT90d7NVRwbysvnlcVb42UmLXwJbsTOe4K/evvLg8lAoaqw8mI85MDww
9w22i2DjJVpq1zL84bgkkE7UW4vlAu8eNXdqgAQGjoxGSV5HI3kkkPDC/NkJaZS51DQGY05Q/JXP
NSqfhF4xD5b1AGycLNoc2oo2KQbq0fh4mOY6gpLemH1nswGzaSkrT80B5Uw+L0EG9TmgIZtvj6da
8qhhFaaOxLtDZWd2lZcBHhR8pid8d+v2b6hGPO0cXlRTef+biwcaABBTsdiOaCOTea/N1uO5P+m1
xwxVePNQ9wYKP0xKpsReeUY1rGYzLEh3LeC/WGnCjknRpXVGzEXH1TC2T6lvATeHE5+buASiKP4i
ZOh3VyCOW242de+vJz9GGDYVdzVCylaluL1JT12J35YmPwy9wQjXAkCvZajhTG4X6wgFyW2K+JO2
8aqXdZNHQDkWfTCjCLMFXl1GLhnFaXmS5TrOvWg01/ztYtL05sjDHnD66tv9Zql+sspvHXiEqzAy
BonMpBm8qkMjHuH7uVWKeeR55vNGf8XTWaqHPaAA+g54A61bQ6g3r4+dt7QFEtSBxZQwlC8JtTIV
NLeZfU/grgZ7UX7ZyXtOe/3Kd0M7C2i8CH+hG1X+mMS5PXbcY0MrdozlTAfiuRkbCtQTTHdVrtxD
Vgog36GmXeQGqtRYm5ELVsSWc4Qdkxx97cO+MHT4f80mSnWkj5zvstNvYGH1Qz3ADDJSv7/PVipB
1/JkVjA6AlAQbN1tq2Gnkc9F2Rr9a6BAAhdFt1gCbQK8vgWLVl7E5TXcwwajjez0DUljoBB5V01Q
SMnJvxAPA1egcm3QX9kiJ9JofqaCSDXyEx9eYWZ9xsKedUn4tPoklnQDIMcKwDBWhI3UH+YZJTaD
qInwKmWqAoxdQdfBxTSPxr/3IuKRgZXYvYdTsICEi+Nssg9sUvhFV1rHbk0LutMXexF7rRjB8Tav
0VlMnymI59/gfB+C2q1ZQhprVbYXyNeYncvJA6XxHj+c2kz0kY3VOyYcide72nH6GHTz89j+jGrr
VhrzkWlQrwpmkQNghTLQcx5xZy2Y1UtXfTdOvj8pNzFqJzSpjUgSnk18LXyw0jNmbnCsb7ut1px6
Hwkn93B6jlcJKs82xFQvnKky5xaplOjLJvq0HVDlVrJpVGgtO0ej/fqoygPxvLHj+LyWRN/r6iwh
MsZ+1rVzzpRdPF+2Rha5lPKY4dTyWumKOt1bVzn0HmWIvtyCtfx14Boj8wZ5TC/ORDpsqm2AYj6f
vouLEx17vl9JKpjzP8QkmEABCJkkegfcZ8NERPp1xRVGhVWlCaBweJTSTCA4v/sTseRyabJ0aNbJ
ZGtXaS+YCKq2cBJmJyBIMmMUs7Un45kaPnf9qb+psEZs4jBfivo9Tb1eBmUCGyeKNI1jkdsHTjA0
oFExMShrfXF6eIKMhjV98yuZB7tFC+MxG0W43syABoZ1+6txr1+xMbLbEUCwetOatVwiM3mvWD55
rGOkaU6p2/xWAE1WY0Jpbig/8CIDm5wikPY71xW49WAbYL0HIU318aOMNaJYAaUIrqkcnzwN4R69
Qh9B/hGcOkPFaUdFaqDpL7p4Qf9spsQihAs9DsVyrudKgJOzYeUNb7vciFtA7ps/aqbJkupKT0w4
ACjSVoKe95vwbj0ii4m5zfOsDXUt/Ath7TrPQ4bw0spNWDAYnHMwC0pjIuA/y1PwlAtPxIF0Txv4
JALMIyibnxPRUKhXYYOVO5mQk/4rnsJMlMZAXEQrGRwtgCN2cSWB8QkgDVmXqskcD5iuQ4pq+rfg
Y3Z0KG0GGkxTG0nPuwivLz5QLKqG17Qpdoee+S359k6K1O6zViRQSgh5C9b4JKIt9CX1xDM2sJup
6aPXJjbXUinP/v1Jh9Wixpu2q0j3U/ytYGUE89P4gPp2CZltPC/5SC04UwCelY/D1SUEOW9Rc36K
a8slE0lejiCmPmpJ/yrtnTHiIg8mQ7HqdmmiM6T4dyfeQo9qwYpgpDvSbDGCJuG7V6TkY4T1w7/S
JRJ9dwAov5LA6ei4BMes2OYtAN/AXGjndTr4t+FK+qsOdq6pMiUPGsf5xl5m2G9PdeFT/PDn14Ox
GwQOJeBY+gjMVkVtYVt8R64sf6/ZI4kkuSKuED0eeWM5h0/awr5bhwhZ1UxkTgm86CCQiZNo5cQ1
blwuhHMHpgdFtb9COpHpw8NwMHHENUa/PmMDj/hMP30VgM9+7hSVjQUS8bTnGw6QHHXc9kXezXOO
8tG9NHhZ2CCHL80gVGmdLwCtrBVZTSvUQuSynRi9O56EzaQ+3laZjyGCAE/Os7j/2iJ/WrwOuBAw
yeocz5jueoaXjKTyhE7tF6+F6k8mwSTJLfx2l4DOuW6nCIZSBqVOvQIQ6QKuy3acBv4rr/a2fnr6
LoXK7hToRygvVJpYA+3huV9CdS6QnpajLeYcTikBQKo5KVuIO9Zfs1fPvihbo5gbQwF1DmX7j5Va
z0TRzSbeTJNXrOBzndeJMb46qoE+qRI789WPfrQ4bfHFuBK+FqzvbTn1fnab6/j10jmWxTlhjILZ
dklaVMRyvP0f9lDSzjtnSn6GYnipg+Wrdk2n4igy/25bQtJO3pcnfu/E9GKoMSzcNhUSdIOqgiEA
C8KouSSXmCOsMs/1bIGVqLLbOVSPmnnuHXi5oY3KXf8LsaHvax5sVaIGsLMo2GKJ/IkpIOaqQdya
XOzK2DM1LPTFtAzFh9gW0bZx9sDMIiQiS6VzuI41kUKSpsnK8++Elkyg8cPK0ddE8QJCpyg42w7c
HgZkCSa3gDSsqznMW2Ptedk8DZSecpkClyEUPtllrVkVIk5eGWDIoY9d4m443tmT6GyZ5yAQgEeh
EBPTIHbrNbcwZIYC0IOM74l0fDXO8NcBwC68lEzcofl4SASuVeJWpmwBY8fdf/GpZo+KZMCbQ1RT
AjFs4LceYbH60a5vdAnbKlDMBE6eDQlIBUuMk7Mg7xb/DE5fsU7pCWW2OD4BAIklF0KCsdjUXhRi
RvbzfRUmLnA5v4VEFdHGf9vA1Kz4e0/j09SkzDvwxdHcw0F6Pg9bK6qaRtr1j3Phwde4T0ME0Di5
o2LvvsX77gsnwla5W0ufSz2l9TWAIgb+Abl9M4o2XQwr54GmCC4J461a6D5/wgfTSr+3w8/l1xHY
T+l8Dhn9bNvTLZis4wqrhB3IPVEKdpTDCIvMP41CwwnmnRFVWpPJfcAezogEC7U9UZsXReREaiGH
4YA9EwX03hNPprNh81XiI5QUIo9FWwf/sytjUPukLvaUJdnPjnwwa88f7sfpvj4lP2reZHCQWN5I
odEBq4vGuwOzGf+GNqPPjCux0s8tJapaJuJM/4Ks18kJ3/Hl8aZvBAT3+eoPuqgrS9OW+o5rVsTF
WGa5essGzcsgjX7HntT8GK7+ZEehIHqyowPRfxnCgKSpzO5oAJpDQOAYq3mHJUCUNGHS4vArPn51
z/bYsi0S5GieVMGX7JO8R/q07nKwa8qZQ8fjGeHPLKrBX6urw7ISt9jMtRtAwMMsAnvXVf4GsyRq
kIszV6miFrGEL0AqT1qx8KcOkM+ZJ4wIghbEKN/YKTa+DkHlEJ1k2YXgxi+wj8zJcqnXcb7s7s58
0pRPF+vC2vXSLwJmQR+9iQTLNir4WIR+nhbUHtXw7v2TpGdw3qwWwVWR4jebINMrsHm3XQx8l9ax
t1hwkspERcrHvLhkxvqy0HA9i8or0xzCOOGs8DAwcJyYoEWcRHXQgxrODVnAJnDsQaAWubBC23Ov
50kKwUldsiq+WmJWdlio2GhYX6NQNIfI1q2HL27/6QdLts76cxJlVksWJc+e9sM0ABligaX5la3y
jSCWRoZZgBCnwucLPe6kg1XZkBXwZsDlhg9jRp5FNkBo9yTuWOICkXXYVYLdHyb1Lr4N6wFVhs8u
liPSvtHzmhq1w+FTI+J9/dNT6CIQWPLVe964cf4n1ALSxI/L3/xcSasQ1ihE3enCfVcK5HYh+bDz
QPjpkVlSxXoPo4D1ymN7uZwCWAzsRnZsMf8ft+HhVIAhL1hJK8KRBOpN1RkWuHnTJlbcX3dsYD9R
u7G2WzNPIY/flXDy/KIZAVFm50/WzLKIadlf2r7AksywX4uje0gJm7nfsJjyP0PgUtfs3eWYQhfV
TsLF4aIW8nd/kRK2TPJ9WtKQwTHim+F1cG9rYGAENOYfqyAhznYtUw4428NQ43n/NzNjBYM25i0X
B/MqMdZjZ6BbciiBe89iIPW6sM1laY3JZzn8fkvlLPiPkSA9cIA3wYuGLE+4n6xnIdi2PqZovBvj
gBjL4ZCNqL2Z9pjbwVYQ9rW/cV+DbhN9d3fH+pVHcRrxFHJvkXBc9OPMJ66KPQbWl52kSrtVBvi8
8dlV8LfMpMeS39HOirM/KccDFEoa6GAD7AUEpDYUHHZgdIgARY6Gdnj4H6Zd9R7FiOZOZQlYFLR/
YlDhDaGZP4VlbX0e/HG9TLEmlybAVZDFoSls7ijVt0pWUXA+vTAtTZQR97GzcDlb8jz35TExXklI
zAw/Jxkd/1WylZsQIU7jzMuz82mK96JdLjaeCLC3F5s6PUB8VFMSQKjVBEFD6ilwQfUaOz4k0FyT
kEQ97aOzOlcrtmeP40TMo9BoXuwQjyqki8v0WoGyqaLRJriIk9FLASZQDjKf26bZol232kmufmQd
Paf9V0qYXDhE4NFcqNYz2eQiQTiXJPd4qrtDd29ZwXgJNwiD2KtRODDbCshitjmhbVkvojKHFW4f
vPdZhMEvMbyA3XESqKgP3UQ3i7eUWZBX7l03lM2kU9cE7q/oXCL51mnizLguPBH/ltvAs+VML+43
+22kuAfDqxijCUhGi41/U9PIIAwecvVNFExd7FNmLCzDHRoJu4fU/lAwi9uJxL/S7YvCfWwMXSH2
9XJelPdkFn25HvNGzej4MpcdRBn68E36j/u8vzPTlJCxCRvAmP+zKatVlWuL6yS44KeO6NRTTSen
EbjpTODqW0nv69CJCNBWSD7NySE3yI4JfptQ863qVRHNyvy6ONfZxgp4XLObuIb4HnSz2hrrDe/J
Rp+vCvg7G4QCWbXiVnHaUvkc5uH6dEKjqvBo+C2m2GLSny4Znhq8fu1zVTJfUhqV9y9oQGrhV+JL
6FcekTOIj1rJdEYwx77fzXpoB/oX/2XZIdQCU9IYN1zPjEh5SpJmtzsmZeUFdtIItovR1VPD6hbu
y8ULJLIht/Sk1A34j8QMCnxY9deP60K1Yopmw2V1onohN74AwsprohHNbZOoG9nDLLT/Uch3iKAY
CZZAeChd0oiAq0/atTZ+suWsL9huODenJIymQrQmd4APVQSeCcCf592aZQiGxBPqxzrdRCg860fe
C/80HcUAkpvm1fdidMr2C0TWkPX8FNLMqtR7u7Z3/VJOIoo3mx1dhKL1kCj9EIh2A7BBXPJ7xwvK
WD8cjlwAp1vB5Rk17E72L4g0yxIM13JcjcO+Sz1gNyUEmk0J40MtIjxcVprFAtY+Pb4fuRyecyqs
iu49FK4arZaAHdGkAV+lrPJJD0U4qXu/HD3/+KA4JKTBkHdUgzXJt8+a7QgI9/6rV9PtzEZjT4Wl
fFs0EWWx8qm4bqzIboSInp4CwOJVHHv0Xvjz/WfhTO5mNxw+9bmg/vm+RfEAnz50/tKGoQPJXrUH
0n8DlerBVKWQvc8gignT9AzNmrx49Hrq+2K+D1aFp7eosaD/H+SjSimkIfMDjvfeuZGOB4ID5I5z
+KmdQH+7V4/bPtEVF0oejmMRJOV+0wZoB9+eUNxEA8xy5diuTRkIR2ZtsfwZeqsMXOHR2WQ8TpNW
q+URFlewFQpWgWdABXtChoZStzyFMYceYE9JBkYhFv2XJ5EdiB7vzy9TjsZQS+9BX7e7EsxsSST1
H1N5443AvPdQR/y6P65hyqr6p/b1u6+wQgNhOwx5rL5XNJKlu9du7vmtgJJUORQqr89qe6s0pfvd
fut96vMjRskYGNY4UwKZqzF32YTnxj8WXoZpgR0mQ9+l8gRNzfKlXnUBWsi3+DDCRWwN0IIdoMex
kLdquT0Rp4vwV4QRt3PfXNpFA4vSuhaBat9pFuZKkIFpAnnaJNrgFbMrkq2QYoHr95xEhGBtICJT
OvQWWM76U2ELdFuFJkdvBARzdiCKR8QuvKdfUlW1GTeklLrBI0Fx6Rhc4APf1THoHGOndMyqCerh
rJuwLt/pvy8TBowizh3q/VcLsORjL+/2xhBEEFeZRSdXQMcrzLLtzXV3nnBIZ3ExcvYUJn9sDPGq
xtTYXHuZG9mFNnuxObHvItZiXLZCzjYkxihRcCeRfC91tfavedM0BauLmxebXMZ53kk5DK88NCrH
jTiSF8R8dgFQqU/nE2eU+uTGG8eZJkI6xt3VjjBMYfx1w1//FRygCxlKhyLTz9ojZ28edZEeFeV7
/OAPk/lRP1QeYTRK6LxHjRRTFxFKnSHKRph7W9zpktLYC2E8DY+iZppHql6OypobqBkiRpLLTqIu
EIIGRRpIPFMhjunQ29QbMkGHa7FHBQGsxrze1WQfMZoMsb0cEkVd5GvRezkT5SYVaeS0zf0eZQHh
JGdm9xbkD1O/zoMoyUmMoEbc7MooESD5sEzpnz7Kn4FhqS189SQopvte2eLRQN6S5eHHL8iE+UVu
E7HBIzno9mopkcNZ3HeqyNYITo9YO7irmaTZv2cuJQGEQu+l2y7d7qvENTggmuyaK1Is3c/F4WrO
xya3wUq8es3nxvo1H0ohCNtmbDV1mcdelVL+zFgxgjeHfAbGcgpUQMGMnsIT2EZA3dbPB/TbtxTD
6BMPy262KVDlt9RHZndBk5JInqcDN2koGYE54MrGVW3G/T/OKUH+k0IB74g0ySDw+lHoB8hB16CZ
uLKLilcqMnZ10Ynd7DKtxHttJviVQWxmIr9BlvZtTwt+cWtwgyOCuG2wEc6brQ2K0nBN71ZsNDm3
k+BU5LbxNQh2rIMy55RKsJ2qUEWOujF0MXZdEdVF75GHzkUHq1iWOxGkXUacGqmB5z9ywrwydPf5
Z7RenBr+LwDI6kR7amP5z757e5JCyOD1JfAqif40JRfW4fymb8mpnhf0BYWRu5kU4Cl33u5l0crD
MipnqGGCSGpIZc0o+H1JcLRKsHsZPMtAsfc5d9QeY+pAbhCsnLXfZzAnwNFDYpY32AZPqP2IFip5
ltaVVsC4A7DpwxJ4L7yHMpXWY/8SrulhQT5rifLTPnmSgdwZZiUrnaYrUDguKwhTtmyEoDlqR3eJ
No1/lx4J1z/RaCx9LDNcbJB/889fw9MuYipTuAnIftR+5PvygpZiR/+DyepHbmu1PA6metl39FR3
6WHp/uDz0dx1INu8zKOGl6VHFAOEse1yoxI2Qporfva22NEytwvnxkUG/DNkmnRVjlwrem1/7sN5
DnIftO4T+CumUbGvFqIW4UTMsOHz2qls3s2iBgVlk1Rrr95xBQQTbq2M2S+emVKI0VysMlEJss5p
fOe0qWqflflOlLs4gS4UYLOQ1NeaSo0AdPn3pj6evDtP9xh5FTwgGIgWDH/GHvG3E4qwkP6Zl/o9
gIBX4/uFP6EPQhIbQ/JCHL6jtc6H4EyrdpAWx2fv4hV6KJuFi/ODgx42Ru1E1GWye+94GrlKDYzf
39y2iH25+EOlDedBZsNxkT+Po6dZH6YeJ5bzEoE+QLfz60Ncnd4CyyXsAqCDsNAPbRYmTCN1r12Y
Y/g+e6TN2T0Brc/aYMQO7sBF0FrUuiYkHkbvKnsr5e9F9qTXXBLTF3Txs58DGdByNHKvpm5glUt+
BUp0woWen6ylvYsNBryT1FwOaTsqhgP0+uHdJzensWZVtluGNPQugFDNdtMVjtElVvWcgeN2JT2l
+4GIw0AMEm+pP5B6Bobp7XIRIoCJWCtygmb2McCTgPyrpTqNQ9tbjAekktJyLwbaKdorLfsf04hD
Bpbzq1f1VVt6iWyPtWhbCDHsFkg0eNnhEPzd9+O8+GTENt8h4wpY5Z5Lg1/IpigQlufVSJeCnca/
PilUcxKHubU5Skzm0h6BMPFhCOwm+zF385v5f+umSXs0cuyzJB45LIdCRlNVv+YNAlvUlTzvJy6n
UFVzuD43QuDO+9U8EqWHVQkGrDxWKp7/g+V7ak3wrEOZy9Ucvjhkr6E3ZY3N8+5B8j1NYWAKKZ1Q
ioM5eySYJ72Uztx2MFYFpdLKpwm5JWg0+eJWRvqZHQ7kN3qeC8hlKNgM71tw4f4ims1LX5Sy5whP
hUsYMg0xlQvE6yTrDN4iAV6BO/KBMflL7ZQnXQZ7XccrHLTbQwzis2Msp6R0QS03Z6HUdB/q8+x2
IyoOJgT6G51lkfSBVzd5zio3AoCFm+s7EFLYbuYzks5cGwClCsoxj7ANe4xMRuQ/pCaa/Mbseld2
Lq+oMc2pv0OpSEnQtcOhK3uaXnYslCpe1c+Bcxzs5iJtTYoM0/2lEPmPoC4hB4mnCVoRaiYAwV3Z
rH392LsXKeAvo/r4eWDpgUnDM6fXb2o2R3ZudN5YmFb6v1cD8HH4lNHpoU7K3WIbgzlBDBkXbrvC
uOHYG+U4MxaY0oIRIOp8DEfn0RquxOsvxoGyP6fJvU+jlg4otYOKoebo16ydx6VX/8uA/ANj+oxc
yTTV9PiKfSJazKafJ3u1cCg6mPQ7T15vOE2OC6RyWTgVSgE6Qtnzp7WbgEEbdmyAK6BMo3NrPX/W
vi0oQsy/8V6moDOSOZmO74EIw3pAZpaukynYaX327GF8D301TDmx9+WUDIOk2bKrjvyQQL2Duy85
A4f3ulWuEQKLmEPVdGYn86y/2cLjlaITPc+58tSJQA97w707cXalwW9h9Fx45621mdZQ5M5pGOvS
a8PB8YvcBjMq+ZOYJeQ4yEJzFmriHJc8cvIXmyqg1HSqN7n6lK4pk4Qd28pTaMhYmkwhjrlgAN7s
GnZAW5m6vopolXpr9tbAB7SX9Do12HlduFyYtL0Aqa6JDj4c3Ir9/33TsZe1MHIpkFJklBc3nAUi
Muj776CRgH+UZcZwM56fFIF/lAnRzkvyekB0lArOCchAsmSkT/vcbeji9JIbV8B8DI0+ogsHpwYe
na+XvJsfjzhmVIkOpT7iKXDLprLvPrxBzqHzHWSog7dZ0uitZjFQvYLLNPCAquw7d4wwzypV83dI
MjsaeGVC27PY7hsHs04kxdty85XS0yS3z/aXXtUgj14RXNmnicki0jVYx2G6WP7MSPs0I1h5wQXn
kb1jwYdOdqe09c6Z9dYzEReLnhwcIl8Ksp91f3gFf5JQuEZcgZG9zTiDaVLukCyfTvGPos176UEQ
FjvQpjIRjuVEZjXT9ANJJzfJg4Ebryy0SNtJ4XXLA0dv2JNrSPMpQW1wR+f+BuunIJvaWG9eZxUc
e4yXpgYFN8vzSDerJGuuPmFoGv5lguNzAH8vHZvC/WPtM7xtkpDqxs4cU+OLG319l6fDgk+GHFWp
GSi+vQYF4NEOXyC5d3/2rEzFKZFw2DoUbjT6dK35FGyZb/TO9hYJHO9iEqrn8LvjM+xvtDl1LMha
fPDtaKx7f8aUU6xCApU50HAGhJh7qNPEicVlRDOBH7g/jKr5Gd3OeQiwIksEPFrP0ppVr5AOBxjb
hdpa6YMsdKGa2iehXP/REdGyiM7B8o4fNAKBwTOIveXg0AHQYtFc/GlS71xwBS0MuptDe8xF9XUf
utgZtp1/yexIWsXfjCri2qbPF4RPa0xgCi35O9ubcNYLZMppinMKktcGI+R2w3RRvAr1lhRMIdwm
5+/nlxhQo4VWrDB/xrTv9A9iJ6RpPrnfwAkJajTOZmgiCfAKAGu3qQpq0AQ1OqL0gGKswM5xyw22
f6DIBk2nS8xoHURjXj3YnHtWlK8cEv4igHJFkosI7xd2M2kdtGDuqjT/vTjlggvk8PM/kb9fJckP
rh4xJq7NQ+ZvPjpP+o0FJFFePKCT00uG3uqWFfmfuAhz6FYmu1xuRHNCCt3IXkSpqGgeIHUEzMTI
Zf996OFBngHpewQprKU89oo4fBlLsbvv76lN5KXByjkZngVJPfNXsg6FnMzNCSWXtXwWbOUecGLF
U2118tvSCWpXR/qxjzRjSGLJSEU5TgdKcg2xIRSi54Yh0U14H0l8RAvsbKEmfK679Mu5sfm6EbMD
TVs/raaePVZhvTTAqqgzyQR94xKpWWdD7jdnnRWW7uQ88YHMrdcjWYTw8FwHbjB/lwpD/PAqSBJI
v/2CrIkSNFe9vtjHJ5B+Qcpxkdl/Stov1cgoQfx1MmiUJgugf+Idz2r9x0dqkygrFuc+AEBBg3v1
1mmGDa2BcUPMXwLhn3jouk7lYgGoINfAUIWTq/A67Ee6/NpcbvCr0PJ1NWfwZOCJB1j6paL2zU2d
fd4q6etO1VkHsj3LJW5ayeBefVT7pnQwlg3MIdpiBK2NhuoVQKdaNxpfYbhUmSpIpNX3yqi7oomn
tjHZMfjc4P99XFuqcd/gteB5CuAXak8RX1bdD3D9H/kGSxjpsRSJ3DM7kBj9xGpcGLdyxdciUiWn
SSRU0iwgQxmU+zKnbx5UQ3QRmr5orwQCAAdWTFeD2xwx2XhTHtbPEnSCiWioUEcOK15vliTF/cKj
FjNgeOOMgeEEbmYSGl+7DBcIzBByNM0isZXWZoQ3OBzn/aF/U5u/21flLXm/Gu+CHy6qfT81oSG8
vgxHZFR8dDL399Qbc9n+AzLJvzn/xYxEdQKYpVBnYJ/cHMvgV9lhNG66OnbRAvZMUi5wKQ3nTjP0
gouDYbIhCALt9Z1ghmS6oNQUxZG8AJDsh5UbADwygo0i0F4GKxs8kGY4IcxbIOOZW4MErgmxRyyo
WReRR5r75ffsMILBbRLdWbvWmV1z7+/usyZCc8i2v0KGyVo9/pVpC+P2AYsUoj92Wcxt6i4f6Z9L
sXIQs7RTszK+vwi56rFwOVNM6UF5NFZG/Cv1YkWc8w7LahteLblWqoBT0YNXxmp+TpCYInrl4s8t
Ht3NYu/cWlROLK8eT31elUPOe0jhsyQFNBmD7AWiKwH+C+4UVCxTqrqjhofxoiSHxvxacrOuuPLF
G/yE3GKLE9BqSzLbdylVPTcbPwE9CgGm16PvIAf65DLdO+t9WFd2GcZLsjJEcKb2Q7uQlZZp8FZP
DFGSWYfwFQV9n0fxq98PtJRDgLx/kCrgvdTayLggVMSUsgI7qe0lpj4gTKH9lbU/T73rJ0XAn4/I
dWQ8UkwqgkD7bW0YZRijW6fPj7E/BG9POKrwJrnsGNMeY9XYzOurtFW3hi4xoUFM/FELhnUGyS0T
OYUrLF4j2a6kzYerY26+LCCf5srbW18PV2fR8n24tbmoRwsuAiRql9edw1m1PFFKuFdw7Kt0szGm
Nn/0afkwurvlY6eIceVi56r9S9j0KxNtMPZES4IEf3DGpvl6uHP7gB7ocss8D8JIPx+VGiMVwiBP
NBnxYkPxvcEdgf8JpYOqaapGo6RmI/2FhZaKl8hGw0+vrbu//iSXGBXj/6SdEQNgWe7gu2y7Mgg1
O1JRmgzFL9k5blkrfaOw5ev9Tl0htuLZHpHKSJ7IYMpEmf7lahimN0sqZv8VrVDlIbLtUlsU6fF9
sX6ciXTCiShrhVt81rs2UryNOH5BF+IF9FuF3/SC3VHskH+rKX5ywmjhIgsWm24b1UEcDdzM2VCE
a1uI11CzIG0e+o67NF1COUCkLoJAlw6PcxCbF22kL4XHdCSan41fqaZ/3Bdsk844+mg7Uw6Pos/M
1emkBwrEd5EYI8QaLSgxSU07cIDBPCzGK5sL2aqLnVirveX4TpTCJS+MKe/S/7/lfQhMMsPwzHs3
nw3C89FxiZqqcPxa3Dgt1YyOi/A7jX2bp61lqdwgaYdX6/262wknhRjOW+M/vc62o/K33FKZKLfh
2s6hAEFJ/MAQDoCZvh9qeZYi0fzMG6zi5rB42qRVukTEsh6FVB0R0uH6CF3ADIHgxi02mOQHlf1I
5V9cy65iohWdx+vED1RZK/9+5D1x9A0HJ7TaQtIQiknG0Z3Rvr0a0U3ykzVLVx2ZCKF77OwRNR1c
PpHTEoaQ2pGVM13FwM5tHGE2DlPAp5pOrlc/IUqCa+zLPRx7eLzHVRQvjdcal/NcYNW5mKgjfZdy
5zfpHWnA7ulpKIpFoNejM2cYnmBNd6JNQSA71ToOmwgtk7IO9c2Y954X9y1NgpEuXZjrGu/18dob
zvDSS7QbnEEyGIpkQsO8ZL7t3fuAmWPY7i2UK0SeqMCDecX9HiK3XOZVF60CMbLAG1zuv/3atq2t
z8xhE/+JVRr6S+WbsLeG2iVkJe820aWFzc3MTYfv34yPJEjwXk/pw70sMzOD5VYSpL1L5IfwrkJz
z7JlrXGhGLUN4/qxnxVi25YGRNx2et4THdEcgSnXtAgm7PeACcnFp1OLTSCuFuFa7XgK8enGaHqo
FsPSLkjSFxfXVj5/ytB2vF7yXFluR7+1GiVVBb6cw9VuAemlLsihKwvl0TWshIOJLg22viVRK+jK
aeQQM9jkAVYIitEIX73vN2eRyDL0xJLHMwqgNrEsT7bAWDfmuUHwEznmFVkPjGlk1r1x0/Sslgjm
2hOPzItAvsv1NJUUQXAChYQw+0O2/RzfG45EMGWkN2xdQqRTbI1qILxOYzoxN8km7sDLjl4H9Ydq
R0iVj7lRmhCUENkm4J/Q7VYqSMpftgOFQeQO4WNwK8itHDStsKZcOYtOMhUH1gkNcuAyQcsalQoM
fSYEyELwVvrfgCgT6Qe8nSAe0CC/ZOYeb7VB2s5PdtV6Vlm2CASXsjOFqOHUmHE3R9WyVGU2nwQ3
edbJF+6wVDAV+ETwK5MVAP0bGN5Vg53nH0Yxbte9d2PYevx/sAjJid35LHBMdd0d/oYy6xtrUqOq
n/bVQgTfQNGXunAfgm1Bk4bEh8fGb31lJMxd/v//nJcne7lInK8n//JAdcZ3RGnVkWQesBFxNKnG
s3yHcYZAjmuabDJVX+TIys+gJ5N2xVCPJubkll+FiShydWrPrPlIs3YKk6cZELH0DB1fdYUTpSFX
ajPXgi/KuoWsPLZiWvBFDXQ3ERh0z5C5VmKevpUQbygc1/VHzlPWSHWP70RqCM3I/1AkGKXTe3FE
qPDAlqjAl7EWnNKitlwx6oQ3rsMBY8NnJ6h1/8PMn53UExtc5X5ghtt2Oilvzn56zY7tf2V8Obc5
X+kuZIqsFuGjUaZlpWelnEeDpHyC4jVwuH3tL67mGa/crCkQBXLas460NRU1BZKjUnslnS4PwojD
CC/o02z0Bnxs85h5GPv6dVKlrOOgfUZq28rgcp2XLhrx8zrqe9JZ1QBpd1a7/H0uaW1F5byrM6A/
sVii6mAXn9ZvKe1S5WYYpNHCVbIa772QKBPbfnccgHLME0f/EW9PdHsuua8DgJy9wRQI6wYRFSJG
OV/Q8hji3H+QHUAzzcnh8VM71XAJHT8MB2fdqOKZ2tx8ZSGEOIcKuImw5BgopB35a2n9VgVehIgc
AeA8sR7yNXNcz+C8dlQjZLl/ELl7l+78KRVtNWIf1+8fiq2lA4xfkir9u2mXl/4kS2HlHkwqn1Jq
CsG2SUs4ZbPKOWCTMpM9qL/y60x/n65uBaAz05unz5XYkUpldiwe1D1CD25uSR8XGHeBsF9kIO6N
+x/mROCxGZcbvrj1UjvK4SYhv+U2oRMCTCLffWvJbjl+hlxPF7IiPiTl7QRuGCtbypuI+Dp5Fbx+
ERD7NEfZChp/ffEPVqF2Yx92dFLcFY/djqxLEXTtWVs7S7CHaPCMXWhDUMZlU9V6uaeFiCy3Vok/
2uWiQJK38+dxl1IalzQT0NAJyfOWq3XGPbpVDNZ1rpICbGZun6N//gz14menf1vkaOl5aLflFOXe
l4yd8P2OiYHDF1eG/k0e+eYAADvuGBvTFxuONo/182e8jVdMYvViZvlEXMyej4Tk2wxZqNVLarx9
GHaJ48LAPw7oROzP3pJ/kvz2pE3bnDXQm91/ysTp+sCo1IllHxhv9KQ0INqXUCEYORoZhHP68zQd
0PHSscFjV9UMmuikZ6TyAG1owxNCnVX6ZxiI/a0qG16SzvxyreMqiXlGVh+cZIIdzpa/lLr7lZ7B
T7TzsDgYQ3aWJYdq0VAN0hN9VMMaKQFSOIkhKrYmYwXElxSU16LbmOmWjrRIZHCsYpWHfmB1yLDu
sNVvMbTBRuD2Hb3tN7CZogP5FdyqUHRQIwF8GThU/xM4Z2xBoBwvKlCm+kSL54o8MXZp0AymhFuz
NwLXu3p1e7SYm/B+jeitOabwcCJExmWPEnEDR2Ak/qzMa0iyczB1zYUWCnSmp1oECnEpm565lQ+t
XYt+CA+sBTizCUUiN8EmMtthVWJfxbY5ZuHa8BTvd1xWIMi4VBCUG0sddZDoBQ1DdJ/fKCD7CZjS
m53NtGmjkzSrpGWHEKb4CMVzwuVMGBXIy/5H6f/uv03PzC72vQILbu6NjfZ+d2vRTGTymOwSkiuz
vJAqz9kmIo4vKGLOwuke/ZZ2OQhRWfS6q2E4zKIuEKuD/ItTjzFK3J7iNz1LftEvqxI8Sb0xJLsD
xkY5FvwgwcRPewzw3QltuCaGZaAmiZolyqzEvWv01SEO/rLymlvlBGXTvR6hMQUR5cqixbWhF26G
OpQwS4U7+6OhT0Phn/lvDuLm6NJQsRW7yQTslwZ7ldREtbnW6trlVxiuEAgLFjIKdXUUWBd13Bxn
RnPPRH5/xXa2TXhfuRjk/fUtbOtzOT2diXtFKWtyPemtt2TENjWvomg/fY6+TLIR92xpldj9cNQs
7362UaawiZQD/8gJE0F8Ak71ChBShlKDyhxdeze4wGrPGI10aKTNzvdQg7yClWjFGrPFRjHL31+E
sMbeT+yrzXaCVGzmjJ134VQpVxMrjgUBEFOyvuXAFv75dVZIGA8ZCK+HkBgmo0p+gK0A7ddsu4mS
mqexW/CUnkzfNeEf/Sn9+CS97AwXKuLN8vJiUJ4hA8VEeKuyo2WBbWfAobrLVHay6gnjBjOoQeBR
6BGStSpUDKPcNzE/4LBYBkQb6pZyzLfog4DBp2gCYIzAUOtXLWFSwL5RScljD68WozWpAKfiHaRo
ZtWvRJMMPwl3m1ZOLi3nvPLJ1SDs3pUKyqBa51/r1KsqfTfxFMgZx3BcTaSflHwYeFeBglRIN60Y
JYvdIix3IrRj/1RC6L4otr+z1TiQbSuNdtgoB7QoR8kEFUZ7l3QiEbdrNIc2WlJtw28oDsyGhwvC
S7Sc3S6B5GNgmI3u3ScKIWg0zJUo/eQLznwnvUPH6ciVQ7aAcC4bMYdD/ApJuprzbpoTasmJmz1N
3uKoHZy5C93+aKkes0YvEPhH7wdb9NsqnjcvBT/j7BkyXWDLLGrMkO5WiZ/bVIdDV87QXa80q8or
aQtn5VldWTrHriOEkklPrKAOIdXD8rQTuBVt1JVSm4WxPp6Ye0mWQ17gPDC7M+aqe0N5OPoXFLMC
TiA6SX+oOoc8Ehf0Fd1l6/uikPbLOvS7E8GgNJP8VpseUSKwz87d3wzOmfPSz0Qi/+dttXmehdDb
ag9r/ma96nXwiaGKIcVH8CRcj/rbVc7rD8l5LskE3mSFYpxUmtIXE7NXWxbbTc0Ow4Nl2RIwSO3t
SVoAGQyJK9c3ZNzxWNExNdkgu7yMGppHAigwjfr9ZH4Jdrp+/7ElNsrk6DS9sD0AWsP2NgG+KNEF
owoPzRz5lBiWinIr6pCF4H76KBXm6ZwCu0QA+BlUYw81OFQor7ym4q+zuruQuPunxs1EI+UkMDf8
ttSSQVOHLLphstR9v5A13PAGqJZe4gVkdlCWE+7vtIoh9R1zNOQnPylxztcETA09BQFVTRx50g/L
mw33/qoVadYGARSTanWN58yu7ot0nb/PwStQ9hMbeAmJVz0I2fhrLukTA9l3kSvJSbs+hs7YCg1X
Y+YlUB5hxEDBJPgNE7DRSIJ9ws3E4lYYuBDJeBjFffFn7+1X00v2cKPdRc/eJJipWqWId6/N825z
NT9kOVDoX3IkXvwRpqwL0K1u9FA8GcEmmkq4VHmNzRRgzhKrKF2poBZYlgNuB1DioX8oomtPytxO
p6/EdNnjsfZx+Ny4e0uWUACXFutJ+U+P2JCb8XulTrLd/duhNKd4xNZQRCZoI/QxO/juiUjdU/ug
o5+fekIR/2VwEN7x3LLB0R9ENmAK0QSN/heT9RMfkbuyupKrdLuHWV1VRgaMbcoa5pNrlv/RPCb0
+GhbiuBuSJDNznKZxkVxtk33GBXSlqyPZU0npgK4th0Nn6wqoBiinZHLn2uNFIAhJqAj2nmWZMxG
u7tIUiFYNVm/0qF8JRJyKB5FDkRNAmKnW5zwyCBxcXfnGlD6KVzYXpPaCgy1eAF07NOVI01u+0ZU
bbZykJYxJXjD3rNTeF8dn7ZkrhY1TOvl3bnBjdwDN8Putsy+bxlwiAO3Qk6Ei5lADNOQVgdKrI9t
EGmHmfZ9VHk+iepq15rBhCYrNX1mdkAvbKvBmQBpZyLLmJBOigTgWro9SDR/6cIDAD5XeMLcnsoc
LhZ24w1iUs/yOtSoF/HcWl9KougFd0VTnZryTkPs5Il54qEIodgjKfh7iGGtlnfpAaZ8NCUJSGFU
V7bDDs9ETJ54AR+l6HnqVMK4RYGTrrPtahvoh2S+PFwt+P/9gTWKb/ApUXtYl1LPiFr2dUIBZwI0
yJYFqXjrgmO28T9w+v2apySKgEaW5nR3IS7N3Fa8r9wTxWZDaYF9svKlnA/oBzHk+azsDkpC0vP0
ugM/cj6WOHAKb12Lb735yQmerlhpfOgLkmdMu8sie3U+PQVY69CBj1nnORPVZ+AdA+9hCnIBhvtZ
tG8rEarLlf+5CMyWO0DDf0mVNwp6vT1IkFq+EwUUZJgnrsb/v4pmVA4ZviVAUkDd68xsR+Y9ODic
LyxZcHGwskm8BQU55Pt/e8hxKnjXI3DA32KdwAjUrluuCw4hcMlOZq5lV/qCGI0rTb7+XRWc7q3v
48MM5nlA1oA814RJ+jqruvgYAGIX9rUSa0EmOq29RO0oJP4nFQ1K2NfsN6LL/V5HFQUokE5x/Gsn
p4wVm+0iiAtucsSuzlfgMrTCMyOAmKDE57TW39UWnsEv9GUDr3OOg1o54IfSEDEzJmll0NJ2dWs3
2w8mWfNOs7wH6OU25VfxCr+51Z/jjBaoie8tZ6hbYvhd03OhbXifk30BOiYfKroPUrHQfSGmj7Nm
+4l4w2knVJ8x/TcQ6nW04edf4AVjD6o8p6rT0koq042UmCqg7p/Fo6pB2LMtWp2+tXmuBiHHnvWa
6+7wy3MSdkDszPD8krb0otz4VjXFpiDzlMO3G8O00Ar0buqELXo6vIFP9dRoCJlVM+wdFF27CCjT
ovdPA7QwZYZ+BSoB54We/pcm+LFvW2UJrhYbQMrCaA87X0AvvND1uGuG9TMk25zrIGhvfODoCOLj
fhmHPsmCjOljfo8OjkV2iWxisnyPLEbO5HB3fW25nyKkCw/bWVkIXrYtABGmobQ2mi5LoA8tCtz4
6BVT7GU1BoM/iqTzSr+E6TbEWbb5IYuaQBXnk08L/3OUN3/vqLvtWuqZFcvSM8cTPuQRGmfmIEKp
JYWYneokGbJ0mqnKRx9SyrocrEa5CUgc0m/hdgBB2DOcXrLrKe98tj1phj06GRMk0WAI8iscjk/9
jsByRjOEYR3QrCYaXR/Aa3xPjz46JxkFzrOIzJK1c7I63G1obYSKH1+uVeI3knWbQKNWbMrr2Vrk
mNOOA9nyehU6bZx2zUeiBLCy295GK1SX0CXQDnStMY1kn7V5W1KJHznZGTrVExUy+3GyjKKJwHoW
WVjvOfFLjutha2h+VLlozOorIKws8XbjwQY9+Su2HMVnhyJeUv2fPh4YQboI4YJgc054VZT9NOis
qRnG2EVjg32nsBa1fPhsE5NkqDT8tbwEge/RxXNne5YXbhAg6cwS5qTQ9K8d8e53xNjVG9zgr9Ed
teE0zHx0UZetJOvLkvsvgEpaZE2OTnmIB1D1ozwuI0dnEROqpsl3U0d5vEswS28EgrGdsdEZoJdW
HqCKEXDfNxYb1nrZdrJ1GF8ybK5oeo2Jjaz5rzI9MdQYq3TeLOjDtRjVLbf8ymvwPENtAt9G4m0H
ZmWv8i1t+fR1D1dsUiwGzzZl4c7YUPggz8w/xhtwr8fHNUBJGuTR2ffJYCkyjW1e8oGq9+jfXSas
Fi44EiNhqMdib4uMSJ93OJhpaqTwW+SvetVhrjvwWnbuFJFUSSccRORngaF9fBntiO6rWQoDBXIt
KawFNzqK2Xc4pfXN1fMGzhmT1xp3UMJ6kPAzNd80l7ufW72lYWzGggwfa6P/G6rw3jyRsN8Bdk4g
4xMRp1Ag0Zmpkx+wYbC+izuDBEuclGwqE+dVPfh6VXYc19+YGftztW6yzKf1E0YjYlua3NOvGlSf
XYERblqNmNGbmpSjFd+yCKDaZR83oxMAYyC13qIVw7/x0Ug8bl90fk8/um0xJB/i8VuUFEOe9uwf
HuBfK0QB0bfy+qdGqWHkpBd2FhiCUndFDd1ksIDq11cslZC6kv7Tzh2BannMEHZR5NdcOBf8uQev
xtNdMC74JLEL3p0d8lGnByQJegW7FA+Z6SVdaBpetX+al4QjaGZomHqWpv1ZjiICwdj3IX604/Ns
OGY4nFyonvv1w/DtzLqlXSBoaXeuvvHK5JqvSZp/fcqKp9WLVh0HUQBQV24gpHjiMlHmzz173ild
dMPxuEIhVubAxsM2N3zrTA3DkXX/XzmxzeHU9ySRef0K8grzBcbIxRN16NEPYWcJ/uOmsuQ0orRS
aMUojHMmzUO4R54sS7OCj0jgZUZn4H1Nn8i7UVhDeCS8Oi0InOebFm+YVAwIPw77e1HGW8j8u55z
ielKl74VMDnAXtQiyZO1Z0jAR486dL4KCM7hQQ5UB+piVp+Pd1vlcT6gJgomIAf5dDe4vIHIlZJV
CfxgYQs4wyiadmpnphHhto40TPNoLqI3wH4weQ3y+q/fPphN27xe8YAsPylIwQI5EgAQwdfo9jt1
PDKXWBzAqZ0Ce5gPrkbfC0U/IWWzPqm9fcEWf6vzNX2e+i8PoZnJCtfwszTFOpuMKs8jpNhUgy9/
1Ki9xqtL95EI1Sg6nH0VGWH2Lva60UD3nTidzxtI3N9V4vyjFN6B5l5w+JEDUrYmNUZuh7h+md+i
PaouTnohGKpV8rznaIiXV+GMw3GnLK/T8p3DOLVRxaawUUxH/sjxDcvi64kbW5xgD95YRtNQi4YV
nO/82Kj4db7SKCTa/HRcg+I+mmOhogNQlkHItZNEPUz0pgP1cqQgTrQnv6H2UVNsZgCEsOC+3qMZ
MGdrAbB6Ntl4LEp2CzvFAAPQfskZt5BNINntQSAchLkXdxMg+5/5NxsqQo1i/g+2ppj36s0SUlaT
/qv2uZKEl87EtMMKsZEeFVAoYW+MagjBJPpER045xdToXr+IrfYGR0Owiyl6yDXsgjb2DjLJTxP3
5z5rDXlsoAnhfXzm9iBJTarWs29qHrhAk2edgXsVhh9PWd3sppkJrE/cNMizBHtu7qcHCQuubNGf
AQd5zJdZ6ru39Q0A0aCKezjw4d8mVH3IRN9bFuMYgb40OFwEjIiOvp7aavrlIIXg1PeR68mVN2yE
rys57IKPCe9PrxjB717j4pKK9SiAQ5N/GTdWd+NaDlgmV4//Fk1BSLF3ItwqIwENFFx42O8G6tGl
vJAPtCd1LnSi050YGU4jmUnHFMehHBziqp8BCHQUJ8Lbymfck3WqGh4PVal3wX3p1C4SzsDSj79C
0uhvDfC4vBW6LRHELNVHjaVY3LbBYhJxO9mPEb+mPyQno0/zBPiTOtxJrXSGRjr8maRuBkTMpRCv
I8VnEZ6orvmfcVdUd6+5jSqSsFQqo+poyWGaXtL8EMy9FSr/bFtsXzg0qdCzLWT1T4B6KW125VYU
cAft8EfRuEUxqjRRKtWRg5F9NOGxeOLTxLkeWF+U0EGHAS9ByjKuVheInIWNuML3EFWrR/B7Qox8
oXzXm0Keq/xs+zfpd7LyFvXCQz6EUxBOnb6LPOwc1bPLn8YYY4KHjZ/qcxphj1zkpIDVU20zQHCF
mlN1Z9G6GQEad36tsbzf2GHSImKUTNBEBZJ5/+lBt4wKr2f/XlS/X8IeWGU5GWmjRYurMmGcRjqj
aMbC+UOIpaQjjJQE63qftBCDeAkeIDaLMRK+TYKMCiKJdT2Kza0Qsx1jgdaSvX+7vII++EdwGlys
ThFghfNsCHJS3K/swS2iUzYd+RjaAQ89nuyTczFjlOzmzXUmynKHTtIQF5utpsDpmr9hchlQ9Ai4
ZOX/4PQhQi3JorewViZcQ11n/BeIe8X8yodUYUYlvKTS7cIBDJZiB/4p6AoTiOI337e2Fbg8cM5j
B/ojwAqr4nYnshonrGkm1w0hm99AkFFPLhsKgmJEd+OBwrlVk0dAtDpd5cFWj+7Ey078tpCKCyj2
8wVj9SZUTxGopGffQoRF0a8ac/KLDJkFdD4/0RYDVaTZQMr8plBqWfamiSn+W6bAIFfc8fZm8GLP
3iD49nxyeWs4rXRggmKVTVndpZYabhYJ7nyOn01rOr8Lh1/idnSPMTtkI5CNdfqosDAJxKLJoAem
GQ9Q5dH30VUmUE8JemZGhumA9LjhRBxqHgbMu7j1VCDQUSLzwS/CXrGnNsVnT42vfMhhdr0RT0P9
K1XHRGPzumQHwIYScqN9oAdCy+OB3WlawMCschArvU89yQgKOuLic+tJqyLi2goz4rlJjWi+oHw+
YKX604Qnmqyl7xzSN96UeUi6nsfK244KadOToLoxPrnrNq2/hHUq0JQ50bCUNWqx3MiXNXvucIC+
gfoqzQI14UxDpAfIiqb4cYkVbybhIbi1lRJC8nNg0GJf5GgppLULRAZc1q98q3DuUbrwbW5CWOSO
PlgNUmZLtwinXdlGeZHDVjFd4k4oQ+tuAx28eqCBfAImWXffA52vl139UPX3hOzIp4WznPglTPIb
0YOmgw9jKmnGTMivCoeszH01LippqsHDxdsCqYoz8yUDXtKouL1H7VA5oqnL0HmoC0g31rJwIks3
MywF8IoRwcjq2mmC9PtFfzimJgr7p4pkphFcLD2JRyQNxTfvsTEIjuzY4jZbXIhemlE5wJQXfgOw
0H3wuZglTg0MrRJcmXpJcqLcOoIsZ2/aPTqKJXJ+l1qCMbfOmW86WPwRdzy+J8jKn3v0QOU4Td3i
+5xPHZLrraGqMwKeBlzYdJH93Nfx7TplgOIgOVaW/AMtM5t9tBT7sAs7hl1E2NhmQyX84GWbC0RH
8Ssikbf9LISf9TThiuhXIrq90bpC6eq8SCZphFdASc93tfUmrSBBEQYqENdW+bpa9dWVLy5oGYkS
ZTw1abzFpRJQrQHSWVDoRgHHbjBLiToAZiLsbFF8N2Ado90EejElBXVv7q345zyT68Kl5D6hjoTa
HJA6W43GyygB3Ip1JCN9PJ4IeVqItfO2BVWQ7mSgLUAtghAx8IyQzUytC0PdRbyXrLRaRhch7wyz
kCr5jiypLgXjwdSBWdJiwxJXZsBM9ld4W6r6+TX2JfjRdMqhAFGQOuTlOMMAI6bYQ++55AwSg6Fk
yxFlSxe9X6skbvTIDn2eCBbpVVwrjKjcRpG2a3H+zL7wNTvl3SfGr5rvcj+6Kr22NEN+LQlzYf6K
AIZJE/pRsP1l1HZr2OFYSj0vRJDrvOzLNbeKxw868UR99amwvHYJKbYQeETHzLTnYrl/88JCJBU5
BS7t3rdOAKE9w9so8BOTArgnZqS61gXCLpSoUb2fcoUU3RM9DgML+bsZhn1F2qbZNej290fQMpg+
HzJcqeNUW6ProVqYsCairScCA7OBydZ506FYwn7U6qpMIUIQ3zmksKURK4AfL4AmgaD+dEyoiaFG
Uw1Pa0Yac0b/h+mAq5i71CfJH79ofptXwh5DJ1yS7dO1+CflXMxusYY3MYNWPlq+tj1LWJNi4Ta9
O5HOxX1/6npkywv1UuFe/Zmyt6M2cpTJEUNHAT4aDQ9TsLsFtDrtYXZsYA2JvUJv7rj/fAJ/JjEn
Sz4zyRJOIKzEPv70SfU7IrDYAwQcSFC6cblj8Ae9nlK0/jaQpgFkZQiAz9ZMl9V72aIZMKmdTfHg
BPZWW9b3eyFVqzsRU0BUegjUnDHe++/eZ37SJWdXuZ1tkpG1hIKPOCd3qUWHv0/B3cuWCEgZwU/q
euMHRTUhvZ12Ex1yX+i3qNoVtuhsBES/aXMiqVHNABSWcvduVar2sZVSVFJl6kCf9MJvd0PlXVob
WPkyAuaT/Mo0R2bOXlFgkZI3JBWE8vwygKs+1rs2KAqk/aTAg1lKRMhdvQPURoswOkzHx4pfLIMi
DqD5BZ8/Cs4u/6mLrohMOBzZU+lYbDJgmQmnqActmABOe7C7Z7sOnpDEzs5EYiE1NgvW34EF71uy
MwzOjOQv6bYjDSBV81O+sbxhoYmchKZpZMHohcmwuKQ3SnA+QGFMRmj5+k0OUBazr92unCWRcNpc
OkssOBkdZ96aXjYkn8xCU1G9kUAv8RaSJCPh4STq0GvQnhhWXePBWd0Y0U9/RdptPPDQiMCfvw9l
ngsCvylQVBkFXexXb7P6wkcasGul4HEg/pSUcUyT9i5zoqz/WMifTfh/zpMYARcT7cu2dxHImZJo
A6MMvZ2hCDBassZb5rSANYCS4HCJCtvI9uxuqSTTZzkyVmt4HGnPCRn3fWPrf+u8d7Vy1JtGV54w
Rr0CbLBQ/yEq1l1c/IKBJMQHkAqkdklbd4Xn15KHSum/WntGhlW2HIRdc91ZolCxOy8632f+L4yb
Vrvo44d2HNHplQzVj8hv0De8ssnNgaQ4sL9vgQC68DF87T6jzr3bWlMHAF8SyG+AUGGjTIWJSxHH
sZ51QKZ01mGp0iR4YKPihJz8ppm+bNnput2NkzafxTnIXizTMZw24JijfLH18s9MdOVfY1u7bpAf
fMqdN/4IaDMxnmPCau37dKb2BiHIxJPgD79YIv9WILgSGkbDHq0dDN3CROnQnJtdfaPGryCJ0zZX
/ZRT2l5yEiR8M+FCfFnF/xQAcB3WypgHegPq88MA555vd+BXmg52iMZj6mENuz33kFsmEaBKAGwC
yD7JAuwCc21RXCzEl+iyNJHczAP/sCZa34+f14dpudokeql04Dl3nuBNyRQv91gcHsLBiJQYmiIh
EiqTiuUOwshK6hbkffrEvpyqQ/cmiuelYtsX5qJW0SUJyVxn/yDaJaYC28w9RWd3tfqxLLF23lgk
ZcJdmeYNqe3cUeQmF6q86PZ65WlPzl9Yj+7CmLAOwPWiqmFjowjgRz5BEBK/gCWFMahqwNLvzHQr
XgMzgNFHwvZfWeaiva88DTg5tj7HEm6oJM+NpKmDZgOgDewA1LDkx05ZxbEqnBaxC537derfKL5/
KnVZkT96y0bOw6DkxOVTOvy0rVSDJXJcXf3mjYHkC3Sm98CvgPMbC/TLCY0yiyNw47pfAthR2sRG
Gx2V+SUm1vJuYAJiTWjXB2Ipq6vMP0RbUn1AtOpsNkygP28TVau84e/ME3DIjxINMfHVMG4SQnaG
JNKX+9POpCRIMcNk1OGMm2Wq6MxPI78Jy08VITDHqwatcnlW6bdp3FEsX0N4hvjnvLrqsDiRbWWH
Ucm15l4uZsN9naG0CjMkWivo5JJPEPvaBtz+OK4iQ+aQwhj+dqsJy6JkfiwVasuktBvb0KzGMqOI
S1q61619BhJCPPtRs4GBTBdOwxKU+xw6ab5AXBlpuhf6u89EskBGS4ADIoViVJ7uDjaMZXhxpHux
NiTjolaDB2kEToH0nSyrGCwdz94hhvhLUzWor0hcFVPTR5u7caMnjSb0DERkaRWQVUTsPIbmq1vB
Enk12iXKySM05DLSEPVVI7aGg+MKZt9KEkA4d6SM442mVwWK2GN72lJvg0eldUq8PoKZkPXdNS06
fA4Y2n7gu7PPDwwbXAd/npWnWj7f4hkXlKJ0gAFkYuWZeDtP2kfpJU62A0eI9KCggjhNHLeRmpCL
jnDvjrXIiG8mEKBcJs9zdK0E5uHF5WHZE+KbT62837qfD6L6+uChK6cbbTrwO8oL0+xnzzedIqui
iGHFdpWPX6/GBhXYkziT1TClAMoaW30tcdC0k2vfRlSfL4//BDkcnASb+31ssSkNQHIPmpZIOWl6
ZDgYuYUcG5PzvAaIljRJMkrba2YZV12ryS36yf60WmihoJCd/B7QM+FxCGnJaRrQu84A2X+WL6VJ
GaovdDb2/vVUouyNCIH1p3aKkQmDG4sCj/k1G30NnoiEQaNb2M5vRJMEpS/P0cEznqxWiITZyAuD
dxudWj8zSJds66QCOtQJ+g6pz8czP1J+BcJHWm5tmjfygLqXQ54BMa1zekcBGWmOCNqiNdV2YLP1
eeakVW+jHcLo9Jm4tBXPlnoWM/DBpGrZ+Lm4YMOHEihigxiY5c/0w9lG4F5hIQthFf3ZHRFnchpk
tySdaK5mPMyDful6VKUeH9zLnc8ZMWXF8p2H1IaweCz2WJH5nTdiDFvcbTGpGjAlLlHBukimGXFb
sUmApTQIozcYoy79peRjm7pejZfG8888oLJ56pTRV6lZL6pwxQLl2fwyKTVb2J5vRqVuFjLz2qlK
uEjK6IBVjKXYcstHdMBkEEuq+TwT2N7XUH5xhNl56iKWpCjRMzQ0mmUV5hjd1EEu/sFTjn7wahK1
vnj5Kwa/sYHlXySO0F94+ei55ovFYhMJSF0MoJ1hH+lKOSMPgSx4kwGIGqr/YZEcmYuBnKO/aQOY
h4o9D8yhW5BkDkv14YLZIjTAVLFHcdc/fhuwBapChnd+lv3sTVjloxTLiHf9cGbpF80s9peyaN8I
Aqhys8XUWdxqOhb/icsaGHrFbpqzwQ/wIeRpOWyCXBSavIUGNKQr+raop6Nf7uINFIzQuBwP7j5I
sX55kMCe77K9WVZI8L519bf/MnsTsoPGS9G0uU87XUhXDMfvWv4I2Zu6Lfx2RPdkwgm5VhFOfNOG
U0Msuazpv7W3IfRRi8z+CB6Hme1MVi9eVsZvZT0YTMWhMi04Z0AHHQ+QIEnZ2XkQBIBf8DCrurBb
RYMaV4r3w+n3brk4R1eGHvIqEoCWw28GdPozG5oV1RAY+A/KVgfCO1OgbNWkL3WeyOOOVVgM1CHk
f9NsIrCi7WelxWUgij1rZX8+tyEgxdcvFXgpUi/arJ3SjX1kpc4bMNlyyku0HT/PUp1PKIbDnsTT
IRSAUdcKDIgPIPrmVDIDImXuXKv28A2/fUvBU4jCXJzCqI11P4bVM9O/lVaEZeIsJMRhORYXHMVK
6H4BoNZqkz8kP4c77IQDEpSxPB7I5wUfe+LzmL2dGjUvzHZH2+v2WU5MVXyiC6fb4fMMEiWT7t2D
UU9lEE3KKpZTz0TlyyfaAI0hPs1bqU2s+M6sw1RrnI5hHXrmrsDdrrT9ICR9/kxnvg4c/8bABXKX
gbr79xvujOKipCFrIkXzugwkmy7oF8XU0do+u+VwJwwiVYBJ/Cea4Jd/Q/Q9vk4XKyxEOx2cKwrP
ax1lugYbhNKnYJkqtyqAEgLub6HN1GeA9yKv4c+7lrS52MVF5dI5cVG999JUbyAYZjelN6bCQAk4
L/Z0wfhEYSZ3zHTglFdbxcqZfBuZAB2SII+dymJxZBTgMHdKG6RmlVcsJlH2WWs+CSA/zMaxfPw+
TCFjxGrDBPfiEqu8sxZ6Q2hqjagstGLnjp6LJg+YtFE8sNEBtesxcFT3mywSgh+8LPrCSg7Z68mM
S8EDdcRNG49ukzFU34DGZcE52Tpr4sW6AhCH/WWDrqjGxbGnw4EWhEE5KueHHx6KHJFL/03lI6pZ
6+xQJElKa0NcRgr+K7abMJAXNdStBfVLIS2JYDZzCgJyl0Nqq/0zTSnUAs3MXZF/NqOpNHjXsA4J
fzJdffED1j1WXxo8kDBTWL5dXZEG1/Nz6zRvhrTDHEh4MGwGPgaF2bLf6mdeQ/MjuNUlQGXPNfiv
NrHmyweN8ZWnStgo+XMk1YnbsvhXT515py8eQ3gA3ZD90ZVnZjGNAFaERVa2/81gYQimU1uZGC1w
0CviGyVRSk5eJJFl/3V0MXT0+ZaQ3sl+e3syrMAHVkU3QI7tZ6qsfVRKrxal8p7lnQsEuNoKkpH1
j/bMX2iizj3kHhx0eS7jSr4HnO4vDSRcSvaqcuzOrAgFmuABcM1DT0BSvUjpDnye5gtPGNRS0cx9
noznMcUcSsNVZsWZtm7O6X37rLbjOxmkrvNIKXAqljFV9B8Qr9tY6Ra8pryyJIuMQszFHIdrK69U
A+vk2O5hHPnqY4z4v5au6Y+8i/T22NyG9q/yVGHECd+6dlzuF0MRz4HF5JOqSQ941w/E25leNxKx
dYkPx0wdlqWueJxBJg7IgPxXh3n5VBMKQtbjKxgsPNrIPLgcWxpPJwK7agKUWMnAxF/u0KJaEs+z
gPKWp7By8SgsTY0r5OsmTzPGSAm3jf5eZGsnN8D0Mc0YJQ7bN2L7rc1eJfiLd4lyg9kZpRXSOmVc
WzPiqdJuT4L75DkTNVbfol/rLy3JcxIZy5o0KozlyFUQkgbMLnohLVS3y+GuvxQjGBQQRWkBCrhM
LeoyNVXakmuFQMLzho8Faxn0cKrIeHS3o/lhZQibQDld6M+WDzh08M2DZAf+aWYoHcUPFE8LoPqV
+QvrqVQKSmqjlbVbSWfommDyd9klCQ5DrIurLQ9G1Ya/TTSViFWjnzYebz3UtmI+ypxtrKZkgou9
1s3CiJrl4L20O3rPMMIQXmUv2SmoU3S7Q+OQ/gJj3D5tlpUzEq7Enkw6lDvOLH73KnEZjN0aLzkY
OuS/GeB35w3L7kO4aVdDwdBavAbKT+RQ7inwgT6zvWTFuWa/uo00qDXSNTkJdNBOHKRH1BjxPSh5
wvmB0JPz2NZbaOuqo2gdm9g0WeaoZ8nErfj2FmiywY9bdcsrFlH+JWavM+MwdvJo3l0MbOIZz6yr
XSesZQ/qAmSCPZMSVkE5FwU57Eiks9RGATvru8xQ+MjAfsMUZaRNG5G9hAyJ/cdJfYvPeLPbvP3r
3I1bDnPhqX9+qAt419e4ea6VldJcqbmbSinaNRRXOccqqEc7SfOxA78pOkaXb17CcsRts0x3Eq46
eic2trzph5D/sPOJz9XQ+GlTDQcr2wj+qg5dH6M6wzo54gWjBTx/cVuKlbBEiWJoHjIdjMgduRP7
lgAcl8DPlKs2uC8m+0YTBFr1b7ROEDBY1U7vjYDgyqC18I+w3Wa83ctkK1FxWFI8UzKgynSllq48
a1YKmHFLcnVoq7fiTRtbGL2PZx2QG2Nol/5UIWIbt3JsaSwXBbs8QNuCXuSk1sHIayRXwol/FW4R
Dx74CGsr3uufhGbkv3O0Tz55DLCPq+7H3JjVn1WAYPCRvHuyONNx0eqQJvgBsh2/l9X/sCBBZZF3
gxwGUhYNrzeyLdqjGrrHvvh2RM88qC62Fh4MDl01VAHyu3ljfo1U5dlLA/YDhMdx57WPy8TzF9rf
KtMFFdNZSkeU3Vo3E4Enmk+ZdjQN1pe+of6GrHfLl4NLHwS3NNMToD71qg7NeBuQz8Uzjnz9rQh3
06iW6TLoSFuNzZoEe32AxVcl3WusN5cPvhuswkHePpoJkgMqevnW41QfRqPWP+KAq+0z2sRDVxIe
effL4DMWD92zRFuaqmtw/tj8vyNRjia0qhKJlQQKGFNKKe1WRZmwe+KH5DQcXKnTwm8C5y5+qh75
rxWcNwJ2aqufFzXeZmzndalUmEVor6EmqwD7Skf+0Uv3OTM1bizrn3Ndq9KcUz/WH9e1oNtcn8wM
aLdQpkEhgwkrW7+dnIbYY7Dng2KVacve4MPdWsnz345K25H421HExmS2F0zbHzN4/lLLiUd37+vY
UqWY0Joa4VgV+O0TZtMj5w8WgCmi24VF5X7fOLzmFfcG/bbNJNxH1spoGCJ7/TUMuXHq7UaQeGgu
AFKBkPuCKe1OIFW3/y97VBKrYEqfvsk88kepC5speWFNUocZtsQwY06Rc959JssJQksBfaDC/qRH
ZkoaDvgJVJLUG9eOMkA0kpqaVXrgTW1+tL8d+xkNB2ezG4kVLeZonwcwGPatTAUuFVkG48c7r1WV
3qh7FIL8rNCwE0sFKayh7oS9PJdLJ3Omg2oQF+1is9J1aQxSNaOjjZ9mwRf6gYbrik52F/coNF/I
PsVdEPcq5ku9I+/1eLulUIMamBBAeIxZtUN0TckedlcgMuPPFwY7ijeFD81U6yPJjR0YkkpaE/BX
9NLqs/Kd+who4uJI4ML018T/uK+bapyGA4ULkK04YzNIzlC6F/pfTdYSrAt2xP1BBbMomqPqT4/Z
TZzTM4Jz6aSI+hUyIABHNRgeiAODvOlSqenKxSSe3HydrPBAjaGOivgSIHNfesRcorPK9Ee6bw8A
jvatN/npWM+mEFheXWMacfVbD6p3t0NoT+dVJVYnOZH187UDu158gzRb1EG5eO6p8fkLPciDxjMc
U4pV5wz5//soPIkSWtaY6mtex7HItisY1/lzLND/Q4snEUv6WUXEnZTNoCsItTKZMVn1laIosqj4
L96DPD9+rouRTgZt1tdF8dyJF8L2U1rB5BUe+bZE5X+wBIlSXlvIo5QT27Oyq6dTayEyrWtdJTqj
DuecvfpuGmlQZnKlMUFDwVSKn1LTW6gVuynq50wxfnO+sgDDbqQWJblWaUHlwRqQbdQlOPBjZCeA
jr98IZNAa2A2kY4BqpYeKOdoEXiWI0Qup4mwNcfgH9nFPRtqAwuoup5YWkM++FFRs2i34WLXg+rJ
6KkAbZV4LA+0qUGjY2aP4UBr05nkjNZkxCV9FfNFa5FtAAXCdcEtAyco9wigfy5mx06KdzH15A3t
6XY/vCmWITKtoAFLAtADXxdyO2JBZYhzq9hwQOpHepH15qrvwQRXtE1DmcMKFWrX/zHzsh68/N67
U+k97AvPU5WuXgzaOF/kceBAbUsS2HVpfhRck2RVQnvbPBNkjsxgDLZ3bHU8iq2UO74+MKFld1Wc
HahN2i68kh5O1fVWeVHBQ4DmGqAk/+AtESxhJWxPdhG6DL4YaMJFNm7xdzlkKgv4iKYX1E45bgo7
qu3qvPP1zR72h9F/Bl/JR+kfMFnOwZ1XrS/7tRiaKDf8ND+8iw5I3tD5E7Wai9kIApIu6xlGs2IS
M6fyGSlsta6VKjeE5xSm34xCSrQhnNaA1ek2UQs5aWXwjLk4gx5ap5+whxFcLqIVLQULcVhBwMdF
5f6JHupimN8hNDLq5YMxZPzNhxvI/cHi3cfJW8KakJ2A4k/C7znQmOewpEK1rbAYZVimbpGErCSo
S5feGXKmM4DYa3qCtt84dtVEUPMN+w4QylNCmRqFeQqtRR6gD0f0ZjHF6RY0KwFic5zZm5HlLO9t
BZ5LI68OuXaXNBUQh8ysifB79TUj2WcwRZtihVc/F4RqYW7xZx6UxVvMm5UImfkU08vm5nXoMYTq
0Xt8ZtZLW+hMCSAX5Rd7XPmKJ+uDxG1kAyYDlp6AIVgzx+4hqvjGAZk7IpF7TME1aj4a21pAazVg
HzkcGoc9yPo091pkNFryNIgYbQ1PCkMJ3ZEBcghcyOk7hBtoNJcr90x6sToRfD5iqLxE3OrJJuEg
fzTJZOBsNCYX6aGILmec0Cmb26ow1GrlYEmz5eOAmrYF7QkSIYXCqUcZQwCaBdl81rf+HPmvVjdO
yyg93wovU6nJU24HyjOIY857bF/LyhbmiFoaO3DCtsLl7hdz8XdIPdM6rzY1klNs9I4lY2PP6KK0
WsGKab0zpUj0O57pbkhJeXxTNdts3cQ1KTTCVX5/rAZLURNAvB2oDVXzbVCa+TpcpYe1+emzMfwr
XsTtAZSlITxMENyRNwZlQF+KAnAJ68dso8JD/wC8i4gyuxYATcjIlgEZuBLS9KPtqf2IXZPibS8c
88UuBgErLImy1CxbL+ahBKpRRNJrG3Lek1HyBEA35ax7l+7gp8TssP8PmVcraNGD54DROoYcVkC2
SBM9WP3hrIyn56oK6MqKAjiWDybGIa/YwUerzTBm8tHKjVy+Fgg03XJO8CZLEg7Eb4WojRcK0cd2
C18ffz5J91ojAuHq0qQH3dyyT+TOqGW+lIjdNwN/z3It3pJsnpdoT2NrwUMzE6M/3DKrDaZc4/jC
La8lgeJa8D/INH5SgqVIlk9I+6C8RsWBoK3lZv5ZI5A2/9YKX0UsdvR9rOfD6qE9qHaL520GptEx
xxSjiVgFOIQAVPNfWPZtdMCU7vdpjWVYT+/xGUTNW3FvOKsXkAMvzefriwKl7+GGtBJnlzXUTZSf
v/hNwmbmSB1ZrbLc7LGYmyOWQBzF6CBKl4pkfPbnuzYCCQ/zoPoDZULRAXEfxqvZVIPtFfzHUEZO
Vl8FSiHuo9+pACPRGizSifXhl5QtcLuGGDiIiJByClNMvI94u6qOCs+lh5pyPbeK9co3H0yXv1Op
TGUooxWJOvPIZzFV4TCbAhjkfTMDcvOBLIV6GOT1vx2CbFPw1XXYhaoaxMLKsqB70IHf373Nja1r
QUcplf4nBJ87SqZDN1gRzIl6TUFNYodii15Eg2dWyNHnkjgUSbnSgVgknE5s2rq2QyFqUd+ha2iG
vyyp1Y8emA8YYfMLEz/dzmx65NyihD8GZg+ycy61IT0HQkZC70S/qZCcV05CIi7xf7QCBc2CHMef
NlfcyXAzyC2GVJrsFUdCeKBjymu8h21SYEdhZCo7cOQKbTySY54l4/O0kcGOmiwYBdJiLrkcjOAN
BDEdk1w9u5jnhHMhySFEm2DwBNxmdBapG8yOaG4iyW+cvk4u+LzhSQ+jgNGlh5hhnvyNc+4xNflz
hFzodYN23rES6FIGN+m87EzNVhLZ8M7mNhX3XC35q8w/37oGChJ3TyVzvaoftZX7n8qvQxK7GNZi
bvj6Vcz0S9ibB0BvBKVVBOmKlJMpgnnyWPi1uPQgja6RnwpgkOcLXCVIsRFxALu6lRmJdTflyS+J
M3toZp9wczwju5zuj/vdTspaYP/4VK83d/oA/gQ2BD7NjkzA2i1/a8imxYvg92Dlpm/hA4P82/fJ
z1fAGH4LmRcEcoK9CSNEn9Ze8fR47ywk8hitOmjNDAadVm2ley1jHnHhUmGOE2shqOLbxpk7z7DX
ZuzgWuY3WAm858wj2xMvQuZA7SA0XsnU9mBtUFyQ0LbHpT3xSLkaMvaRfPOrvc8FkA1Wd8o1n7rK
r0coCgVx/Uxd6JvOFMFNpecqjD0Gvh6xi+F5mAXPxXni51vcAfhm2eyKeggf3UKANR6i+JZa+Njo
JY4IJYqoDYKB321GoV8A5Whde/b/bHsgFrMfMMnuooIh67n+BD27tpDI7Fk4RwCgBZEw/Pq5lOS0
nG0NFrdNNA2IOgFR2HzcVywKN8sA/RLDiqwMPS0Ysku4KWojPLBfC5wwQkptt1t3CL2OGsDCwinP
tPcGCh06wu5h/wNYR970xyvJWouKKA2RxBY4FC3jMExY0h2J0x9K285ViAMvuDm4Fa641fr3B9Pw
Xu9SaT53PVLLSWVGM6zemIKRzAgjfPUXPxOAt8JUEiMhr2PhtTlRo/m4XKG8CSx96BX7ljBhCih0
/365N8CtrsG37pMicDlX8dHJ+YE2IHD4jnK+xtlXwo/xs6af/5h/p1L3OQTYhsaJQ6iKiUwy8RQO
F3OmEeig8phJ6fcO0UYlpAYo3CG9xAhCdYcYwDtPZXAvSSEaykfaolHDTfFtjp+2rFwLTtizGtCX
Tgk+TkhLXRsUwrMtYv79soOy9Y5Ca1arPwe4Mny5qPTTKEpCC7YwMeGgHRzqdgpiYY9BaBbeyHcd
Oes3bxE214vPl+YuWV2YOczjx4P6qq6DhZ+lso3Yh0zd/p5iixOIDmp6cFID0gPBPBysc7DYoWlG
kh7jgvY225DWWjOiymDUtqm0HoIi5XyhgxZGoc5MVeCkxkwT2f7/6LzgzWG6g7QwFnZ6hZhG0NSn
1jHb81VoiYigxdf0DmDXpD2vGxsUg9dPglFfeWwbOMPcjqpUmh68V2uszzNPhfPTJujHhd0G/CCX
62O1b2G9vx2z3rzkUBOiOtpLop/fw3JO94YfjIC3jBwF7M+B0bL/F5lODAgqf9WAyhtLlBrp71p1
/ABXG0XdMPmj2l0lBy4QfBxQaGXViVI/dZESJCUzX2Iebae79yWIywr843OtDdLRxBYdOivLEken
B2YAWy63HkUV6aRqN7JnuphnCp9EC+LNtbp4FQtGP4LGnzkdh/4i4e1HtB+QV/NyRjj1wv9JIyqs
JZm+gbTqxzqfgEfwV86b1WtpNewbrX8Wh2a14OJFgbzdUOe75bnFphdUHJaZ0P0EYGmpoG76ooBA
vCwERrlD5Q5oLMjTjUppO00nPoc7uEBVeEfJ0JBozulerttVrIIxt6d/JC1iEL69xs7D4id11cut
eKzbS56xo1PWSMW8Wy/0hOhttBp4I5nyRQNvBDEOsVTrslU0KdrS4MBK198pSwzIQtKKMYW8b5dz
v7WPxggkUUY0vyp9IWRlRPY3JQxfRnB3fCGMEMhenhxDnlOkn1i+1XZRhIWIafBmLKL9slSh0eZC
PKyVW4qECy84jnhdCd/cH+KIKE3glNd3wFS7pQg2F4yhdw1A6wYshBOHFOcaWlG89P+VfWvEwF+q
grL9gmgpRIWswhjk/X8dAwVXb3i9bWEQC6YBSM7VbbKqlZyc7Qh58qbBw7uZGp8Mr20LG4EyvAc1
y0a6Yh6Ejg3txke6t+m+OI1/M+Gi+rBnxWTRY6BMg9OofKYui8j4alw3zkHNI3HfbVbcS4E8t6Gj
WwqORBhgONtowHTNkb9VYZWUoNIAG1N7PFaCJibjZygeg00t8BE8xOSPPGVZKg3jk3TLAcFOs2Cb
eHdRTBE/6wAL5sWvmLULNTVS4I1zY+8AGYBsxv811LmzHz/gHoeT/yR1G+/NlxsW5lXV8I4EdZ1d
fwbpT2du0ZSYGBVs1UafvD7zBk6OaWo0UfewPvs0my4dpCTGmd3hHtijvN/ECdNDXQaieTaKCisB
SZPd6bB2LQV5IjoR90TYUnTGpEDWBiPeZkHWCY9cHQF+/uq1S/EPmNDPSiXlDPzMo7AWvk6wSC2P
QDzbwKBPt4dmpPjujqD4SGUyoRcVrmH8TtIIilhiUiLbeNK/+ld30++1xQTbwazfZx1yPrCps70O
9wqFGKt/f5WTG5YrgFct4oxvcVbrws+S7T1He7lBohZ/7MThNHmrG5T79JNH2VwgaZ0rV7yw6VUD
r3d6mTJ5Y7Ss/32AwDCK3YWNWPXtjhKgUG9B/Xfp8b3H4BQGVt0qQzg9mNs5UpwkBdycWiKKHNC4
TbXadndUP+oiwfMHP6n+eO7plnHftEjzY4Car7tyduYDBCTV+fhZYGPTt1Z2zYIAWOwbtTC2Zv+h
rdHJ9+YC8n4VbT6xV+UCuMOKDgR5/7z4m68dwfwbHbs1B30PMzpA7tbRVFTLXzb7nimk07cGwa91
ltnBOWACsYrVSV4jUT0o3heD00v0LFSX50Iud4y2ltOeHVvb+0mV+vNVnLlgQaGcYa3olYBt+YJx
8D+tcTLOSawKWcc7xaEwMLe/xJ6lHm4Vjdlm4D2Uu2LLYVbsQC3Mzp8ygQ4f0aQ4xJCfq8c4/FBb
cBSSHCC9spBgkmGNHD9jJ7T07JotDZj8BBi8tb/UsvUVhQmbvxIJ6AZaSNqYjuyNMMgS9yBjslLf
4ri4Q/HeCo6RmJVytSVsnXcZzQ+M4SfBVQ9noWvG4GeYqE6gjdSnQYWTFTkowd2ymiaA4HXFamEe
KT/B9Zz3GNaUpBqJ+vc0q5m6eRJa5ZXJhbtZlzDCZVZS+g3dqPGHRCYBPSxAM6nRmaHKr1NmN5Wv
1BV0ynF62JVsJlzJaQhzlVv4+dqVf7mCwtNprOsY30sWJWADqkWVllBlwv5CkWSbv6Z+PN7dkCzj
qwpLXoAfHPElsLLxNywtLjUecZaVg7A1mkNr47DuPMZ55XUtsJFaScgH1pLHSnYAtYJRXWD5CXI6
gUzSQlk7Trzqx14/WF/iB2h1pPQut6JDiBNmPffKkaykI7jdtsvoBuer3UxDZXz2sXCIzmC2APXr
zuAmEBoeU7bwLiNO4+mVsCJBRM9dbrhtZzGNJ6ptSHTkZr5F3bNVViM7t4NKQHLyCUct+ieKu7ri
5U1H6s/+tpJzdzK/UaTQYcxBzbbPTnV+lBttcXuHV3JTpyfofWEo2gZ+/XFRFSx9GT0bDFRyrCJe
eH6Z6lZWiqqDEP7W9lC9gQZQLSjK82CNUE8nUOncAu6F0HzDse1+D2TprMjCgtZ/hOPmbcXFf/Sg
vIPhU5IyXI1Obhqn/tlfyp8aE+ca2/ETcjlYJ8wK8lU7IF7/OleoVOPGK8sdNBLVkS9v8BQMZekL
ZLtyFbynoP9t+R7wnkt3xx1/UezLaRqGg9lX2yLFN+ByTMxZv1zYOWOroLXqX6I0qI6iM+Cs3TTz
b4auiIb1O2t1XhotADMnSZxFQaqyyVAEALvUi+OUEctRAU9weJrV/OSE+2ZnoQjgABgGD6iavpWJ
yfeeAwmlK3zgI/Jt0NkwZF1rE985/utjuFpK6CmjyxwticFBQ8yy/xc4Lu6V4cba4jl3kKJh0SM9
McnAspoKTC/z/QKHa48pICEqvPAfYUcyyLm6qcrip3SJ9h0ckuAPgnDs1ZX4d5mw7+q+oI8N5zNz
+ifH9AuT9q8KpKJtygJkjq74QWvz+sXuRWLAJtRMP8dT+WQ+gE2g3t5VxMZXyH675gkyYDbB3qzr
XicGHSqyXo9kcE5VFqZ49uqEuYKZQZhy01QgJtjQL1Il1W0qr5/bwo567s08pmENssx++x3CpqNG
dqAt+BHizSDabeMIZFwm/5YpeYsRXiIk7WQwkbZYTlLf9nYAmkHxMj1063Wng2WlTkDC1Yloh2Q7
2TFtJS5vdAA2A86Bv2YOIXbsTCy4q9Q1OLqPkZK+bWEaCmZstQ00WNY8kj6h05ZXZnkrHO0ta8tl
Clvd01QYDuQtGHpCXNrTdFVR26ucfKnjNzZHiEZMFRsEzFJJTlB/aOtNWBi935TOIeEk58V2Ccmm
k3TiDAuTn5pqP/rm7NaA943as8QTQlar5vkNVgBOHW1Y5lmkAFPqBmdzbk3w2a55LzD4jCdw6Djm
8TGT23l9a0jR6IvJSPqKrAKcAhDmvrQpFzZcM3Cn7ClY5kKK3tw1gV7v8FtKK9XC0ARIwE4TSLPi
K0qTSr9Ggt5LSHwR+u0V3TQuFEA8wno9C6afvNUE5UrdjRPA+AoFDR4rt2Lk0L4HNcGkURIEFwk/
iyMgVujrJSkalxlNjd+qzBM7Q9wbdkwcz2cFlEQqnmEgL/dwsU6/rTYMTKIebB2WK8Ei5IEXCcwj
hiJzc7riB3Nuw9XObNvmetqN9dnnxM5TEvG3FjchAxNk3IoIXc9F7tQ0rvgqMJmiToaRUkU/KmG3
ZZJZXhA/+sct27PL4LQNd9KSjNXk/uz3k4aDuvHHGL6b05LXuj1isMZ8APDFDRUxp9SaXGINFD50
Dg9P5Jth3jhwiA69J6CAN5GLlJlFPqsc4htDTw6EaZkVpq/gXNxJiSyWPHekRyHyMnOS82yXYHKm
SFt8BSW3mEBCydjslKUHZhPEoXFr4c0+WFc+IS1Qo/ivi918JoghOSYkZEahy28CaaFpBg6pa0O2
KPpFLIewy2bQIRytazGy1G3yih5PRGEuU59643p+/cydiDexoV7pUHa+KKQncN/q4Km+HSz+y222
ukPjXqSyJWAoCVoOwTl6u27y6umv/of+PgnWYxpak7W/1gJ9MM52cq4JZWMa1UrY3JILrqM2/HwY
juyHMKFOyv4cXp9RH4ddZ26lRkSDpvx5MO6dLD9BB0XidEnhQG7jrPWOXfUA/5ATLorgqhNEpO/L
ZwlNfY8iCWfZN0vBiImlt8KB5JMQHB4d66JLbZID0+J1s4uH+fo4/XgkFMJ1mzOGfb/hMS2N7PAk
ybRzXxeHl6UvOQfZIU15iSOgSigoH/h2taC/vs9b8e/j19+fX4v8n+DZhsMmrELMw/QfYyG0hOuh
JMJt1/lktyyKTV69Z9ra3feLCkPnfUObecgKxxH1fsPhj1O/TIKXEk86K4GbpjFeSBjwdGfAxi7g
y2WaWmbZEkFNUt3y42Vpozm9TED9GQ9vjU1OFt5Q5nfMg9doHl+4fH6C95fXdjLmZz/1KOd9c9xp
vo2dWILCmazEwZM9+kx0QP9gUo0Dy2r75D2lHtfmVCHg7AGx9ShMK+kcgU2BlHwwxlb1Ncx08mpa
trhsd/zlh+EX8m+wcxW4GvT2iIKNyK9ycGTNI4ypzBwL9gh5dizppvRlv8qqe2xieBK35T8SAAa2
JSeoV7kLVBKmLVenIa4TUVTXYmzFxTf0s0w85fHRPLqKk1hybxz6gdeP+RJxGgbQJpwqYvJHX2Gf
wdfJMk+D7uCWiKHtzu4IO//PIQk78Fe+iYQ7mSeOm/jaj39tDzWAFdbYVaeBUEqpNYssSjbiSoMY
9WOwn9AZqEvSu0M4/jQESRsgohlGJjJMxvsDeHyAlfifBGWPYOtHQm3GExTQY5hFOojmzevZ2BZF
U4prbTQP/9gAeslHpmSToxdo7gXNMmhxG4tMsceANdS/vow5PDOLicgEilcZoWrR7MlsPQf5eu47
4E1c9Lch0AvtQnu6XtSwVtgdzto8QDhlIOczEVUWSb7wPbQcN7ZiLowLrVXPlFHkJGEJnqkOxcb5
tfkGouINpVpQyCFUZWilMX2eacikuM4OqKjxqtJmIGF33a54GiN7ATWaNaAC+JukwMmlAyV0cnFy
S9jNpCu/FhYUOHPL9zhKv0G2C2v5M27J++xPfcgu8TccyJNFenKEh3/sKo89gbqPIg1JPLLO1ECQ
lR7ZXLOPxdU80YOQaU/O8UF9g6N3MtpA96sLhnGuziooFUjn7b6YAOZupUyNb2yUGj/UdtIBOm9x
q5WscTgCx66+BXYHxd3cYn0GWUiPwnW0PPoiZvg5gT/N5m5Hy5TmXifCO1QNzE+z857DY6QIxEkk
61V2nL8ec/4/6VtLkYbY/dCyZLJ9dUG6Wgd4o4YASXo5YIFdxB8RSp6Hp0lffC1XiZ+RecIcgqdz
U/F6GEnCOjrQUEYnoaFhB0aWw60yZZkVeMt7IFUrNi9RWGGrV5kIzZZHHJi4GcpiemAVMaA7m3ZP
b5+jeBmUXyI2u+s1rPbCYD8Qd+ZkfegHvdjMxzcgKZB+hoStHqzlF/rGAdB4+UjutTYiyNpuSbYS
6VL9m35axaq3TGStaD6o4Zz7/+Y6lTwBGs5N5kXvfrmjgpsTOOLeuCZvXEgshq03g4UGNKY4/8xv
v2EEkP5yGhV6qMJ6pGdHujqfRD2APgcr7tzazGzmEEBELnlrND7P+pQokiNs+cjUh72hvRm1rLRv
l9eCYhip+dcApD1Lwtfw9Agf09lGf1vRVjFvn81mlPZ/DZFdr/+ZCVOvBvlDi9GmKcAc81RQPIQt
09OHYO9ulgAT9Tb+3WZE5xd/LlKceaTDAoRO/iNWqTGQZUUgRMAr3xLsUcZvXEljuISGSXNV39KW
26GtNZKubmgCrlmakxujyBHXxzDw4hoLG9GzRlwKwdJRkg6KS85yd2d6xGsS/3wveUv9IEkqBMu/
6O7MC3PFsKdNbAo0WOHUlhMS2FbgCbK7vmBmviHESdb22GsZiJImwbCUxs/8b3uQnsQf+BSd1JaW
/vLi++AcfD+dFQmsqDuEvytqbFJYRHsi2RzOmrVLZDBGH2Y68zWQMSaiHfLiZeyzEJB0VrwTbrQn
NzIXABYnJLX+ZzokmecegyeJo0xBABNvhuxcqkA0bfm2cMRcEi5g4RWXDy02lQ7nFqxFGXMFeh17
9ar7+gFUOO+JJRu8bttlXP7WwmAuN0K8vDbiCXpsRpKX1is5nXuLW6U+3gGuSph2A6sWpSCgqYcM
ih/2R8GR68AGZ/4PiZSzc6ayBF2OKYJ756vCj54sJYw0ts9wCeJWiJUjAjPZk/USXpbaawzqhihA
UxbHxgzm7SHSvcCvOlw3nIhCsMenhPuEFZgr4ULHZ+I/KUHqcaOs+ybso4jrai4hs/ruvEgv0mda
VWanxPDoBHwbHtS+2EF2rSe+Pz1JU8YX5VVIl37kEDG6niI3JMZ5EcGHPbdx1IMR+DLgwhaKwg0j
dUmE93EIziGZ7A+xkijWcGuCScBpNqjtNl9cvruqXjD8FDxEtF4eCpJmAPEVRkQrbcFFQZ5Aa3uO
Sa2Hf0Lg7/EliYRSFqg9c7fF3Nw448gAfAz0G5VLS0Mj7fUIGnRfSAwz7tI5nGpHkfxIq1phVNf3
0cFaEkbHH48Rr+/cgl6YaYoyk3nWaBVAPINXY/SYMsKdWu+0CfAcgzwk99Lnbe0uRtKvJXG6WTIu
O95XrG+fooR/N4zV2+6EZ+1dXJItnCfrMvv31woa+88aOq+GQ+sLCfguV5d4u6p8pHWW7nNfYn1x
ZYnaNu5tOEXY+DkI3NCTjBvY223KoLCwO2HnEsV/0qlrSpK0SM2LhVIOO3SrkJjShOlXtLC5NgIg
3bohgMk17lj5AnR/sy10x7OcE5yIqA2LVPvRXYM4Vt47I9NGB9svHPGwfGTNeZfcbN79gqfndj3U
5p87c2es9Uhrrz8APAA8EJ9C+gbocm1qGgDIbq1q9savPo9/Cwdvp0ORNT/DnRIIZcHs/kvLOVJY
9MsLSGHBKm/2ZYFP+UUotdIVCZXKx3iUelW8alZHcBHMFhJjGeWSm2e4EYznEnWsWDLLORYyrqxh
gDgfhTWtp3XdOdy1r9fKflZbqkkhfqrhMkOqQK1aNuRHAW1ev0TZIUQR0/hNye1ys2wn/Va0gp/a
hJUFcCakjCFSlPgPXjRzj8Z27a740yaL60EJiGM9yUdWJ1R4FRmSoFwN+iGVkC+jBuRFa+loNZBT
dFiP7t+Q91s7wpJcGNHp+vyER7uFnfgEJ2/qeFVMsjBMt0y4PrrCRfaWeWZLS2ujFlUqA9QmfKQD
VW4hxdhZydv9YEoFwZxYeBTli98IeRrAlXj8w+LgSM7l2lBelwSFBtfTDVv/YBQ4K3UHPstXi/OM
YhRNPPVBNNa3HO/d2iiyZwzX9MaahggnYgEzHDytxX2cxkmh9pWq/QX2GfEkAS7M9qDhYRmbSsaG
t1HoB4XTpFvzVSETafpD2JO0WkS0LKfDSiK5TU4w8n+qCXofelVOED7i68IFo348G6XjIdhY97EA
Bv0/CPxoETe7obdN/INWj+EnvJtK7zq5uT9IDchPKhh6NJsHkXJGf/5i9WCy4qcnRuUCthIWfI9B
axquWnKV4wBA5usGj2g5yqbR1/bUTFlaB0pj+8yGp3UPkg6wgsf9C2eSSbo5moBN2RJtIOQHw3Em
G90U7x+zOnO3Q2fci7b/4E7pSsj1E2ctlSAGwWPRamZyZ3g13tczkWWKQxsZZG7Kh3/lyFwUwZbU
wjSfgZyPTFCggPlqocXKcTqtffgLhQaPnWplb0WKgBieXAw+Zso349XGx+TeYjuLlWr2uKjxeZvX
dSLCLae6xr7f8P4FCoIz2BzKqBbO92JaWi/W8cvho7kCVKKPffyt0ArV0QUwPw4YmDySatVfNQBf
QxJG8MDu45zp/d07AVTQdD40cPKElbzOZdwBwX100ABUPik+a3xIBKM9yx3V1kGokGOlPeZPnysH
bodKqLTVrYz5wzk0sO5aW/2LlJ59LCZwVd0J+DeuFPnNtnZ0DwGsZb8sOCZWHi5ARpIjHlgCVY5H
ZQoiehcdiJWC4lfDYtXVj24LzNnuE+xSvMHVCqBT9A5pyokPp8lNTxUQRd66wCliLCZAgMk51xwn
LW0fnDNN/uBE+pWy6kClJqtueGJB8Y+gSTm3OlPFhDqvJQKk2DTHIoKa5cMUiu6TkSs21lyP8rX9
cp1oipJFjZHpIiNuQ9NwNsSZitNwdBWZMkR9c4FUOBffC31ldXHxIc66DygVww3tGVhoFDgSN0Sn
zF8f1dmmvEth4InGIYG5IP5Cx0GhzBQCh6lQKtlnS7i9RefiQZIkqJp3X4E4XyePV0oO33DqaRIx
fErG1391fAOHpI11rq6mQrCLko2kCvduCi4F9xKTbZT436hNoZmgwZREe+KIKPz0uwI5kiI8jCGn
Tzbsg3ce2CcBcmNMYbf1WOm1R/QaiSnjXwajVs2zarn019G23O3KO7nbh3Uo/Ep+1/EOM5yGZ8du
7Ij1tLB5b+lR1fnZnckk7Ii14ZaZyIv35Y+TREf9rTCTb+PSLg1cfYat93JAgvDfrrbs1aor4JMP
0kgYeDeJ9vywT+1qbrrbesAyav+tGoqFBXO0if4DM3aO4cqearumB46J32U9wwinqrSQ5E3cMy9a
vReFIPa9iyvNGxkgrkyokdO3xEIrP7ZmjsXg0k3qtpUBPz0xZJFv3qLX7EPsUYR4wxgj1vLYryeS
6Oj55I1Xl0uer4idBwf70aTpPGFP3eacIXaMf7bzSek77QSUkdvmLN8G0BzqzhDVqxUSjrPjuqlT
bbZQwQmZDMSGI+iUKemnYkMQLIzRvutaDCJF8uCY7cCA2w7S+PjN8YLkF5AmB16uUXWaGx9dmSBZ
Engc2EBLKxbH60nbBM2KofoM/+avcS3B+08qiDT2lMawOakb6ghFlNmJelyvDhlEE+cCcRvgu+DE
2zxU/r4vv6EDOasp2SngeKfclZEraOvpYsL8r6DI+Vk2BCAJrgXqGWlW0wYbjnac+gOqivYDI0nF
3ZUX98N1iaQ1iY4mMuPri4uieP3GrV1wfYnV8g9Ys7PgyGn1to6bK/wP+fosiduBxWP7k2p5wfod
iP+T3pQiXiTcala5IW8L7JFZTGx+MfHYUWJ9fo40VQjFS2q1vBrB73Xfq4WlLN2zm95VGjpUNghp
Lo2qhUgGPr5yBiiVES34YwL1cpWLCajEnaehiASS2mqKSUekkR8+sShz5Y/EERYo1AboT8BUut0k
z7oQkSm3fMrs57O71ukAdkBJfAyMKkhXFEKvZGkPi+FnRwSt+NUkz14qgJno5PN9B7VkBvCGFPNP
GQUJAbqbkjIP85s2LUi6y19jZ/tt/mkQPauk9jsMf3Z51kWmOCy7yv+W3k2+xG8t5BNxRCouwhq5
aT/vtMFG+6Wg8hpHVV59IOv/VfMhJPDLSTzQ1QL5Xj3gc7jcvEYWYUpv0AVHpHF9O/wSUz2MCrvS
/dyfvKq+/V0F1AWy4x0d8zWk0O5Fup0PVPgXEaaqb7cfhawu6L5m+kxxvAKr4DDRoFwqDyGfD1JI
stShIN5NLfPkwJU1NMrM4T42pEoOwEE9O66Ezc/fCeCO8pdLbCpxiLQQwOPS7YFwe+BCCj/tpd30
j12YkZDB3vymCCQyd2BvzsieWAzftWGjJvL8jZPw/OSiveiUnDQ/TXO/PPpZTAjRIZqEFArkpwn8
+MC2k938ro1vvNC03UiXpYnYC/AfcFdpxBnMuT+V2MwDuDXxbNDBSDsBZ4zoOVDUYjjT/obXMuOe
KgGPUVjaeOfFPvxW8Hnn+M9rgZbHCyupMlU7bAZZYgteD9fzqd/nRNqK95bJ5L4QXrTl+TcRyyqW
Sj21vgq8zA9red/T8WR3ZoQ2/jvc2MHmJCce6vr0NNmVS1CN/ozqo4vHgjOztJ4zQvs36kybC2p2
hktScgxTG6yvensvjC4liARVUtpIA7mc+dNz/O2W1BtV6H3oYse6LUfa7fsdg2c+m6VUvnD+Uv+U
WExvz7OZ4x30ixxEIKJjOalh51BpU7DEoZT1EMuw9SePYfCJXdB+u6jNSEWyfVgzF3wUkE7IfMez
bRDQ0KNFhzK3ed6t1q27e1lm21o1OB+ve/Gyy73bHkFZ0RqJHeB7TI1z3m+pF8w9kIKmpsOzm9iC
NKVBiF5MfFEG12rjq2rctWZUIyeu9crYgONhzos6MHhfz5w5MBbgNAPcN0WCMbgGK5y7I+il7poQ
ihvpqbhWVNx32uliA1YV9YG4rzWGRFHOspw45KV4AYY88D4zK3WngbRXDW9pcavDWoe8mbeKX4fN
1kyp2PyWTuQ1KFbC7Z0uN3Peb2jDd3a3VAytASIZiyiH++66WsaW9ID7LlMggsFE4i7Rb8y8WDKJ
QyTI5G35RwAl9q064z+oTa0R+ld5EMGgnTb6U8qvEy7Rk92ApugYepvcW4sa34UbS0n7Sz8CbvuR
0D/0VEelbZ5EGI8NZWa5bQ1OeR5PSaDxbrEhpq7K4WSXDKRjguSo9niOdLE1PbSt+orAZbJUXmo7
vP2TBD4GxwsJXQzB1G9xcs4YYCzPbT/eFHROSMJif1VctAxFcpRWC2X8m5NNCZ84fStyrU/ZKgEw
epm6Tqzoou+Jso+6phNSpAeMjMSpve24f+BgOQYiMFEu9Ud6tmm2/CTrSE6YJr/nlvtp/bDmQCWJ
DDH5w4p5tvq+yyF0YQzZjovASxYABYLXMO/Ho54gaRhdUXLPUrsF8/Mnt+RQPuFJk1vSGPc67oOY
w3xjrxFILUlI/F1NlFPxHDS1KHGQQmFc9BcIQEirQnXEqxaJfcD8fjac4yFW4bew3B0nPvGzQ2jx
e88PXSpR3MCZJL2VfT6sQ2tSy9NyiFuq1S82BbVKRO/S/aXGNF0Be4PTT+Ng19A15eRBHF8B6HlA
ILv62CMsQif70QYuMQmPXxBLDAWprOq3muYcihXJY7s4erswcu34SXYmD7mM75LtTiNVdzDn2Ax5
SjfWKlimSUH+TBfv1qd2TDqjneVkC/lNC7s2RwSJRSj74hkeb6BvtB6+J+mZ08coBtDA+Ymti4S1
Tv9HhYQvrbZBI2FBxdrsOw3GqAwXxoDNLsd2+W1MgUPwJqTx0hqopuvTp0cWG7Hx5h2GT2RQ5049
DtVYpB3or6YUAIjZo35uULbtCkkSoRzfiA0zlzyk0ME1/85WB/uhsGhl+03gzAl02G1x5duePMrf
31xPu7Bkp+erSqp0s9y9tQ/GrZJETYcEISTyO/SPUxr30oFrIi548h0zueV/k5jVLyQO+BPYoHOe
hfVTv310kiSwIhF8Geox1dce2gsl+uGh/LEUqlY8kUkVlUL5pRfTrNdGUOaUBDng6ltoGCWrKKp+
tlrJ7KjVT7t5gYBFyXFGLc/5Y/kDtKTDIdJmHxiPVmsGblb6DOHp7FRsefRWiZmGndyAkKj9ryHQ
cE4lec38ztEAKjitdnwi6rnk7A9G0FiGvbllhSuxJJkKwVzeCjhfRugPiB4bRt2KnyDsDdVEvU4K
FMq5llApdZJSQfaI2Zb6Qt8jMY2TdtwoYOfF2HkXEY2suN9kaQ0q3gTYWXQqOFPIXgEyc4sNS40M
jXUMLU5T/pP89qavg8oQCWQYH6mr22LD4D5X3ODVvqmX5TIqGrbI571lKnRx0o+0PoJHjgGUoh53
EjKGAJdbXRH9qhSGVK75oe/nWE4qbi7a1IpuNaOegL17kT2DE8y9QHnGMr/y5QQowANDOb5tWDPz
+AMudvyWxXbkrhm6SS0mVLLc+lM26CZDOqvTb0bmoNllSXtOsiLYjXWuYbaD63J7axSWs/3QDyWE
JQnNDOltmMZSCH9z3Ab6US78SslIP3hsje29EWtqR1rp91+7994OnIU12ShrgfjhiNaR9aEII0rw
YC8fHGJD3oT1cK5J+JGuI2syn4RXQTf8dqIRQD1V1pTwbSCEWybf95I9U0gIxXeP369Nx6nTNO4u
ZzAJxJqhJ+Qc0A9TbrcSGAWf8zUc+yarQwu7r+e3+RD0ks6s7QGwf9+Q4x80aQUoxWVScLAhYPzv
tYOlWxWePgWkHg1lpyAxDuuEMVuu6miqi0BIBDepqksZWuiSPzZKJKn74ETrcoWZ4+9ZcpK6ur2N
cRRb/KqPkIcS1ILq/RYD2dN/MN4lmjYvrKp0M7PnEt+Z0f0Z05i4UgOH6tzakyEBmfZfLbmeNRsj
9Ylydpi1ru+ylXnkoIJSi9kPOc23KMkrmPauVeA84aqBttUs9PGUB1M7wDjf4/jweJltCvyvwgtj
mz2Wfq8bpwGSxCygaZYmd/x5pVtYOSGrA8h6cLwCgbbcjCMdOCN9bGLs/CbcHv4sdeqtHZDKLsCB
txNOP3Ro5Ry4ObiTx8gaO6cpVpMNerHvB0DHo1CZ6jIGsCjvVpVaWt/G6RrWd3nU9CakB1shqm3V
6vIAyz85fmZCBMzpqIRepyGFAfOQ5bGwrPX4M9aZ2ki8m90R8quD/YjlEhUXplozSLYCMUvQtaX/
q8TH9PfDqjgGxgrLncNGmdTeeVnJ4qnJDB9WFTqc3TLHjhGgCVVEMsGyT6rpPFFZwYpA2rR/yLyB
TIiYw8mqmMRPctgzESUA6qY1SvXL2B5Y0YrpbKc2IC/+Onrm/y6jnxqtxEdmNmh8tgjB0PK6KXpY
rMzlsrOJICBk2d8pHBm+h1xaXB0O3/Hf2fii7VtRVgnTvfawtoT0Dl83jhFoqkk+NbxISK8mCTci
ohdJxLWJOohI9PiwVqPxdnueZj7M/SdbsRM7k1eDgJ4yV1zTr7nhlTGH9xVst0LSuTVXg+uMnBs1
wTTjsamf4M239Q3qPiMpA9GTi6lJDXEbsgonCFJGTz21J0e0YzuUqRQIsNNKOp+DLt2P2YyDjEFo
kprHjmQBfaEHQz8U/Bsx7LpzC0whQAtvWNVhB/4Uwry3xN+02qlPclzkEV1T6xRvsTKg0jlCyp0N
A6DFMKv7Rz42A9f1NlVmSxYBXTh7V4NSyqU7WplnQnasZ4KckWk+1Wjm/UfS2cbqFpbQziv/CE3V
7CLRRITIYkQMCTmv9xy+/ZVBWrXEwqFwvH5FlOD72hEWwqnfOanHwDCgDLckPj7M+DRbWSRA0Ekp
61jKJBt+ZsCnUWBx+XpHOO+3IBbV79XfL6YyLyRQfMmbbF0Hx7rnxxwLoM2zoDIaN+3n5+7B98DL
DZQ/mvzoEBhJGbxodPXwLV1QGuN4rBUSph2gzK9mmTo3Sd9skyudz5KawKTIORA13KwA0LZFUKmj
Sy+6yqW07jrCblJ7L6Q1idg/3vk6/sX/l0xE4aoE4hELqMRBDj5FhX5Nys/dM3VRgnu5TRfkFmC3
o6MrdvWmVO4/fQ78whDSN6ue4M39yiUfksvmf/dUx4QA/8ZsNvTdto2K9wPS3KKehQuAELjLh34v
EPdMwoSdnULgDT5RKEdcKJPd1XKC4QLLwqfkuKWYYlEdeS7Ia+RlC5Rwor9seYG8qFAk+GMLM6SV
yqgZdnqrOBRz9Mv8KMegn8mLobEcUOi3r1YzbRiXZl3WkSCHazyk/yURbMYm2Bv/G16eX5UXam9n
w2knbeAIFVgGwzkmsZyGLfbC4ZP2Liq+JoxFa5kfXFONl+kXmJyDrCuMSANHq3HsgG8E3QRHsm4S
U4tzcPVT/yOSMUXz4lbPjRYGVFN+QakYQzBNt/Hve7x4SHQkAUEJkuvYxu7LuT30RAbgbqk//f79
nd1HTEtU8Vksim5tIAJRXnJWoFr1TXaAB1cYjZVD8aO4DX80CczX/Sey1S2liDBJ5e7xbgVN5rF/
XdSBlvDJCpCbrZAWOaYT5nLsgspiYeT9WzVmPs20y2SLwiAvNfRiI12MbrcVPzlGhePR+c5t0/+c
A4BNArvoVIx6A2QScc+c5r9QHT64ZQgY9gaPPlGh9X5FHomIyiKVeo47yeimamu3R6yrfNmmJWY4
Gp9yZu+NCS/7Q86q4rCQMYsLqjvZwNnTM7BSN4crlOl2QgAPdGZ8zKflUirh7E7EUStcHo9QWyw9
EoZJgTYH8Vb2QKToySUl8pueT3rCfjE0btKANDngF8L6YUWPAT08wgXtpjsU4f1WWg0WRF4qx4Fq
RCpHWKXcDZ0LLe/iuozu2ptaeo6smACo6Em1cW/sd9R3Hp1DfuRy3b82MWmRUjtMdWQNdXzvo5P5
Mn+FHvsTT7z4izmhnixzNem9LacU3xLjx68r4cStG1OsKSSkkLvbJ35RCgm3zlkWDXv6UB3Mfh3i
U6nzZxcx5IQdMAcgr91SgVwi6Yb449dn2oqIr5Jn7qomqIzuZN82BDJo9GLObE5pMzD/2ArGDz98
Xj54c5+H5dTUJXdhg+QqtGHfCa1dY2oiCkUwCk097pLwJc3H71Ci/eqgzVqrJLp+PYrXnlMRBe6+
PQnvG+P1faMu/Ix2RWPxFRDwVwb8ujGufHpP9dw5sucCzMBB8U6sd/66FZoLQInMajxKy99An/al
eW9J2r+E8HXidDl8/QfYysBkHfEwiQk0VhW/WpkoyPJARt620g0S6k/y4DrsYtYxndyzt/Y3mMm4
SjXo1I0jaIWW/LRHNA60zhopCWwp1rUo07pe3odZDZdCbH9kesjP0Z5oqtNnld4uaZFTc/XxMcuD
8UJbKYwUErfDNT0d+VSlP1SfH+squoemeLpoIGWI9I2X6codYqAW6GzANpPUZJuAjhJdk5GrvEC7
vUCLTk2Th6Xn4Udu7e+8sYx2m+xZecojwAzc27V8WP18HsST1aKo4kXf7bkfuWqL2npqV5uN04tc
/0Kb2ox9OxA35w5RVGv1SGahvC+h84vlULw4hUQD+3DKQgO+H7Wl6fMMUsR4Es6TcEpLGe4TKt11
qKdoo/db1ZVgGfRuwPeM+CD1aGg0R/EDJf9ady+UScF7bG4c/2kVKYgWN+N6xBUaQ0j+dT8IlfC5
uHSt7wVF/eLze02dzayVw/T7bpq7Z++GO1kCoBpGTFIs3YR4G+H76NNBH6Pu7gcKPNoK8oz8aDd4
2PTGxE/UTnXnvKbG9A29uhLtApFriBGhm+DXtyexomI0prxCxMM42WU8p5DtZotgpaU78FixeYKP
bwTnqpMN4xBNSkkLF9zqwSIGKh7vR14S7zsc7Q3j/El1x7eNCJZo9FF70dCfpHhXhSCdWIpuzwW3
D9GfLxaF4AjIRC29YiDgeWcxDkHhduJ0rHosYkDS/yQ1n+nFVAFtIzVYJIgQg55D9oq66jfWb+oi
L673Izzclh7z01PrREuxrZW46nBVNSfNwjNFrlBSaUFqbR7z893AJI4LHuFNILnmIDJb+LbnU7Z2
2BI5UIhDCDkSqML0D6+UHwOAg8twna/n9tyrfqjckA3cnfeH/36n5tJ/3VM9Syx7hThyDNXLm63u
mgEdMGr84WTV/iVYFfGq9PR4TyWBeQ8B8sANX+tzqyuDg3/Ttu53aPyh0kHoGTVYAHCfpIqoHeu0
n6BuQLo0kysoTC4PwmNRH9sw6wRuYn1eJF39S4HUJjwusp7b2NnjdM7HF5U0KkFXLjA78xsFqSFG
FFcj8tlER0T8SOphdix4HJmrgidzCv1hWEM21IEE5RwbVfdkpPsGK2e5tCgP2IxG420bt8SbhQof
ELbruk57AXLOFha0dO8daDlRdqw08oeE7dEBSR1ayDzmSvVS0hH4JZZVByOquJNrIjOggfDkju+M
iRcR7KqZN7zh1gxf/eP1jd1nFqLsEjA9AVKIvsrscsOxlmyfLNccjv3eG2EDvcDSyVCk2XAhq6Wo
EdVVEOFxaXQ+APo6xK6LLNH1SCPKFRxuejyUNFShqncUA9LhQxq0i0Wu2il1Edk43e+Lev2R+iov
HppyWkFPFycDVnmmnrIqe1wcHKhlY/TFvpswU2xw915qtmzEVOIxoaRTKOBrI25WXdk3Nw+1hLd8
7RVet9FEjnrchLSzhfyr80C4ry0dcEZ/o0xoagXjXjpzMb4yg/Fwa95TQldYLZmJeGhFExfkZhOI
7UUHqJHsFDv/WW53/V0t5e1gWUjYit5QT4Cyu7UeE/Hig2ydOInmDs9pnH/0PkuzwR7UBv059OUh
YjdnEHDYn4/mOC4EqKWQciLhQO65iVxjYfEXZRNgp36q1C+8gPZQZM7bvDcZA6YNjE403xcGvIHH
qyW918wTlRPV/oRjp4hsA+WhkCh10eAzcAK0Ms2geUc01sb+ZILFd21IbYmb2T0BUzXIDvA3tc+r
KiG8b7D1ww8YqVqJirNiygphnmVzlrFv+GxoZMRVM4OKHm0VJraQyIqCZl+xJm9wv3DRwC+SIK6H
8USaKjfzjJk9vywoSXT9KfWFEb7sd8A+9MsPWeJEPZe6XQB5SNvU6kGCCG86H6SmHFD3lAGUDE+J
0D1xZNEbtCP4m3ARsm1f8KaP/92eH2YYdw9Nly2E1YmvyIEeIVQLtihRAyTcUxO/WSfjjWvobcwj
oRjS6l2qS6BeUSEKQNjI3FBYn/I/ho56LVlums8AGVvPMd+ooIwelaWLP7o/2t0Ur/rkyl3Y4LJk
wMVajJS1bACk5yECY8REvpiWuS0IPR7VLTPe3ZvoREZ5Jq5bG8SEfkde2L9C2diuE8Tng67f23NV
hHDOX8tIIDsM4YMX7IZ+V4+6N0IYPMDrLFjuuy7KqTcLE3OxWQjkBH6Dq3Ou2mNmS52ASCj5PCq2
8pwV6zB4lG57GRt4mwyqnFBcWipTJdxE+1lg7IcSi+9vsCVdHW7sCVuzH00b6/fUnVZBitXArSKN
A9fHUezv//RFuJAf4bKXBlZSihNhxlpqMGeof7rFRIPh4tDhNq6YZV8Cm8EkAOqgF2eb0jx67Fkk
498rzjz1YEGhBnfTFAuXCHxBRt5e8QC92LRsvepZYFAvPQhYc2WTAu3mioDqaz6xhIkcy+MJU66q
O4H4KUT4KD5+2DlbSz0l94Ybt5s6LyUUJ3c8biPJxEmz98JDtpwJj0wLciGgLYi4a1n/EjCWz2io
Fv+X9NhmAJEa5zlW8cIc+Lknz02Mh49RCCg8kQ/MaMGKB3JI0eUAEXSGS5Uvc08sQ/sjYUqbxg2H
gAH1L/jl81P8W0Q4T/1ZYxsNpYjX3c6zcUnUWNnXWdeolV79ev8WcJPf/+n44wYeK1NCpQfY/h/G
c0Urh5kxwLHJasXwahUM7/DmZ5aZ9SUZWX3TI+w7U3bhRvfctti4WXCLyi6ql3ZH493UWbj7eizo
QJ6CQUjY3pLiqzj+dZmmxlLpu0Ochw2cFiyv4aMStp6SmRj/a0AnYshoo1c+ydRrl1JpIKS/zYoa
s4rZYTgzytOAF+B9ulZcDYnMB2XEhWohUYjlgI/IHRTL80wNQRjP3loTaropFdaNHrcc+0MzaHI9
J6T6naSVkVSmnncwqISug0FIuKAD+AZ6Wll7iijv2l01DSkJ59zgJG5Z61x4gXToKPiMJW+M1aKj
Sox3BC9AJ74WTdNggfSV5+pby53o80qDQixiZ5wpOle4ZIlaY2LjjXQ7Xlx0tMCeF/xIrYfcCsf8
I9924CD0FvxSl3ErBW+8FPnitUjB4fzV1Tptn/az5EN/38T+1tWAhhPc7EIpHAhqR+hR1yP5Wwf8
fVxBlUUiXqDrgBaMC+2yS+2I02CrG0yWL9OyZzOThWZfg127X5lUl1Cw0qfrhhZ8jud46NMBcRr/
Ru5Jb4+boayWgydJX0MLdXcDSRm0C0Guml5lJXEJ07YZZ56k6Yd5j0Gso8tCh1yirdhiBx5S08T3
HlVv/IJXDA+81sf5fQOVX1W4Ox7bS/VTBom6MMmzwWXR22Kvx8ONnVJD+Q+xGoyfdDRU+6XNBq9F
GVwdHwMeR791/VOX1Q6ehvZQryGF+8veuyiA2b9GvMTwITEgr6VyAm/o+q/3yJXRSdlUtUYjYmth
w7VC046sE9WKxX5Os0h1uS2KEV32uDtx2GD8CqOgJNfDjCZ1co+fENj0+09wv2Aw02ijuonwP29T
0GJnBKmtSO5dmD+VQx9WEGrrzEwAO7MIrhcwNMQp6D+hy5zoItIpJd8dvhbe6HsUlV2CO2gN1Pj7
fZJHd2RusH7mBE9wRFeXNpn/yStr+7icxiT9eJbp4KST1hq7xZIvK2dQFZsIMdTGaNFCkPcrlHip
h2gES9d/rPmE4sxGBQUi9DWEcBwp0isJelVBAwSLRSX8IJW6bANSChUl5S0sNPGSola8/aClio8p
ZOd83xjYF/qgCEyli+gqe4WRr/pzyiA6PDk9/1F1WiVCkkTCVbTuq/t72EZ1RSWU+ILb2xzpgUhR
7gSCn7MScyG0gNZqp3BJXnpaLEdHksV2sGG7QQq9NRq9o6fqeFOHy75g8SNuy238Xx4my2KFN5jo
W+xDASndj4eEoARH7fSr63thDNIoPi3D5csv/YBLuOqbExd1SkfzfINUfvIo9IrhxANIqc3/Ff2q
kMmSDNX1eOLl4iGcu/VSg8lbEzOt82MfiRxNsjwguYGWf4bGGZTlUw8N6TNiVvPzJyTlnh9j4/5H
ccjYXUKE6b0SYwQSSZcTP/gASj+vzYmuQg71vDwvg3QIVBQYoUzhp8NgcLt1K8dpC44LRbSaWJVQ
b3rAOxkeyKOH8vKkJqyfeqv8SWL72auE9iAr9xKt/Cfb3wMDquIESzyT3yp0/00KKZSZVCZ/95LV
9Q2brj3ujKkCVFsdpBm9m7tnvCYVFkwMymktmPv2GJBp/Ru2jQrrWaGgc+os8348YbPsLc51WIyO
kFvZ+avc8EI7VqfIVhuXl30w2ZFd+Cr2Y4153XqSMiZNQCRRdjWbvtKHLlJB8CnFzeb/5O00jtFr
sMZAGw8H6Q+KU+DIzVGCJsSxW4gvOOe/RicjCFrZrqKYXMY/cXXrIah+zKwONfAl0oV1cXrOQwAK
pEtt32iPzWAFSeU6ukNctm9UqZy0Y5cO142gr7y2FqelWk7huBxe4STPD+9TksIl5qi90dWwy7Dz
HyvLn/KR2LTlqNxlTGTjW/iRA/AoEHwInNN3xdyMZfnwIxv1uJE7tHMPEd70hAlkLYhvAbLWNvIp
fDp5bCbqSjrP3fqGLbTKccn4tyf+iGeE03c9COKo72WBgW2bVjXXz4e+OYVEFN32NaMqd6lHDP1U
N06Fh499M8wr6g13gXz+MIZOx85rIMaJCg/eZ6RTdhcRr9xwQWQedKOOwHg0aJh729k5+2PakWd5
A/nBbTezWqQjYbYUupVkd/y5mN0WWAlgeGqwT270gLUht8Q15yGXJkoOYH/IoaYSwJ7ap7+HZvzp
5vYKGuuYe9mkV4aI/BgnFnGe2N3BrRXRpeIkqPrqXSdWyIYfidhqtaauXLJ9xu4HLJbsh1MWOqzm
mcnWVOTrN04bjrzlAy2TxbheFY2i8nz3EtQmv52GIQisw2UtZ1wFwBBV8GekpGvvT6wfB/zlX8x+
1Jqku4QyCyJaVRmwrLgw9iotUUaGJRIUm6Tf4I1pXjumeT8DsKFCO5Ydgla4pvpKwqCLXRRKKrxd
1Q40mcDvz4LlQi/OSuj6oW7FHB/UerB10HhwjMtE3maXfXkIgHzmIqv+ugMgbHw80rnNdDbGYBIU
B9szAy8AsBlJx756ZwM8hxP2CMUTdQSkkflrfAC0in/ZBrB9XsYlz4/z+Tkw9fN0cE9mYLF50HXo
2ND8sm70jmT2pWsap2s4KuQ8QSTbehPQVLlW+hVH1Qb8pLeL0GOvsw1GsPdz83pTjyLP85/Lartu
r64fylKbzs3sx2J3oAK5QKxzFUN6OMKqTgNle3s2AYgILLaYj8grLf1Fb7ei1gwoSJlhSCAsZoZj
6adu7wssoIGEdewqWAefl+jakB2BbucRKCoXNEt6esI+/+EPXJzoQkNIOnxBcnAi8WRZ1UDb+FlA
pB1Elb+RY9iMkZmbW28h6xrYmyyATCcAf4oNevj8pBnAZde+fdU5XYsvYvGHr/JVcYxMRQ6Fnhkq
oeMeu3s9xTNpa4f9shGdwHwcrX2V0+qTKdP9+mR6mWrHxPKQ+/LSQsgVoW6mHGXKe5/omBcACT3D
wNGT4c6AvuL0Xfu5sNvkaC+RimMI29sZdnCqgKhJKRFIAhCaJUU0Y9JB64cb75nP/jsJRR72CWsU
UFeoTeNJ9BdEqsNGk2MJ4k/nSYE34pz6B/zoyl+aqfdFOPL+8CVvQfgywS/kqgDR2WXnvMkPBs2I
HPh7EXXlMPna5deifoLzFB3dAAEv1BgN6MJrwIQWZCM4VDGyMyaWBpgTeYTy+nl0HCZSJFURUasX
Y7fNPf3faqicnCYRz0a8GNH0CKzD1AsiyM5kJEL+1QJ8bAIo19OSeQkVgXdoEKzO4NrHbsOOAMzi
7XPxFDtvI5XffOmN0/bpQKJ8/6i5Ldj3l0lvHqHZD10sVmjDgRZOOPp9bqf3GWFKzPQJffhFdNt3
eofx9/t6/SBhu0CaxFi+H/hE0q9fOKHxMJKyJ1vL1LEtlT3pWvfd8bdivErSYywNDE1tBj3bppq+
TQafr73NHOBT/VTMm2ECbsVfXlkkYWZVUgfUJ5hUiHbFbOw/qQ4mh3d5bTRfIUCHcYrdQLRZXegj
SoYSEC3WBCVAAbGSxfJCb4365cXd2ea2DbtvacoCgpv0PdefAVdT0KVo1N3mLiq4C4QlMZEYtv73
Dx5VplkmV0e/QSIKaqa6qu9o0qzgDDlC5FmNIX4+UXaxmKQ0DvHNTjuNfMMqaJssHi4taIlfeIUu
Ihb3QUKO8KSi1bfpCxR9qsMOryfw06PIaXfNpfYGQZWjOsq1y8QA4AVkvuUhz+bUNHKwWfzk3ckH
4UPUDq9dNRXw1XrPuNlo9btWV8EqK0NjPDU+hBoqgxiztx3Gwyx+jPmgCWHqKi6cuYRm+akFkfgU
MY+KoZpWvm4yh2X0YTPAdjmLDa5bg1tfxMWGFT9NnMSj0OVfr8jUhdCIC1OfwhYa2R7TLA0XcTAV
QQzrdDh3NdJItEQo7iWL/VUOdqtX7Uly1rKA5/GyJhpV/Z/6Lc8Pamvku8oqtVqGx4kACGIfSgrn
UQWoMI3jI8AUEKMdwEOPBGCCkhu4+RxfR/+bfW+X0VwsPxPxqn/gBpCoOe7MgiEg6m3CBDbkOjJC
khMIRkXYuzwNq5Zn5w0d2UM4DztwSxtK6eSbyjPFlS6eez655vnnRcx1mEPWSun8mn4jAvszw9Q2
ja8Ks2yLIhqwVT4qCyn6Xjw4ZkcOc1/LPVrJCBfrdxkwGv+8HmBjkWNLKXi5Yox2zpI+TUcFCxUH
DvfgOm6VKA0YNnXqFB3cp10RiZcxvdbm58SX6JvrJVsEyYEnzt0LEr2PM3UxZq0Iu9YKR8X4cTEh
OmaQzLwlNeGelu4uVTrefz1srKtvjKOXbXG8RI8TlP80DgN+qwBHAs0TgSrIUSkZGbyuSZQu3bBJ
+SLk6/j0iA2sqqplJIPDcq+KE2Vhqc0TKlSlFdRg9XbsyozwbmiYwF8A1R2lv5PyXJ79L7dnlj4Z
GtUJw0GFeC7iX7MsIgB/ECi8FWmta85M5pQS6LlsIX2vDBov7jFITnxlqebcpNst7P4lI41AcLWE
nEYTBpsG5h0WwAS9dpVkPshRIY5If9lSwwziiKaOSxSJYkbdKVtCC9QfZVQ9SVa9GXNasaMWbW3G
ypl59kJknABGiWYvRCcZsVSwO7zyUxSSeW4JblLP3nZlT0hcTZJPysVGIosAMnOhba/MB8GHy/Ea
Wmd6gyupL5jv7jbADjthVr1x7PQNVG9vAtUZJIva6D1gNanYNYW0NGb/HII12FuM4/ps7fL6ef/R
CgEkEFEybRerMWt1BybSHsxkzxEodjNDhh3ACloX13Cn9eezzO/EOXF0b6zRlIkeXBSwf7k5T+wI
pGpM6tgJK3DUZuY5rc+6IVOBT49mNK3zqr/TPcJu2CHNl5QARjN5GtoJRwz7d5aHGSAEQvzfsdXq
4p+tLVFVL7//Mb1fF6c96rj20AoQ5swiYlQiXXcuYQ66Y6HRzVraNBpJ1NNcmVKN2xJy/jtF9y1C
GuzTYCtEEA9g4bi7LCjuU+l3dIsq536MNZg1Dx4R3RoiuOeeB1CIiRXbIMAJQpr9BmVNV/StkBLH
ROQGKf2JkfidnKIrrU4Nl1VQ2q8sEIqtO8QI7hTuUJ2o7hmigw9UscSoCEBuctT0h0EQQjtzxWR+
7toOojX4t5RVfNSLntDuU+OKcws00YWzB4xmKGfqHGG+TO4abSDifr3HmljAQxZidUTPCgfQIkeF
/P88o3ElAESZUg1gS3qXRswmrRfQ7mTgQHfo1t9uC93Oq0uLCtFBC6KK+UTa+js5hvYUCSBIMssL
+uSCavoHnJuKZRk8N8L4OuGhQs5jSLcIfJm61LMvivRIXX3L33fxFAx7HBaIN2QJuOK4Au5U+WU0
hhlFOMI/84Ttp5KK0mDa2drOejGsMCUy9l5CxV9tRAVIpIefwds5myxC/ZCQ8IjRNgouZmaDRnCv
fJpNUjoI3XNlBcE+GOHxLumq9rSPnTe0sSw9T5RMA9AXvh/5OrK5+fXOo2t+Fs6qHhQWs345Mbfb
uAmBdafID3Nnf0TrRlJ656+bIeWa070WoyR/LmNwODg+8xONwl5FzYGqRvK2l1CLF4BHHPm7daM9
kEFeoHvfrRHRNjA668KDPjPoJc6bI01pzHdU0MPhcpEFVr4yw3dV2l911nI+RpePVO1lxgFpWing
vLmW+xDq2xad0ztCbv/B9DrVUA9to2TxSIAVViCktynL9mXz04OOHjKCDqWnoA5uij0TvWBylqmw
ALo6qqYQUNBjBLalOjldtc/yF4yN8BHese+cHEUruKWQO8/Bs9+vDBHplaNa8szzcTJ7KXgYEQuj
0YiBwWtO3y8YZObsC3u3jhHtGEC+JGbCn+4D7oHyl8VPFhZYmF56Y6lYKQ4D0F6KlIaj32a2Z96U
rs9FJIOdSjOBKR3ltGTQhQ5mr7Ff6BRG80d3fhx8BcMSH1JDofEoaiPBL9GH9meAeGzh4SMA2mdA
YcG09vt10duwWfvbDJWFS6EkuxLZVW10XAmx0WcpMsVGIfySYOHZKMjbS4DOTgAefiTz2oRVtFof
yWohf1F9+bAVENHMH7jKlN+5OClnBn7/PSoDzQx6IhSw55W4PmL4EMqciJP9M9Q5uZBnyNjll6j/
+i+RF201a8s0Rwpk5DPDluNxZw8h3DWKkJ3Ke1JVW8/uXM71FEacGc1Gmvk04+CPVooomdWQhsTd
UJO1hN4tsZk+Oqeqb8lh47PIIGL2DjY1FE3UDliDS1q8fbxo6bM3XjJ2SkN+MJUl3nnB+fnQNUdl
+wZ/Dk886Hl4edRwH2D0bp88UF551kZBmi1KL+yK/kZbDC9rUoBfMW7xnWq8173BtZ+VpijJ+bha
N1mg42dLxSMN7dQmTfaq56pLfXMBCzkT6WCfWmgeLlW3wbmMRBZM5DQGrAtnOQY7mgc7oyP4OZgI
PVsfMyZVKw8j8/LOGb2jA5U/0cvUZlxbNjx6NBYjaVjmLEr6f1qgBY8NQdsoZlLkrKG1L53UU77/
fzan2Yd9UyfaC03HVUz4tXhfA8FxBNQQxv3qQabH1yuw4S8Qc63XmsL+e/us/SAyp939OmC371Jp
GL8gRK0z0eTVmD9XNhJ/VP+V8xdZBjRx8uie+kg6VEtUh6akHcqh6whbBLyuW+GqqvbL5L3atZ/n
F4pJJ8ZHSeICtFsnxXijd/u458C59QAlLw2kwDK24CtG7okOFLLjZF+VW0st+WJQBehj970QFUDN
26TtnUm8atDYUyHMRvcOY+JxJFgAUiRGaQLDpL3o3XvHEUC9n2Z4UYDoKelEfzK3uBxq//TjcG1R
NiEzF99zT73yT71Y8ngxZfxVRPVUMlGEUzyFL/FXaSDULeTMl64ixAV0YUGqlOcL5Pssdcs3zn38
Z0DpgQjgCTo8PEjywZEXDzevmFNJ/819TxAuTFvRkI3v3SkcApUTsvDQGoRBumBw2Blx7utZpHg4
14l4DWrIRuPYxb45cEWdfWZNZ4dwc3xCCKkNZ6jHjFUhCQYhEKaGBX9K8YQ0saH+5/dGxALEY1pA
3qviIjZBTyyZT4XnDp6/nT3Y+mGRKQ54BhM+RO68JPORiCITPimpfdjtWr8NLJeygsjk1+1pr1J3
aVGthD0wu+7ksT1XMNQvcZ5dhL96eqlRVqgDAT37AlFkeaA2i2RJg4FMr7Wpx+M/VOuwhFaudQB2
4e9+RDfwYvVCq4E3P7nmQYl/3pJjmwXI993Cy2Wlt9ucunhbSl1c7w421NDOeAp0WqcgJGl2ukhL
N7Whpoe4mokTSMtmz79y/GFOFB9FKQNvdEmpv0DDDcaHL7ZQo6YtXh04sWnC95a6QIUbHIfkN/pB
r+N1TtEgK3wX5JVUlXkrhIzrGOaK8I0heWfzi6DyIXGSpSZ7D8Mc7c90vmtMA1oqNXInYBedd5Cl
hZoUIbUvx8KBmY7WM7k509UWINLtHqQbsfhVDv4hip2EfqnKQwKkdp4Q1L90p9GLPIPHJzfimxLX
fhgZK6mj+PqKuzRuFrtNQ6U5eZh5bS9M0KUJgRdw9PYgUeinoCpFdGSqLeysZWeFlvzquIBXjVcx
NrHJSbOhTeZxBfyN6Getc57SBJbmx4BaS/FtaAabr7UF9o7hDqyN9Oaf1cLAwVGlh2T3dq7NdY18
JpmIheerh9a1oVHmdCCXsTpxSDs94FjZg3sUROO5J1y+7amTkltSRkZzKAAdE+GwGoiCGI8KpqMo
Opzb10CpF4yr3XhDPzeaOfI7zZZxrZsoTuu4BZ4832GLA+2u39TSbwjWcWLJE1XIzn43o8IjgpS2
bt2iAM09/zapkvFvJYn7IibpmZElYXx8u+ZADNmdqUGECq+ArKY6qulruoOWLDPP0FK5Twmp9o5/
gikeLUzz1SRrZiZZCz8kgnl1506I/mlBxpWd6l8pVs9aZOZ0BK1q6scTTAz6EKALWu0LZje9dpBt
XQs2YRdGLl6I17prnzZNq8ICuGOlBxDCU7MvxG4U9PIc2ToGqv94Bs9yYV218QxJdmlFqpxujmfo
KiICu2tnUimqQykJ+TsAPH9SeNnBJj595qy7q0cfy3CO3J2+Z3/KdSRYLElcgJet7/OqOOqBe2c/
WJzeQgkyhD62H7eFmSZepHMUga+w+QCe3huWsUkaJ1gbeXFEkttpm/QQZvbIcrxCo96EvYK4fd5p
edvIRsGJLCGv58Pwr+FtCrz+NTC/LM1INyrTPOAFxsTHRl1T0THJg9c3ongVy8b0xQ5I0AkqCXLD
f5VRRBN04m3K2WpbyTt+K14aKM2vropU+eTCQAOaJASSKbozn4ZW5CI1ubwpbr1uFT9J36KhQtHT
a3bj/Hb4YQPaMzfECWywclnA2Edofj35X5tgxcy0PCLYNgOjbfJ/ig6ZgBsXEWag1yf6+3Czxaoz
oPFi+vBXNB9h+Yk8W3A63t61AddXaWln7mTbgwIiW8uSfqRcpMz9zhAfLLVUgwWlFeRqJ+Ul99KR
TwBrfQUFdGLsQ9nAqxlR56I6EoneoqIaaRGybY3f/fiYqF5t6MDRIBF7O3EsD8AGPNLvNo/Jy7Sa
yMKj1XITZB9SM4+2vM5pCdDqb/JABwX0HwG5MOtjcaAzLKYYeY607fhWas4JVjVawrsjFWGYNays
M415CwZ12lOo7Aux43Fh92d9jIfGTiLTQguSztXgaDSGEg34EzNL6J85GQo56szPCzIxnF+5cr/+
vaYGdpc6NoRRE9poBiU6g7zl40bb3EKyaoR4ep2EfgS1QClVlEDNEgs/j0LwYCKAVP9vFa3GU7zV
mQp3jV6RdCQLcJjVy5BKHLuLx97iETecx6KNzA5AKaDKrc3R4ZnKhq10E5TgXtauqQf+vR1m/1/N
5bxHO7Ndmu68uiO2MF7m52WCo/vWUcCxF064W6I4FSis56EYDdLv4kqNMTKHG0z+JRPpTDOG7CmI
6X1qwsCOifn8sGxlvibhZcd7eAWAFNZPY35NudNIkwHE9jj+E3o+FCRuZm1F/FT5Md/ULSijebbW
+YExrQHU9vZOidK7KSN15GhlVZ8ddSE+fkuq4LzgTCMUZONb7VFBj6gOUzDyaFNp90f5oox3DLXW
XZlmWxsU/aSeLwEYu2QQ2I6as/uXvU5EH0u0ecA/uXUd12KElyM3h8EKGlXA5B0mN5IG+P7SCLz+
/QCCR6H41KOgLaoIGyKfD42t9/zHK6unYk44a2mhvvc3wLLcx6W73uK60HsoFYi/Y4HOT+Anw3Jv
LdMbwNSRn7bEtH657Dez5rFWVlvZpRZV0DCYvQw7cLvxGnZTbht+yn95NgP3MFpRySl80MGmGpyu
6OPSTzIO0LL9ahKFotAGXvskFFVr2q+x1I8wxBNqaDXy1O6TgSN9U3g5XziDHJPkgIbSlIVrwTHK
wvDO81iYVEEd+7SpJTE5VIEGyWbymNkSyTW1IPptpbO/5eBUfmkTF2eTUGqgYvxggtZsHztvBOEI
tEvvyzJHBHARfk30S5t4lRdmCCwcae/blzZTH/VMEZDAENOzVSeMq2aYs4hrLY7OJO/3tHHBhIYR
ZBFQwjVsOfMOTtjKa61FxdQbBVyR/ukL24muNxEVQf5SA/4TRxjNx8LJWsWicAPQ4jWEWp/I/qjd
hT1EKUSEGfdPm7LEXhBifFOu2bbx36mh/5UynNfMyHUCuXJiIUJud5/OhzlHbdk8lgDyfgABJQBG
2vlTvt8wGLxcjP4SgC+7UybCrPYrbrR2uXDJroXCYh6fC30BsmRj3Xbr1RvI4qrRKJLbL2m0pCr7
lLISIfeVuQNAuqbDeCfMCc3uexMxTgp1cu2Zfb29WtpPzgOik3aTZ1OburpyC5LM6OQvIzPSLZ4/
UwR5r/AMhwWWD0+7r27lO/PlEyJft/SuM9yLrRtSZOXJWe5xD9yk0z7kvUJjnqkeneqAn9F8O/D5
paA3cn9ceLndnz7cI/eaFm8qBeSEWv2Dfxm4Z3qDkbwhL+9L9n2B8qLkP1UGDO8ONYXyfw4ioYHT
5xSU+u1Ce5k7dmaYQwFrHU6zrxL0gY3UcaCsLNnW9ET2BnEhd7rQqskBQjyIted4LgOb920w5tMD
ogjgFK8fSaNWulCNLMJIEbO1rhL94BMQSgs8lnwddzIpQrmanPLrnY/U3C2K+YIeewpAZYdIyJhM
AQhAua+0xMDSD1+aGqkf+UqRzNptB+XzgFtjAqkiN4ZJ4yvxZskTIUPYYr3AEkMSICNZaS/qcNsx
CCBrnJIG171Zp+Veu55+IPTmAUK6BhWhMUsR4jcWRdF6lkU8FXezYvVd1QzzFtjg6Fnsgiew5WVP
W5ZESb5KCLATmgsE0qbAGtpSgNzafcJHqBVtDGvHYD+CrRKMNAB8Z9Jr6wJIYfPQSkXzxaRPbF+g
bN/GdjBboVIsIsGiI3Ba0eVO51YPN+yILm0kpkPFGIIWefzVNPMZkkZGEDvP48oW93sJMm5pNs08
4hlBgNvglnpzGyf1d9ZpPIXgn2FVTN84BOF2JuXZy4iYbj2qaQZFKmTpZk8iD3K8Ad94s7yWEcSx
eSU/H4JG+DrLE1lnNWMsVRCicQjEA6SEiyfjbowpGDKn4rXfxYCLRXEpmmGyLEQ2fZS3YWkYi6k+
no5XdBkZ4m/DZp29Xnjya/A6P6utWiZEJLEVhA2Q1HDQx4uQejMg0tsHlwS21BaE6hZs1BoU2heo
0ENwQzfa3OU30jJudil6cuS6koCfjQ4vBDRIngX7XSFGd0x8/VJNptCjHqY6LJZwdpLczZTSX20f
hoIY3GILnW9xOrou1Yl5peW7gN72i5gJ4rXe7jDYPMg4NI//hdxtSsjdReChBfRXoPql0CGkSdAG
JzCTF9kHcng+w4f/xIU4LRK36ZqxDbcw7o51sn23J/qtmSwquike5vvWKlkNt7PEm0qsDhnLbJ1D
FkdiQJ4UP1A5VDLvviYrcgYP1gnsK4BU8wcBPG7CFgUPn25o61pTYyONsMOq/dXu3UUsUG9kUOIT
QpZiJxSLAhg2H/s4IuTUEy5EPx4P3opwe0w5qlS0+p/GrFDcBNuh1r8fyZ8NUJwMxbno4STsjkBL
KGFendZmxzx98RG+95bVFaUwJdIc8A49FwLuKJu3yA/pE1208D3kHdjF0fuONMfkAX968IyB5/Oe
mpcOLJpGJViBI+JcWhMFFYj1s9cjofY0Uf6Ogb9ydVckF0ZVmSQudIcVqR19dpcnQM64NFJpJXoi
BQo8wZL6iIhfnah5SLysG0CPs95PQ88PxQZ4YLZg2uMSD7TfOEJjgWkOJ0k4qh9SFuMkwPqvguBU
76lCp3c8uLOneC8rISkOHA0mebq+0f4LB/oLNWbba+dZV/NJiT407qDT5yL0zLE+FHXY3ktMpn4y
hETFDCB3CM1mv+aqy0h9TCgD/QGKE5SQPyjozH5ZokzRFR8woWA6J524usT3NZEd/GI4z7IQM3fv
B8wMlImXvdrNDQpXUcHBgk3F7XE1tZxawKgWxQQ0m+8Jx14Hr9sLBDBVT7nVAPx731aql6s/S/nw
tnxXxqUxC9FeWMS+DvEb8kUNfXsoWOsvDHS7pQoGsh8lYavRPq7oxlBJwNHMX3xTSvQyEM9R8ujD
/pSO5RVMypwe2tpNRMipVl1Hrb0calkF08QtdkTPX1MS2EIMqAXXypO9jdB8aVZzZ1Uax/heRNQk
6VsKs/ZKI9v4nOtX5yUbfTgrdUShqe+CBiwDbLu+KLvjiS7QDS5dvNhFjtMI6MDVSrZBJUyYmAWZ
nErAYi1kcfFW7EVmVVA38ISTlOu4QDH/CtFLUHonQufBlJVvi+6R2UGAbu1O1hNFha9nPgNYZlNq
yBFpJpHYjNjU5n0DzrdPl04Dy2hM3BxWhKOlxcqg/mnA+M9Pbx6AIj5dKwHGYCb422HhlANxhyWr
W25xFrTAmTWWoom0oKpKN6Fd5Bk7Z47vPcZ/WoKgU2ufD6OAz4gnnJLBuykdzBZfxEgOVQ73U/r/
3WsfbTGo+RJ4xkWsxn+z4kx3HW5wvQ5PHA9JyJ4//un+RNPHCONBqbccp+hFCv/yvrj1zUAstV2/
XqIGmu+wxTSnWj8Z++6otUvbIzELtPn2vilAGvWNPWi9BHzIwfJeqgWnnUd2w3IIjhspeAOSAPqx
zVG7MN4kqFRIy1kseRrI3CYeQMHx9yhDowF2+UVe8MOgUmsx64rExIvbKKmn5zoDICME03NUGWqN
Ok3dk51f62ftuAg+I0VOFfJ89cfFfGpgAM/hAU5iIqxzbUOVdLwGtsEMuwuQo3bjrVRw+gwFSDCY
w4RiJq+TEu2rYbabhuOkG8+EonOjPpWRDb7dqFm1B6YPBH5StEcHzyn5sBDSFLGpjM2EkE/pXWAJ
qIB9wAcwn2P85WCsjNF9m0NfyLuV8w++EKCtTCmj081hx6jXuLQtmkkYHiqo5VX909brtPvpkxvk
EJ2SJk1Y7RS2W+cnkZ/8yY+tYOfHA4SfL8HG/L6ddLRG8Jbki1zo3CSd+bACk0qPt6LwdGyQedh4
LToyBF8Us0LXNlbqdBwElKv+ykogd0mR6Eyq8os25JQEMhkIc1fqjegRF7Ww3gLOoFYtr/z8+0oM
auchjMEUDvSoYOCEWKHkCZ3S28f2auUC4tNudk4I3mlqZ5W6TJXzpyYi4JSJRgcfu+Mn1U7o5Xss
u9nq0ksSp9Gsm+kMtF98nDo0MyEXBNntehk9YDXTV/+/3In12Blsh/cINeHlDnaE/pLR5auyuH+O
beemyFZlMJb6V4WqL8fe4USZt61A5ygm5zbEaSKviL0MuNHf50A9IcqXjp7JuA5V3Cdw3IZUTw5q
TRsPxuX1CJ7CWVeiee1piv4fnpZk5ecMEkiapXfMIRRuKdNdLmrb+1oSmMAJW6Z/KINlL23YK4i4
1y9K9n9a0mWE7G023WxNvv1ue1ON/h0fqhgXcrf6ApA667ULcHU3UEPdB1J0/7I1I4ZaSHQPB+MP
hs7vZZfvmJ73xapPVdBXGziV987BwPj8HWzSakJEdzl17VCX9w/dI78sTINFbSMHGd0jSljG/t03
mT2lZDjn2TAzCqjGx3a7RWcEpuApBeu3Cuc2B+FyV5ub2VlQEe11kl4WF5tu6xRbslclfHBFLHtE
Dc2/Dq3Kw0XdPmdaTx6aoj6HeW2SknnSUT1Nu1+xhZbpLNUwedG/8+M0JXPsj0Lu2oDc5IkWfw6+
CYH/TTqxcG59CM+atx/30KLjGQMM8VmgoJLlKzPlt3mPod8kLsQi6G0yt34o3PGwOhBxdLttc1Zp
6ODplYzSrw0WEiOItundWXKNzF6IhqdNePuhqbKcfZWbatCgTNcL2wr0H3BeYG1VTXctfpFmgrLE
Gh3bQElCExXed2nFZjP0hPOPxKPm2hETPw/ykp5GPsmHL3QZMjGYt7rhQEcjLLEGcyKnShQbqPRh
E3DzFyEJOyYNCq7fuH5OqfAltjCjx+FfJtOCNwfiEP9HfU+YazTvPninDnA/UtkYZDtVSxGv12NM
0HlDb6if3+ALZKIJjO5d7aSj2vh+ilF8VKJSBaD8p/Dt2eUWkwhB0I4aSbLFIQ1XuOuJRHxjpZuj
1it1LaJEFtL8eoKDYrj0JYdk2y6pEO4+nIaZxnF9qQeUUtYcQ1HhkSYgtIFK7lRwW5LL0L/IBp/m
sWB0KUZyTm5JF4T7of6952qIFR92yuf2zoJ89Dxop2m5WgrmHTIMPyrqEOv6oZk/D/+P7wJr3EoQ
hOEljzd73iUcrnDfF7xFriTFXi2rW5YerboaR/PhK8TcqMI+tVKQiDQXbex4W8Q/LTpzghUn4959
EVYRe7wPQ8mfzPBk7c+lxSSrJmXk7DjeQ/jP4CByaoISc7vjPVhxwfw9CkZgoGxy5KcjfCE917hM
57Ah1wniziqc0gMqrg2pDuqqQZhM28VrduEDtz0AeWqqhpRq4DDzxW9gJK9fPJViafSp3s4tkap7
l3DMLm/2AlpkceiWQdsi9Kh2uwzqV2uLcsD8sgAaVICPztlWuFSahsCJ3DnXKnWxH2vtIOFtOZQA
jY5+eLm8xN2DUpnfKIAuXQ1n0SkHV6nPt0Gw6oYbOHfuA0GNAQpvqSK0Fe7JQpzMl09f+1WAuk9v
VPmdscFViGr8iazL/sJUSpcDoqIJtMhHYMCvJYN//4X1FwKLnlATGHTXaBZzS+tI9dBMs+EeMCWN
v/10ND7wyC6MjO9eZ+r3H1oqeGrzPXIVh0pAj/NZGQbtpgyTrtrVG6UTfz30wbtXEXClWeBTPsiS
WzJgf0PLUlu6cf9lVBcbXI4t5hkQUj3GIz6LgWfzaUeuMecKieVWSpvTONA3S3vLm+yRwv9QhlQN
t5Dem3g5s9FkxEL9b89CEbZtsv+6aLQoqVsxqCDdTI5Sanmc/xWtNjCo4nQD7Cw4D62HWDSusoua
3EVRvjTP2i2VsjAfK1VWMlCJCMByUG10kMaUapWdkZajkBVX6zWeGFC08va/73K+iq5J9+NbENPA
INkVh5jSjy7SNXahE/aL6zqG/aq5I3/bj9djnoxfZ8CqR9QAXXI25StxfGDkFg6zvk5nvfqXoi/W
bw44NKL8zV/SiVnxNkQjQLRV9PRVEwTCXoDUgq7CsWp3S5v+ZZiJjnKwGVmJChsVwJh4TZIduNeq
sfF7hn3BQsOYU98Q7pTfjL5tq8d1cjM9cl2otmYlgsk3m1E8b6V32+u3ATYJQCGTZqAKr97uaFOS
d6TmjzqtHzjS5zdNyOBhPIvAGcosNdEeCcIqUlPlhr9Jul2feWqsdE1cDEbS7vx/VAhsksy/Ecov
IIePHlm5Pf7v5Q2IQdBBa8w+HX4+rIWRHMo42RYhY1nskpfwK5lQAUZ5SCeQNjhLsECEepyLk3Hg
/9rBdY1eKh7OZ8+e96o0FqJM+KCFRWOLpetcS8xc/TdpmJAk1K2AIWMRQbOeCPPWX+9K7s3ckaxv
i2sbTtvtdMlHvWMF9CjffJ3agnfo14Vmh74VecHyTL/jZ9RtbdS7nMGY1n9XThI38asx0tZDqWmV
LZif+rqbF2wdHMwU4j1LZKpi01soG2KF9VuHHzrEaDG9oJyqbkp4w3ov30oP8C8w7FQkH1XcPdDH
p0iTOgY8jQMkjn+3QLqXwqzUHykwPsgWh2j2EI6bzHA3PVK3qVjGUxJPH2bYJ7W6DyNFs3CSB76a
fRrhvnSvHaBcHjE/hCnO0qFZvJeuIbnd/fYv9FdVH7bIrx60CaabtpaL5QptdLoF14rNzN6GuFH3
eO4XBK+ZKDgSxpjgvCAPjSlvYqYeY1sHa3klcafweU8LkGvvbxkIAX7/PXe3aM/pmLjGYi4Py9bo
ufGxsVTieZl+4+3Sw/gzA+5uU5tM2+WN7Bp33RU4HM96yKhLBCxJDL7qQFVxAklirGnqg6eVCrSD
TOC4j1MpQwgaulndrd9AkE+BlOZIz9WIRvkjzTxPht8TLUK0q7iXuy14IyOTvgAMXahZeSXoU1sd
bac9AoILHNdEet1Js7YEo9ByOuEu8bHQZ6D7jBp+5hoLbCW7vb6kygJIG/LqzXlzaHjTL9qyAct9
th8PncnXAUQUgwWBx4vSpjqbT+9ppGtrjXY4+cK/r/ts2YLJntbAPHlrVCDPLNJsdqGwhvcunQOZ
nWz+Kv2yCmBjZs/V5mKhztay75FtvlR4jVzrO0ahBNDs72OXjK2uT98f6WY70I8DRFqxrfqTDe99
3wCFIQwAKKo0vkIaU9XeDjw5c/khYREKAp5KuLfNMdRaLrz4aS3NimCxIPtWXpwsboXKvlris0nb
ddrXnAIDOYzd9rb/w8lPOppUmOB5U0Sm2oMfj1oRbd+OdVplV1a840Gb5NpuXMnlqxlLsAwNRd8C
UvaEVKoCipwFUVCkvXAgHKBmeMQAWQ3GH7YPK0/hd2xopyv30oIXeQY8lWrvX3EZSRaPUoowErBc
a/vFenisry+kwpKrIzZzeeoxIkzMI/S/JgebTyv0X6cIqjPAyx9mSTwMxurAwPNx8zdWZmXX1dy6
rz0OcSKqh5azZVv8iCFcoNMb/zjlIZOrfj3gs+ThnSOvC5bOZVzUrx/mOLxsQXDMzny7e3qcVQB1
3Z90mTZGX34cp6SEVARwQnH/DDBH4yzmjLxpyRy2aWqdKAMgAHGYiMNh1hOsclB2Y0Mjo0zQmb6K
a4v/wuw+IrJ7TCFAbO6IiNboj/5v9P/TrN+tqmT3lYqAY6byK+t2aYooHV/6FuKxKeYUdpBE7VzN
2HXnzaHAzzA4BkS2aCf62e02ICDyCN8+vbvvzM1zh5yO9VoH8oRQePVT3rOdr0b38yCGRviovG8n
wpRt+WfC1mnFMp3Ba1ab0WBy+uZkk3IYxs/SunVtXHQzx+Xr1/zfHnGKf/iucVoFxexN2GIITwCh
wbincfOhSs+uu3SnBUWElCcZr16Zf4NmooZu3rM6LCP41XDeAn/sR07xcS39y7YUwLfDxRz38mmV
Dk3IXc37QiF+6mPkLHAdCQmL9VWkdqVoGTpsiHDbVAqOagyp8clhm4g8zL4d89djVBJcGykov5QS
TBSdvtKkNul9N+AJh3LqbKa+NJE4whIfxk4f/bk8uphOMXuSySXJa0UMWx5kCCIoYWMGRvn291i4
l0tKtoZQQ8Q3osCIXdoAky3MRdAjH+Eq7CEsccGOfb0ttqm7GSxvquhEpojz+YNHlWMVzCQvPWKk
TcuaavkQYIWViEx8ADTokc2UCsBlzlhTWEjYbuS5F9VxwI7Nu3QvUhGMoYn5Ol/AEe5v4rSsJCW9
3vYU/z6B2sLDhPWIjwn0P6nxLUf29gyljjez7f8Gazyyf+ml8mKCRO/Is/2xjhqShjWYyt5cRkK6
aAgyQOF0qIrgoOw7y5DkD++urqS60X5xXXarHxJzxkIokSQBhOYSGNyan16wVhrX1g8kwaQ4CKg4
1JlZTiI+FMWtN/Lv/G+AVXiScgMYwWe3UOVmZIMIQtWT/PKAe4LeOhl+W7vJ9atE6HYLfk2QO5VT
s+SDpKMwNz9qVHYd+IZGNXf/B5UfFMMlkBTPTZAbggzANpA2OdEKjs81hRz1hXqAlkMJb+YJRebx
SNOTJ139fFcrZ9wigmV0JymV0yofTzTkZDsFYAwV40t/7prSe1SCR1thEVYrn+Xyr1PmsS7LnfFy
6yeZsLKUdQOU8KPLd2sHyVoYBUCNZU2Af9FsBEY6EwY74JxGojK8KdpemAWcXLMAvE/53UxlDI+4
UQDYwh03W7+XXQa734Ae4sUvc8YrWGoYevJHB8+TPMA/8pgbopCG6UmaT47yxLWEIlgIGUOoBukf
W7TEPM2p1z3sNBPONXKwX0qvXgU0ZMTXUM7bnqCtRtiMlgZoAkDfLI7BTys6AcUSfwfIqKzP2omP
UtxCc75jN1mu4xkV5qTuO5+ZxvfBMClexJcwRNe37ANZoF7tAyFdx87cKCRfwbjr+3eF2U89eAs+
FQdVfkSajUHmt8W2O6pFUhU4YYfl1wj6vZNWJanECwL0KNpsCougaqJ0P7qY62GLHaknI76VGLY6
oKMyEfv4OrI+IKEIwg4Gci7ksYhWS7twhcnkjAmmHT/jJDczHHXOC194VGjtaOt4emlOcUpupbj/
o93pG/urDT20FUdyD+hpTKRzeEdfieIBVW8XSE18hM+EekZH6fu0trpKrivCdj7mvO0QN+NSL+c/
RyfCujk0hIXeq4vrXjziUn6z+378/GG2YyPOtlrUPBMWAyB3/ICB2S7h0UE2rJzyUnoDTTWZc2WG
XG7NMqFmaWA59BOgQRyHj/w3FSqHt0ZhhUtG7L1/NiSHX5hfDMnjWJUZts1pzPRBOu/MniXXEDH8
3alFjo+tIOr3TwdPRT+Zy0FCBggJiFQAj1xcGjv4ZZcueKFl2P/q7ULBcfEVtvg4ySt+en+N1ug7
du5HnKmenY1lX2vW48Zqq5FVTJ8kVqrZuHWIpkCsMibiEbuRLey6PCYbPWbjR0oSMlm0XLW2eHPb
BnOi20TmEBSLDzae0idpiyFtolQUQ1DHFrL7DFKXbkprnVorPADRsbz3AidXpAUO9VL1M5APHqEf
RxvKG3Oz0MrMlWI+AyjwS4BII17d7Q0lkyI1AvUZYPHmWJyW85VxS+IR4L9+9SFbIj19TdawgmWG
OJfzdBxHOyKz7voK0ph1qXGpuHQD7GoDCPQy5gNx1uYKz7wXkSsJg8tbenGbr3eKRqEbU3pNjDvQ
aVeoeSxcAOdP3lXl/z8FstXWjqu8Xy9FiFzBrwBZtD3fRkqUvdypbM45qxYpJGKDPIdtz27/ropO
dtT1J+sRgfc6tw5ah/0Ehg7SLb03OIzIJY7up/D3B2PDh90Ro/FCXD1yrnw/k2wwk/rLmJYQoCAz
HtCfW5n5ce009IyMHKiy0B6e7iLEtKG4M2ZJ4Xg1AHMEauJK0km52QpIkTH4p97yOK7gyNXophAG
wmlMLRl08SiZ4pa1htDbvv6bQ6hDO74pwxMcPE2N9ft41wFxcM1HBTeGnAz7+gWHaXRC6eEBhkeH
YF18MqF7qLji/Ck94DazCjFC5M2OtFcvQmkcwxfC6FnsW4zEb7t86Xvgkg+269JZOUo/zZK4puex
jMdL7FAR3kqKxKBglo08f+sqJ7XkC3ZLs60uP2fYqwkusWxm+F0gbdAZoh/tf/2xOqlTXWjIBHLy
rBGurv5GK6rlP0hH53WqDCPNeoGgkPJGKszwFtwkneVEm9hkLROcVf/EsIcxZRoQwaX8Z/72oSBb
rni6GhsJOCn1udhLl0gzITowf0zhgnjWber5LmhoVRCMmkhBzvfzGJGGGY5Hj7O/OjLBH9VRZMdr
Ej/jyMADgYYrF4AizY9/THe36XNIWMFunmxG3LPGQoHKxi1o64ywYmZnG7HS8uvMJsoIwf9qbjVI
f7Zx15BfdW6odRcGqXe78AsghgL7UozBSMA6pew5DPJwXhHxQS0+fHNRXeiZiKMAJk2/mj3mZQcc
SMPvPUK0M2bKTqCuWNNaB8QBK2ni9KKzNnf9zm7Hi4Ofs0opEGJll/q5Lmz2bkidj7dWuvL2luMw
RCHXaB+h5BruyvDjNscmK3l2KmnB1Debv6U7C5uEBlg8vw1bbFrhUfEr05LZvqMZSh7lFKVAvI3/
CXyH31Wit820R/EYk65YeMDnHYv9b+xCrsK/Iy/lQRmTjT9u2aSGThLrp/Wz4OSZWj0V59CI4YEs
zKR2dIf6XRD5a0mpKCt+64/HAol4+htZ42NstkrcNYX5MzMWl3AXRv73eSxpvYjApBs3RB22fBMn
DsQ9xwWtVru/H/l99hC4w7INdQDMt+tGN5rmUZvunkwDfCF3l2FRX4xvmbYL2VuNAN1tiFmYFNPW
9uubZFaBZMH+7YvIMKbGbG9BWQWx0em4I2GxQLcWi7f5z62gGweNaExAWfPr9YIf/Lcf5AI566+z
GfTkzsPX4sEMunIWOYwJtRrqlW2y3uqCX1YoVOSM2hHSX46dcKQ7bjbHXEj7bX7zpBBHkUUiUeq8
YN2OgOp446SdxaI5ahp05XvSgbP2iBBq6UoCHKgmNBCiKgFHzxlx9PHp2EGSv98qXUlBNogPG+6j
n7TxpdiHvwrrk8XNrMQL53kFoH6cyLgQ8ioYxTLOSGgvN8ye5T44bZqt9tIsKP00JA/umqEhYQSQ
RUgaoWdWxrjb5KKpjWnHh3sLifQo3CoNR24Sirt/8n3uUC7Q1XSy88cP7+t/99AU5hkwiGMyipDY
OksSUHP9IxLM4xIybC93ER/+HltkEdr0569TaE1pPu7qB5c3epV/6OnaYsxZZee0jcn0TiLBFGZn
eKEeyT8HD04R6rCzZp2v9+rFvcyHUmZ+tcZECopgCjvImpsztgblLVyFW9VaLtCNFiIjhIaUIssn
NjsPhnI6KwO1tcGwRgCsorEBkPfddQN4fLAyNqpjC4IwTTU9BzV3PiYxOZx1CXoHK6UZhPh9fDZj
8BvcG18FRYHfNzOV4n5n714JrrK5MNX8mbYsH3byhpsWj8b4c/69zm6ZntsYucc/1+53FENeRJeO
TpyKwurHIaypY7qStqLzipcmMsZ7SXr4FiFEdauEmyehC5e2CrWApC+efutxfS/wj45eWJhOaiwg
XcNA7W1GBp9tQeW1rdrJrXnvF1bdrlSUxYPmWIHmVqJjPEbDgMVE5DedzBL93CN6XYwSVxoj/0K+
CoY9WaHsddRgMnFFFsC3xF4Ut8lnWtLKI/RVlmNAfieM/E6+oQ1WauhyvhtzX+Qt3qHjGFh9UU1H
KxtjgFNB7WzHPjdoD1JGDAhOzk7SAbPE1I35xsveVDcB80frIHdKtZyKAVkltAB2iR4XgeinHF2Z
dpxWdM2jUodKfmAsPXGByfuyNWcPmGnbnjU/0hrckQdqLl2F0L14N74nt/vs8jTalZ0OUHO/uQ+F
jxkbXm2wvwLEXNzBQiu9DfyeDTcxez4jP2/S3DAFB1QyQUxpwFl6qG5A56/g8GenkrZLVw4PN+O+
Hp1SPZ54SXsm1nI+PXY5t+5/16A0QhepPeN1ztRvKqTC8knOTA889KsjuBIm3omnRYpmc8s5rzLO
DtdiFWQL9m3ZQey6KShRZhlpYS2HejwKE4dHgJCUKNRpwnsMdLNur+husCBd3v6nS3XYlqjlXzNM
qiHJFa7h7UdFKQhv0Kn6u5/Xz+GYRaLPLvxl9/7eZ0e59IoLLeiQJyvv1wWplLgEZxk/TiPPlYEP
cP7R2OAVGPLEv1xd+zB8Pit+WMewRE70hGTH01RTFJ/ls8BEuRw5VegAMRYouRtW6aFTr/rD4Mo6
fVf9LDUrB36jwfJWp5AB82ke4OHj4o5p04nytstxRZm1WAvbTxhPyYnoFiaCIK6886uwlJGdDN/E
c0pDNwMX+Am+2IEAc2LJx0LVOznTGe163O/yEFsQw2PyhYhlwKpMz0gPgUUD7m6cc2TQHvSLVVjh
eYZmQ89GhvxNQ5268ab9VqCCPI0os297KBsX6/e7jjCJa0IeUebhDzuA5DBR1xtVdcW/w2R6rBVt
NpqNUmYKC8qf238O2OKnH1TuA/E1CzTz75Jxj6Xkf7eam9+6VCGLhV9eb9H9r02I8PIhdMclYz3X
L4nk4RD/1DA0G3e55weV5lwqZWLcglRnGqqiyg7shqwPLfy9VbbuRs8w7PL4AkQuGhk0PNb2y9nA
1E5UjwBTR9/GQKo02rtqYeYJHn4NWyWFyQiqM/6FHMVPvlTb2vMPwfVNhbr7GOf89x1oJvIxquZI
KOmTfbJRmfDwXVK9aVrSHFTp5bWambJiRXHk9XQMwAWPQoDiaA/2X7BcHvMEvYoqWEYN/pXhI6ES
wQNMGuJKVWYVk2kzBF9jGS7pNO1xxL75etiDEkr8I7GeX/zuXfhRR5ORKAeTPsUuTIVTzG6DO0p0
nePiVaUVVPyHoGDbhyM5rTgq/fIbhTZVygc4kceaeLA8FOA0rx88gA6YNkdI9vpxuIlsjRCat5T2
ev8LwLcoKFmkJ7skriri9WJDlmSsKq7vdVGdQdBgD6nKV8vxfoVdNHkJbVSXEKyUIZkyOpJgbcuf
/Kb1PpWjJ0+euyci0ujs2WGua0inMZjcEtE1I3cVlLkcLuzNuJuWwmwJ7Dan6Q4Kltuvsou0YVZS
ejp5/+VhCDaHEOCQCXZqexgj1YZF7uR4ZECwqVj43t2Rrkw/FtdyoJcy+NaQcyyQiNnAdGabA0XD
f3Nt9ncGe/NdnKcseRdSrhOgxIt9b/B4P1/VvVtcf/N54qSspSwMxOqFi9EenpHsFBC82OjQhfwL
jsLO/PumZ9fCepy3uFfduWzPf4sPR3WaX5e4t7+z4YwtoNvw74MQ7m99vSb3QIMq5UOA8f2b3aZD
kybBklaX2AUZko9WP5/mt/o/9ATp1ZRzf6EFB11vKNotqW+isi8Zh+2RI+Ic/eAPYAeDxAR0xKcl
eCdp6nkVwuidQZx9csWzHMX48bgnu4bLJ28mVOWTG8sDKQAo3TAwPASNhDOxK9egZQTui8rMxGwv
BJ+bMcSQgbx5BxL+F5/qhSXtEEjJlVeDn64GDj90teG8V1Oseh3RcjY1gmNLdYoYy1qKSjiRWw1O
YZeOPDtHfZ7kFZWz9kLfZqHn81l1Tg5BS27q1VCl0LyVpY9fJRfkc7XSAUMS5tzMiIHaFb4zbfkh
UjGmO4vbCHMkadpQJYbFvRz+D3C1rsE0Fq4/ofc1aOohwHkh1uTBICRcB1qOC3xZ47BLJ7znPCZ2
RlcrPBvzwsptA4cnqhYOrbYDZDT6G2FVY7UmAaaY1wfIQBOr6zJe4m2ylNoq8RERsDWf8S4IolKU
GmJdC+2ECk4LFSpPGqRSufB8kGVvMlZoIXWsQXT29sBLb2CM7GscpHtzxBekgu3IRjRc/bmUJT1C
xoaml/cY1aBXd9Lyex96RCX59ERvEr/DYzlfHoCdUURLwMrCSgiZQdRc1w0CNVMmDiw/9pnLiXVP
NCK3G5IYhnZuHLb0TVQAtBeTtTZbg175rUb9N3ic9ZyXxUeJbLkN+A9rPCO4tL8AkDLDg0hjR8YB
+8SImuF8k+NdRwV+RPZ5YhPsnw9VoCu8n4xIbqQRIi8kEc2ujtFSTAuplE7vllbNiFFgX8pLmOVA
Tgi0MeX3PLSlG9bpfPaSoWAEcAWrMRIs3WoUFJN4wKCP+rRfQOdbYIVNxdj7L3yZb47EAza5iGRP
dyndPSHzKIk4J4+unQSo081hCHyFWPvzCrjdiSzqtPddIHgrmClFDjdNBmA4AEbClhSuO5cxwGDN
e/9TbSEImAIjt4qBmEjpJDt0FXVYTaci370QO6VQASrtbF/ec9trRMceX1v65RA7r/FU4B92TN7L
k7WM9otDw4hPT2abQ1EN7P8Uzx5C0jhfD0v7CHd/kUEalOfkNzwtf4wGYC4mJ+vQMvY0GwaCFBlX
WEel36Ef0WkrYJlm+1Q9lIWItrpftW5tQSb+KPsgpPJLP9CumbfiT+xC2Fa1lhiJO0hKUA1+N6Hg
xAC5Kw7yz+VkBAzqAUksJVBPATvP8wwF5RpH05iGnyEErhfONFTBFP2xQSHeNnV4nw7Xmvnjx06l
lSLbL2jr95jFQF9KdFoAtEhjcQ3BDTPoi49d+zaPJJNJfJdcZl3sKNndDHBNwEJoUZxz5lplZS9y
B9eXSHwg0uJN/g/bqz1LG1bY3+02uXBT80g3EQOIb7jSDHYhgbGskYJRyGsisJP3OCNU+mYnQf88
uN1DsDSoZTSnWKRhu0B5L6expKL07i75EnZzUI9MtPO8LSM2c41CbToPYuyYk381faJSWM1MQPHP
4XD4/FpdcALhPtnK1MIwCUgEtjGP/nk9p6wg0Ps4xpJWBq/2mQ2gH4Y8qPJwKRLep0a+KbuglMXt
gZfTZo99xMYfCSi1Mk+xOEVOecte9OyIHiXbSvf2Dw3pTJS9Vf9OwiW8vVk/S1LNKpsFv15/cIK2
lGkj76kQvfL77FDpa8wNfAlQgbXnlvxP2XasXIxvEUpcndG5DPD7NljqyOvFQoynqRl4+fgiFtuL
GA1iFrDFZozwThOJgV26dAY0qdx11JFvfSNrGkWFaXEQ84D1gR63d5k3/fsLOV3jWVHcwB9H5Fhk
/8j/GRHRUv8w+Qn7ZHpkKnlmet58ercT9e6QAblK5T6egU2P38r5jlRgkiv1/knGkMrrmfxsX6RR
hJ6YOJxZq6FXgBNqrWgGCQU6lf5t8ASwkEEAxY0l7ZzpEEenyFj046Q4UE+PyQj93sxrZxuJJkhf
a9kd6/vLVxPPCDm595HiAoyxF/u+SVr4ZGDe2ebmcKlrWp2BNfmcNK4aJJFoK+rnE+MkEzKpntKV
0wp6oWM1jQJMTYE5/rW9iogFWxbNrwLlV/c4UUvAIiRAW/3JhfQnJdiRhca4XMXYuTePACZk3p88
COpVGqeeP/yvD7yZDZSRNjL0h6bhnwOopEj4t8GGc4d1LB8eWjVaTX6U+VS6lrOGpZ2dh+CQulpx
LQklm/mN8UcB3Ni8RG0iIAS2hwJOfuW8dYg1V32EAWV6M+uTAGxosHMyGapoauHL8erQd2diwXYp
2S9lm6eBbG1n2pyAem/Arcp6fN+27+eAhYCTGjcF12MxgUTV6dtP46T2I21O2Tz7axCo/PFkhrf5
L609ApI7CyTpetRR5Lma7eBhmt5FJvy97KImvbl3O2uYd9jpR8xfl7s3CR700B+NJ+tgjunnXlzb
T0HJxK8BjKNKrmCM/JDDY4fz1MxtzH8/XdPKin+//t1ifmoIeSPvyAnss2k8zu05+ssjgeXzcUnG
MdyrKDvlAiOoXSL+ZJejoD6ZJtPe5qgh9i7DVSzKZwOxBDQNj8W3uh7VAMmRyUYgTUsO+59N969N
zFqp+zY/SNt5Dj7Ex2Aezm5Vo5xXCcpOA+XsFxagQ0DHhAUMPBez5T5U37nbDIvhbnVge1XkDU+T
F1PsP1/qb7s+XEV0xtxtfOpJKTFTqxdp1+pwzF0HY74DwrEa3IXYny3NrKyEIxtZ8V35S9S3Pw+j
okXvN5/5xIPvWyk04BMOisMduYJ3lugGs82UOn3MHrGaP2iS+1EqH1AmZcxjdIU3jnhU9ZBTkKQ7
5luum1sI0E+b0Qgal2+t52mKJZQPoBS2WFSQkz3b3qptUxGamqgJBCZjsIXmVptfh6zWFdq2sYPJ
9vvNLlJXKshdA5ADfvXWFTV+l3/IY9MUzatgP4IH32izkbERMMi+z6jZq3wvoW55+bqN5IzOILVf
taO0YZOI+6VVxuuCJLXsCvgw4rZ7IUD06lxsIeRtkJV18N9gVOmmCLHR+w5W17XHNO4GsQqCbU4u
aLs3ndjxsURlQPPvU/408i883dWWzYHc7reL2MYEjEluv6yoMd1cZL/tB2zpEYi8Q5HzUJQ9qAFr
DIZKuRNjouwH9Bvxnyln7i4fj1ORTsUzL1YTOI3SNFcXIO4F26QRKxioO62+41Q+9MDNEcWgznjf
tjGMFLzsqTFgGbzM/JyNe07nemHaF2Ir3mps2JKOTmKQsGi40rbXeF6WylGUU9O9jBWsiOe2gKhe
nR5tctPc3V766wULGiT8vTYhJfJtnuqLv9CqG2inU8i2/u/q8OBiCiGJvNeZ6AnPimT5DO+R80Mb
iBRd0B1/wZotxx8qqwS/VmkTVMPo9LlQY9v7lniZ0cLWKOAb/4WgX0KG/v36I1VGiTayDRP/cZYx
rKQ7f8fF5hcvD0HR9b7X3J45ijIR3WZRjD0urMZa/W7ZpURS0FAAc4iSUtUSgm4pSMVWs3ArZ8h9
PlOH5K8uwE2te/ZnGXk+z8WwPFlJiJtkKU8R83egqySRaclGshcHKuo7iN4Xt8SE8HZQF4Ljp2xE
vWhE4aRfVtuZvLgijBQyBNuHCA+rgbAZF9m9OigytGZeJamiy4a1E2ASFrsfQVyfHAxfVanzMZot
vFOP/SxNxMzLSgFizxQDZ8JulrPrlNz5Av+oDwtsRW7Kx72VV4K1C004RHJ4Br0c2eJyYReOPF5f
V9GNQjV4NogdeOyd6B2fqplrwz4f9gmGGeen+81lnNOZcjpg7xchuzLvaup41DWfMZFLu5qvv/bz
g8e5z8qShk/L1x2shl2AnWiPFqEyfftvjUDolZl4Jf1L6RKe30VNXZW0gXVgBJcj6KLVueFA39mH
3+7UIqhenJ1dsRTnFQRPQfq8vTJ2kxqU2vJra+DgORlbXluSjKqkGq5hI7CV+PD42UMWNul1rCyr
JjvbZxQHCdqcP/vAV59ejk374m/Q7CsWNXYRdkxseE/Bj4dmrUnR4fqXurLgUu0pc1Mx6DGk71rm
+Dbz31VET9ToLfXNk1JveKd18nVM2VvR1WtkTVHZHpB3gPXOt0SyoMJ1wNg5ATm2THwjPmuQ1npV
31LNGbhuOhPHkFCo+yEDthgjxe/mYHhcwuN1whGj3rc9he3cnXk4jeIQgX5CuppvCihKcbmclwGJ
e9wkUKHCFUSeSx+OtjVp1xu6i70OWr79v7QagaHf+bPvBo6TcfMjXGUIazHrAzXG5q4Bz5JiAOmK
/mM692iMhfHwuS3BBJs+wisGlanr46ynxScu/wHqoaCpz49PjMgadCOAxBI/OPLkGLrZc63NwjZc
t6IbxYeHRIqWpySiorfSCLq3b+6v8K4mL7BYBcWggAbW5EYg4zeg3aEuM5rZgolXw2HNb+u/KKbE
2Glh5SRNTvbw5Sx3SzXfdQQV4eRq7NXu0qM3OHf2r6gQULA8Rh4jJXGi36h6EzWqAxs/IAmQo+QM
k2LuMssEbnbTxADy79Au/VRXa5+SFk7P39yesqSEMmbqF00Le9ePA445J6wN0jV6APW3A1om96i2
/q40Ro3LQFTpUqdjffLlVIgIYG233ipDGM2CZqEeYp7qdoc6u5UfNWwrSqi6kvf4eOsZmk3xkzeG
G8aOHqBR1OyuGrjote4F7E9pFfGdbrAvJ2eF1SNLLitrfV1Lb1w5H8AZq1ITWZbyfTtdIEGfDenm
KY5Qe635gCqqfVnYqU2mLbBzKKjVx/kiHMyce3ecgukBIi+8nd089iQXB8X5ysf0LrlHV8+r76gZ
nUpQTJ1LxjX0VeKFXAkivZ21URN/oBw7ku5AX5NOrcFBoTw+lx3fB5E/Au71vKKiypO3XUyBSKzl
FUjRtyakPowwKu7VF2tYksWaapWnCSukvB4q1hnHgQ4Jq1ujeGt9bqUq431UUEiAlKqcV/foGmIN
yv0qsp8hMdKpflvNvqa8lWjoZ8yO9m99atDj0NCTNZTixqBzTI8meCWuIQ664J7/cES/N+yOaWYf
tU3tQ/qeve11CfvG4I4HigbzUW42IQXAMluHA7tiMT/9erXp+Ptp1m+vjHAC2VUDmUqqdKIrDTiB
4oQmSaFgGa0cgAshVrPaydrTfnuFuNAvLth7GVLg93GcBJYTm2jIoAaD7umzVisySdj8QuD/8NeI
U/88vwtXpV6UqNOATmHReQPCpejCzUA9JgZCmRU6tRkons/EW+9XtEDUJuhEUGCJmMMuwAeyfXBL
WhGw+vj9hyk1PIzfQ8jWObDDj14UJV01k5bUaTJhivmLYhpDD1FwqCeCA0DbqKU3VHYqYO+qRrNR
Qc74IDENZRGVGtb7rosv23hA6bIDbiIl/gUPMYYjKjI8wriW6SFTZnZj/WMXKYZUxyPVLGAzXBEW
B/BsR2oVUakHMwQCajUT2SD9X/gTNiTdwqiSAFlTx71AJ2x/Mju1um6hK1yEqxOsQsXEPGrtGBD/
RTCBSOqP1+/CQpfWyDnI0SSc+fKmV4ozbM2M52p60TXB4Q92UZZttRLAu164ck8IyINYkSG8cuuq
Rt0AYtZM7/3krWZsqUlVfLpbLNCk3TgAPNTneyZsuyUhk4ELmmxGUgi9PtLn9P5F2YSJRWIS+MuO
ZyMb7UIyzEmX+ZfZV8jXxXUP+g4xxPie4xdt/LzpMH0pM4MMrkl1e4Hpm2BR0hHBdHYbfs3QZSk1
19Jj1FgYYpTVDFWsYeYD7H7891m1ogKwu98jvdMZXbF7liSTZkT5vOOZbxeYgwlaEy9TDDugC2rq
OqqTO0IVv7byBjkb21zopb35z6v2+YhB/vOcA11WkClzwR4hbGlsNoWS76UXoTZ/OyEAjzHbdyKY
msQQKsQR/E1NYGHxKuSld221EKdkeRZpmzOVUDhmF/VrFu1aZBUZ6Tpw1ig19MtrZLxk4rzsIf1v
3hvszZMBL+RZNbRPPKIDNWdyOrGit/jB0ND4qWdXEhJPc7m6RadqpRL2YkYzz8i9SLcj7HgRsBYq
10VbBMkOarnpqdWAM/XBAUSbq8oeYggHeNxtRNv7vXRBrjJ8PMCVUVmn8qDKOtjHkl4zDrS+AlzT
ro50kyGsc7E+TEo0QJom6AmR9tit9MeQZrpvOmfJbAVXDDSLE/Tva9nm+rFSvokEnMTBe6aGjob/
kjA0clMmaUuJ/M7FJ5EIeY0Y5lLdnzE1zXTCIi+Z3pEYXGIbj1yo4iEzFgZVdnGb+vkNpMcdN+0p
+mYEZD9+4eFztX7LvPW4aw6WcB/wWW1gAiqMXkXh886VUU5vli6uLt1SCMsOBllMFGYorUS5E4hj
w3Kpz1nGV/f869U6ug0H7Raq44UakX/ELGlGixBNy2UEcaETSVS8KB1I0ZYCz8ksvCSrZOjrYCQM
uuevIieELtY02YcwfvpuS7Lui2uyPNq/gFikOZxe3Law4MbYVFERgA4L+TWAkKWMPcgzsydyZlE7
FKo/Bo94Fj0kCQRXM9n7DnJwdvIDYgdfIsEzwil1n9R3JseeFLRkHGGqsFdsRiMHsOMiv44QN+J2
AeIOOn8FAWPMx8WHyB3UH5lYLNxX1kTkbtJKKpA2MmUuqrv4JdNgYpnHQ61WwzzHYCejfRPeQTQY
+HB6TRIJRPa4KqH8BUOvd7f4D9B4W4VQMz+W5sKeAD53dFiXZwW2eQDl0wDCt94/2jVQtTuvM8Xm
GNkr23Kn/yy/aAOdBnrcqW4ZczWKWhb6nH7vI9I1Q0jo0O1MjLSfd4McJQMTh+HhhzvwbnB57ipF
5yBifDKtE2IhnmpdqVBGOvD6oTuXCjqxFsE6e/W8kxFQ4G3dc00/M2pIRy17m6YqRVRc0KUuguRZ
GT+Zi194do0Z/VTIe2AfwElNBpeW9e9/vULQgeXeJs21nIijOyDKoZkCnFoyVzpn9yrW7oG/MJ2h
VkU5umsqMpO+yYmZgVw1CYJEztsOV5hCVwrcI8O7tSyjzUINoRdcMsmv61pbrNLNgHhCPMUKz0iN
vMsgV9kGmLOZNDr58e1BMPpXBELVOsMPJ1Rv6bYnJ4BmxBz6JX+m6Dv6ftkeWIUah/xy2hdPigt8
9QTct2mnqt5o6w794rHlKVXhDz759+8Zfb61E+xLIfSnHpNOw7+UGuuw59VCa3n3vjOmGgivI+jn
8cRaPhSt63RTI0DCM/uJ7J7nGJ4OhpkjVVslA3SeSBSD4fnYd7MtzDZh8cdrninb/CJwDtf+ocjN
9MIufJdFBuUgf584LTqfCfXEilgBRORXiZMszyPDyzlfPH6kEll9y98aCF8Bhhi33EXQIG5eM3/7
dR5fRm2ywGPHggEY3NL36gH2OHaxXrWJn6xtGy8TnfnGhLmcRkGTSs76XxMO3x2Mf2QjL9OsjDg1
tTmDwNqSh0mKRlzQyelmnVN1QywK4FL7eM3e0/nIncRqyrYMsObfx6POxRHmH1X/MH2ZhQnR1fhA
wxZ9u5IoMQ+2IHucSoghnirfIE+C+qEASn219x4TiG8NFLRA6wSTMLrtxEIkrF9gydKM2Re/UgDM
mNmzW+vHzjsmv6st2cftOFABuK0vJKyjbKV2OGqNv71UP1LT903YwDovcATsnw9bYyFiVjP2Q7qp
svyQZKSozuWs7LUSbSaS8I8FXS7txHh214zRw4YyB2DKoWVElsShab8PEIZJtJ4+Xk5MNT240nuB
oZKQzLk0sQLsVJswRHqLAqfPFYLyhZ3d76irAlzuBO/i/STyU6v8fEcyUpqT1R6bJgqwXHAjpBMm
x2+C6hQ1JAbZHnIVpQ6QJ8R3xuhN/wwh5QevryC0zxqRs3GV93ysd7Q4qp0duPB16h6kR71qeXQf
x5U1AzEeBNuhGr+1yZVaX8RvBxPaxj5UpwUD55/4lpsAPPKzWED5VCpalAN2Tap1e36NXFc8b0EC
BOiQa80GTI13QXGP6/Z7yT7SGmgcBwm7ElsPqRvMtOfvnIbO1Wd7Ll8jxnlMTb2NPrTgD9/Qvtqp
KhWwrLtzFwgpBZAqQhnRJ9tNIeceQRDbTQoIKQ7jBugSKtLApG024E/F1Yy8U2hMlp9lgiNPLEil
Ykzz5rAwdhpXGCe0iEToX7QnZEKAmn25mxijAXLY0CNGMARnNU8v84qcaOEN6AZSL+kvM6/GVLqX
upp/gRxHggbSKU/6aZDFTg+LM/Ic7SZyuRH6dlVJa6umOEB3gFVAkPcj+cbt2MZ7exv4noi/0dHY
5GWb30jJKXveAqjC5opnmqHnVqlswk8FJzKlcHx0WqSJHtnhA/hEfZevIiitghc6QswCQliAMuyp
W2rvsJjxQii4HUiVvceoDRVFV73MNkd6lOwIDlMWvIF3IrKN2QiHJ2qAvNpk2Etgm3ZrK2SXpWpb
4drt1XWnpchrYxP/RcfqNLPy7oUIQtgoJ9AUi+25KAWKlBBsBnD0ieMmTXiTrC8GnEON5h9mDGFx
cNA78lH7e/A5RS8B0QiKDKegWcwFMOX6eYLpe6WMdK5cOeRna5g9gUt3/pfxyI86PkuvQq1WWy13
BsV2q/plmK3DUFlTHzGET8TMVBnjRzLgmZHF4PHl+i5vArQjo3NIR7+Bd8phF/CHlhYbopJNsBY2
M15ilSoWhAN0iuGDrYbssXqOxAWUQFqv5shzPelrwrtZrPf9q6JjUphB0uDABSB8MRUKJxSs9dlK
UvGQ83/y2Vq0Y9N+cdMsQ3XyQ63XxsPUNPfnd6jmrpJkaCZ8CSR1gBhCEhXJ2B9jqcFh0VhtResk
y6HuZPk0Buyu/bODnCvQIiyC9bqPF7siXu3BleM02qJS9FeQOD/hFwSLNE6i6vpHXoe3trfz1IC6
DWx3BZIB+9Zp7yVhON/jBJTsic7D3a3HPuKMq7SLekN2xYDSMnWpMGk5e4wCFM+Fxev0CMFMvy3P
Uk21Z/o//NGjiq1wU9wwuu85NfbhjRUQvI9FoyAoZ1dlDUcgQHQ1c2mFcb0SKbBRJY7UnhISlGzv
LEvMecUMLqU9gEH377NpDtDEd77l+SV9r6wdTrwQPksD3Ow/fixy5gyzzNqyBpZBiBWsyYGflikj
hztV2iuiQFNH214iqaREs3QhHZRXoKfjkfNUY66dm8mTwqB/cJ47CI3NiRnDhojH07ghicQD54mp
45OGJVRlpVizoYkQfxg+R9925iP9XvfKD+iwg/YLSgTTe6l1OiB5NBoE1xrRyfP+C0rDKOSHFJ7y
OXeJ2sn8eSj6amrMx+ymD7kA5fhpKrFrhcD9kB9pxZ0bBSOhhX1yQaAy+sx7v0r7pff63uhRF+TG
UuqmLt0OfTsbNakSKYGaZVMvou6yhdP1mrr57UNBekAeTTBdsSuSrXh21DoEHODkDBkiow/KzBbP
ifuYgSEs5AgxmkvUuU7uVQUI1QN7cYi3AnOEJPrMSZaS0zc2I6tEcCjpzbgSnOwRHmfVe2OezVio
MIcCU8kg75nPAI/R1MuHA8bIIaun7K1EyYHEWsMyREQCOJUjt0565ST7fHPFMit6ulnWYxfNv4di
PX28Bbg5nelw9KoVNEeylU1eiyh19vDmUVyyUyeHg+oKlCWZL8IIJKP/Z8NjbuwgCwXAWospe1lS
j1CUBk5SI+C/yAn/FKX8r2i37RisifnIAG6ARkhSCm5tDuF8GQ9IYWVHK1IeOfpRjs0bEoUFC9nQ
wSpJmwiDwLm2fw/CtrsmwEH8vEW9PxAaIHdfNVOybitRFr/hLmWMLv0U4CsN4PHJAKA/UbMH56Ak
iCYyTXgs3Dqu6NaHwwpszM5AOP4z7O+jf/L8gkODCxoYaeQHII93bgFZ3ihmePz3BRO6KEgTjh6i
VA9yFmt1IFjlwCtf0iqZub8HGkj7l75vqcoKfYSmGFPWV0Ya1mwX4isWprUo5Fo8IFEDahQCjW2M
qyVDurWN3sdSjQzwt+ENoFwdMa4VoXxxREiEKz/xp8n2b4BvgxlkwzKxgOecl1XpE5O+JI+wCxbz
H+ofQ4o7VzS1c/s4N4eo9KYt4KvcNJ+NnL3vMYkS+w84vmva7iDmqdTT2bquCQk2pG0oMLJ0vWmO
/GugJtLnjEXoYnS8gHSSSnp/Ehu00K29QLlbk6U16fHRNRDShmKVxHvqkTQw3ActNZjCEspZS09c
ewx6JGSorplG5WFGiRKSjDTqh1NMUm+owwlmVDFMc2qnQAUOrrVXTl+5zGsp9YPrc8m7P/qEdtYI
m+xy4Hkado4ambs+kUxjPLUFUBVcfAy31ArrtiBVkvEUVuHT4exfDIWUj8DCz3+ghwF9eyeeiawq
43oy7QOv9eYC0qwUZe0Yq1QMTXP18P7dUQn6ZDqLq18xQ8qxDqQCJjZtNiU9YQ/J3ONTk28XNZrO
KEf4LFWyd/UuwSm0Otg4VkjNFzF5jdMs5IXb1SKTyoiXXLhpP78a0ATxJVR2yFcfVSMn52Jp1hsP
GeW3LxR/ooazjxTcm6lvIcw4m+8dUMBqj2/53g0azR7N6oFO2oGAQSJ+wWvzb4eZtSAh04rqCYII
GIESeqF9d/Knhs2X+4wMb4emaXjFbCiLPdJXvNPKCYiui77atv5zWIiCziSqr2zjsYOL3bbaMPvi
p2RBvNsdmc+YqOy4OE+K5ya0kFsUSeXB6XT0ad25a5oGVxZ/soSCZ8yxm7XgSyQA69X0w85Z70N2
nJPUOilJ+FGPtBEF+Ib8QiGuRv/8iYbtINW+fAt0M4x1Uy6e1PhFAGRGs/D5gkFkhD6OPaackm15
hKm3PSsIYLLc/vNThsh5wK1ylforKAKgPlHTxtDSO2R2j5f6iGk90T3nQ9dsgUvRf0ksxR5YkHP0
sXv1QZ0VhwHs7rKoyMEIk1iUvCIgUnGvfJpgEG1GWRmTdo6L+X06fSdsp12xKOBOY2ktsOEV4PJ9
cHi2w6xAyJMYbNk+K9UQC2E6E07e92qlGmF71gArW+RJq5zDhwTFt5vwxUhplv9aK9C8To6woksX
BZP+7uKuvkF0MecSx50FamANGE2JFYuGEFTSdHvTrXeEGhczifmeIsnCLqNmbyWfNHU5OLL1gL0A
Iq/NBnOvohMUqJJPsTZubvoMys0V4l5EsXwzmi/QWU9WR/UNes85mx/jTKHD6LZ49ulyGP8IaHd5
pfQ7YyzrU3+fyF+ElW136uvlvqNVEj7tC69nTitgT6L2r3bUuEXecsoc3D1cBOppuSkoYMb+6uyp
xLPqXlAf1HUuoWHmKUxAqFSBzsSwVPD1+Ag5SVkLvJ4YGVoBbOyZiJwZBXn8hsGABi1CAqIC41UY
jQecaosNb7w/+8QthNchVxU3El9WremJIUu0CURE/5oUTjySBHCF28Hxpb+RzvTv2Lpfe7pbd8Pt
3UN2P154aeVZ1i1f7cHsBxd9J001bgiWNCpKh60RZqgRGVuzl1q6fNDG9LEnx3oE8cHKaoHKTJzW
YhIzOjV+RhYLaySSqLr3QnEJzuj1TzN+5cAxG0RiU6xKXe2790B1KjxKHrShtU5d2rk7i1lX+8+a
zWYbNihBFpz95cUICOv61u6lCH8b5XNHqaISe9BV0D7XzNX3RzcuI0FcgLgnIkLdgmS8r20GB4Kn
oIC7eiq3XddjpygNERwTRPaF3vT+6sUwBpSxwomft6EkuZpK0DNqYd2T5BQMybTXoFaralIia9k7
qR4a5fiWIGNUo34XUwFzHCeOwU/hOyIwFpFoR2HMCS7oAK4mujgh8e5tEMRLpCma+iUgTlcmtXW3
CmjwwFZkItkU8cahdDAFwjuUCoJLd2F/jxMoeWqaqNPRdC3+8XZ+6ChEbw33KwBwOFA6ZyzSE28S
JkECAV0vc81WnX87vfWLM2AygJNNKzqh2tTa4x77aDI3VTFZtL495GMK7ycOeBPCCoI288Pso7gM
a3ra+uQyLILa+/W9AlENUGJwFWh3Ha0PVaGzUR2Kkk2QdAEnY1TPjObXg7v2MGNSzP4oE8wLLkhR
+iTksO/uXT5G/d1h3OWUJGBiG7pZUmLGUfeU+FmWteiIsgtjpHoe94Fvw0AdEhD4KzZ5M3uwz8od
O7polcDBlP/vFCF4P7aS1ZcyjtaLj1o164pEhMu3DvWHfIlFCg9t2dvwJDc48TGtJmXKmBY81F3O
PIYuU26amrjN8jWwOmg3rmHNa51hNbSUOfgAsHscR4BfTZ0elri9dl0+aI2c7agUKdOsBFUnspEz
7U5QzR/Ehptk4UfI9LvE5AUYGQlcBorGONaeX3Te6ZBqQPobN2PfVfrmvjZ7wc7glu8u2MLkB6IR
hgXqC5NGlQ9+gLs49JHH5rXeQuFwPDqQYkue2LrsVFY112y2WRmaiIozOidPg3O20kLAzsmxvONe
FSUq7x7OPojuHMIQsUtQCB9StB/qnbS74G1wO0D1ZPowPHtF5Wn+MLKLC87nWlY75YVKe0yFoLyi
qJynf5IZtVaCtcBjfadbr8VHz34Opy6shnhCSfkV3umIMs59JODSuRgI2o1nTcqZKfxznysTbC13
ynwed8nZdM1cFdjJCa5SaJIxGt38hf9/n6ct8Y4VcSpUSRFUuSJzzdNdRO3fNxz+ePQuFkECvHNO
ew+GhzyjL5vVKTlCjvxXtefgNKPv9XdPBEtWufqYEyOktsiG0M/e0VTS28wQ3zSpALLaz3uB4uFl
1Gv3S1veaWCcGSMOdoCV6xFeqM4WiDrIbcbRkOeRnDodYoza/qk6YDI241hBbDbUtQGzDDnNu834
TbQ/UmkLAE8tPGXD9I73WZgTPZTJ3fRHL/67i95YwGkShw1wIs7KuQGGQMFcK9LMRPOHL9/pU0Mc
CII5EU86J5vTnpziiYspLch+0ehpvvGmHqwiKJtrTCCcVjh850K4NGoL7pTF7nqZrz1Vl/rm9S4J
cQQ9HYw7srdIKcg60UZDleqT7VmAOkxjrYwxxQFBJCmZSaoxUs9ISlLj6wSiC9W4eJ8+iZhK0+Rz
jr810ruHhQ46BLM/XP9xvDqxTmb8lpJHDpCropWUwQt6/yFhYGlA8J6DryqGTIFWgRlf3tcntPhA
h/SHACJFkICs8d4wLamhQGY+2ja5rqINOZFWbGGw2Ee5ceHh5388CURBEqxxokfYJc/gIfR35pFy
terdPhRH2XVay7ZkaaQ+U9C2mTeMny6+jNGvOMoJPAJcFqpOpm2pCYtUKCzoxddSsAPG3GbY+3g9
cGCnT5GrmV6q50MPApPij2te6uoShyk0bGVxlSmhnU3SnctfZZUdGcMJL7C/utfao9udSEmmLwc2
vkk+7zjQ0ejQfSErtt6Yp8z2iBsEtlHStW1E9PpLdez9XX/pFcoxhE98Tr4yuNQ9klhGrR89q6Gn
DDIsYtaNjLzCOWqTe/0IEhEMwohJoTkg/IJcBrswR6OtDVHykxgoncnmdjOiPks8ZhE6x3XF54XX
c8lHrvzl6Ola20cq5wFzM/whQQeReauCbSFmKouCxYcIIkhDdGbCQRFwR++0ZOeZKSN+sX53DEBE
q3zH1v68zxB4qpSPycE+0fmkUUZLTHxeeSZYDJBxoOWi2IRF2OFh3e3C2t3MDuZLMiGd0zGb1Jit
UQevKNU4xrqMYukyjM+cdBD3IsniZcEucaXtjwtN8zLeZfAWfzdPaYV02DfGG7pwYLydZdXKiNxe
3hvCO//ZWkSc8YfHyk4iAXcvQwBsSLpSg+HT7Vv7T7heHqOoYszRWW2Gy+Qj9jb7ZxkEu59GaLYk
M1cMkFSBjcoj1zeWurTa0cXlxYnpF+ePKMWJge1eDscUWz1Ahyvd50/O2H4BWVegzBLeUneWsYhT
mfE26Q9uAoTMUGsJ2UUtfdqMWPxuyj0uutv2c7vx1jq4YdFeClxJFH+gns3eri4Rdxh5ueOTrFyz
qlCo0vsNsegVVQa+LqI89dY2RmMGOaetM2KNZuXww2dqx0tUL6sNPVtBWypulH6Lk2T9RweX/ETt
tMdOWQZ/+3468M9wix4ETOhSjNxTYGnEnDigCXRw4Fi7+hjOqgjDAIPisOj/eD1OIMnCF7eBAx2n
mkBmCizEnvmObqSTyGM6WRau/bOxI+FGN8rB9q+gFhb/O6SjWmjR3SjhLo0sVgJ7i9s/OzoKfFkh
4I6/82liXacWERUOaKMplCyzTjAE+/ktYJGBkOIET00bT7VvbfUDVSF3TeXsBfuqwjJld/smxV9f
ab6PAhA06vD8mtWDYAAOm54XhgMM7LgXMI05J0GdZsRkwhrUi33POofQtUtvZMWDAH7h5JeyCOyM
cI+5ghoBBMTVOfVrvCm78jvkwTbD+rXlPFfioqoQOuLIawtd84KknyOxJ+PCq2P52weLI9qZMg2w
qLI1rmDmuhsVkqdOVLRiYcGFUcT9oXDH9tux6zI3vZsBP9ef+X71/yQev9dSp0LqW0hIXQwDy1ts
XWxhp+4M9ErtrPBZ6rd/Z/dr0RZ98ZNe8TAa7YeV6OAg+kWgebQ4G/cwChM42jsPVeN/7CfkGCNr
gP6CDhrdvL1yp9xP+5MPgu/YCA6XdNCTDyGTBCHT2Z5GdgLm9FWHjosF2HH8TWwCiRq873dN+G/t
e9v/156oaw6Gv/E5YCftkSuq8qsn5WRh8kVFbWNDsVVAibZZ45dK/PB76/aGoGgMIP9Uz9X1eKry
T9q6p54+s9aJutx4khyM1GWMUV6RgYf4QDdKCiLJ5dhpalQLBb4AzDkLCUMGWzbE0lBrNG1nviIA
EhvdIRAAjZHU594qdtVZFrqbYupp3vzz6op/0E89VkVBRmBBAre1NJwRceUEiuDGEQd4qbBBtLUD
WvIsRN0ywSguAt0DuQETm3sqg49E7++iFC4pcKIO+FCpyP+XY+SnM0zUQAwLe0XPUVcT/p22iqPu
7b88Xq8cabH+H6uRrjGauxFEEFZhDZP0i2OijTpo6BZstWqGK02xWSK3lKhhLFvQQO+ZF17wri88
AM9qxCogoOhtx+XyTmq61wQyiq3Fkf3j7QGOjGho3ArJHureIYk7coP7krHLHr5kfPngpfqvPupi
XTyX40e40SIVFCuJCacNOQgYSZn7Cs3j2c/Z4roEYH1XuRay4Kr4Lh3XxPXC0HnfzMshDBtx5yKz
zvht/Cp7LHFSkeWmln9OSX3/0yK0zoWw0EKcJZXEySK32FCt/qSeJXDutG8IjqkCyotLZle7O9X2
FidChmNbmDMc8dFtE7sc2OvyMFeT66f90Q+0orEs0S86Wj8WMWOuTydX65W+wC/jrbhtUDPiZC/n
dEZDof1/rXGxfqPtDl+gJPqrqz1sFh5jX5PMJK5W5xH20Ax35zuHMPBOMZSlS/Yy6tknTzdQyCH9
xK+A3KNVJL6ngr5ARA/4Yfe1ia8o7Df+rP9kRDl3FWZWPyIZzQbHBAiNE7tsm2hoYtxvL7jnfC3A
5RXxoPArPqtcf7NOrxA3f6fGZjgMV4CmJiAUeX3fiLu536olGBX2GlxgV37y0dMl32TksfmiGHWZ
UbRb+thz6tvV82dGak9Hxx7HcqY53R4I/gm+Ce1zA5Rr3fF87DIt3nQzNz0sy20kWq79b/GGyTLn
wCYGfjUrppiueVX6+ygpMoi0qSXNvDDeJ2wOripB0OFvIfGhJl+UyUWH9tUJB4yb90yoHNMJpZz9
jSG0YbDN/wFwK297YIMjLEPJCiR8fvAh5JBmxxQukNvys1V4xoLnKfUHnbgd5QTOjAuPWPpErLP6
e0PIkpf4R/3EXLF8Bkr6JvLYOE0sEgI/ajXnV+4zVWrzMMNy1j/v3qC/8b5SZrmHiJ+U5aarLLRo
+7T1tl2Yup+tZqzh6hrayFCG6HiZFw5JZ6HFkPbHxf+31TpkCC7cK5SwaFc5ryIM+EqryM4Bmz8+
AB8o9q2uCZ1/hJ6ud+KIjC6lgjaJUzth3PE5l+1BANLgLNuO/UuMEz/XQucDXE4I1p7B3hmKswIw
DWiofA7WkNRN8/em3nXmjD1Dg8GALcVIgpiKEcPZMk9Vo8wgosCArtRXxEpzRSw+++DLlp5OyXFL
qfqcPBO2WbbJC62n0a0jdLOY2UQjt6m+mknGK5xMG09DoQBBI1Q68Pz4KAmovG/tSTs3QG6Rs3r2
o1uyRd/eK1XjTA1/Qiu5nffcokd0bQEJCZ4V1U8/uvnGbJB6Wn60vSm/kSK97wN5eq+kIB+2i6hm
Sft/3NMBvwfSfr+otaLarNd6qJ61DlmwHC1tBZvCKUpkkEi15cQVfHRD1GgUAyq/wOJYWJvY4/Fx
3IGC1i9CAeZB/5t2mKMOmWOlameQimg9OWMPPl9Gi+ph7dokBH9xmNkGpEXko47AdNWzAy3EzTkc
EMDmZU1/D6MnvS4pILrG6AhYs/CsBu2zOwmSXWyK3WXpv74is7j0wTb39txSdiHyO3OW0GzcQbb2
nrAd6R8s7icz92hDgVg9IeYFvKuAJ3h5e/dGe7zke00QMiUEaI8jSQy/Q2FGbGcI1KTUzUr4yrxz
hCQES6XOOgJL8Gkqo0YQvSzWTSFRN0wkeeKOpRZzvbY+ldTGSso5yHPk4JLuqGR2ItObOhGmHf7f
XYkEsPtI0RhWUIVzxusXQoOb0PRwL//h8/coBYhFIMZR3LcV02uSqO4B8igo7hvtAN0cWrXBnCqs
++j2QGEhIV8ae66rTNzi1C8S3cRE7Eef1/jZyKCIFjsg9OQol87twC3pb2Lp+NfhjDNdzwLtidi9
IrzrKeriJa5ezZ/RguaohaX9ypMtO1s7hzTeWcGXPlXRKxxJtM3tuJkhbfDeNUC6Q5zh128h2x5w
iNa46qWji69bIMq793i+p6NiRnalAUSynf+pV59Mp/AmyuHVb4Vbh8/E3e57SLVQ044bIRhITwnd
4/NR7SvPuyOt6DcWy/xFSJnDW4h1XSwDryG2yCT6HoahhcBgFVcUH6YtNhgoObJM3q8kaNJyKLDa
oAB7SnWGtWyN8+c2XNOxdtZo17JGe4AUC0uQ4JwmjzfjTyn2uNKlQ9fLsg/9JVDYuEvX30+oOLvV
qdEloEo/dCETC16wSD6B4yLstrYMLL1Lv0HWW7EPIHqhOhqZxEqy2FMB4shQwHT7M+BwcLWtpdED
Bzk/koDMbY/FC4dlfim+KBLCtTK5CXja7dG9fZcdsXgE+foRv8EuTpLJ8shoGHkRGwDxBmivoLqo
cyqr2K0I1nRwSsKruXrI6cId9SbWOGLo4mgDMueWbBYXmlx4NYAju8e8vTRgCFZ5IFzWLRNv6K7D
OCCuVzJ0uIVMgCGqcZbQ1mkuDZ8NQZ66/EGyZ8MWalWjx1zPvNn2nILJ7JnrDtyeYzbxTyWI+EDS
EcxcV7ETDaMWLyuIz1Ye5L3GbJ15tDe5Ilm6JJDT+FttRT3DBZZJRP03PT475muC6MdPkRSrEwwB
PFNzSrx4dUk9Kmdlzcj1ENjXuWTbmhwZVbf/+JfgVJ5yUZ4lgk4GL3FFLOZznqR19J7XPp8sYvug
kuuEAQUx3kjyFHZ3huAfB6sNgwxpNWloLlo5lIir4OO05NhybMK9nWqvEl7T9OIGwznC0JWrrDMi
2nTSYCAjyWOtRJXjqpsog826MoeBRpzHpod14XJ0hw9L3hrej1Ka3D8DUjh7Ff/aFt+WkG2znWSC
cnAb49/67/MBgai2PCPkRm4s7JCi67jpXX5CKCAe509hmGG8FbOKXAYXikCwyfscXKBYoN2/B97O
dUJgSSamDuKRJfuBiZq7QDROvilzcqWaKCz1dpT30F3o9m+B1DeHD/oHc8U7//iwPI0qgsdZSu17
QyUvBBiMIJJwd1E+gRc6H2qOl2tReLHywBCLxUNN/MdZRNMvwnloiKkZqGAqjQTUTFw0oNIVcd+T
FsgBod8H96Sg98uvgapqpyA339JT84VETLkWUSozXjexODlTDXyqu11Ep2l5yYhkJIatzTynipyc
gYNix2ulxhjS42I3HK27ItGJNlL68paPgqhDEuIIm+gITkNLO+uUeX4dZTI69pBxalz5iTlpMGqk
LaUheuMMMT9f/r0QJKj2KsesxVE1FhlKkcrXwNZpJvoipSdaz22ejx7ZHRBidv98eM5IVx5yD3XN
WKOU9+cd9flU7VEYivIwumdamebQUgfoNUkcOIfbaIJlhciRykotNar6344vr0xv8Y5VR93e8cz4
uooodXgJ7B1c0JxJtjLhcAxRByex0/nmial2NjJW2MlbOw5ywCE6E2J+0tnvfufScCvnoigY3sTe
tU1X8wxLSDIl4k8OEF6z2mYgmiy5T9nD8MGr6x5Xg3UbU1mq9+1TSqjHGFw7u17RdwhgIB32kiKJ
rEHnzhQO9cbUc6poLDn+/poPBhSlAuSjQC5ub7DqR6GZ6jWkUBev8B/wH0lBNApqRVwe+MgChYCg
nyIITO9TaCBm8FbyxcC3kC4hS6qb2IbPFoL7D0/SO0m/apyZxE1xdPac1qhxZu3GMn1XHCeacQ/c
isABPZo1UYolmaggIxpjOCCXDijT51139fvZ09w6V2tAUWuhiS3Hdsf9VysIGGqIy+zR8DRKX5Hr
xr5t+7fRAFczCAAomGizJH9XNCowXU4+BDUNa+ugLbeeAj28cP3YfNl6BAbAAhueDAvh/4t1mS57
eU6QlKeryPNLCTBpPVboeb0jOf9hqoTws3yn5+3Q/46EydQHiMNjk6wSFwQpYA2KGxq6IQ0jtj+t
5PCMcCyofRkvVyO3fdgSrnWCbk6+Ghz0forRy6tTZql1IXZQnJqc7VHoxGgQ8pfZOZE9nsDqxnNO
vZQktl2NnxsNXnMkS4LjB/yhAYbXkTum9cnEviZMaVENpdXR6vhCN5UGzN3+PFEBUEp7Ak/Bdi/q
prsAUNJLbmp6K7bAtM+i4/Lx4J6x0x9WSYXV3SODUO6jcvqp8xYZpd3kLY9S/OrW+9NhGaEZgH18
IS9QlKkzXymUvwaIgFhqpJrfvUk89YgGW5Pnfg3hQe/WEO1YwiZ8NWZNTBlOWj7lHmwDrOfSpWBi
QEzOBTmXW9swdBGcbeDPe//65dmlcWQsK3ezBAKs9ZI0CsyeNu8WkMkar+JKFKIrnW2a7u2L0MUO
31gz8Oyv3mBV3gtkD+KS+8IHlXJKqJmW9VkwzuRzRNn4Db2tnSz5Gc5PL33CmtIj8tgPinnSPAcg
TBhP6lpK4X5OG/S1f7f3mWhy0PtteBz6Va3QxJvMd1tOFjRyGSj7zfYNRRxrVuMzPMPvN/idhXnb
SibSf7B46Q4G94rVQDZQXdHgeyRGlrqO5NgiX0ZBxSiEW+htHImQH2DdgSdzelJuSUBL8t/S40sS
teEPUGTDxuEvppBX5BW5Pw3tBVYshoGxUs1DXXotUfKmt4sJLVFsLAeJ8ERSAypF0vssehVeuLsR
CDdtYsREzQJEnqGQcDe9BqutO9RNZIveJbephjgobTKWxpC7ovhEYkXn17RPKL2pYXZ4g4hw/Wqs
9uDK9LkobYI5rubVh1mcVpzVpLr6C9HB+UCX8VUgREKFp4XJL5geZk7vLOuDDiaUHNsU5YxIL/t2
sDIkZM2gt7s3OMQ98z1b9wztI++CjRxZFUIIoZHaRYwAzMfUz+q3peCuvNuzJ94Awg5U5p49nop2
bDeqmVdzt17i9Fhrlag1E+gDXnuThWAd1+9g7UTWSMv5nQVtIs/TSAFgEac+N4tNEqsM/vMttqIS
nf61Xxi6kTrgIIGaQPHfMspJZqPxh+fGbmiTGns9YXMBWTRiktlo4V6zp69Owteq5xZBcz1zfPq9
qtSn2reCGmjEiN/92Iyat2ZFh+vC8UeOWOSrLOQt0Nc6CCEy8VplL2gnzQ/5qsw4pXxfWUguBzR3
265NPlXaEQdMI72RgUpsQMv5ogce9muDz0cE2itsJZMFGkXQpP0CCjUga+w9GIjNwGTST6HpWKgn
EWdkkoaYKjHjJzTVXa0NeYk40XwaXzzCOZm1/Zno2z+QnnkGOOGJkGIrfZ0oitdSqmpTVBnIgYzv
pzYbLJrbYfWJUoBXW/ECfdCbT/Lv1kKwvbEXrg/QiFZ+GYjQ41hI/OMt0HTlvVL1GuVW7xG7DFL/
kfNhRpHvKgqsPo965RU8poKEzum0UU54AX8bBr6wBJt0z79pdE9PUiYHKc0zqgQ85ozpvANRfltR
jDH4I4gwQWb4K0N4aS9VwrpJeLc3SFX+RHBqwZ6sr3W+A3x84me8ZN/QlrWLhHFMoUVRu0TYDaJp
YpikqeKjOC1U1uM8MkOF6F0HQqlx9VTqLRFmyrdf0XStAzDH79O2LVX+f9LwKIeEaS7Fc5FTDjTh
PJxJ4ZhMeqDn+8oN16BMosiWDWTSpB9xOIv8wtHRYq0LdRlT9TU2l7MWYmx3ZgE/JtH0RBBgp30B
BZj3+JufNbOrhlaiRt4e+uPfksq5V3spyz2ruGiAPf63fcnRVKQJ5KT3f6D7DprcE6A2q8Y3wCW4
xdBcSgMSJaFJzusq6cQN0VGNSnxJ8Si+YgEqhCYtd5SdNvKkDuMFYNcI6pGAqnVKx+HdF7NigaNs
CjzqS208b3Cha3ON92XwXrZP1V52YzyEdj8wx1TU2BeQa2wOI/TcYe6LexdgHR/knF2Go6h8U4rZ
95fFK7T3W+B1edKrYOnful8Iwg6T/Y75G1reqER5oSVFdwHymb6M1NmrnailBooG+tSqpCodNeyc
VTXv4UQIGPrMYEyYo7n7AmpR/7zTugKk3F3kveCi158iiel6xCoGG68bri8EsuAzRuagmHL/DNP4
ckQwmssXyy1P4I8Dxd/l4vjfuVlNpdDkw32b0Z0d5vY73kSdPDVGMrcWZUrOQAO3ySFskthgX3jV
Fi73zEtqT8yaZxGTxXVile8xGCefPgDc0v0SnCmhk6aHAHESQV7zYIhl8ueke4BbOmd9ZK6d0Kc+
stQyaq7iNdUtBn2GjTq7+Yh5/mQne/laBsgCrGTF2SWHXcAHLjClSI+lntonwDrzNIc8FYOuVpBG
JgsObG2GSYDJxBYXPZe6r1TWdA8LuChclmSDKDddaeklcT9EqeNd31ud+olub9mkghp0tm9ogo78
8a8UupKZC0Va1aAJZzHf8CLPFUscouM1brIoHtmcWyOrWl6gDMYBJ+fWIgGzr/xtm09SCEmIOE0B
FRGSYggngxgc5q2AMQaouJP17EI1+G18us3Lc9jxLdjcbW51M4ImlnSHq/w0OwWiiu71NUGTVEiR
eLghYaDjKWCOlss6pq33vw2Vul3xlqsAgt74cxFgEw9WeTi6qPMG2vjhrrE1QL40N4Lc6ziEUUJg
63FKWeZQ1TAIjf7ArnoZe4UlN3E4NVWdq4pPYbJCl94c8vvoZpM4AKrxXC1mE5lUkUOowwemrcgP
bF5TMhgloN7Ocf/xg91VchEaR3bfr1qwybgT2vthdVvWo6dbtxRc47aieur6uc1BB/n8WmjCKMHH
VBygIlVSZ0I53OiY9zsGF9ejkfSSp5+PRr1Q62y7sgM95MdiVK2289eokCTorbhWZs+Ypy7O4uPR
MiPl02yycpuOQ2I+gqaPPyLv8sM7XjmR6UEjUf3Dzj3zS6sRf+IUDPN8/kUBT4EDP/9Bc9VsCX2F
LFzYuo7tJXC/7Hhm12EtKIzEfu8vC9X4w8hhJiikPrKpMQ4SVhu3BCVIgCfOr/QoKG1Vax+RwHfQ
YvjXm8mpInhAH5of+rvdvO+J7ENsm2VxLZP7bE8IPsNI4cAICMKiVlKd9YEsMojGgzZXBgpI3rSK
XM6B2+2WWkQM1mKT+gzR3lA+wF+Kv+aNwuX+LhHSsBwYBGiUuAbfDWA0vPOJW89I3tAZueEPmZD6
JlklX5rvO5PNbj9PYxfPFaUSAp2UJcFtPxEza6YWSGb4Wv6X+i8RzfmQTI6CYENfMm+gpV54+Mj1
8QuaBroCphg2XtYFF+5TinxriJmVYe8lMJuf+ChR8BxpL6RfdeZgJOqcapDNVC7AuVXs2znGWlvN
ZFW8JxFRAlQIZVKfI5SwO5WKtFEuhO6WHi3eJNmtrT5maelMExjvRWBk0+aOjBhQtS8fgKEfxlXn
ByxYD1LeZZ+2jntXSJxMsu1eNGMNXaE+QtjRfl52D8kvpcgqHKflfeqYr7YL4FlfHLY9JqtUoHFI
bkJTcXYspZQ/9GuGNXQjQGH+il0xxcktuK4iCVMfz9rS7uIbqEItAZPTOh632WjGCcI2xSUvmgWl
TXoHZm5Xaq5jWONGws2qihz56e9H1096YknXcAFV1OFU+mfpVm1uIQoYbqsHwNuw4Pj+TQSex5LG
2cY3tMlTRRwFfrnjzro9uKK36l0o4hrmnirX4kuNVaba5bF9zyw4psw7YQT29/WTx6l2TNT4jqcS
B8qy15cag/1Ap8kmb7kTdPCoYs3kffret9zzIXMTj4x4JZ52tuoGpyWXACepzyoREeZx6EnBJprh
wytQ3CggxRrYEVvHnx623vad72WQAO7MNZTDAu8nub0wm6pUtFDKOqUu+S8BuOFqGGIB/SkuGZIj
i7VOOk0nHtEXw7FyMaM79eRCuX+HaULzXW+5juEVIJ37BQMrNqRIv6112BtgXj/s/KbEjIMYpE8S
S1WimTWtky6QQW16hbW4f1+FU/C0MgV1P4DT6TCPRXMH5EnaNHqQdCZjH99ShGUbbhZhAhiDsN2T
0MAYoFwOcfhJiJTXOJcyFssBXGaXPy6qaG3Vwr3iWP714arAtwb//DrYX+iLwspSM24W5owqLb4E
Rww/7iIEhWuiQ3KzEVZ8ZAHxy79bjKe34cysEdORnARGAHlypz+8ZPUrYim+hDxB3c812vxELq9P
17zR3LKtKtf1xjfLSEFlNacJN6oZC7WeyOaAQdTzvEevPbnW4+CjPIaqyCy1bGDEWVGIwe1S/y+U
XYTquWV/1PvrJanYMLqXujLT2RxvwWSzJjdc9ZyBnBQf6GmLZRKlG9bA4eEkb4H52esRPAYNmOvJ
TgAauW2FJ/peBY7YhNUIaPnL/JuGDp/XzIWZmSKME/cSyAqQK/2NnZemo3msMeN78QUmjVedLxsu
gxlWqta4v4Lg/BVbrjCXhCIsyq0gcgZwwSlSsATjXUFWfXD0lL2gKAfEesn5RIJk33LbA8nJxptn
BAuo9FJKAi76WkmszlPewfYa39gPgGwT/a9Uw7mPgw4QY9bU1v/uZPHKOrBbKeirxOFJ0fN/AaiX
1QyDHeTLrgrUrJHYnzEbmqWffB0FwGuYMe60JYd2TsIIWSt7jiSjCHnpEt7RJAdJ5FO7zX+6Rtl5
DnRQ0Il42A8CJg+732UtOj8HpxFg5VrK5v1KwbMCzT8JzEwOiyZfA/euKoihXHNYrlzS/ELnAmKx
RcNVMmq+UtnIGUo+1PqkTKTrRE3/kgiLA8diFzDith0CS2X3DeYSdT4EEmfxvXmRIXi2KvmObXRD
ZNTcyLCQDtSlZsIz6BS/mhnuNJkWlgEqHZaz+wmbtddQgv1UMf4MHDDZqi3QgJnjxLaUrh7Ni5iM
0PxecqqSojfvYv4jiZuGgRA5jnlkUiKxU3fT9Py6hNyQuwyCRq0PzxF/ssiE5ZAdk9TxyCJ519Y+
oxYrJVS901IG6m9JlJKW41Ff7V0VspEW4sTUkZqEBWJSBCOkPPY4hBulSg34MtzQ4iQgyV6oSGuU
6Lgi7VlJaNNl7P68eMNm4Ott8WDvhbTd6xw1luzSYVOVPwJt60at2BZBX8vZkE8uqi5LSm4eIJGg
bples+uZxuBaej1dSBZXJaBHTHYOLjh/uLB+XS7Wgg6P8dAXOU5nnzazG95LMWOUAMZ4wPTT8SfJ
MHHw8pcyNSvGth8qdV+1zUVgGj09ITK4bISBIbRRTnIL0t76MvQYVpuXPCK3yzEO/If/WtJu9Waq
Wd4S+xgq2LwphyLW5M8C3JWQjcwNiBphaqW9c7jHcF9OWXQKH37E29rsAz8ZBKD6N/IURo1RfZvJ
/0HBf8QxMv2SuH2QhsMPmlC2U+W1bFwJcyMgJtbbtsbcUlxp24j/5zM+xKvFKAmEsSYjqJgweXzs
nkVUsKmHSotB8aqXKNMdMw9JmdX/uXZUg65ieldkCNEjlG4BcsG0Tw2C+3Cm56JWSV25/vW7/RMg
PFeUn7CWQaiK9vRt5U+PhySICozI6PcNJZvygSI4OEtks8m+Cm/0sdXELySOlz/39eS73a0pyz0v
4tlLNTxzEy7oJ2enb7cfSBk8/3+29SxWzYVZC3XY9WEsSOnLhazrbG4vKnMNrgsPb4+8Olna5jsz
uVUQR0P3+nEglhnglAF7kIPvLzsnju2vUZhGe6gzK50o/qEcSrRvGYy5WmemVuy99G550T2ua9ib
2LfuhqvB46qkHEhNn15sjBHYwfcvBfznfc6fq6XV/W/vh4nlRb1CQvwfjFBxta9+B5JjvXdcnCMR
g2C2MvhyyS0emdsWEQ5T2V8uz5rubM6qXF7yvvlLNoQTft8ArINOwkuePlJkv1mxUZ5Ae8zEwr00
EhAvYZltqRdSiSH6XM+QNO2JGcN0TgGH7NanXGpLutvzaWQkYXi6uKg98U3cxMepVKs0IBur8+pA
nC2iGSmI8xQPmfY7LTkYeRJVhBzDWiknjZwho5qd5xGUeGrtPRASUOxxl3RGbffJEC/9r1OGvqxT
itybXgsHFwjlUzDJZJjmvEg/mREYFK7EsPAHrwFtwMeyDbOZAat9U28kyV29gP3myCkJa/Zctj/5
+S/8Ds3rdqcDQC8kx57Q8YZEY6bcf4Qmt+j3Ws4/Ja6mrRZ/2RWfUKFgo6LX3ZhijBZOqklONn4C
ywvJA0mU7/dR5842C4D1Xu69zUHxSUvADqmnPLVQbxgU78uS2SRaH7nK3PeufNQ9YP5UOBNWrQ3t
YiCXM6lShAoFXUuOpx9fii32jqiu+JD8epNErHPKSFGWrQ/bbcY+O0dUy2zBlw8G9E+FdiOZpGMH
fBVd+6PD7l5eVXF4KKop3GAPx9kLcJ2KOh1gi5LW0G3pbmW0iw5Vo1XuWGDkdW9pa+gkPfY0o4m7
JTW2+YLMfQi74vgaM+xUZg16TuVrE2fs/2OSSo6JTQqoFNpMFt4FHweYcoRDxyYUuTHEDS2cviLl
Rwu/bNcw8pKp4Uv0Pzin+zbiXumku564+DX960+ZtLJH4PADhSQptE1DBMieRWx/vUnfZXriwjBH
biKK9EIuFizf/eSUWkil/dz956pTUt5fn1HU/dAqrgYjnlLbfVAc/VG1IjJJTIxuDuljfOwUBVi4
T5z4vbJODQ/KB5Q/SZlKo06m0FZcDbh7jf+M7V+yoccI/vDSaiG1BYQIEk5/dsk17VuKcb+5mOtk
26rTF10oQ9kgUwM3HeWnUjRKMTfUBjQfzouN7bou7dTGE2qHzUKMC7tRTywrXMZejDnDgoZo1xDo
QpQrH4QvkjP1lC5BFDwsGzo4Ho0nh5RAyDrANg+p88tq/SziPxDTprc6Lyoxs+Fih+JrFk8w1hoA
paEf14zO7MBdflKa6/k5NYscduhZJhVRnMUh9+2H8mecZixjC5zUVc4zIRMCVExWaYBSq7ri6uMe
Wtmsq9f4sSOAgqbfmFlvjUZK2QXHMNr7ZAJEDv3vHhD5GF1lNnKnWHlEDdQBsGGSW5iPsuvS6LOm
Ld5YzEjhWoslVekGObJS03Ssr3UdmMl3CuJ8o5BrLTXZ3Seo+R9oi3xQqW45OIeMy81vWmCI98+L
AH/Qh64IHMXvIxPPi99wD+7a7rLwrgu3fwjIhgvI2mgYfAP1dMFj9lWhUoXY+njrADpbvUE1or/w
QoG/7UJg7E4uAXj89qjuQDhgbRGixPttEkxZFMhadSOMNL8KQTUWhVe463r0R1sOljOKYRTcEmI+
jsQc7IuC53hpxZmTHjeS3pAAhkpigkmbzVu0J0f6ZHziYT/emEIqH20GBANMMAR2pZAj5HKxUmeZ
YHZNxCwAHuXHDgDXpicJFNIH6rloV/6R8VVfjiVdsUu0M0F6ANG/vAd8/fTOEsFV2MoiKQqZ/M1a
uluZLHMPSWVNJl3RfKXEKTCnNYiqTP4oi1f9/9lSRhIxwk4AsQl4yeYM/io9LCDDga2tI60lllP1
/oTbxErKM0L6esC5hc1hhFhLimKz7JLOz4AsWlSvuqjtvhvZgdirsjRPY7ZQoQveZPuyQPDr7J99
9vNyGvr5aFheqRjDsdhQBoErUeKrVPVaIgpGJO/gk6LVJAuwOuV7d+ti3FuDAP2AmHY8Z8d3JfGP
8VXvEBgikB49Gi3mfQjSGcScRaTaQ14G5TtSrCHzGC+GsztweUoTyeRitjkrC8E7Z787MhN99Fqa
YWARqmiRtD0+GuTzctgFhxO8MgZfGiG3bFso1SK1lhOrXY0gmTnfb3SSaeGWYas4Bklic4lwP/nU
edbm075pfd1wA+5WVltzGwlGrz1fTED2GakVypmMKlvPiXRCNCqFR6f84KUNy4qezIsa0aOZULcb
uZdIo6hhORra/KrQD2r1I0VafcT9Rmk1pXegFaq4mDqwesfaALlXbC5Q6ZyQed+uCmYfnrJIy5Le
mXrW7lBKmDvDzed2WnsYccRxbx7rRq97Bw8ZOhqYq7NODmYGO8vpi1eXXlrXI2Z0oVANlyA6tVro
/LpDrrg1Auq9HyeRDQp2kvjwPEmp5NwWrn561ljOAZoUMHfoKhu1OxpDqHlQWc8U9iKCrLWlTr0b
TjrAfvu2XitQEUMDL8z+YGD7smpujdbvecrrTpwlY7c2nu+wa/Ax63r2465eBC+DnNAXbQFv5LcF
WR5109r9NpfAvTiIazkFrNvb6J8kgEE8Bq2Sb9qng+sYsFJ4J2dclT5TmIWRG8ukyhPPdKEi8dxq
fYaId48M2yPcOMVuV4FrpUZG/Jckkb+A8byNTQSQOrceWdjuz30c8bpO0WX4CZMmNBYb3FBcvndX
OXyFHh9Zh0vZ5gB/c0znIKzvSIR/b/Xu0Bz5/7osHEnCJrIwjoci3L8woUvucEpgcJFwL7CMHlUe
O4pxK4YKfYLoPFgq9ve0CxvRLMAFk/rshq+k+Lrkt+EKE554YAleyIP6j0NGlwTQOndtXS3yWhW2
YLnAO555VamBUYLrAEzDMVVV9vh96oF25xlrH8EOGCis9au+rop2EdxlVZGjGn1FGEFMZ1xfW2Ka
anImdQngjyees8pB9AaRrA9GaOL3tGPHr2BxQO9iyMsd+oL3On/LFgGc3NA2KcB0a2bOletRSKU0
tzy1qw9cy2pVGgXuclZlnB9yivL4joB6JfMW+nQ0TS4dwQ1Qb5Ndn21iDaxeBIZaiyvP4ghOT7nI
f07svlxVhNlCdQBH+yTnLrQ+O7XXneWSpof/lInFDQVj63F7vp4a5x6ovsH/6KMExg/wr7zuAJD9
NVzmH9MMsv+Pp/ME9DJPLtkbx1uUSo47l/pGWPiNa9Eu0xqvJ6d6DMzBXM9V/e08LQO7Yx/GG/4j
cyOFCpXllLBgTreZrhDcUrvpekCEohupWIznaSXDSIiqQGM4c5yE1qbEcwXV6jh+0yadtlNiRSoH
KpIxH551me8/LJDoatzVY/UWqR87f42ypCnBjRBWe80LCVUbA5sHTaTlRuyCGY4djI4LOjD/7aCE
BK7y1XaExUs6PI8mjnnXCUCT0ft/GntBA/Qc9Yg5K5Nvag4+/8NHvU6wQyQ027JXzeN6245ePLJf
9+BM8oPhgWNpo2o4y3gtZ2gqrETxTYcI1xTYjtT81O6pUlafI5IQeeaa7IW9JuJk7Y8/QzCk9Y2A
k9RXYhoQ9Wrb+KSQtiGiOBoB6MNwgzSeW2GBiFZerIBgz277q3V0x/nXPMOUlEYDkuMPPSXk/f9A
FwOYyo92X2XAOOQywaRtqvzKVqwo8YvcgUuA8rvBSIl5ImNldpDfH4Lfh9xuUYJwrHLEacpK0Udd
SHs34hPnEGnjBliGjKJnPPQ0BkEUnzbVWmECoNggAYgldYw6IUklOfl3xgi6I5n56nW94JIOgg9j
5hc4Q8ktx3hWae8Z64hRdQG6LZztqTXOhCuLu3l6IZ2ACwrNd9xg/1gtyjwlCIqlBN6VKrYsZ4Pn
nTO0oDhKcMnCOBxFdiJDgIJte3LZ7VGECKeVUQcYwVgheAKVQEyRA3r2HhU+q4c8CSGB6n4Hs130
u0EFhQUg2P0lM/KDWUSs8wQ0ozzwNTgq9Pmpm/PaXmPYJL2veITio0FcKi9son+fiIgyGGlgtcdK
Cq9DzJUZV2FtSwyje3x7o0jhZSCea/z97hSqnF/cxNHhYEfydQJLBTmkGR7jQNah46F/5yeum17g
lGuHqd3m1Ah9AwlFaMWMqJrUdmF1v/pl7uu9yfpEqTiR+VicZnYFaVojcNSlYq02+GGHxE2lRGu6
9GGiIpiztJ9RSXwcwOmaj8mmBvn7fXQwoFA3FKkfhNQY6VM3fFmwhUwbvaZl0Oe1teqPMjj8zyyJ
hes9VUuZ+HswQy5Ob1kVVzpRxTY5CNQrLh8z8NCVO+dr+Lv51UoYSPcpoun5O0x9pQh+qgiY8vEA
FmCHrR58aseABttySM2BZh3HSzjsFFPxeKYfNPyMriCdjfuBqjn6boiy+Eiwp34dzLWd0qweMNvO
jOppH+TNee7E3iX/CE4Osfax3BQiVjhA8NZl2xAzIK5y4FW+d2p1/vIklJMooqo1pZeeWYLNaJNn
9MOUCpqQ1Ss/RyBV4SV43qGwlm8yCCbDZspPhjqrXZ6C0kMvgmohiq2CiIZ28MVXC0u1s2M9mVM6
t2cVSitfVDZu2EU5IVr8ykS+K/fHmq1s6pnOat6ZbcDaBANHrqHvpDOikJyn0w1csZUJ6It0H6SS
6LYJvCW8/IjyM41orGXx8qRGzMo4Ksg0XMUaQZVhYJLi9M4+vQkordU95T1n/KGIUuZ7TINvzu1A
moKFF7G5edps950oIBzXJdd8naON/fSBBsf6WJsXVn1kA5A5Qiy0EqMhMxNLYkixMb67CyEK7tk4
GBa0mqdplQPBGG6rzkQEij8wo7M+0cUcCZVJpBsfGDdJiFPJFwPidfF9Fz3FuNngOviwDw9WjPsg
DLu3NE0vV6aoHjYzs2buL7yPwK6Ix7ggjy8zcGwDWBR81TlKWiBqSXcumVjqufxPQ0gsYs681gHA
NExlIULqPDeKxPu1Gno6txkJkppjGG5dUo5ckYlGFHUR0r9UYSi5MA6cKIfyr4bAisGP9J+oDijp
BhdQqZvMLsQ1gpYKWQBe7aWcDghQWN3Q4iyNH2g307nq+okAyFp0jb/ZfhaxF6nLCWclJujEwu0U
sACAezuVzCS+VueOlRORrNByH/h6M5WNAXdV+TwoFPDXW056FdfD9yF0aybXUzXKtG64lRRcIskR
RwXOBbOtc7zlBbphY7yW9CWmbpMPPdd5A75Dr0RPrzN13VuO9gyAa+LRCdBKYTC7g2E1SAUk8Xzg
LmvVX/CXFe0Gd4fa9VB+T7+4KXlWuEXNJgADzAVcey76LqRu4WetJONRXwrnm4T7Vf+iyPEZ1EHp
8sb1xA32gbYFp49N9KCfpOpIZx7hiU3d81auZ/4JjTqCbwQwSNIVOpEFNg2JoliRprNeyzUBqGeA
hhTR3ttq1GZZY2KjAiZ5IswvNys+5rNEiwLvDLgYoPfp5gNxjRvoqF38lEfzAaTwhYe3DoucCV0V
yvVRa7RM98gc5ARae0QLpZ36qgswW9zcpsarjs45BJ5K++VSEE6B7hcETlBKTHvo/zOQ+hH8wvQX
U5BwwT+73qGxQp7C7qkuWQhDFjFWRKYCzK5WH4zETeoPlxtWDtYaN+hnkJWhZpHdT4iqAhS+9iLm
5nvULtpK4LPeu2L0JrYc+a2FujTohYhWmwlN6YrwRal+gPrCwO7FJW/jDzELNoO7KzQDDZ2aMoMa
WGLN3/UOkBMSdOXkV9UPy1zY9cITOQVq2dhmx1TDQX2S2pTINWuP+qijN9lc5NvKTk3pCko8K+tU
SeTSKlbmTqVi0pDKtK02bjF/hMoJLhu0b/fjvXr0g4gqzETAqrNH5WEe/AHOx2gVQzfwDf7sCeT0
mKOd7xfCxkxno5pLE6A+dke2U4vLOrCUtR3t/or7Qkxw1H8CP8XMoYSZoxePKlTnkMaZoGQ/D1Og
uQ8lvk8Wf9pkIUvx118+9ngeZ0GI777/ZNRnF+8BzY3iqiK9ThKSPzZymqo66yevu9sIAYoowPSK
kWCBXO+j4EFMcCcdMLGA1YMULSoViTf+gS6nNreD/RbCVJ/7vEBi7tvDUd3+Fi2CB8DqlNNls6lA
b3pKgngOEuaLsYzCsnr7rva1C7C1chItaCUKZuo4Mh86nW6csea4g66HI/NBgQNMcq8nl3DEt3wm
innNJ/Nl/Z6nAWhHmtF2Qmv5JAdQ4G2zaDOxRfJnLvqiSpRnh95vE6/zos00Lws4bQQ8gHfn9Dae
87Lvadk/JIG4vzSnwe1rgSXYcF1EUNvNQU3VI71CiyFpWjLvbJMmpmZJwVdscBxR+PF9Nr8ELKoC
hHes9amZuep+ZZVYTDsHkvsLgBlxKdk2/U7PeVUvGVNzdIVicVwf7fNzeEmapiU5Ez0TBl7WDa6J
l/FhlfOzFTooR4I8WPI89ukKvbWUlmbWO33B8q/NviI9VhyiDjBz4by0A+FMbrFcuJc1eFsXIaAz
6lXcYTG2IRL8z74+3Hf4A2ykrgvUGZ5pl0C0cYHk9Wd1Ncq13kigzPk9osS6qsNvl3C36orfEyG2
7xmshdEsATtZoOloFOlF3hx8uORZI9t/4P/DUc/bTIvZPZKjPHuyK3U0q0ucU13MNAarSTbBHbig
QELpurYQmTPJ5EJnqeb7ldMQDTilNGGVF6wBcII6cWpfMT4yVXaKOpP2K2bRxbvu8CVcfNMihTeo
xeZFntkcBP5CMOYFRa8ud86W30PeEUwTUql39PKBVNW6g79DuA0q2My9H25KRPg1Zn6B56RFZWhW
E/TqtK2J9WvYLdvZR/iPv52DnuxIAtWoJvIxLlFDnx6TPfP9ytiCYfzKJSPGSfl+hYK18cXkZ9ze
/gnbgcMHOC+k6JOloDnbhV+PAUoMFHmw0RRE+o/w6Q/r2tYkzSE86HBn8qJ/Uw/drKwSrLw2F5aU
ImoKjNrBYdg9SmG8XbEb9OfvV76oczN60EkjG0qy3+rNUVAJ0YcaC5igtkqHoJkNnUgPfjOHTKgE
van30AHfggdlW9aqVbzLZPiLt7Cr6PlILKZt1hLAP4gUE8XpEXzhVB9CnlyibmSPpnZnaKBTDlpD
o74q20AOKIXaZtkoR8qNo7Gt+7Yt0vebWMg5acdYe8xuyR0gdouB0aFdvRd66BJVdXyJ0InZs0Xa
P+b6L9X1ToaEL2Y7pGjp+T2hHBW7Gi40AUihrU5+1PbwG66uc4+RrDLQns5oalFJMgLitHrFpoeG
kqm/NxzM6+hcjK98+qbZfm1rN4lXfOUxEd3mempzgimYKNn8Zzv7C5LIt5+EmiGj3xrqX38tz3j6
45V2P8ftHkOwGUxKDsBuljGycSqpYVjHKs5rga6qXEzqdX9YotXE+sTAPt0F0Gbv8rFl3xjW61gW
lit8hhk7sEVA7W3dXOOacLJrmqSn0XJTvSTOmXk3iPQd546OJXLF0FROrbx6BeSLkeN+z33lfrZ2
Ox25L2FRo6yFLptJi2yHzAAmFgexokvQD+A/GtMpwX7j7D2F5S07svSsW23dLm78xz81o9x87D4p
ViV2pvyrNRT9Ljc07vOdFsDTTV4kqVtHxJGst0xMMwvN3QdNG4qDgoxPCJ7WLzoIosdyUFM9YHU2
G6pAnQWaNlcv1+s4korQv3j0iLfqf0RQrhQUH6WQgs36Y9EAb2e+ITpEBdiilJSpbBB/I0HpBYcT
OedOqRVrTgrlcIF0G6n/ooGo01C6S10guwah207BEFrz45MlquLnEv8mqupRM1YYQSSH4az2Loex
VlXHcfmX21/CBBhAx3bvs5Wh8KRbEmRfmySw6k1lMf/WdhSipa8wiAA9Z3eDJ8WauTaBbstF9WUM
61XG73OWLgNIwWr8tkfrwiu3o5C67qPD+rRlmfSHMWylnuRqbmsTVkMU6KSkxj4TqI99w/QregLq
ObHR8RpOxBa9tqP3WxdHazqGBtkLi59HQXlJZO93GwnkN6OjvqmHb+YiZBM266+1Ei1Xk3KuuvrW
0vhTM89cxXwRrLROW+GV5KsUoFS0l3Y6tU7C+HwGCOZ5mz8JTtFHIicWRYcLf32DlMPlNYvOPzL3
AcDIQ59ZVrHIFSCNNwPo4OrOSzhpql6vv1U0tYfgHDPJxw2s0IlDh6Kdd7UfT+CRTouIVfGRER+W
F2jY53+2HB1QR3jd5BTIhfPtu4HfRuONFRXDQg+zuwnk57B7EGqGeFh/Tq9Tyzt9pOvAGmdQOKyU
JlshzLRLx0Cnob35Vr+orfA7pA05WpJTvCW+/S6PkdZxidYvj4F/fee1t6yZVl2TB1vX6ScWEFnz
RGPQ9RA77rgeKPf/Da4OlbV/Skg8P8JWeU5xiQTH3XKElPTL4mI2586uKpx+Wj9auZxW3bBqjOQ6
ZM1k66scoyTfXwkiTS8onudgUylk37MX5DMNyuyFv90Cl849GCfhpCBfCo6YEzC4dAhUUBUDXX04
+h5JI9sNVyxULZpNmxczm0i5jzNMltR+4zOfZw9L2CwTYPRYTQbbW7SWeSqoqbMX9F3H6vx/O90d
5l4FnxWgt9zzFUQU1b79RIRo85h2EB9MKUJr74e7GTYdA9a0JBjLRVbiaGB+S7LIEdYz9qoZaCsn
GsjL8xDvNfmQXC0hqP+iui0/FjmOEWCdeyuLku6QR3j4wXV+1L4cO6LS9BT36jpEF1BLDcf2uqfy
dnij4CBFUnPNgsstHxbdzPIa48GdZCxamnPNxuJFxDieZFrzC3TkvepPmAfwO3QEm9dC+ItSbpcN
1QNH0a4IxBg9GbTdXZD+3fw7mKzzKM/62mUeTXwqy0PRGBzyPZfgEwTbCtOBXiioLCQ6ueQuFbed
bf/n/yYXhWLZD8mMK8IBODvVcncGra4wImXZvyJp4nO6YOTLCiW0/daHkotzKLtlxaqNoWwXegQv
VPezMpxaqTCHM1kOV3CmWhFjdswICve0//7KKnsFfa6y1T4EQdE9890TTLz5MiaaLRy/9qPf5Yto
wQPmNUFiHjcUlCMRoNDSh2kIY6liujUEokUheKZlfmHD0U0KJgYftfNRdbbNbFLsmX4KoNHvmVm7
gKu4xz22geanqZQ/c9Kxb1lyj/KNhbhwawwGyriPcmU3c+LOG1m3Wqf2ERNEwH6zJf8gTuL1Qec+
gtZznS/h5mUH+JtKVElsIpPe9p7m3MANhL4KcMNzLwTWkHTSWVcbwdPkBB0Z9qIiBSD6bzE/CZY/
tmhWekbv4nhaV/sd4IFqOUNU8avxNdSab+44HCRa+N/3o3Hiz/EGyquh7JqSCXzRK4jST/J29Ory
qTYY16pVB/uLQF9oQTw+BdvfgLrrIqh0Tl2o1x7s0P7W2f4JVXmDwHn+Roujk6uZS/aCoqhqzOdw
QIgqe5CyUkFzvZBcfcYWdicX65YR3om1S5q9C34Gk7yVf6CML85EsTHmJjnnnXykM9vzCVKEcZio
QFcAZfONFg1xdLbn2tkYrZOWJle1T+94cRngDgMSX0LJb2KlyGhIxX+K6xDjyvartK4Ns5ZoOw9N
IPtf6mPXdyEwxdvkfR4eZ0ZDL/psCclXyZyeYjD7m18TOFN6XuMk8k4SP/CFzptonqvKhHcZyi4z
cPTvMQH29YQA3OLmSyi+g+QmYp9k6fT82vwdHOCLSx0VSqqhe2CCPp7p2ggaN3Ddg1bP1b4uB1/N
TR1ubqj20DBZ9dPs5LDokYSD9uDamdil6nAwCN28FtOYgu/muBvjvW6XxUHK+wA6nJASzdWIcqqg
rdurJoiHRLRfv0sFOkDXM13r/Bbn4cWLf+6KOf9bogY/Q3AIOXUtEpflh+tMbs8STkrR3IkPVeqr
swfG7NH+WdlYgIkULrPY6oG+meY3l50v2Vz26Yxdewe5RaqayVuN70zL3CZuk2NvRU4mRtoXdAtY
6wypAV5phuqVHA9woS3iMTmZ3ZtxZw0dpi2x+dATd5XzShJVzTQOvxCX09VkLCx3IgL8lTfmFz2X
PtZkyBsLSRq3eY15+GS8XElqXaLfmTGkhQ9WocpElOZLWKuUb8Pi3anclbJxFJZDqVtpxPQttWfb
UoPtOaYS8Byy91yTPcXQ0yd/v+oPAQfLgsHe7OUjgzB1qXclamcf3Bctw6TS+mWIEy4/26EOOoWn
F2j+ZJFNW+hElHZP+EpuoChXFNa1mxEkvEU8SXgTPnCpuNPDUblL1IKRoxcmBirO7ZOuCTpg9Wco
WNCPchzCQsWVHZQzgl9MQuJi+2eqUpafSKt9gcttbcKQLRIfB2ZOSN/JacluVhq8RXzwBZVcfL05
hBFOx0XxVZS0VDLeEZojTgZvhhYdFPGOHxsOmlIZQZ72x1G5XKh3nWMbOopkBxbg3BvD8Dd+/f+2
OVtFVDezlF7IePWJ11QAkZ3Fm/Y/9SiVRIwFlL7CggiZOZKQ1p81slejfbR/fzsDUc3NpsAQNS0K
V5ls/DQ+SzoMygmOHz30e43kJPScIHJkMWsQrNYt5KzO6e5cu5T/nOHWvzdBhjFHXAz8icK5iyM5
lrlM3XS+riT4gqfsYWrp7JMJryoYlQeZnCEBc6djUraDBbnq3Xk/+hkwWhU93qGhe27zEx7rw3V+
+Wj5D7r5GItGd1sSAlcUonvImXZ95KPXw/vkgq6g5I4QSmpRRIH0dHsBd5ZpaNLj4vrLzQ/ggLVC
5T8j+6BDIYVMFmX0HkRQHgHHzKDzvQhMQxiKv0PrVm8xja27nnfm/1cQ3UVHRsaEeUzpHlaqDwqO
RuHZmxBTG1GEboh4+Qaq/KHpydSMrvhYVH9Of+4MXPy7sMDXEIBRFWSMeEYKLM8Aia+Ep5iHxSng
M5x/ZKEV/MkRf7orc1j8bpGyJz9R0CrJpa7+oVKhYcwcdMjShmuKy4bCjGlPfCHNe7u/QQ+e3mjq
0L+7xlM//Qhanm8LIxUWKQxQtMlIDlajTZm8pSWqNIxnhiWce9hVgbDj4CbCRaC84kR+rsf2DCLU
FgrvCCD0GkIwWpqXoklOuUx80c3mNejpU5qx+y6GTnjz+VycY/E8FTqz4O3pSbKXcodeG4/Dea/a
3ld4DtCaPRMbwdH7ny114ZB4LFWxmVpyStMP6nnlyWL8BMCfqxbrn0aZkcocBXwx/iEhXlExSD9O
DfJ3B4sIrhpPmED9ZhQRv4McMrpURMRHMNa1TAjvetDZEnBmm5DqH6KdfMwdYJkJMrw1DJNBlykQ
8FBizri3gcc+EsVTu1GhHcLiC+pDCF4E0z4Rp1p/aI5uFIuggkEUXG5Fs0Wl7Ew6NAjtTktOvCJR
W1zAGGV36wsHjGF/jP/0UgwZocB0XLb4ML1Xd5OXPVVBU52CJSl9sOqfvfGfVBxbarhgD55yb3DA
FX98cLibyO+KlZFqMIgn8AtK9MVcJVaElFWSoyjBL8+9mgTto6AcJv7uukw/xKUohtsobyHrWwcW
Oyj3czfEnvO4++pQNnvwAKuHn7WAuD3MfSCaaefhhRem5MlHzBNq/54fszyyh0wY5uigW/zSMTNK
k7hq+nbLIHFmX5CRPuWhnslPzI6fwUXnCpRuOkKZlZgwqiy+YlKOL3IzDZvIBHlLyHCYOZnL0biI
r1W+eYtn01hRoe8smFV6yhpGyrMTCf2nrxEHQx8LCcBIt2PM2ME8PvqNe3BE0ap70Rb0yP04afMx
QBKyw1ZPc7xENOYa98LKpN+fVZcASDpdRNIcKP+tr1hVVYTDjZELtKxBTRD3Bv6Uj/PzJ0xFgikY
+sJ0dWzELYFypkuyrWP3x7AqeA1+9MFi4bl7cqAXf+2VZ88tL9G9NnUlfqrGcAh5UNfaR1lXvwCD
Lz5yQua2ZKQ25G0zPw09l8rsShhWTAYeG83+IXq8HjlIgIv6IqRGhYlV5Gm0bbMxJSLHnOzo0a3L
0yyfRwnAd8Tbu57PiGxhmKKJaopn7ryIlwSs0XjHUbx40VnzPQ3UEuSjFl01CZVKHebY86Xl3w/1
2lfCCrRa+0YHnCWoYb7yQU4FEyU0T/0icqe+VLVqYBWmeZdq7e7EY4oGUS8aLF36tcGQcyxAQF9g
tvR493L3nL2X7D+N2aU4f0b5IJMTPFbUoTfWVo4iGEuiljWv6OJAtxF11NKhs6gJfWAjUqrTAKhE
zUmyrYwfLVSNp8yyXmO6Om+JVjUzTqstRvYFrcxrtzLELurMvlaK7fBxUyvCRko10Tr9gBy3hRcm
d0cEqJxld662YsE81Ue6kEalZnlj+vjY//gp7JVlrKaFHP5pLqEA4sgnduizG8jJg2413aQdRDvO
p5ZIOQD+HbeXQmF87VLuNnXZjU0d5GhnFvK8nbUdxuoier9FxMZXvw2O9gWtT5KDoOy+jXovTI/E
mnlecSfL+/xClKtG3cHC4w0/RI7cmNDMYuKAnouchhXO8J4DYMuBdHTpTNhtaJp5S0o6KMq/uofL
P6CCjbqJl/Uq/R2iOm0cBSMrIt94Sv3nzNQyeDu07h7S+0ISSDC1nefJj414bxfpfJd3Sksm5SSO
GO9LGHidXPus4O9Jcv7lZPhH1sJyuErHgr9BdAUkDPwuCgQ237/KYrLrcJCJggIPUGst9+/o1Pdb
9p7piND66fZnVZ0Ls9dRicjMVmejOwO1YdDXxluLfw27wCVjcQcEoixZCy4F81bUysnNwEvpNCfM
aZ/lbptNRDtV8WcMpRg1XClYOmtHpqpPOOyhv/4mWgL5Jl8if5wX6xzZfosULbcv+4fapL+7V/+c
jNTJCE/694l/AdSJ5ESF9mVsY8AWC09+wra+eEvSWF3v7rlWkmHkV2EK617WMk1MsLnKfK+W7cVt
QYIQFQeuLCsGpb6V5jMHHP87Tw6JKzqRKwB0ebh5IFG4JRJFJt3tlBmzGZPD6UVfuir0EGkBvyYd
VWCkVyi9qh/RYXbtjVV00oEZZiTvfmyP8Mi0lkFRxZZC+FPNtjmh3TryqQa4Wino7M4Wqu1kt5G/
57Ysogf48x4YBkrnAM8gyEC0U/JAd6FtbZow07c29SncX80/tUekR9UGTCanLCNY8R0+OjK7krfj
jLjhB979RP4tWeR9GJvlqn9D/x/9R20qKr5f/uN7Zt5ITz/0a/WLJ7zqIgX9+yKcmUk8piy8Q8po
IT3AIYWbIvlUaL4jp/HFQ7iRySkZGkzXDXZZ263FcfoKGQjj0DE/Z0ZbTCjJq7uPXSVkVP5FyDVc
dhWYROdMfPz6i2O/2po2RGnisOiHNkeMfhwJfIqLTamqT1Wu7v1PIGF5mAZ+/Qph3JoEJBp1+347
/Xo6cODWFFjThY8ihpO83/6hGotoXWc7Y5Hn/GF2ZfSdcFciWJhFnGeFill53v7EUqZyAZ8SD/II
eCqig7mmgKLBSON7B1hjiC+SFZozmqNNdeIs9bEfjEU8OxWBBGCa4umoHkJnixzRRPWsTt3k83LQ
9PQ7XQGYmLyfV47gUBhTntiv9ieB3lW9Tpz/65+NbNeobfxTaKy3zmYCsQaBeyGrJ07hmR6esZmQ
3KbJu16AxiLEnOhgSnmQ9+wC7JY3G2p7blkc9XIMWTU1QwtPTNd7qSXY6Btt1IrNMf5dLsObRcvb
K/OEgu/WnicGssGVOuCJytZ8MytJ637mCbk78KoDTHnOeHkOiVKqravLAgteSLHP5vhHaEvseacW
z5LJ1UQ8Zlojl7tNauy+dTp7/g3oWoW5ZztU4txlqyRNhyPOzNHYYV7vk8v8r6WcsI4RlFusgf5E
pK1b4GUfFNRzhG1BtFlny9Eqb/U0FDAbxFHKvAVRmxb7/u24toKUbaXh30Ll1k9Jwd7kT+vJoyaJ
goHgoL11NQTSlOyT7rcKRuyXMh9oS8fDiatf+s+ShjSJl5W09mEPgU24J0E7vKn7mshAXEaScM7B
pSrgORA7E6GakHg5kW9fABgekGvT9xHX5YsAa7ryc25ZdfgKi7f3YT5PBYokCj279vVdChiQRVVe
LTnRTgzneF1OU0pfgXhBg+Er6mrvEibJIQXa562GIc31OcikDOpY5nNbbs7uHstu3gCFJsdgqEmr
wyApV6lGifSYCfNUDzp4ocom8xynKw7+IX0h4OqhrtXSQgonZK/K8huWQf5tbQQ9inp04BAdJ+9I
WWlyrtG9LSsdXUiypnCCU44LQ9OGwXav4vi64aOZYOzV3UDewetY4LXiWqE4kaa3woebNSNtYeQv
JKCf2KvYtkcD/xQVVz+YHBHrnQ3PIhtr39K6eLNiOcqULiOtjWBc1Hjql9gbY79whPGFPs+VAj1S
3ZSUy0JMJBaIHyvwBGV/aw4CIKuRSb5VOdDeQsCZ9ujz8EioceRh1+VWbKRHH0LewOaGAbnLV4/f
4R+jLngrcoyPeAk15/pu6d+xqg7V0XRAFCKCVlTzCYPHh9fhjFayItqFAwYS45B54NArSiYDLR4R
ZJWLaj+TT75vhcnNfZHRawZExjLQbe6ChKSx+bXbR8NHViE94cO8phXIcEeQ8m+7+hGOhGIcT5c9
m1CGlz5VvpFdP+8Kc2wNddsvCRmm4CD6Jr/NSpRPPPPoqBXCbSDyzH0FOPe+YnqnTUUuZOXBAMi7
GVmpWekHdL5a6yAeGi7kN45xy7lD+TYfjL3zFUNGeVT61H1CmraQWFv9e2zC3i7hyY/C0GBP1pdW
r/9Ir+hqUEKH6BcvAX87CcDQVYV2ylD0c167fWq7ACBZXZyAxD+b7lvyMF3RjpNbFv0kHTAtAoCk
weYKjsXyOU117RA0UpvUiqUBWxHYiqXrxD5qNrydOvU2v7ydr7LVuQuzGSy2UPhUX8P0Upgw8ncN
Ki7Cxe0NQUNb+Bf1AiZaP6D+B1/WCxJtWiQ3FcxmefxeE4rvuBBYzMW/8SnBuhURL+K10LbDaIHV
ApJIHPYg6Oe9CNCBJGTuyQIrc2w5McHMa/HNtzoKFJNkVQYsIgJP2+ahUCfEBR2iESzFAmoeypKr
xoQzYf74c2pPcj85kZCdGqrEmEnLo5ai0gaR6VDbU1XObEjmsA1O0PYvgvJu8oMtDF4BCD+KT9cK
AWSCuOfwBbO+vUMWZ7bJ4cLdG1shCaCRm1Td0+S0tQ7/mc8R7/R2J7sT7uJzc+TZQF03+B0WCSMt
xv7/W3Tj0ipEWqrJeheDyB5DDLlwi/4XQzqEAKMz4yBQKijtRw7IDnbTXLsCaAfnp45n96dEHBQP
1tbAWptE69su/944Tx1w3IniHh2KMp9zS7OeijIcCqNsRAUrwrQquEaYQAx6SWUM8x5D4bdrVGwG
/hGhefEwh2l1xmhmUeDwjEWqoiDQLZjQt7f/tfKnPUxa0DNDLQTyFhdZ4bZz2H/cnEPB+JGFV3l0
ayDe9vkHkS6ttEwjp7J0kzZkmGa3eFaiJK/LN/swTSGH1TzIw/NpTI1IS3hIxx/m69ovZjja0s8+
A50pGQEwm/TbTjSVbEbIqYn1g1E6uimLJ0z44chby7D9NHdfCCZLUAoEax4XPMUdxOMk3nqdPz+4
6mR2GmHeRkGSYpbPXYJ2S3vTXqP2b5ChbH5lbGBb7VSpH5EZKI4kR9vJwumvPCrrBlkoGNuAmxSt
EmJG3scyTk5DTh99WW3LYguDBRHQzHc90LQxoreNllt71d/zEfatO6+sTLubiDisqGlIvQvqakv9
uCoy9tC5p8DYi3Iqk+YNFqrpkdODgpuJfArLA+P4R0WFntzL3DwIVOpoiu22JudyE8RWLsYbHg6/
MDgWgY0vSiMUi6U8v27zDD6HIHxO8Djf41oak4yY5mmZwkGsu885+iWSfLKZlKFKzLvDIjavA4sy
VB/NufMSqQfgkfWu0SZ/5sZJc/FCHiUmkBaKcb34CMj+qgj/gAJq5kF8bRpvUa/Jv4iLA1yfS5Iw
zp+Sp24zK0V3YAtLpZncOiY4aHRKSw0q8nZC+qyyYgW41HE7eB8xdQDr24KiHcl3ITFAk0hw9cjL
bXTnMvBA/qSsvGF/3b/Y6lkbykSytunl+uLqxY5PHrosVYBgZ05UnPdGBH2ndN7ofSFDS9Z5e+me
VKKL/6pdOcsBuQYjNbsRjnocEHYWeznAxKLF6g9Z8UnFzX5wNZxcpIFRIcA/TrfjDXtZgvXYaUpc
VHNmGlZW8ANv6bLFzUi74QddUw9Kox4Ko4URSs4BNfip4o5JyChtcQ44d1WekPfTnVMXFmVjqaAC
YgTYgSgB7cO3E6qcSTS9sUXh0QY5VP7MNWMfADKGkiV2Vw2tBi5C0/c1hfEgPWtFk3NEHIvgde5/
ZnBAEg2/wg8cvbvYJcsyME0LVDR/A4WTu18Vow3GpeosebjzJpdNRJGEgRcmZxghk08+RarpfzBS
LKaQsofSrrhPWzgEF9UATLGpWDNHSj0PpoK99qStfGCuZML3CtLvW1TBdVLThNrvxdK2Juc9ebif
Jd7zNIip9rrz5HMWMnkXUGTsAASSfSXqLpXl8R/vAcjaSzYfhSZqYGhz0yX4MQBqRqMWv0cYHVdN
u9p+4Rg+//FATe316lIfOtJNzp+mNBf4VMvdsN9Kvd/xaYVVEtFviBTQZ1VU11KXyfrzCzjKZJTd
djNLbeMOw0HAN+isUGrd/WbdoNJvrrz7Q5Ec6mxkeosI46M5aotbY3dH2IFpsM4EhBdzbG+uCExS
jErzFpQI9l70P+TU8C8kylybZn+JZPeZRoQyp50ERjiCOCYkoBlvIusUFkoetR3eU+xhA7D29WxL
jjRUwV5YiJLzlaTm8mpzO5pFSlhdqiBRWqxwWLJ87ct7+T8EkT0lmJZdUltW62OOz3SZMzaEm0BP
eOVtz61w//yUOYg+Af0V/gug1jhMLEevAedik1v45KweTBvlpByD2HKLJqQLvp5cbyfE1LBUvU82
58DO0XQ6EZeg7Vt2vI+c3kHAdJZ5nKMtGK7KPtR2nKuqmPPCW8TbktAbCtA08qHuycEhTIE+ZSq7
zteamCZv1mcqh7j1r/Hp8HvgoZQT1HDeJ+y8Oy4Z7/YMpUtcNt9vR+eCleCKOKl/VxNd+Lvy+oQR
9ugNo+sDZtsWjzf9QZjl5yroESvhuy8+oYYL7aC/KVmYh34ofd+gPtFB7gROStAAzJUb7X5dn+eT
glmnP3zWSqhJau7fjfNKFGCNOj3P+GEW+vn99levYhLxnHolGypRomBRxdTJitoqBIYnfoafWq+4
PGDpPEgxquGuRCSQ7Uji32zyjK4GdfCUXkEJK33e7LcjIZqwKwU0BSlj2YO4uCVBma7wwMa6i8NR
ozHxediLOtaBNwflI7n0tuxX/UcYTdU/XaL6ERf5CJGOcctVvlWpPQP55iURmT1XYyaNbLfJohl/
Q+No3KVa0KUF9vLsKKnq3D3rtF0ssjxryppWnlQLpcYJRU0ApPqhifi9+5hcIfoqF35gLridmdZV
EqB3NGVUg0M8EOFQfYSquzYV3Mq4fA36UiH+c5dlmbg/o08P+0pqzFlz0NO4FMNkMKUeHq8U7srK
QwO+V4Fsymnah0INsOHeULs/pYo7woViE+0XYKVwAti7glX8Plr5izqx3WNfl6Ts112vF8iTqEkH
UU7W5yYovWHTtkslK3v8Wy52KI7+g2DN2KqUD1YJ2qes2lluX8HqAj9Hn7IaBh4WdVU2KlLfd/R5
FQo2+iQMKQqvfkIYfGOMjixTB4ObW+IoStKHxuxdKgOozBU8xZzy6cQJ3I5h8wiwLoa8HOBJrSZW
3JCGIA/Ndk1nNN4gGpNBfJEGyduZebbrxIHjtMOUVOBJcKJz9C1RfpRgHj4ojOU+dl2l7uB9mSB5
a7V6ZGTtupYDZLbk8dO9xEcurMzJM4Dd6UjmiZ9WvbqSs0eDys4mnINFQPgzPVf8tEWfL+EjGgNy
ubsksCZdFJbzKsdIwEhso42U1N65Wh9XvP7nZ1aam9PXVxejY7WrGzDD8MFMZAYPEqryIZEN50Mp
WoDvUec3bWfxZscernLDkaW81CciSnILdGYfvB+6qWFIRy6vEm30Enn+RPh068yFZqcyOv9H3CSg
XgfJ5JtdtpQD6UN+/FAGtF6Ac7JyxKEQjHv3nudm0mMNcUcw8vbltBOQ4DA/ItxSCtGact3ltr0r
Vk3Ow+qvUFizRcv5yAuA2/ty0m+kgvToy9P7GKlCpDHV8/dlQ08vvRAaV69r07BVCJlQEWJ7ZB6c
0mNXivRQnN12D0s004CX4n+UAg56IzChL0leV5Z9TGFAYtsGCIy8oDQvFH8hfiv5b8L+ixANIkYk
z3sDrOU7zTtza0sq8gr+gh160vWPSrk2LrU16O1jd134Nzohonj4E7Tsy3aVsBJ+1OVBdq59PKWy
LVkaRQIfjajd/lpXl0r8zBz+7tYildNIsly6wSeu+mcbeg0IprMxqBga4EM3o0xb4zALlVzqtpDW
rYEWiL23rmehqRHtvh3K5x0CwVz3wnghIXYgtNxgAxIenHEiDTwrtQf8b43sUABNgFi0TtY8OYxc
wtwqcnYG95pwpNQ4gBgvV//gvN18zsL01x9JFGwtbVJY2bEV8+LnqdhIKqpigsaYajAK2o4HBnK4
56ur1sN41uYKL4VBxp3Aenk6YqcsF3QDMuLxgMIykgL67OdOtUWFlrZRlLayYdTmRWryn2y6ojKH
SnidAEZ2XqRnS+hNaKCfEmM1a4vDT+AASLfCIsRD4A58xIlUcBSNTYcwC4bwcmdJZXf+4fcSGfsh
sdHnD+eOek/5ebu9JKdRj52bQw+RxlBhLGfQ4wRqZkMaeVjJcv9Czhmlgc06Zh8Hc2ibetxTHy5S
S5uc8T/faLc3jPSID/3QBX6MNsjnseDsntf8++rvBHrutPL4khVEsRIDhtXiaV7vBc3v4kIthYTA
WPYv6HUeMFFHb8ML7GRY5Hzr0gNOFRh+DekXTuJerCL4s+d4/a1WSP7GyBnKvUr7aqh+kQlVgkbp
PNJ/ebcWplbf2xhOp+Bqzw7YAdqjQpdtDV9YiqG2Tk9nqQqugi7aIPEF/sOAzfCBCfiNaqVV8y8R
q9/woahDT9aZyY7XRk0s/Os7ch9Q9ZZSDoZ9qOGUyy9BcdVsuXTQ8hjnGyOieSXo+Dqpl66u1xzf
WXNlHio2ODpQ/Pi43U8jRrh0yB74508gUPeUU5Dejq65xtC+trH1MeGx8oLcZ7/IFYboceWug0RR
nA59MRfGydKB+DS6vbCzCzZCCgE2qale+kPrAkE+nud6mr6vlo3IISJ7Ba1PR3zxGW69cjkRGsYi
ZHkl794l3m0JE/J8J3ohyD+qvSRKIf0fwBf1vK/I5jMWYIrDOGZAjqhiBkzBDvZyXQwPl8VkzM4Q
M+tm3o6fymJuRj8TO/JK0y8mnq0eSO7aKTOxmofpXm5RIwM7QvLTk/FG1St8TyXuOHniMVQwLlql
SqHvd1ajgGgMtm3abihweCnHs3oBy5Pkqf/J3AWfMA+pMWn7xC5c/dK//fvvGDJEmzDsStCjQclb
h9kgGEBTGkwVVHVO64cqgubvJ8a1WdUoyTivqZHgpLPL/9S/vgz3rdX0O/lt96Rf7EyuJDASvEHm
F5REg1kPTmdFkeMWujfh6vPFrQ3UVV6zsNFQTmjBqSMl7t5x/MW78QJzLCpgniSZki4aFyBvgHWr
hTIzLJaqFD2De4KjUq1mh/zS34goe99TQu7kHRbKTHZtbmzc/NnInVqkqxFbiTXxfgS3eyitCipF
y2Tzxr4vrX0CpCqb7k8u728g5Bttsv8fYOgiqqi27dbtlRQYLdzSqOeNJknZK2nyLkIb//pUYepw
0D9YS2++nppOAO9InOdY1pUH0jLXLzTUhuesZWkqlwiVSMmyhxU5NYTad/0aikcnQzEmhkCzYOkx
w50Ne2rdDekkHUyoxgz26a5E8iAB5e0PQjsF91ELVU9LULVyEMBxJzckfxyQolwmnHtH3cXbKDHo
NkVRb+bXCLzlX8NVQFSq68xh/x7anrmUbtXU6oF0mSjk3+LLP1EsUEpyLo//uAp0M0boX33q1XAW
wr5vtEegds/5EHixEjHcAMVsvU8N1b7zp/Aik+URN2+lSfF0Wp/gYzRgu3O0iuDusi/QgPtnaB8R
rAnxcZqYT+vms8a5WkUty9qBoYxAPAL6V1JePl0k5DkU6Rn2eKevyUx/cdg/kmb4uo5WsbGBT1hu
n46/Y5b8jbNcTiMKFC/eH3bMZX7Ezf4b1cTqyqPiv73X5pp+ec1ZC1dtKs0Wgoq4fSKamaVOXuuI
WEk3kC1/BEgY8BLYDADgpJge+uQQxYa7hZ2LV5kEP9S3wlIsUPth2Bcrs/eclk4pqY9S5kX+xMpi
9DIXylGLJ7enspkpipZctrFENV5C5cRp8tpyo3N47QBv5ZGKzmPxbtUpnxlrctcdvv+W5B/w3n7T
xcswIMPM6EwgKzEngyEErKBH4U6LWC2I4HLTyE8NNsgK1qVAOQadF/IL4kpqP2sC0gnurquIHyXf
mIqctSp5AUNxPEjgo1Zbn5RP144tjjhVjQ3sA4lyJUc4+2dB8SJqWUSSqZPy5auqiCGIo8ANlGGO
sW73yYEPOD5ygp/KLgKmhvC+RKIUSO9bVNowgR1S63KoEYc6JXXOJqciHmkHhf67mY927OFoLFkZ
4/sfyiloE8O99pIWphcvl7GWxpncQejTcQDM942Ke9wtIjrX3aYcC0wg2RqlpcAEOYSPV2SAhM+p
miqGfUvTJQZw1s/kxTvByv5vgbBW5tchH5ZMH+YXDreNtVFqcr51CiKSmYzLfl+3jXUxS/SrQ7w0
oqSUofWvgq01HH4IURNOtU+e0cfranmdm5n8Yu3h2TUYRHCtaj4zz/5p5l3dDBgVY56TWOMpKnF9
IOK/MpCfhDIQWtHyxibQW8XQ1NGkmcLpt6HNp7YTEjdhHpiFmF/r1X4eUd3EjJ922G3+LAxtvTKI
wvkuSd5yCgBkZ45++pLWG8eqtsAPo5RnBE4tBy50a/VTVrsgD76aIs41ksCVD7APYuEY/dsD0b+F
FBt4YaT6ZJ2wc1v/XkqodHYQUgL35XJxNZ1ExZ1VLJ07y3hEcP+fcpsMpN44bXMryme53qtDK5zS
Da8pzz3yxLPvLFRVKjSOoxFIQxfe5JMUQwrfkusK67rCpZ++9r99T/BnE9p9TDFJj1q557pRPw4m
fizW5PZ+TwyibIECtji9Q/sKrBZRnfef2TxB2sxryfUNnR6DWK8+y0b8Rc70WctkeWNSDXse9LXx
X34kVqdvoS0/VhAFJDBCfI8vS5fka7ovoUyd4xRfJeIFiikq+ssX7zJGy2ulKQvVkkYcVTUZQXMf
UbQ7gFaU99DMIPm8Aje11BuEtdDSB8J+xCtJKyHFzq/b//3PaW8UiJVe2+yBfh7X7gaM68lSkjCW
ZSPLQKX/ePGFr/xM38C/KTR/UAFgGtOkRz4PJYEtnMpkYCPn5YzdGHKKutW6/32FXQkefhRdHvml
ygfuRr4IDiFEe5Hyz2toF4LbZDDjRdRY/mG3gpJ2QptQ0glu8D5GVrzqaVm0Qf1WNDFNnXmmyVwM
CLEjiiwP1lwY6ujcQWrjhMpo3OCMcbAGWTJGHolixpoSX+6bZ+lpSFIRO6H8X/2uYw/fN0+etH14
qJV6TYC4ueFeBRAviuzYIlqnrS/GGJ7s0jImgNHjI3FxBbwU9CMeDwIH8BQ38ZPFMPE9EuWK1jhm
IbUh6icG9dDyXPnxEvJCaS3HnSrdYCFrigCVX373IMbVeWuZYcv6RyrratsPV7YMvmOmnlAO0FhL
D3qfTyACY2QXtk03D6KzDMqgV3BBQXTHEyGuv0E/TTuxpsI9+5F8+zuJl0VbeiGk8ohE2zh14XUl
h2xTnhOw/bfstIw/pXye8gldxlHtI4SmILl7yObQxr5XH/LJr9zhTy3BrhKSAhn///vUHJ8krmAo
1Y7WyuXKPiv4afqXUo5Cn9JXSkgFWiuRGXhNWW3sGGt4qoXG2nd9pUPjnbu/DVPIwIqmeE/epAdJ
njyanEiyeM9G3DhUz2zbM9ovfz4Jb1NkGq97TGlo+JjGsm0jcQ/2bGKDpZfUd7lVa8otya4bZb6+
LiL3V7BjzeGb5pSakhVtKhNsIVMpvM/uO/NdouDt1uEMG396nmjVVJA5CWudeLdDoP2Jzmuu8zwC
hoa5SEkOUmhx0ZA1KPwP7rYbW0csft9dYPTKx96zQ1uua3MGYsiOLhZWAF7em1iVcHQlBGtEzc94
eYMIF68wVBiB55r3xribV+zimhwyPIkIXNZpNV8xr0FEabIwNf33vp2q0ra0tMThBbRN9Em+pzL6
aGHM8tdIL7Nm9NqF4gJriYZPfg215jdK4arDVDrAnqOnOByoD+npj7RaWsIGLUa7sjUotSKjWmvf
fg8QwsCqhVswOaMNxat4SMXH+sP34Sseo0e4iM1LBO/xA7YncVdv+JB9OumCp1xLSadppQLszrah
9BH4Lx+/s0/hoLPicroI6PJ6UwSeROVHWdUUBaLH5ZEJ1gjeG9a9+HZ13diQtx4vLJfBwKQ+ATUM
7JJ15TTRK5fYpjq4n3qqRXalNg3xPHoqJ52O37H3TIISCwM9K/xLFw6txaaqx9+yPWJ4/cJCWM60
9x/c7quePMr7rbfO5ap8GxZQ0skiedQiQvFVk3AgVAzQZMS5KbpFjaX7p4FAZMg+R9ZLFtY21qQN
p2Ul4QdU0o4H5jITPa5DbXRrD4kWKgST3xrzCrHYNONFbeOojSDAqq7TkxyeMeVDnwEXAS1UrJ9q
N6RCnIDcaSAvj3PsGNy2ucHae8MqTNwh2r8R8+e5HsjQlQMPftpO2uN7F+nLBxWYUcLDKMPRZZIv
hlWgSimXNgeibu3kKWVjHNTMaD+vw6/o0EVZ2hRJdBBq5sZhRRyYpOQXJwO75xxJnl1eNuo0/t67
zTwObuDJUUku0KwBypZLmQfql0jvjfZLdnGdXcbBapBkmNcPXhCwhMbxLwXzmoDYbtKWbgS3QJgg
KJZ9qmLPdj/Rxam/xFUo6S25Kcf7FWmSUFT26NjkrABlYzwpkNRnglXSfZB1XsSTu2ndoBmFfqhL
AuZVC2uTdYG9Mf0bPrCYYwxvijoQEetdGu9JhxmKBophHtivomWaXvAQls0n9vffJ+iBkwuS6TX5
tqMp+D1LGI7i8EOsX3TlxDr5KhiBVeDmvnz4PhgNO/8X5GhcFI+Qs+FyTQdiUOEOKWohaOYF2qP7
3cGDEqrAamo1WrGPGcsokeE1NZaeJjkZsX9aPVYH/enO6UhQrS8dMtjVXIjDjUD0UeNjs2mf2Ewx
nBj8qh8luIfUOXkCZj+PcxC2pXDA0/IZ/QF1rmubNoobWXvbLAXiUwWG+LWovSdqCH7MnxOMY5mX
SB9RIkCuMtqvVURpA9EgWZsRL3V6E37mFvkXfVq3eXHeJB2szmeKjLjZc/0i59Pl2dNtuuLVbge/
IYvSQboF3zE5myv4f1JzEhzGTfgONsMrFyVsHKLQWS6ue7S7AZUBU4CghaMQSOvQm0em0Hn4NoLn
ZowHPhiVbxUWqdRTDZUpWgHvAuvFtbREOHjDYbAQNR88jR1NoKMwU3tvxvnUX0hBlWAKK+OUuoof
d/OmbCTjP7yuLXh9JU1qjblZO1nM68U9ypoPn+6v0kZcas4Srcc/1d5//X6KpDYdyPl6HNEXlrs5
tee82wCMKUnOXrPY/NdugGHT76s/HujX/jZ1UFS6MDsKXyUOcIB/yxCJu2WxSbmV3OVTngBIMT9x
1SmBuS0P7KNmzOwQdGeX4aht/7okSZqBVTYKTuqoLx65hg5hiBcnMQI3mvMSBU7jLhVt9JrXb+xN
WA/xtep1oHCj6IT+dw2Jqilbl/nfSefXkDgBZ4nUIJrpdOJ+kucxe9oQ67r2fIGv7cgPNJD9vOYT
aZt5H7AD0BfX3dlZ/1oNLXNYXYlrrRVh4IfJzUYjFdM+M2rokHH6ZH1FPfoGcZCi1VdPAUIu9m+B
dJhBycGQAb+oczmjeURSBpaUQWt72cfgTkimCBvQ8EnvP4orCxCpLTYdSpMIwJGzecvFZfh6KPkN
yQEXB4ZN191cnON8rLcY/sFD5eB9/tDPh0XdVMRYcpS/dN7JnsKiuOyOcHOfn9GYVq5hpjoLVTx9
urVctQAsYBZQ+udcuxtFj7C0P5zUc5W3wbD7EBEZAPwfjh2/Rx1192p/F1dw9vvVWqVSCfEGru97
BBQp9Q3+5OLigA1MEX/pT1LJ3rixTwi9kQl0oo3r2OMM+lPDcskdAFmD6sIM/rEWAl1WDZKQM4YE
78dtPVs/AfnEGz0DDX24LLTnF2h1SOvMcSN1jTY4AQ14uZ6QY1123FOlLCX7AxEsZKvNThrH0vDj
cg5oP0cLTV31jboAoGTUelJHAaI/MP1ehSaMHm+2OxR7Hn4Su89TQNhYMNmrsyt3gCdoEVWloXZa
iNNfSe2IHiRCoJ4f9UdoAEKEMZaSKXrz6/UnLMu2B5egG6+PNfcCu7IZ3OKQJWGIYM1ubGdu4xaA
fECvg+eWhLSiaVGuMon9tgV5Q56xegVBciPlI0a2reEhA3WHXmWz3jxKGWpfBJxT3VrOM/9ac12Z
o8k2QQIj9FqkNUDJNP1PCZapXp21PIS5ErVxAxxJZdovYNnTynR0NiiOHT89+5Rbzyj/GfnEIdlf
Qy6fqKU7TdaUbFUdGTB84vE5u1Qh8xc4iYKtmcqiyBoUlY6SagRCZwTy9TViQ1tnYk88nqpHblqI
TwpaQe0/RDls8Hwb+rC3Cmjdd+S4enILTW/WTpVrLhEH4F/8F2KhSXn6Uf2kmIshOpjJYz/6TFnw
jGc1BTjBZTzPG/wyDn713MS+W0OFu21xBF1K/EIYvPMT5xB1j3CgQSOe8CaaUVmrUAZMQ9/4iZd7
Q5pP02zxSqSg3uLNWPvoOdW8Vj8V6jCjWZb1wma7U2CvvyxmReijaQM1m39/1+3bxlNs028npz8X
t7tAQzpSU38cnL5a3p51qj/krfTYYdxDYxOgJ+NU/5CC7bnj6aR6rwCdJsJXZbqLNtPzooEsNzcN
VkWxAXz8rdg92Qnp4/eTPyHU/K6sF0Z+9dteo1UbWlYyBN6nJCIOCizz7kPxdJN7wyJ/MDiAlX83
/JLeMFAjQpxa4JSrAYsF9QCxQ5yQ58k3twPXyJlQX5NP4mMa4b3w5BLpfVqiccUfgbuNJXZoyqVv
Yn7bftdcPCbvNcK8E3WhDZAcyVWgA1YKHCWUsZkbyz4cc8rOuNquv9TKP3CJY3VFY+LU4tEpKxey
kKLhL9gO1bfhrYAjGIMJKKUTmlc2Y1oUXV94amZR/E5WxvsEwPiGdJ5yXjikTIufqV2/VnriwV0w
hrw29vU+IVWn/ZxSYrjh22zxdYd3jIz4n/iOGsckhpVRrCaG2zPCjkydXyVP7RVewTZ7CXoAtRir
3y7ChvODJNwzFMzqzcB104+0KriE5LCW1DzyZF5EC0Lcuhmz5Yt3vKste3nl2Mi2oYmDJnYE3sWz
iTj5wWJ7j6Bif/YTB3qRz1KSyDPSN0IO4DB1PoNhadxmsyPtEr4kFJQdQOAzsnbg6ZbWnONH/aZU
DHDfy+6P3MaU51muCwlh12PY+SkXcP9+o1jTCdb2T2rZDW2mkdWI0QLbumxEf1IkzOs4mmuflmOX
a8G8/yJTpFINddTWLoWDJNPLu/g/T7xtGP9i/hLvevqYUE7+a71NuFbQTlhAoGN+1In7t34uRWG7
Huw41p+YWmSqQ77wHorcnT/Wamp013gZrwI+hkxIKkehJFB0PawkecsVR9dwcK8ln68yl7bgjI3/
S/bTcZ2/XLAcbschj2Yb9LO2FhL7WAhsL6bNGQaMD7L5bJxiXiUCjdR8YWMDi48GQN+0PybykNdC
apyMQVcTvhkasfS5KQ5t2Gk8LB4OFe2lsSz9b1BMoV3EOCwTEtARNl4i2oqJRD0/atAEATmac6ln
u0ZvZ9GNFYTIC9MGLHTi6RmHE12U12NJLw/015HGE9tQCdV+v/4vJb7wIUZ43rXvuXn+YOkR5gg7
FVa28TjEsCeq+wfGuNMXE1I9wVfnUnZaALyZpc9FCMZD6OjrpHgnfPAibr+DIeuMqD4WpA+rha47
/bHpQ7bk5W1rDGSeoEPmwDyeLJCO8uyvOErt9OSALkfiq0f5P7f+HPYnWN1c9cPQTwgT4HvubC3i
nW5+F1qS9RboKilmZyFWrJf+PMjJccGpJI5BDayzsqXdrOdiEma3lnJJh8KArQcSC9aMyWGRmyUp
BuAQzItDW8S8xuWUzkz00RQOIhR4IYWuqzfDPshUpBxY20Gr5NnvdQwIoMRhtosRHboNGy/+xAd/
/G5yz6Xzm51QNDl3Z9yMhd54AhgFKrq2xtf+6V+jzQxq3FTEVTd+WEdLw9ty+R7p+apT96aYRtgQ
PwVygKuy8x1KvCqzYSzCken6r2VoDIsIBL0qW/brlYpwLLlkSiyZSIsz75xBhWyEQ/OTmg3VVZWe
oHbDkJZmqv8mmWo5iffWXWN+/PjW8d1RbxasEIvqRrtusWAQzlxhX6ZWah4dBFIguJrL4CzaIqk7
69U6TLzgG31m0yxVjHamrk3B08odjQ0VoKeAddTMpD9AafwFfpD+exbRmoOzxFJhMjj33X+Wmln/
Q5dn795gR5z1t56GXqFFFa9CgZOBaw//z0PJLSGTaeH84lNFKT8veUs+BFEr2m7YDkpopWOoXbja
LqEFLU2RNlcE2EOgzLpsa1rO+7p+d2RBnC2zAiXHrK/WgfjxY+T6ZLqZpXTh4urYnRhSBwsmcr3M
sLURrJYsPKZSmSAxfCAT5x1Gz4VLavD5r1+wIfFfr+KUG6/TEankgFNMr9cmQX0HZxs+ZoPYgSJY
TU8JgcpgnqwNQWw8VbbI4sEY8Pr3JGQJHVpgAdJ/dXc5O0KADr0SO3FXsU5r1eAU0obdg8txmYIP
Z4UhM5S9o0g5YpPZ+bQml1OV2keDvfXWfOvSa8z6ojqrQ5NYp3DJuX0nqi3m7kMuNwV2LGNPpeg1
aZZjuAuFv6uKi5n0/ZH1B0lOazYvlkHOsn2rK+WtPNqb/sHS3DfUJeVRZK35idNw+BdKZfl8Y8Wl
m/D++LH4eXFknc+ZiE55rvBP2QmMahC5YwU5PrOjxcwy0ZWDBilVhSL4W1msiI+pASIFI2yhxzMh
VkHouo6D84ayyVCUHjegBB+gVthEMUvnDTPeP8VsQYoyOt+DdrFkdYEeN+RnKIQ68sgP+NyrzUMm
kS0NmABvjw4uw0+jd/CzZdxtDXOmHEn5wyyhz6po+bJoi3ZpC0hWIopqT62du+cMtHZ/BldyqcZo
b9fldZ7cQ0WLHPI2z8k5YfL2IzBKBbs6M/Tge8MByAkW9vlZshxyUxVfwTWs1bhGsgjAzv2GNsy+
LzLUB2PSmbOuAEywTn/I4JNq42x6urKrcqcucPAiCV7ohPcEHi6Fr4vwTShgW0rhxSZ+dsoZBXCa
0K2GkUoh2u5aCyIQ42YETWrWRu/kJavQe51CxsQ55OnTcj2K2ApVoURBL2cYYivgIYlda6bXdKnZ
CrJAOuaMUf0YCfWdyVCh5LHrG1z/TciYV2CFUQwAJgafF4fK9+g0GWRPBcreA5ondhh8+NrFgBYh
PL4emU1J7heQmqqqpG3XNnZ+a3X2yy6gZ0WLpKck5kFLgJpVIzu4ArfeJNC6Qf38eI3ZC9PolkFK
RKVGXsIP1DEnT1YqXmjpVFbtyIAUPtSkNL6EwlzAmb6IqTWTi+ala3es3hU31BsHHncM3L7wspji
lRzYqb2ruNRU7jgU7bC31eQuqq4wJNg0sbf8AerAGfN1wEayEUabuY0VyK18hp5RoPF5DcLHMUyV
bug8xZOLmW3vk7vggAzaAyRmKVsxqVqgO58oMoG0pMFNsdyc/DNVEt4VSi13qhbW6w2KSHjw11Ed
M9QDwSmy+PY0dL3eQy9Q6ZATwoYMu2JaGKJ/6SxE+WlEShhopuiq1HBl3L/ZKo9q5JCCU6htSKQa
TbuXEg6ElHQgalkL94awDafErtkBpqvaIQqCMkcOaT5YoFS6E6R3ck35b7ymNmmkpjdZfdCl/NBp
ZzN6NkmbH1uFCoEtUZWYVlgg6lBUyjOangs3jRMOImtPLimXiaX7KZ4LtVOgts5C5EYXECDHVfNs
YiF9V7wF2Tqrky9oxtYfga+9Dy6Y7i9yZXM1B9jYVgJY+jeNl2LqltcS3Zmv8R7SL3n31BoYNI7J
1dKi1/Vg2f8hsT9NR8yxX83IAELCLVaFwrg3xt25DWwhc+ao7G8fw0w3mu73OgxeBfpJiaBwiioB
9CjqcZg1mpieIlsNfqp4lzORs05jNUSjCIto445AksMjMzYxhpTi2V5FtQxhlU2DK5Vax/aDl/lj
K7E7OccSJg4f9EuoI19/vh2Nou4hejTCWUtAN7Ulx4t+3OVV4FmGwADniVhVq94CC26R2PLrzr0B
+CK4rLa79c8WCzD8YOsY8RigejQ5JACqi511XzjztZlwqMAYWQs1SrAFWk1KdOTbgMUizPmDArr+
52gRE7yui8IfvIsHDebD6IYTcgHjxmuYxVMPE1UZm/VXAEzaAvw7UHoFbdqWWKGmTGkFReWmcCDt
23leD5Eru/Y1EDN51fAzf8u/EdM6SFYXrC9B2IClz4AqHOkgzK+kQ9KQVK6tMM9HEMKBasL6funU
TE5JokTzkB2L/75GoV+q9BUkMknP+YFqArCCfybs5o5D0E5AJl/v6lwoMtSSzYKQtb2t59vpKdY/
n5gPbbvTreKSk4c5GqHgwoZcOKTGzCocHrNV3vcKk8Mu0N8mE7FkQzhlbg5fQRPAmQDyVHGGmWpp
CCc+B/EYDT5StfrfMeEGuz/TJTs1xpHhI8kYBY54/+tE2r/4N2fqtV8OHbB7gJJIBBsGYZDiI/5V
M5NOVDhTPgMMtpu2nmF5n5KKTN0Pd/qWFU/MEhrP4g3dmmrq552wSnFWLSZ11bfe84CakXORFiak
nfQy2rx5jC4dW1r9RxsRs3j2xC+Bsj5+IkvpV0AX3s96cfTuJ3TE5QIcUv47mWkG1W2SRO9fKHq9
DpiBB5I+q3RpxEIntVeniO3zOQk3txHbVl0VgsQOysIHafcKR1fzJepyCvBf+lR2XdulRipWuJc+
mf87pYl3bhMyQpQMYpg7GR/LMxTkqWaZcd1RuIPz2zinMDLrS5YOgBgqRt+tzIw/xJIOahiwE83y
MKSnCjxSgvRfl8t4o3gH6kSpy9J5ZVojzR1R1xy5UzE0YNW9V6crKR5VZc40wlMvlCN9WMmm7QLu
H6rn/VWxLiPNavGpTuqTov/fxbae5LRzI75L0/1CRZHtAN2El6/UlRexcTAUWDArdX+V715AWRIF
zv6uK2zP7DlcGdBLuvJ6sOvlT++IYe5AMyUH2i1IBlwgvmdfhmkYc5WP3NePm07Xpk6t1jfx4rmS
FozvmSsA7jJbXbVbFzJiDVv2vuujA1/AhIiWKWISHcNH1ftwH66nZNskBiwpsTlAOJIzT+ybBk/p
DvpVFnvMAgjKniF0iqhP21K5HeltTa3yOzdExMN0LqHvI8Vtwba2MtFXFjvEiGAlfUM2wTkGNyvy
eRrew0qLmKKBiLZtz/qvoDdDH9eRXIUmgAmvDI4w92vhlOm5MsoUcgbiE7bA1ZImbZBsadurqUli
qjxiqRADIrHzyiS4nMdYD6UB5bJmCeE+UTnJxkVs0CHrBuFk/T5Wsi4MO3WNhMCd2V9q18YxZTgg
iNHJAx3nQRVj5QxY+jTLH5PDcPlbRlcnpP5rk0YKBXWKLFlNylH1UzYCci+yDxkZeQ0vIa7iI0KI
tDvmegmh1gjfQCFkY84Wzi9POhw0GbvIfJPQWNjmWIFDmpk5aNXBMwwF6W4T3J4HgkJk4FIcZaHg
GJvMbgoMyL7rGi7fZCeeQ9kcH88jfgboBlFUSO2Bl/WY7DvEmU2mACn8k1wmAHgNWFjUd82KBksX
bOHMuAfukLSc5r3OUk5l4cAtHAEaOrMdC9Camp2eWCmEdyhFNBEV50DEyI2mix0F6VVrYiOZxlZH
JbFnSsz4sJSe/xFysJ/DllfonaBdIiyY9/NdFjZlgdTFN8j22TdCF2+gc/LWVaKNqV84Zp5lXSD8
zPLBAf/HB8ga56r/AW/D4erTESR8Xqx1jpBNdzqbGMMF4Mn0YVvTwwLUSkcRHpnnfEU0hnwckmBA
dqJc4oZZpNRNMyIsec0X3pfSEsCarlqM3+Kk/tVHIOpDSzb5ob4A4ex5yTx15RYKzbQ2pF7o/g9X
QgLt//WopaIV4uQyTfRt+Fu2fd0xyp/Yw6ULFmJW4AJw3hfbYQOBNMu0U7qch+102v2eRZjZoBhR
kg0BUZz65KISA5M8JGX3h5fOKHwtX0/oMnaa6bXwkBfz2oxwFn8niKRAkVRIev/TcfWEPMxr+ryC
jgtAY4X0M3EgIfE/Zf3EtD3J1GXB7fdvvVzG3U3kabLK+d0cQDRMd2rtGle04B7IiT9pdHehg3kq
hD6dqxzvurQHAR+2mf9Ry55wOfDwhiGErRik1F/SZ9ruzgvket2XBfZcDZhAJiRSVVUJZinGzsVf
TFnoo03pl403biSne8WJX+B9Xm2PproQ1pJPnEs50kOHLY+YrGiqmVPB/6bbfV3GUnAtq5iYUVXB
XrftQZPniE4AQ8jfGNJ9R+9p+hU30nZ0/h3FaA5KSUslxzZK1RmOvq/2H1N5i97ch6s27MBh+kq6
wloLNFiymQzXVdr7XPXrTGFk1Y7u/joVVlXACTfy4in+/aV6jcnLjpPhxlbLSU6RR1WSbxWOhwZz
qMdO8JhPsHQ7pILhhCbUMEYNdHorm/0N19yr1Cs/pQWiotbVgJxk1QuoY9tToqMAnxLg4DY10Cx5
KwjD7ep/AdmG4cZRwggtf/vVJPyz06vAz7wxH9xdfEcE9r6L15N8/1NVxQSu+TI9eDkJM5Lp9ZX9
SJRxtk0jqHA6w6pYfJtwViEhJscOJLa4wj3EAPkojwIidZNeM2Lyxa020U25VRMPGCDg9aQKE+c6
8Wv4dkfjxi/cmFpSN+Tn1cFt9No14+ZfOjN+uObIeFgau5TJ9a1yaPhd7seRgMeY85NdPqR1Wmqw
ysf1bMxmOObZtWjOkWM2jpfH97DyGGENOqwe4t47KApHBNEM/SzWTcE+tGjAIn9eAhl9UVEk7dmA
mHQ15CU4MI67LRB3hYvRjEEFWaTdHXuUsOHgi2OLofk3XSnscDoF1YIb3HivgBoI8uOZuPK1P42F
95dCZIjIhWGNBBculR46tA4JBWpN2yPVNLEDhm3a1+87xLnOyOooulgA+e3Unp0uXmmd5O/2qSdB
JvR3LGmluOWm7R6otTiL7e0182yihX6Aggx3nhbRp+fd3lvYUt4Fd8xUP2gIqT4N+INq19Uqfm27
O61NcjVPGSccoPeBNRyz5dF6tluPs2Wq62oj3i+Ltwf/ASETd+8iJk+WvuiBJcK3jJ/eZS4BblaQ
uhKnWArUZjvKhwa/PqENOt4lu6I/FCpsh6tosKXL0P8kePnPVGH5I7pafKWrTFECp9tBdH4UT1fa
UE6WEpaUuQZFFsieZSgY29IcFbdaWh0ajmGXvEHRpuAYQl5XY+PtPynyW3cqmW6vq5MGz6n3bQeF
mJ8KVKP5XRZkXrXZhPXNgymSSJ27H9MXTkfCqrENnqS+AGknw+0t5O7mlNVeu9OMUexiI3weGRwx
xfCA0oPZjBTrn6l8v7tPe4d8VBoJKuyji3Lf++PUnu2Ipc9y+l4WkZzttGtanvhmQSjKBwbh46il
McPsTftvfAGmyh2zCTvAjwmu8v0lNpB+2B1lVH+H6FNTdPwO7xJr0ZFc1sCL5ruZs/CFwGSoouBO
JMe2iG095qyf+ZE2Te17Wk7uzvIx5yF9ZxOq/TJCtC9UFztow9/ja+cOcAt7ARejUhQf0LpQMQAM
hpPxP/QQVjoYRB+F7ofnI8Spc6dk1S6y4rsoOhb4COxc29MMUYPFNuPAC2ATocSa4VaN0O8QgZZ9
dogFyMMpAOJE8qtzA/kRDsPV2J6bBJyM+tDIAZERj81fPzq3JW+zHjoHq+p2H7WelTwsVZTnCmrK
WrZo7c9ZwYvu3kzFcIpi6xlbCjguSbdMP2etCJDtC8/ajinfnLDLNP+vN5pfXbnVZwrZ22h14Xh8
YAFwbHgvDCEABLO6KNjMyqPQ8z+qSI8dHDMM8ih5vjkjoiUcYPDt7yUB8jPPNws/vhRh7v4G2MmT
ixcv6ePCW24/s1UUkAWOXw+uxr+jf5ni1HWafdPxSlyC5tJxQkETdyBdjzAfTAaqm4HY4Mh1LLyY
kk04ubCNDgoPI9x6gKih1gux8rzwwpAI1fp/OruCrCwpcO+aN7OCRQHbPKj3fwSEHBTrZP6Kwz3b
A72azT6emJFmAd/q7BlsqNNEfeuQdZ7RQfi+MI4Dmw2Bzw7Q3xm+oj1KBDUuHJG9hPUD1XieAQ9Z
BLp7LpQiyqL9EZC5EwnquqFEc60nKaQ2H5nk9YBhSbCNd6zRY7SR+oNMilsmGPRjnyQNRcasa4Kq
HSipjV3Dznpvs3mr+qyJneGOrnJuA6IBcC0Wq8JXA3Hi33fsAHv0zTXc2h1WbzEcZQIcPzjNc6q6
qLH6ffxJDT4SOT0000f9GDKX/5yND4/oU6jgjLd+p9572uOF7xrk1Eb0hx9BdgYOzfn5XK/39dCJ
9K9eDMvD91d6OGAFIvs0h8z8tc5ZKi7mlp+WhQtFJyiiqWxVJhbGPa/U1MIEI40n4ViuBLsT6v4K
nhUmWZ6ATiGZn9pf3BrCNV4QwZZDn4WHg0AYAv7LD9rm1CJzNskQBbzUHH4HdNijpXACidMJIM1p
SwCEu6V1pq2+Kdq6CVO8MAv8I3BJvnO3A+g2qOYUBKNlUTMyRmfNpPMe9wtx+inpdn/iswc6l3Tp
ECqMeUAa7ofH4OVs7HSknT3CTj8Ik9QSNZMug8DBGTViWCa4p0SylKwMZ/d/DrwAsdAd8bdLG3g2
hfhkgzPAzPHP8X2beTvQFOXcScPF1AowUnkRecWybwD7uUvz7G8AEf+ppoIHMhjgrTNoyM8GoUPE
OAV2aD1mE3eZn8s5VgRiiR7WFbD52N30TKJl8wEog1gleQOxR7X82YjOULevszZh7FFCYbxVdDUy
y7dLOc6GylSlVB+6pjpOu/+S1/EeChhjemuClISBpqCHZJtG7HDc7oXzFLXjMBzh1WhCsAY+yw5c
ycTrYD5sh+Pkb/tHIHVxziDUa/KTtBARV1NIXk1ZZNFpnORHvC/txPzsDV+lB4dgDvBGsyDZwUuR
gzjwwX83oxal9uxbaxTAU8eD44ybEx0u6B1aSASOnpF2yQK3qlrilI2lVpIWKlEY35/BTEd5ItEj
9Ga/EynTxXMJ/wnKYWMIE+f/W5bf9dl+qAKVFPbdDP5Yu5savA7JGo6kx3X9xFZ5JxYcTWlPIIRe
Yl6+EDKXpVQ+TJx7n35gEvUm16ppe3M+t+DK8R7PlqyDS4cUWZWk6yc6/RzdsgsDN/NPDDNF70vm
N+Fuq/uk4QP9RjfQKXeU8x3pXxdq3legOgZ6DdYwZK8T1PhhAZeeJ3MAbuKiIvPzhmrISuAKCLy9
Ziu4LakqTYBOj53G6BrR0XQorAhA4f8ovZGv1WZJ6HODDvw4CS/8F/wLng5BzhvwhXfCXZjqf6t0
dIuS7ESCtdcaWHSTg7QwS8T7j1qjXkzuNh+NC+YuAF0Xieak9bpbPwxjHoiPADCH0v4WoSLD3Uff
i9Uky7ht7+X3F8yq/TJE9w/a1aKgB97aKzyOWG88aDAPbY0lR++8lPiCi3401Pir+22gSaRgJJQq
Rj/6TapSRfPjqD5zlLu9nuGz3ItcoJI3KoVl1GK5tAeCASJjg3t9Usz54jVdffIK6KMbxhLDS+nE
j2JELmrnJlkmK5emKkJE7On7O/Aiq1OJDA2RmdRxNGNQlepmcSzKQomLIvcyq4g1B2HaQXCbl0VM
SWaURiVaicbZn9ZrjX1xlcurhJmyxImIFm5gYhg3UCLJu/Kx/luQH6JatpddU9WvTX1EpxFXZMWm
EDepYIRct2bfUhMd2mpWNQZ5pE4DbfpZf1qXXxV0kiUJ0y+C7dkF/OMuz0l4rzouLoioc95YorPC
X/dWRtseQwpUEUS8iclSpRgy8ujQyYJI3ecuEMxmefJvwaIAkaPXcu+LEtF4EfizZZ8T0sUUWhnL
zDdj4cUM7fb91+JHdNU+UHjjLvC7IR7GVsTO2g4syEmcw/NkWWA9uq6wa8EuFX9Xlnw+c47Q0GTK
UdWf4J8nt8SQDaL2I9QQSqUUmJlmv1hKHd2reLvUQvzC8mXcB/wgesCf7jQCHHaPvBUG+RC3oy0w
qm0vt1/Ndoa991wmHy6eF4hUolfmzsdBCxI3zPm+hQqU/HMvaY9Rs/4DsozJxc2bIqpg1fd0lcuh
VwQOIviMXgTQs5fCMnZ+SWxlwdOQ59hPuSdSqAYUtB5BPVMN2RyrQrGwVQ5wmEnqW3PmLtqb7/9B
EON2UbEPt4/ZyIvOMvB0uwR5ZSG62dQnKa7XeNRSOeun++MKBjp7IAsjkuseCA4zM5kJEd66mRpS
m9gneye8MF1/CtGlGAci8mPDvj6YWL6Ts2GZ8XLwUB1br0kLyVc6OSezZXWRLE/ajc9KuwxLYZ9A
TKxv9qTQ1F/wVVQwrZB7WFBHM7DWls3zyoj/LymTstJx3wHvVrb23GcKx8kYfngnMZ871VpjKV9a
Sc9UWVqA33rtT+D35LL0QdakTkOjddHCWuD7RhPeyy5hX7ShQMl0Jb7pn0/kJjo1+PVpVLSmKjYX
ilzdWciTtie9k03P478fDgmmmVkFWhMWfuYkcuAL06cGkW7LfpqqK5JONGGnKoM0pRk2O6Lqs5kO
34IaOGiC1KmeEiQxpUSgFTrOuHi3NhBzuuIeN9hpJjnqMX/5q/7tpxsFA44TtWn5PKldej0QJVwz
xQSTXIWUDTGPJCom0PuItYpfj4OPLuyng8p6As9klKQTmNMzomkx6g6jlHT0KDNCI6vlzp2+nwtb
LouWnhoG0Jt8rv5EckWbRJVakgBIY8msudvh2GRKoQ2w7qF7aIli5iNxfpxd358Cgbkec1ofKqvZ
cUWnlVL2QZCCnFFh42Gx5XJ/Qq/dsTiGDJjOWNdvf0RSCzjhrRTs4HQKhklwSDJEYTnx1F8h2uu/
17FSqZtlTFzk1GWnUtVeXLU0PTXSNegTYmR+yExeqex4I9t0zsF/biJWwnV2jMMrqH+AdpcwOufv
IZLDIUOYwW+9xGSVMLvJluGDC3rfXn7407jCZVwUue5zljf8Z0kc7aD5R3004S2zYOSPsduzVbQt
nlQ8AdSmyb4VhmXw6FMPF1D9JHj+g3k5OmdVIR2/jHe2NFw8kBB6iMZi+PizmAWVb62NZcxRqXs8
dpbXhA+AjOF0H9r2TciTLxFlE9YPCe3o6xG0hcQyM2WLuhFo13knwW5qJLipV2lAL7VSxDz4SLpx
VBfWgSbyQ955HNOpYPkpdsA/Xd5DZXU4B41ODNAvwTQpNRqAVz4q6jgbrFeGSn/NYjgW93w8HKfI
4eA43q7NnHfFYYRZymrleV3hBpvfObJnFpohR8OFUZLgZ2WVixizPWAm+mABIBOAkl/w6DQryQyP
+OzUNLwC/Rls//5PapLphZlDvJaPMuXaN4yu/hyR66BuZ6fF5qOzIRvljOjhrtmdVWpYIe/PngBN
IeElwScU/8C64yjEuVq0p4PYm22nAF9n0zXs38aUdl4pv+uJb3MjsQJ8CrXU3Snn7kYKuLJu0bbe
XHSmJUzthaHW1KgiD5gtEfLq59V9977DDW3W2+OjPT6xtBwQwin8eLV9+1Xta2ftSVuoUTi9V2px
HmkBbIbwLVSejzMwMp6ZbCQxBzobsjlNknKVWH2uyhhWYKHi6KFkdNXHdPenBp9a5QYIYP6mzjOy
Q2Pmf1wfa9WOlg7vWUGyZeeYCP4RCHvzvU0H0ewGl5QrhaU4rxqXelPQufi22JvT8tfgcNKXIKJW
0b8mMqqB77wdSbyjCBS2Dmdj+FFaOon821ByHVH/3lQf4SNWMlBEN6IZyOdR6Uv5xmUoN0UpdlJm
qN31juzPFxEYIF17ZJY7hGuEhWANXGBtmz5z+tMDdja50Fik/e/QrK2yM6vfKcUb8zRsISA6LQH1
p77izCvT1V3xsoMOOsJkKBFRXVkMuaker9alMGBPHuYDj9ol4T1/3vmOJgbp6K3pnPixIZ5j8U8k
4J28HPd0QrxleAsi6pKWi2VEj+0ExAG+XjodV+6IOJA8HXJJFvlDyIImb3E6sganSflljyjp7Wzw
VvVd51Uh95GD3QajIlB97v/bipnMpvug57WguwNZibP5ZUe5IW59j+QKJiBkKrXwWO61l567zwoN
62Fue85Nhdv3oTyBA/FPGDgCpKO1N1TbvXzy2EtolYM6uVI3OPYhivlcHJzex9xfrrSFi1b/f/zM
rWDUVEpUQzJ58MzLWaBppIDNKAxlRHY19EK3JnoBfAshBKpDIroFOXlYklwEvGjPouwIw+AdD22V
Rxa/BzUK+EnATD+7GVobzofvoHhZ9HdAOzRgP68i/ya6S4euEcDObIXBlf91AU3H+LzKe8leMlac
/hKNyedAvr2pgrqvAiwrAIj7HmF8LdttG0u+CvbnvFRsMOVavPq4QNsNilmJeITPRHsrj1aovYrZ
CgjmBq0fX1kNP+SSpwstJtebAHNKjhPU7hvnC0ZMQXvWY7XZfb7GcgCTAV8id//mVM3XTD0KZQ4V
7ATl+ijZmBGGRnuz6v0fQ7PtSVfeB7M2zDwQNbYSRGNPrMy1+oVL+iTrABK50agJqSmFrJh9bEM6
/PBxXlUgo/fdDxE5Xaph1C6nWO6Za631gq7zipKsbw/NYB0/+d787j3Etzpu9vTgvCWEOkc7I1mU
sUH+bzVMisi7YJASXth00EttHl9ToNQLllA4US8LgwpMa1fMIZN1Yl+vcrG/XxVuLS5TajLgzsc0
88ip7bBhZUa1uA71vJgtFfmpo66VUA3CpOfPCpPynP9m7NmXq/vyV4MJliKvUbopIpG5CC43b057
6VJChPanQoHrK3TWXoyA8VHid1QhorXBIBJCrnJu4SVc7q84tIucL/8utLVxWPaVere0Wvisw5gI
47kQJTxWjSN08sdgYd9XibVs63z+0z9/pVq+ExOuL6N+P0NItmyP9no2GCMBca2MoKmdboNNjqW+
5mvcdY8JeLJNRlXAn5RH9i/xDsjLmroGj15DU8NOvifEPhM7E4HMkPhhUefLe3Z7qIUSYWO1kbz2
d+Rx2hRvD1XArD0I/6V6VVm/rZxQ43k7xQTWoNTjeTIlkDU7eS8oaSsTGqgIsz5fmdyk/j2H5G59
KML7TAucLLmd5rAkl9yQwy3sC9j0jQ9MdMrlZTwI6eBQliS1pdCApl1Yo7o8am+HmmVjWCSdCwoi
y3C1LLGJKh5LlLE60W28jc/WP6rNoeXjn23Ba397rndmiESWsnxajhnOLPqmp7yX6rribs4ZpSWu
a5qeUGTCWK6J+kTv0FziR4uXEzfUn+1O3jhokIyAeeQJBszfHiwkB6ZsjWjQdshR/aeKGxddkTT/
2l9jnuON3yHgclIeAjc7ZwoyhjonNoJMBZH/5N5an9sDxehDsECpVSbx9NWurA8gHtAjW7rL85e3
wKaYEppV9kXtQtg/breyVxtm+ByL4bk+AIt3OWWk8fAGePda8XxPOC9QyH+YqMZnqyeaNawzvUFL
GPQoEhkharZriK81/hsKbmdFbAT+10YXQRqfXkakwEh3RAyV4aiYPx1ATezc46BgyV8uphaWjKVc
CuW5pYzK+Cvo8PT8WnDQPosJHkneN65NXvHUmH4Xr27z/e0xt49Q43TthvoFbIzex2TOX7Kam7N8
gZvvZmPyAIsTOOmGpD6Es2r1hBIwkMcqXNEk6TzU3Pi71+Lc7LBI5pv1sbPOx3O2gJt1+mhpB+JJ
F3LPTpa8rsjpFld0niNKXpWSFl16f7My1eW8SzzqSnS3nGfJgu5uF8x8n/X9sFXGNTgT6UppTkdm
VOhIvD6x3BrRXPnyPr9YWNUxVDmq7zwJ5oTeBYWy+X61FGYShV1Way3PkfazvkEavZkKaZagCjxk
8HZrtobxZ2npv2gZgxzqszN8MF/e4snDy/fMkz4BCiBCf0cUq4FswOTCNp3bSfT6cdLuvh9TeCtK
t/jxw07mGI24pDFV4XyZkY6197/elsPvhU2osxDHzIJzcMLXvY1YhnUzLHfKwC8h+v+n/0NhTyyE
xCfASs+ak/y1NzgVl1StpYSmBLp9h/MjLuXGQTIhroSkUR5sEo3ewD4Uy1rYq5XoYjyQEV7EULi4
lAcPeBHWLSsH63432flFbdaS1eX7Ct35lgiKjcxbc+sGlGTZR6axXG4Xts4A+c7/XGkdXj2Ks9PB
2KOJE9kKRS48dD4p39LrkVnAlfFlAoIWDPZlojJxpVSdzVstYiXgncNQHmouCE0WjH1gk1WYHyxS
42E0oZAU7vlssV4fqPKNIPpp24upNJ1UhqH8EN+zKy/D/XHbysFOPLpmZbwBOCxy3mhh0xJO0BoB
smUzcpgwMk9FKYvyoeZEukW87uP/JxaQFWbRnbTF+XkLVcoEyw2BUUYQIbvc2hLDzO68vLX9JClh
mfmd63mGlIPezSdUJZw0AiV4pkVliZp7UTLb/RfsN91kb41yEH3t/BtEaOX57QUbfNnXN8bkqHRB
k8b461yENolK/zucf9cGyyaH31kmnPvZry/KbQFzEUwb+kp/R+BqnaNaMF1pnemwYpF+RE8yTx9a
mt08f8IcthooqWnza2duAueA7aWKT90LlNISRb6yVy9I1Iiw25/U6LXXFsLHzhJc3O80KCtrF9QX
DnQzI0lPglVjimT4gywunUfphERYaWMoNZ8Bc5V16+fHB16JkkBEAAss+Jwb/x0An7axhjz94IcD
9sJ/1wLOw2E/7khGHaCsOyiDiAJk3xCcleefcy9wLAAvd+aqzYug335bvmhKo1kjxS5Z+lj/fUty
YOWKuJ21dN2hA6XBbiXB23p8lVA8ft87loxjKJxr2F6stlH73zQTOOkeWBAMkYQrZYWkoslbN3i5
Hnrn/4dc5/Ze7aAs1V/8gQVh4ORs41gSUMkuxNF2FfsE07toSIM9aszRxD72WdvkFuJL4sEbp1jn
zhfELDMTnlgHtJYKQy+t4uckE7VVsEpvpwmDk+r3fibkBOUI/pnA9aIXcZvN3xtXOa2WiKhcy9MM
C+8ezBnBLUj264dhSw5hgv/lTT8CQvgynw+UGc7qAYM8qBAdZjdqzQJ8jOHxajrJqvaStRyi0S3I
1tgyNam5IFQ5jcCU7Jaum5SYeHRbT0F/3kH4ACwPY2xTOdZA7lH0tToN5NbnixS6xTmWtHGzyMMZ
PzI4C/URTRC8rL9ZEiwPTa5wnuze/ztycVMDTzuBZEE45J942l/pmlHziHHSJD+ToW07VoERmQyH
b+OBA9XgQ5If52xLOioLpwcjIlGXpoNySSu3uGm8gTBp0itFSlm/1NGhVg7yIZ0gpe513jShPqQK
TyfiOiS+0z7UCIRvm/kOSoLDnL18gCUTufI1y9gBbJTjq9ElBtDwlBjk9DZoJjmA1gCalik+yDD3
ezUCBkM/wnNKhXvyjGAhRYWI5GYWI9TDjqyCX6cKKdF97+ihI+0WLKlCmk2TrUppVol4j1dXY7qO
1Fm/Fs6tuMysSNkz6efzoZE9IuClNYC/ky5Gk6iYrBRyCjaXDJqx+it2icPpPuRwVKeGeUAYbCnN
Tb7bzqrEgxXNnARJ4vNMY6zIVS5TmpW/r2RRyi2T7QThagtdzs0cSmlhU9xkXyIkfOiWUK5e6YTQ
nQgeKiUJvAax0hBtPNSsi+dj3lzojFoigMEHwRLvDJoMiMnBX0/v3AVwQdRSvvDwy0Wyrw00F2s3
sisQAM60ynr/N2eEOTSQI/itVMDuS89qIHgo9Dx89i91oIN6+XCiPlHWvG47lAuOUdFEF/9T8wEd
zDM1eOkRqUaPbBukC6OCKM233A69aeGAXb/LumwUj8GpBPXIOLhKcXhx6Tt/2+QLP51UgqkFATGh
IjSIsjsoh7xasrAOyB+8H9qWgt/fz21JgRRjc165323rPFyqfL+X95sl1Q/+RYBDemtaeJ49Ehg/
1bTWh7UV7dDzPb0pJ2TZK4CPON/TMaAVvhtGo48AxWVHLW/Vd8fMWi5iwsD5BVdt/vMtk052Xmk+
/MmjR63ut+KXnK34Ov8tAssH/Mwni/Us38JE79LmjiaBGjzEq2xAaIUBGB1nfqiEMM502CC5yN00
2XD8wenu0cPPNyNSWO2Rdjs+xbzjRlPRWQUEWYZEmoRfvaU7R3shiD6im1RooZ5c7beWeA96Lv04
Tm+/oqW8eulA1K9itqtZ4UG/Oc/PV02mn09F/GsC29pkQfL01Z2/VdFrI2I5Ewx+JWIKAt5k7BQc
9aNBe75TAH5rqspYsaEwXYRSpky9BGdRsDrJ4RXoc242pE7nvUEG0o3V6/5g/aHKlf+IEumegoIQ
X9Lgsdw944xHGu9hpzm/WRJClXGfNAWgULq3T6V2VHWFlGwcK3lzJUXQWuN8D8oDBBNs2yevGJYK
GzyJQYm0F87FjUH0MKtC/IE12rb3IPfatwyVx6WltLu7I2hFyA7O+e5ktAn4t6lYusz7gxOru2Ap
JSjWxznXif9Hf9v9z8R9a+AqrFD4k4JgDKVVpctGLWOyldbrkeca08Mj62MsqgQuaoP+KRmdzIqA
XAkWYR7jswfvteks6sP68G1TsAdkbErst8y1OgaLtwPgK86rmdAIs7Rm/lOdEn3wYP6jIznXtfe0
djAnqvmR3ljx0CmYGa7hxyPEJlZ49bSQTGudjfiAMP8P3ZVwGb/4UalfMpe3+HincusESXo1MEy5
ovdvYRSYvLqkBLugE/r4f4+jmkneabjyokXm6LTNVIOYXulgWmind9uGtTjjlhlhReNphcrqLJo+
DBUF5y+7b/TZNqdxKA0L23z/jUwFLbI0GJm9XlYRNbie0r1yi5s8h26gcjL3IiOFAjbYwLBjmddv
MJIJjFtpLW4onJCNqzPHpCsDPtsAyHCrW+tXkEjkyE7o0h2x/d5IgjGLfCtWIH/2syIQoxQbP0DQ
0N3rBBeT3qbDeohWEbk/ZypPRPqmvsVxogT6sVfPDpDurlS6D2f4tdTSV44gS6z/K7ht6Jvy/fc+
N+kQz7RPKSiSx24xjuFEb9WaTZA172uO5L9ke9ZQr7fdp44f2EtguGMQf5vQkMlfTN4wd9SgWUyT
PK8dN2LmUaGrZGP7Izq3fLAETinC3801+LQF2zgoG/aT47zqIGEyb/z5HelRJYunAjlr5C9f9qiK
i7KjY/okKtQIxZrnh09blC6nQNryEfw6sCXb2bKSYFpCO1pn0DX3rG/1H5TdH53W1B8xJ8Wf1Nod
xzJuVi/ZWvoRfwydx9p25m099dmT+sOauSAZFXn/T67L0WnU/xgsXcZrFKMj5N6vCK6sprTh2ltX
Pwf9foIdHQ2YqJuojkDt+ZH9EaREJaAzlXVEcFNB45wLISPr8RT+ha5wbTe06DTnBF/6k8pjpVr9
2pUvH2GBv8RMzUGaUVArn5D+6DQ8NcGWDku15LFuBhKdoDbUEhDJBVWqL+f6S2q87fs1j+ywqOS6
BYCYtIgrdeI8MU+5eJur8SHC1Q+/SoDiMGIBeUhSjr+oMwqDtZJm74vmSTkJfgGWo//xK9pqJjIF
1+wlJDljKB/km55vJY9eWFelcyQxebzkJraTvWhuBKQSFjpWDJZKlv8fgf/ZT9p30JpIYW5IKV5m
qg5VKXV/T+5RxxT69OXqabTczQhynBqBoxmDNKPgGKJKG3VYYJEnaUxM4NCZ/TlVJCgqN+pkerkZ
ko63MO/PQvJQpQm3i2AHWBxJ+rOyGK9s1P38s30Yhn1LgGPIh3G4wxtYguOAdHmEmVcO9AfyS0DK
pm/DxNwfHY9/hDamZlf8ulXMlFm4bv7vIk4WZ2hehQjUYQp6+j0EwuN3KxDbHf37bmqq7pmoXj2Q
CP7E7afPk47TgzYrwRyIZ7AFZrLk04PgfS1g3KjkLQwRm+WXgB6FsIqhtCLPMMku3FRPXWFu+eGX
PTP9Jyl0qoTSaaBIvk1EZblcPPGHZvittMU+0h7CVmqVB95YKWg2D99JbhI/nvLCEkqVjsoRg8Cz
l9ddqiYGzW3FzKynhZUhTD6wPsn5gFo0lffY3RMkVdaIJtxgok9twIhYgbdGJci6aAUTwVBU2g1q
mTV+IyuWgCMwWiSBk74xqcy1vmmHPzbX8l9ihP4fzlvgM5mFkvEqcHvgaRcVKIKPNZnYnEWdoh1M
YKaCoVqPGhcEAyA/HzXXkK0Rfk4nWiE6R04rkwnPiHdw59GDKGU/cy3RSnSzqQHFdrQWmDeAmhA0
QTE+AsU+WRbxBt2tU6D/75DlKDC4TprYX7zjT9lMUey/C4OcxVP1u14BTTekFetyaIClVQv0xh08
fLIFnJGvgHiBiycMp9u1xSsKaE8Qd52pPp2a8HPuJN4sr2uBkRj709OKpdR8CAJoUx0Ja66kRnfq
lzIhAFqC2HTvbjFZPVPJGtniXVQ8saQ28748ejoobhR5MLuIAx52HOtoHR1mSwOhbW7Ez7VGW0if
nRxqjudGDZPocCV2RULvfGJL44ZiU2ICbGETjivPk/iB4rDXWZqHwlkTl67FXd3XVtTZzEMB85u2
1HlIeykHpHlL0IwOoBwSK2M+85PFLh6VfcpiK2ERLUInoGFyU0XU8JFofpocXskgKoLCapCoaesf
J+cEDV0ssgIyZNgl7JYOr1tJt+veYT04UkzkeGzug/8ek+ruMj0Gc7f2f8eeu4hps+wIJgenTWLu
+3uxIb2nRyG18nYO1myhaqDTmUq4fVluGHKFQ7+NHzdDXxQn6+pGbRFmaNZxMqnghyoMokUs8vMp
ikUZaZyP9SdH2/CpGn0PayghNbbeNIFksh3jwbjQDD5cWBDRd81iKlC3AQVYxsNh/tM3zg6XCTLz
ukw+6pK02QwIeuP/YZuSryGpZwOav2bflt50mwLywL+/qao0PO1UY6q68z/K+9/6vhKNaOaSLZtI
lU8Dlq2GBYKy71u9/gCOCK9U7zh56DaRaIbppvXRcs4bLWYxNYDVDhyNnjYRegBG1VgeoYS63hUf
/xk1jBtlb6rjjSSrpt4H6TUUXak7iX6rFEZDuFs87wAkWc2M/WUwRXqv50kD30d1H7D4BzRh9bmd
RgtBmfQdAoxuoK4+zM0nyKP+LmUZ8ZJwIaqczLlnGWTm/JesnMmnVMnRuLl7Nu4hWJ/Vy8H3ZP0t
iFFm/hgrHPbMbAqCkC2ZHn7TbtvLyeLWOzIyB1X7Am3OkS13z+RE6l3HxVNb6y4afYhvFQQmTZOF
rqEPKtuwph4WqJhAjL9APda9MiVJLCBaNihef4VJYXCt5T037Bs6d6hGYeeD+xYQRGYkvEZ1ftBr
mClyNE7mUTI0+Rm87ahPzqknA5ofi8LhlxyTR+A4SF0yPQEH61EscKiaG1s47kwwb8CH1saab3eI
kdA/HrO1EjdeRylOmE8yRYmQKVaUQchxQ2WcmxtgQ7zw6+IaLI5SGBKscwD2107TLCxI+KSjpgdX
Tg4QAjaFlNJZh2lOuABIaC/Or4Ep/eQCVnpUNjmm9RCQN/dL2/W1Ql8OOGuGhg3vxOn62F88yU0I
wNUAmqrrk5Sybd5cRGVMIOKQndnD56U49OHZqj5PdALpWX/pErMuMdNu2h9CebkJq3/eYODlSw8/
PY1z/Om3FaBoOMYo5omc1NyGnjv+DrAX/c++sY8c+6Vgx8Q0o2eyqfAv7cQu3L9leBZHqr+PzkPL
86HPhzccueh46zRLXfGWv7Sd4oBrLtOpmclg6kJSR9RXBwDRDzBMl5pR765Il/wTroDIudFA+eIw
VP032e/HjtEWB9TqL/nlYt+qi5Ds1bwOOIVlahkijS3sAwJw85RtgXTIgEnrUQwD54Aj8aeqonY4
kFi9+XDU4acZHxLGqmsdJLUKJga/re00MWnrE/l8ESTv7idORzlvCRtsNXlYNQPwU0iVrZoW6SQh
R2V2tVh8JBL1uQr9SFd/jZd6Qi1J32p/y0t6CSdM0YVUXJYgFpA9r9v99aX2b0ySuVNJIj8blhCO
ToOzHIENcWU8isWaqP3gv90ejCjLTNGTnnyaZ+wXAQHhMcoMT6HQRK3PjJj4hbGXtFcv648AE3ld
/SJZLwvAvRu+3WgxtJiAX633xg2gwUnlqD1IYTjiuMBzaGbKtf8N8z8u2hRBVUAfG/yOUsQc6vr1
Q8hu2lYnDa4q39qPGOQ+zowtpUsbJQVM7V1Bo6WNkka+QtynsTVrxqqKSfmnpWCcv8JdcuBzmjnZ
wPrKOG5QeyASweSzplt9SHcEaa5IhtHggvx7Aw5DGmJMqIJZQmBfEXYk/+f/nnyML4TxUzuyjW2y
LiExsz7jFrucpmk5U3d6/HiSSiw8xZqz09ouw9o5nkzZ7ZPC73pzOBzl2k1YLRbXJj8bpwZBa2j6
BuM8qTIahHXNkoxY8cbG5WMQZt0nTizZ0HMKnl/QQq5tIdIw2r+07G2qV1bSME1sXGxgN6qECFJg
MWTp8iuqfsdZ302NeHUnJQ12oVRXOtGnqqmcS4TaD+dKZ2xmvunOLsrsWOwRktFDOpz18s/nXY+B
Q29ly+3dwB8d1GKLY0fV3Ezp12fWyQj8h2gKR8W44peRIiodh6hLH8jKGHUT5PStsC9TpResUNKP
yMIkZ+0gS5HEAM+3A3mOgwvU4Bq3/WBhbQSlsqGj4Siw5qhiZsHUmXAnDeHS5r93da15TCeVHoyA
7rA3gp/q4VEo3MPt7mJeI7UlajO33u6f1YqgQ0cYe13TyUu4FVX1RYSTRTcGBBUdl1uuOlP+sKOX
z+eZVsdy+/11aEYY0TBB5JXR1vqJoQBOprUpHJ8aExaancG/zuOEMnWK4jzbucBHYvt6BeXsM40Y
vQUQzzn/ABkeKRh+ce/+vP0cGGJRVNXyNd5KoGUUfZ0nRGZC7GzoHcFqBjEcg5P3+KSbu5l9emYy
cO1jZMuHAffqg0pFK1jGesqB1FKeu/BqV1WGEsVGfWqsZJwZWG9MD0pIhBvMqbYev8oFoNdHse0j
7iyGkAx+TCk0Zj/2WbuKkVoCeSiaWOEOc9esXRhdGmD2iLpKXXOW7GUhZrjhD8HpM1AR+pqX4vhN
lD3JYo93gGI4YizDTgFmAXvjE6wg7L8ej10w8EJ70vhznd7DXxD87WzCkd0jy+NzwKORqFTTO4r8
X2sagsP3Yy/+EBP0Cv9/eoYeKoyjBKQsqV7js+Ru5YaBelZUiv+80FGSJgB0MTT+9oYuhH6FzgKY
lfUxcp/6UWy/GIdjo2RuM1C7/ysV72MMZDVQGe04PG1LQ1owKpA+h8S6SYS6YjL4jqPXzN6nMWt5
UNM9xBDihLKNniduOZjh/XvSuEBZniwCsnK+tyWahMUK08cSdEVTlC3qpFne4wlat6dWu7BP+FlE
Inhw9MAZ/XhP2ErRHU9SiEKCy/DCXecrs1vQXO2j9nbwr+r9tKbflYfB2uvVF3bgVeTn4qEDr4Fv
2tobZHLQeJPN1E6HmgvgGEYV4Hv3by87gc055Nr80g4L2iAriElvE+lf5PykiGQpkhlSeXCppuBd
ES1SyggJUpxFF+TQxYiFisL3LhmDbvLqyB3rAN06Vs9LwSAMu2Mc8+KfLWD5FZtssBbdk+bGF1iT
3c4hu6k4CVd4eD/OJWzkl9y/L4G9vmdpuL4QHXKmoCbuCY32TslUvTl/2CO0mJmdrwPVXIx+mtyE
evJWhScl5ShPbBvc8Ih2BOCKXnB7dsJ3mmpqjxPoUZvKfJWOKXEwi+2Ev60xZCgWhLWKH1VS28Jy
TZtHGZBgx30PT2mL2RknEpPVbIl7BK+meuLwYSBz9sb3xbNvWK+j0xuaI6Tj5pHkYODe9ZA61qxU
pXgV2qRvVD/YlvL7eoGpZbtzT0pdghUEEBkCWfHcf556q2JlnBI4pMHUAiJ9fJWsIkuDWNctNA+/
QI1Xn9RTDS29/W5DHk7VB+84b2osVCaQYdN51Zm0yrQ5ybQnuwJGEmAYx1DewAXsoB5V6GsykIWy
ixSQPImHT1dJ8aoHVFT9WgVCGSgYAGrjn0gzEBoKdg/0wzen6RI/G6Bxe287gzm/NW6JG7h/mCol
4dZnCgWN4ZGHBYOsEEKM1loY8nwY6q6yhTa8Jci4SItkdYR8gRXTWNeBswapkmbCBmRFhycnejwe
nJrH7rzuFECbws5qOk2i8floLlS6Q0S54ns5jtprH7GEnOo32HwaA1iOlIfsWujTH8WXjQifdfTU
Hf/K28LDrDnABlFOaetkLACkhH6DGOgGLX/HG6UefXGL9NhgKQ6INgEmbN8S2uYESDbABSKuvH84
GVOR2a2XY65PxDAJRdCGJKM3IwIDuaj1BLFjiDRNSMmYjkGWCVAt2QuXr//v4EjahCqjjEpYIf/3
UCO9f6G2ocwfgfmzO28r4VgDz+ZFzesbTtdzRfoGheztWJe8Wzb4tBmjP3ACTceQuWNwI8cVGmJ8
Cyiv+2kvcWqPaKCgL8dZqWivrNXtSshfizsYJXYPvwa1wAMX9vct8cJLZR6lmIfWjhnLK6P2QWaj
iibQJNT03Lr21pG8TWPm5G8M15u0pmjVACXlc8nQYUcyuMkVs/p0e5Rc3nabnaH09izDKQhnyG+0
JdD8q3OGKE+OXsKY4wrZqp7Tb/UeqskPekGou2EIGuqVRH+5Se+NdO4ZTTyarHO+SUpwq3LydMoU
fXSeyh7e0pyQ1IdFhS5qLr5oGMGCzHg/PlLLuyLjlkCGGKm66QtlNurqFgSyJPUekAinVp3u91W0
VfjU22OHegGOUDXxx7H2Sv351KkT48+ygBpw29s+Tbx8cM5FJLz6UJ7iOdq4CJsl+i2zKE4hQYEm
nyLMaYlUCDiDfqh7Y/kgFxSTSn01fpVZ8Fr+QTdRoV0KSddLC6uBLavlOjjVGxMMi4nIDEGA/al1
FRcBhulrWAI6WdcF/iZ2gKJYyTDHH8cDdHy4BSsEhKLOKNq/nG2722tWGkDNDcc+ivZAyRc3yO2/
er2Fv2UxzkcOuwMTYzO34ALnhmTv8pSn13OvNRELeoDgnWgK3uZoNx7A5N401UIFhatmGjN7NiZF
yi9JIPQE7M7QxD1qDZqHQhoqGCPdSg78cPwodwPMY0XLmaV+2gINKiSmwQis0Eudil4YdjG5I3G5
7Jhsx6EjvLBjIz2lALCBM+yUq/XV1nd0QDR8JcvZQXQz+EV5Wlped1vm0v399ObIY7Q7tvKlb/bJ
9ljnc8nq4xAZBaGRYWCfSLMbDpxM2DRnCjpsY1PtPRC2yOjBLiMz9d2Rzo8RLOBhOGlfXojvYxro
mzzFu8+YWKkNrU3CJNupx11+WFyHxJgbNBtckxE/5c6+kznZ1/PIVFNBFlNbDsziZPmKRJlFCzzm
pRWEQRMl3her6CsEbwbH1l/MWmx9V3LzbfnLlhLk3pgLAw3GWfIM0vsz0cN4ZdV3iz+8cYysReJd
jK8b7K68fZ5S8C/7lDqN6ted6QW5E6V+uenm/HbPtsz4izQlPhv6MtGrXXNnPWb7K+xb9mgszDDJ
TH0TlrxZ+ex9R82dtXjP8TYRdBI1SUXqRktqEPhTNDHvWMCuskE2auwWPAPjfm+rm8Ko6iXDGcFk
F8OakYIZqb8qh49Nw4zwEy6HlH2tF8vjn6KqPkpzxymopxngkduNKRWcqMJeYAS99bwGahQfCY+n
woHnDCYjqD7INVHYFr1cdGlAE7QK/vPv2himj8Y/OR+VcnVBFScT6xHhj+KbHz972K1P6PUUy5/n
Uco0Hyx1AEJFVC3Vdn2OAfG9bdMBNGLxylkdz1VtfV/uNnnnRGwVo6PgNQ1v3iE1wp0aLzBH3sTn
ogDIi+XBdSE46nW2usYGzLlBWdwWRjR8s/eR6AcCV5pKtAoDOGb7v1brvWR+VO3JR5MZDAPfbHmU
OXcgBbBTvgUtcgYWn9jZYUnkVoOwmOdILd+w58JkWnZ1pTLr823HbJeB7ynUTnfZrhjCZApq2kGt
xkqnJVGXWr6ZJk3Klsa87C0YtWHGnbNtXRucykRyUf0eR/nKevFXdVTfXZC6xKIpkKom6ZT/tsDF
yhGnVlwfwdn7aO0/8a+HXcrs12IiFB/PscmS8sXwlIyLZ/OPcwq3Zrvd2Cabf7eQEfcPbkywqTKi
LTonCUJO0xuS1V/6OfAJp5oe7EHqYrIk7gMSoHAqhehgO0NrGFXYXYEXrizE5aXMVlWI98jnJHcm
WypmMGv+Hjid9UL8TnBJ9FFhCWhAW700FRF0gzs3QizzCDjxDdjgCF0q4C37U+e2S1H/XW8MOpL/
X3NpPeL1sxRtH4Z0dkKXZ0pSDKyvpFg9D4OcmGlOceex4f42eTaieqaxkcNsNQOohI4VNtB5Q95m
eFkmBKBSj1e6BFa8mjsugH8ksOaheIhY7D74IbOOso/3qYDnb7+mL1jIa/hxx78TH5DA/s/M7PLr
coVdhbuh3fafE5a4KY/VpQnuJRTibVVzq4SJKElbtgzuZZDlHSqaiW1NtE4z4qfyA7JsWgVkMVIw
3P9a6Rodbn68aNqOOH4+Wdgn+Oah/PcyvqLAKeCNMsRFXAqJU9b8mxmYu3VWqDeZdGmaQIgC1chL
udVXDkU7ftCJg6gPUluPhYSvEdhP9tJqPex6HO0hnE22AINy4E2Le7NNikgTM5g7m0WEgyF8N/bk
OAvR65bZEHNV6HRDANlxP2IeninjRSEJMd3nc8pFXAAFlHzirQpHAa0wUD1beyaQIfcKkKUWbgVF
GuFpy/znydaihGgkMflOkS689uHFDjaDjCr7dJXn2XPf/0uY2pZeACKrbeJ2ph7QzZYmxI/zg/f+
6swjjmLv4VQtvPiUpEb6i8ImaQomkIK7N0fsuKCcCrvZGC3FvqJohKhXs4G5lDdUVwqL6KsiESSx
cZInlnsaMlbjSLASb+lKndU4xRBwzgtHw0b9iYHG7QMmEPnvzcxxkq0hQanGf+Q/4WLuensnShda
LJOgEiUzwXUsKr9JpT2yS4F4wIjVf3POx2AQF8zRa/+u18sWbAEjkSOWpTquRoms4nXqBe5HRI8r
+VDAG0Y7IxZhEFp6rWjtFjHL5Kh2o6yyruWHDesUAkCJ4T62l5ee8sHJXgaSEz/tBPRljudqIuaX
fvdJqn4Uh5MRBnx76K2h3im3GEueYncHrTSINBUbuk9Squq022XCtrVpHoashVZ+XdQYwK9Uir7Z
WdBwEmiggbmNafqcbiOFzdApDClLJIVAS3K+62WNko/PF29P04M5p8FrtJwqaaYR5gpQhTTHQ6WS
XK/Gah1jcUW3OU8sv3rbEm6Tsb3FMe7ZhAJqURE+cUxshUrSBrIukFw0OnQJ0OU+2uFJy5sQnotf
ku/Bd4/mBFwW+3Y8rZ8IPVze+bMUC5bbEC1Y1QMtFdpGdR5vDJtvPcpOoTOP33xRCj4Wi6NHTVsE
UPDyQ82stZAfTmWzKdWZd0wFnKsbxk2VPAQe3jLKnl2LiQ7rAMSYZrzkjvLgswAjcBPoBr3tfXKG
xM1vIR0M+T9DHQzWYismG53ZdoZFRhie/cbbVh7JfhZjp1/pYyczSm3i7oWfDndcGy89Q9DcXIA0
MCWM0x5OJl5L+gM3GV3XJrHb4UlqLCjPsbkdMEQp2xXzPYj/bcoWKWTZmXQhLVPw5OV/MJI7EwrK
cm++S1r7QwoUAQ0tkPg4ZV7QTFcHUUa4rdwk+8hqVOYSCtugziA6dcJxMtNZRKaJQxy4gvWXxxrj
0PgICrTpHc9GbdILIdfrfXIurIdyPyK7b4CNUwI1jb8ZxSVBvNIbaNOkIR0QQYAt1MbpIon30I5B
cnPPxZHLnZ9UyhYl9OPg86bsHjXQyi32OgYv4X4VBV+4Pl5tsbHH3AF/12iirQWqEh0GwlpHTVjs
PZImaHG7YsT0FfqMa2RwW7WDGQ7VaS5EF+h/jfm194z5PyGXW8Bq5Aoxwo6nFTTN/fAiaYVLab75
Tw+aDEo3SAfqku4Qs8FJSruv9IcYuAdjIxoXmi5Jan9+YDt2FDQgpLdqFEfSjK5TPzSGYgjhmn9x
5aTgxqRFrzNVEwFuXRKiwt8oaTI44ihtZDk7HbEWvdDKRaUBGkLvfQ+vJOmlumKANRZnOkECIXpt
3u/J0Ym7cwdN9PHH4rG+ejhzKJDN7KQSks5DwhdZh8hDcyP/rb8yEqs6FrARMYbMBAi3W39AINMh
zgFNs/SrCcB6Sx1MB4CmK06Y0ZXrGMHwasfKh8HIFdTYplY0rEU1/Kxs53+QPtrLHtfpOcUZAkxZ
I5siXwij4VCzg/CFDdcyR9fJt9pYwXJE3RZ1NUvJUsApxV+KfD0y6TksTB3T21wHpk9pdXgN70TF
9P3cpleeldRt4jjReFkNl0kG0AbY1SuLW6xZSMAe2CWbaHCe3KTXt435ChtK2hI1dB6knqRxkVc8
QCv6n/JOpe+K1x1Gj7pEB0RC65WHZxB86rgBs1MGv4Ta/6UMIS+0Dg1vQG57n74wlh9dA4HHLuqS
5DT7X1nBc/y63VM4yNc5j1w/yxc3lUbV1rtPR161eU0ifqTMk5zD08XuxC8Pd1THiOtFXZ2QrxIO
TJFxdDx4RApZDwVVgNm1YsrpC1w1OQD7FwuNj9iQjkBn84E07djRE3Ocs6Z/JOlEyJgm/rK8y2Qo
PPfYrkM458J8pF7GX5uw5RA3Dn16h8weA4CIsZsKaNVGXsQR849ThrNwJx2I7FjCcpSWLHzyoGTq
F85dtVoDrhBUvTYGEXGCYuZ6WD1qBGYJQ93qFB6ScQ22avfipW5P9AW6i1sXKKzjETjuxS9vqTx5
EWNQgysIf7x/UjDlWm1BuMGWgZS02zBxWb/027bXL2juc/RN4oUYEUPckR40vOCpB7jtwrcPvqMP
SaZx6rU3jbVfCuaCJyrqWr/eqwHeUmfh6GSKdHTNx1FzqlnA7IamDtD8w8d7sC4cmXOqIBAD4e8C
Xk/QlpmVn1GbUmr/ul3WpTy84Tqhjgphab0PCwhw5CZfJ8aAg8bL2Z4ZnGAYD1rkFdrQpEOYky9n
6CQ9RDGl+65tdcSRwUSTm4erZFyewTSL/p2/tqSzv8y/tgSPNUAJjSy26mYlYG9hhu47YBz1qTLX
9RULHdKhPs5OHxzv2WrF0ddAe7C1nP1asCkGI0NNgujZW6kzuejMsRf0LFGBcvippE17wPWb5zhH
L0JMLWPHE52lm24OToSlmoFD/SyllrFfFcNbqqZ3C+4K53UPTZ1Ue/uMmv+CDDkdL9Q7Gqaspsxk
FcE5aBAs9FVYr+BpK3W744rB7Bsx8c+yv2AXF9uC+rqXRVAzj79OUzEMYmpsLlvOP5+MRI1uTP8o
4WyZ1R8aVphWRcowcYTjveFkZSadJyGCCYAbCBWPpWnw5XBVZ4JdeGaXA94BXTr9n9zuHp52I6b6
PtcjwW9VRs+VQrxY/uz5fss4/1pmcBg51KU6mnee4tY8dKKYnDkoTg1Rh3L8NedAGag7+38fZS1H
c3OavVXIPwY56TDWNaJgI9MASWXJK1VKuFnjiw4Y00ImwBpg3UXX1/aD3TT/LutcKutbvkNXp463
3gtNANiC55q9RysSzssFF6l/TOkHSakVauO3NDfCbOrvndATLN7ShFW+il2C3TmOc9oyLDvRwkWY
UQZSLj8Eg0JreBU94dVSfZXjqDUHZjkFEL92cEyB9rOE+y9X8pJ5BPuzm1I+P6PdzWcVnR8OM6Ug
c5FgG45C8vbEymI5MKRnK+nVJgNND8MrM5nlATBqNqTvKR7lVWvgg3DlNAf6aKm5qGaWWOd8urzB
bPNqT/YrkcZzby/LbKK+sdXOD2Vit5wndhuBwn1B7kaM5AsBO+BHvM389C0OwA0KmBy6AC6aF1/T
AUGGjoPyEPRW9k12Xg7xnFN+C6f5dobFerKgEJnbVMURJp4EsOk7rTj4vWU8kgRSAhPClCdfoNss
dI3yElcr1QAi04t2Mh0wEy4dR218SMiiP+QdomsYqGwdFgvk1iZaGgq63Y6sQzBWOGbmDawOR0kw
K29Xluh3snDbfXCgAH6aIT+LzUwHTYEScGL4VyAAf02T2rYF4bLFpRUiWBfbS/gzh8TITJb+qEJp
Kx+WAzzhNvrn5TOlH+OpVMZ4NQEJzVB26Xleiyj4dFQlXE9ItUneFvb87GzUIA6fNbiX/krcGQVA
ev6YLNcaVjIG1MQtJxkJhDdayHlx3vQNA+5nnaCdEPJsWI6fU7hD9m4AxMXZV637FNDb6il2AEE/
I4Lppk6h/JWVKvanO+pJAwA5cUxrTmUIO4JyWp39yP/He0pcSuZ+h6HYlhaLQjs2noM6ae7uQRTG
Q3XlZSrPioAN6/RNH1jDQFgfdmJ6PxEkYrgO9Y2qZ47c/orR6XSTY7pRxRsaHE405t0rcKO0UDYJ
k4UrjEruYqYUopNll9jAbtbTHzZgCMESwkZl+3rfkzoe98K6AArERIig0y28rAKLFPvPcxwqexNP
yeLfwJoVM1v+rFFJjq8Njf5YFAryUNm/mTFQeNj3dzU/dQa2/9nzTrcrAHrTuUj9p2/PVuOh1pC2
sajzULG+JFaTinDLlz1BTszqKU1TXTaE1GkADK3XP2FDh+xpSgV20PQ3FEWpUm0ZZH5ta74IpCui
LztDKwrM/DuYcdm2/Pet+vRFjnneB3D3B34rz5vnt6rLtxa1Rea1/bxSI9CmAuQkZAfpa/kIVeyc
AOOQ4m7tH7SQdmkgS/St4rnZQDY3mWBXKUrTCgaRe3EIaVJ82cGaOviWoeSbdvxOabFqAz4mYi9x
rdi8O46ZsPMIb6eLfdEs+u6nv7sdEOkChjUPWwBkejNxXToW6hkTH5feMn3a7gTCPVsFf8vBcBzK
9GaZfDGQYhb4kCGJC08TyJV0ne/E6A59+8/I2Zij8ZTbe3IKHVB/rUi/c83oDFtyrQHngSl6bXfB
q90T6gII59TYFhGPFH6iQkQLR2JGUCXGyBIrNByCTtDqk6Xo1jW0GuPkoQ49hS6duFhN+axvNbkc
7ynzHVjFGrVuDAbbmEQySmMIqBIYAHzUsF43e1JnE9ynWJffQ3agcmjMlOOTIPz4LL4Dk36qOnKS
byFt6/w9LbBg1POKNUzOlw/RuLWYrpIYAZxPCZCxpoGOrxp6c2VGPLaazViqimv8ngWFfm3wQ7My
ppMBuxKRZYSP/Z1pRmyBIzqhAtYQo2Tlp9hVnEiSaDjHFlayCKVV/Op34NnZr5eJylQbfknUYKli
VeTdrwjG30UWlN31nab9MHa4aXeAJ/3K/5FwKYGaQWV2dWb48f65te/ITVeVo2UOhT8lhJtEcbYS
GMdImT3dwpzZlu52VxRRnIE0yctHdQPScjbBa/LSy6lysPm+h5o/tyETqn22th201/OMfCJCloZS
faYLdfuFnrRJUgJ0mE6jgy3/WKdFO2glKCkMWkrXVgX8U7sUynF8e6N5pXkz/Hw2vGmucoUqh6a5
TeIiYfbvTipSLJxVkE2c0WSFSSUdE6Zdg5OObxcu9IZGzdy6YMA+eJjE/3z3dII/81tk5q4/1Q3i
rtv9VdnfNu4oEYWkv6EMNcXMkwlSieXaZwfF4F5Qle+KO15eAPrH5bA1oLhA2KrKbzBPjRgVP0ze
i2TmJU1hnPOHLJ1mH8ODXKielYfjDuC0+4NbNVHnaskjOyGPdSSc4tThQ8QxAgE1ge+CYNPtuCGZ
osCc7MMwbzcu+LF7rVymSJxBC78g4AcEDzQl3o1CojIprMEc9TFPYenvWIxb1Ox5Rcu8CANekriw
V93KEgAzq8jn5ODpFyh/jmA0aypdEd4faEprVsX997qu2/EAx3x41fMXyv9R1Xf96FpPxx/sGEn4
CopzGJlqkkTrSHp1I1t+I8jmfG+g0OBOIQGRQXTA80ywGETLzvQIIPDnps3W96gMtXEUWD1rOlQA
FO3+y4JEofb/sGU3ZGBLyX5K8cg9rrUf/VtJtI6v6264FETk94RPhS1S7L64uYZSKf9u8VHeqNrM
dJKDq+3dAISISQaVPntpuTtGzysmaQULmRBrwR1jPZVH5TWsxG0Ld1DAxcLF+lzAfoP0MmGbAIlc
daAgXbCXoTHdk2xd1TbHGhNpBoFOQvoHXHsy+ZFnxVAKacxHr8zyogF11+mxi1el9VPyP7hLYVmz
90ZEE8yNd2H/orxY8kZUCi77blknnS5BgBVTMAm2KTT1qE6HGYiARTfXQoJl6FZ+GWryiJ55ovIA
Md+9CwB/WwSSrgLtCNUXKs8dbolnzkEt+ZDgwAcLUChPOCOH0pxAFkvX1imPY3PXskOTglAKjP3q
pQLPj9hMcPNOyv2zKfG6PDZVpel4ftS5+2tc2nJK4C1AhyPtA9uBNghxRgkIQ8WA9iwHhaKFTZlh
MKJYTiDb7JWO4Bcr28skseWIC9epasPSsW9Jo9ozkv5X7rmOPvQ/Y2mSiKCN/wbovB6JCoR683h+
r3ggqCsQ2X+9Smlsei1bJxRB1VjEf1MXTjXG5Jv/1Wqym117H3h2Qy4bZ0uuJnqBUhX3smv0jEku
ZzzBB3m/qPMf2vI7xMcONXSufzuSod2WiIzq8X3ZkJrIfkdR/QyDSWRlzz9hGPOvkgVmTsIgUwR1
fDbewvZEjnWRu/RLeHA30ZZ4HHdA7vzlpvDzoQrvRnH5lGwWr5mLmBwScYmDXhWEK+/rBvs6ai+2
JhhNTwuUHp0OGJqkmx8RMLkwPspvo/nJ9OE0dIwXov2wdfp5Agok1q5NnC6Da1b9sB7WMg2X/quT
OtGe80QBoKdxVnqqc5P/nE/yW7Gcf+q2kPlTAGRg3LfD5s2GCMyZmq/Gfxs+PwptBi+vXFJJA6eW
HmDrNcv9tmeEHlRS/GP3BDJfzaGMKOgfoehbE7e43w+7JJJHJLmSlDQH+XDHfToMJzW7swvgwJki
zZw+Jm1IW02dOzT9kXzn6jhJz7cyIta2A5Z5mCYL98GFELNv8lnyB3h729M+n24TFbx7fsNsUAe/
3Mn2oU+kidqdQ41v3vrFlM6qPXj74fls8QfE7yBG+DKj7lYuu58x57pIqiThbD6rA8w1YW8RsZmD
XpKpSSUXDWHguoTyQEUX2Hm1wYag5GdBN4RxcUIXB7mxh7MIrBOF8CzG4klkIxGlPiljMxNKtn8z
yVkMWiIp3QDK82iP7/ynthhG9x/dhrvXMcWp32d7xiA9KnmDdX+JEWbdDmwNneg53TsfktwEzMK0
46j8aUxmkyR6Tm6cPD688EhzuGctTRfpZkdEgSN+EsiUopqIPRYr6SDmTFfCO2auw71ZWL5Wh07t
+30MQ6dsL/XBPm9YU6vM7y8Fr8q2FKt3GzCbSwhOgU0SU7F6LxbJkZQTr0Q1sMcnTO3ZEDKFfhhQ
Hg18FkD4QyuWMijF0pHrkTMcLGVIpKnxIvXr7D0gPfYKfvMTToPiIo7ucU275ohgIWeKdDy0kRgD
kTCqMWI1ZE/soVijat8UwsHfYog16u3+eCgFGoZr7ZIg9j4A3Wie7jFse/YgJ2AHrp5S5SMHLrc3
1eOjN07S0bM+SOHCLCNhyPLCAHODHFyyya0gTkDtI5AiPkwBrs7r6QSRQWKPbqCQpb5IGfYqvNE2
ckJutfwgurqOTL84bedYl8kO0BScdMUT6t7pUoLl5YVasgBdK5CG5IK1tXHc0tj554V9+d1ev+6n
MEon8x/qyTRw6qvFY70jxOWrDSCp90owAUZ/utfUsmHb3LkgikV+Xr8TZzXGWQNWjzD8ZcSTx1Z5
zIuI265W54pbmpOA1BAjyh5nsOQQzCLK5ns/21L+8KHhThYbyQ55oj1UPMMbgW8wH5BmVh6HGOTh
mMSL2+VBdPDJ82hE6/TfLKTmutRnDhL7SNFzs+BnPPBCHiO6pseYiHk4/wY+WUyOrDvh5xM8IQYl
hdQ2h4NfOP3rrWhbpUDbu8dtqsuJmcjBb2SwhVFQIvYxc0+o+49xxiR3iyJro68IYFjQTxavP1BX
99hWTf/2QLyXhZbXLMEijVrSKNQlpWBqSL0hDTk6K1774qeKS0sqlw8jCgfPrJ7yKq8nkkmhZAIE
Thux2hCDaJPvwplCe9yg3Z1lUDRofxxL8iZILd4cYFQqSMnbNa5adDDODzwIXW0HgedRzD5rQcXI
NKjmDlnYMYoYN+oG55c8ctJcCq7skfkAD/vLKE4Dq85yawyfi9vNhoaKRaHxQQrayRbJvRDN4dtc
zFxgooD81FVB1Tb6wK5B6NnbGzRPvOKKUpMP9IATuvmf65VjVUWk3f7jdYYhW16f+naKGrxmS9vV
u/2Ws0SZluuEyB+7Tj9WMb2YW+k0hqnb6BH8sad6pt/QkINnivU9LPvyChrMYI5Fwp38UN6B5x3G
VgB1ShlgQS0/zFXEttgBFb84rcNwRA7HoEu2WK0uAdA9E3nzAuSqd89U4CVYlvmNBO0xqv829Vs9
DoPfOdqS/G7S+gvC+kp58F+RPHUNYEw1Lp4RtrUpBjlGVkaYtkart2gmbs5KomYodB/ZSHXHSSh6
qC+ANO9vykdk7aoKhdWaoZyb6tngaZEsu0zWvm4egzQZHsB5ZbPVNSxlK00mrk4vgM6lvVQlScpq
Aez5tvBTyTHCPSzzUghXNEA08VkmWAobUxnKXrM8tLWugCguwSpiq8RM4uHb9vaHODY/lUZY9gUM
KWN4vrgRRr2OzGRjf0OeRHaG/KkU4XtRdFiIaf53x2uIj+Y2j9uSBMsyTn7xxIx2WcTR5SIsRN9L
gUheGzmMRdC/QVtaf91ooSNkumy+wfvy4z77W8E/CR1cyMc5C8Xoh0NQEabop/OkqYrouurRM87s
/sm/qn7EWumWE5nbhc1IB64l4dRBSOGLWF4JH1pLQitsK4SeNlR7hOaqxzDidQ0pOxHjsNLFfwSs
ukS1/nWnf3zhaSmUi8liLOtPx8iWy9cpCx4QVMMBA7kbGiT7nC7MkuVyOEwa2x9US1dO8ZVq/wDF
te0Kko3guJWn2XgR8bdXC6hI0Kqi1eLxdChA3QmaU7HmSKT2FPiT0qCWieR+FApjmDOPcXa8Frw/
998MidLW/V4GtGQk/3mONbZ4hKnpwoRWE2J5o2IMbFo22Rfqp1tfAfadNJ+uVSWDnLnT9qA4b9C4
aU8/TN0ntcU59HCKs65nwUeaagTWi9aLwGtMXOcVXKmGh6fRYsS0K1dyG3UZUpJvCyFVc/RtiaYX
thOglLQmrkC4KzZN1zYdQd6ffVDSQZ2z9sh46Qei/nZ0c8WJm17UUrkoLKfI0AFs5W343fO1uUvz
D8maZWD6O99rCGXulNuESr0db0u178b+hasWGrftA6e0DflfXQ7BWRGshGi67MdCGPNDpp8a6TDO
gohtkaKh7XxM5ofvexkGhjTK5f/3Fee9x5V6dr2VOpCrk7o6f4CCIHkscMD1iuPV3Hg2xWT08Yo2
QbO5pK4RuO8Of5a2xCWMpi0uLt+x1Uri+q6jzjeM4xCnOt3o6zAN3z0GQUg0kFRVqjRWLMVK3TdH
0r/Qbyha+4uTzHgdnEz+LCRLwvJuhwAej4upoFaOUNObGAv/HGuYXjl/UWwszqOpNoXKKnElDnKB
ZZxtFqwYC6cZAvvyk28MNrmajJ4gaVO8/h0UedG//z4Eoir9CqOwbY7ywlAoQxEgxWb4y/bRs/WI
QAhiV4MX+RnOixUyKQXCU4heYTj9KQhypPy31UlbISW3EyuSbqhvwDLDgtYtjMKIO4SkRo3w+Y30
96rR4Rhb8z//8uprvoxhdHzKgWy5DYj7DFDO+BcLRpoSazGrzQHzlLCueflM9bsQ0dpKjcqbXM8e
ldsvn3puuUIR9qIujrfvn1pspRnCR3n1AFCVFskmwLv/3dr4O4ETXzPcmpw21lYynfGSCJfLOW4E
UgMTfJQhD1LAzxIVgF6QUwb9e2LnlEptl/bFztLHUgGV+M1YHmZdFMdPpUlLWvRj6/gCZfaB66ge
diRbddAnqoYK6/u8Y4n/amlrbYtIeBG/WUzMoHYJKgZIyBawutE3QfeQZYLUYlTxAhDjMveBiKdX
EGAA9rlF3jFCGMoGkSkPVd0UzwkeBPUXl7AI96VYjc7doJ8sM8Kn8CInl6iewwYmesJAsAa4dUx8
cUJzvBaKSWvKd192vLrn/+40CpUc5s8hCyzWSyso0G2T6GCLyshkH6B3FiZtnni7yee2VqmEOe+D
iRw9n9MSPrSIe33RSWE2XJSULJ8qC0LaqZGc/LqiklNFU7vL81yMIYsVcY3rOk9un7tX5iNu2FLD
kPGSVJrDS2skK8PMrUH4rwXP7nv8MER3E8/RLoVTzJOq/7as62oy4vR9k4XG6IvirpU26r1jr1Ir
ZnK5PnZWMI1YJeff0861nWb42j7aNmg5f5Df4Yq7npvOoQB+0ASbBqVW0DZLctTChtvI23rWVY/0
m/N6VzW5yP4QrACuHxpLZHddK5yoAFumL8bHdsfhqk8riKnmacrhWWpmX2FtPIiNL9cCF/1FwshP
Q7qaYPE7uSa89uDL5t3YR2elrSjWanJ2jinm4KXr9mW5o98Hpq6jjepxDWuHzeIl+Pmhru3ckku6
VmK9jJhd8r3Ytah9gXRwjgQgvHdA8EDFG4SLopO8lqCufCQ1fnCqCZuyg2VbiehvogO4+4MDITae
kzzk+JJ17qZyFQi+6Gwohse+7lJK1dIDWLpD7PVHpQjleneMTyDLwc32vHRCL4by0vzVnDjm8O0R
9iBVSmQ2eUuJOAP1LnQpU+7UVe2w5Nt8dIAHzMwg3EscjSSrPq2Ek/op4vE0Y1RuHbsQ7d8TTvgx
Ru2TAk6lWDgfRklhjP32u45cn4zohSp4zexlECAUtOxUqQ9lkeM+dNv9X6xtLPZFvFLOdAr1ri3f
Cmr0KSs50xc0I1gTMy48StOOUvQgMflH7tVXwWr0V04YhiCDG/R9AP+zzZLDXYMvOEHRWk8YEBeP
G3XfivFxJw2tJys2p+ITwrYGUgKITLe4fRKqGU9m+ff2w9XiCkdzS1kGulXRw0SFDZ+Q1/k9yzZ2
CikKcm/yY3R0DUDODw7UDGuTehHQihfc7zy0U9YCkJ0dXuTXuUQ2eT68xu+FjiTFWCyXH1K+PUJI
46gAv+EtXK39WbDo3E052Tfu4bXtYU+gi2pSzEnyVFu0QS+uO+zMVzzf2bA4ZG2J55Hkt6GV96qK
ClVsvhIEodyo4p4IjgbTDHStk6lkbOK4miP2x+xLx1PDTpLsgWy+exY5TnWkRedQhzv3ldczbIaI
UofECIxKlKRlEHX+X5N4DrxwggM28VxtFUpzfRXzXyAJBFrYIoiMrISfFMsAFlsv/SmVfjyj92DD
jH5i+1ww9N7bKLshCEN9fxJbEKJyLrqkrvCAo3TYuYc1h5QXw4JJVZtXvTrB0FVOz0hozdiei8Ub
/49Gjvb+G7GrawJnvhUvnsqylVUuMUxKPjPsoRiS7/TlsYlHdt8PqhYCtoAF05+/c/DlP0DG19sh
PeHf9p/iwMgP2w1bgS98dOMSGyoMU6p9SbN5JHLa2yFeQws3FAo1Y54CekCbHlk2+22FI8hm1F/A
8f1VrwKp6aswsxFzC7pvFpZ4YqdGCPvYtnZa/zCOYOgKCtGyVc3QUKlFWtn/tgNG7kI1dwT6obIq
rbrmyYT7XYYUGJG6flb8Dlw2HDnm+dp40bttu8tBZOXFPnFifrxxYH7RJKiMkKVtxpDrDOjVNmRa
DeurHC+rHhbNFJnhDKFu+/IrwmvgaAWNFSsercUI2y0C41YZW1fnDt8gw2ZqND1qwc23pMXcAo3Y
YqZa/uDptD0NCtxbGQQ0gMPehmq9/468c54A1cmpA5kMUWCoiHLfnhqsRB/mzftNdeN+RAnWDx3j
89NQyzPa6+zIufEhBNNA0sniNNMKwkkYbBVdkjBEMLY685y88YoSlAhoj2MZ7FxXkKpC3v2hNibJ
AMkK94Vx6eK6do4wWSBdO803nuQlGIWli5BOQZxBNPLC+G9TYSl1zbCk8eavQWc3GKsbm5bHticp
dwGNCg8+UjxMJV4g7d96bgAWv/Ncr1/HtOsq4obYY5yNG8jJA804cfxzBpf8v7f7Hzls40dcpeZc
VJs39SSltm/YgJG0qpxwP/6fWpGhEhArbuAFUFmhcLsBk+Bb5YTtBrIxRQsCQam2RRmbyo1wyLuy
+El9e5XjSOIj3etBJfUjW/O5DwNGTDDlQJCKjZ7OhIZGdHxLn7u4sp2x1WoSr4T/EPy+0SZIYlV2
kOEjxUHt2QN8jSMLREz+0r2ArVNhHFvfiCRZU8TtMYkRXdQcp/tVLd/VOznu5azYmgoHof1HRzzt
oq6fHNoBgzLyj28xqo+qCdsA+kzGj2Im8ZolpnJpsT+qvbksU2lLOLlY4nPnYAtGR41zzpugQasR
wXls+wzOw8cSglMBKghTccsYl3pREx567c4X2T0wtFYi/x9TdG9FqitenNUCoOiTE8Sf61oio4hu
AQ7SbVxFP10WUyJx6j3KYWPu13mi/a0EhvLE0lmnLjuSf91gzNd3JyXM3PBerc6sAauOG8F/oqmq
1mY2x8TIdjjQKGIwQWdRz8sNxW4NT6mKxFmLDab9nhk3xbzE/x4wmRT5g1jGiNjvwPhn4vGZT07+
rziJgfIm02TUxe4W1sIKahGQjT4yZfw0/3smVFCY3IKl6Oo6ayEYNgla51HHQWHk01zkL9/iVB33
Vs49X3As8A3l08GKGLQ3gxqqVG9rZUNG8Q3/1ycLy4g0jXWEwVsSKeTBZRxF0ieLstv8szDIRkzb
UH12MkNSv6q8SbfrM7RYNKGTelEqIbAQvSWnoGTKtMdQGOJi9bSZybFSCzxG/qAeMvMpyDL+jjS1
m/RTjv0UjDLnNn7XDS4AlGKuWbfKSNRu4pXM5EI8WuY5qqTEdFYIudnccoVN7Fbkz1rNSs6gwHDQ
pKDB/lGYZVgqL08A9uCzOW/2OELJnJAIXgQs3D/QKx4t5Lqv6C7Smxs9UPeaxooe9ej50+XV2cu5
FdaE76xUPddySbUWOBkcAd1L7sqwsGMAK+iHWVGPjXJHbgQr7j/1zsI6gPdvBPcr9Khrs0pgcodA
hj0F4J325R8Tk5fFe8PBFnaelJRWa3sFF3TKgB7b6kekqMIROVI8N2CmsBZ39LMNQHsfhkzRJUl+
iia8738Dw3TA+rijjAMVemoHY+eATdKTlrxjW3dKUoCWH9bZr6ANnlCo/v0Rk0WvVcnShqf5/NUI
9AzfoeeFK+j8C2DiNQEtzNFakLbfWEoAB1vC4hBF6K7csZ8qDWMYUP+KAmvT33fBCqCRbo6G8hfA
EEztfi5YIPQkaHAmXm+bJhZtO0B++AxYZSwsq/+56C6gOX5J7zfMizH4+PgH/T7wzo3DkFP9eG/X
Wh3L6PTZohAiGoxV0hL+tEF2hHe/go9iVFs3CkbXap4V9/pJur/11sAxD+YIFoUjpzEQpVJrdSwJ
oerMYSTZ4r23r4Kh94KHg1iJP+eai5VMPzYCH5ZVW9+7334hzsdi0Hb5NzWcdhscMANO0IIB+YIT
i4QsTx7wl5HP7J06E/ClXkfAiAXFSUnHcjqtF4+zropLijZbCgTllUNzWJh4Iwul7BegGVbmfqfY
BkVFrTdAm6i0PM6rgxIVSRbOAGcXeGnjPmPU8dt7LPuu7Cs/6AHAcJzZoK1ZnfMM9LbzNm7uZnis
uoLIjjITAzqj/8i9Wu9HYvM16s0GlTbwaiMQpHdWLfYutmfbXB3Ka2fBbfwRXUCsGRY6iKA7Xo3e
mjWnDcuNFMSMDsdnZ5w4nn2I+b6FOs4beI0/bcVDaFmsozvXmcsPFk+xBsWEW1pV1ZwZhr5aHJN5
zFqoGaqBTCTLvi2PO3oEuEdAK8PpYtLqwM4VNsbpQWJejCoh7rTLMp+WQpLdeOEAFds05CUuxnUj
DWOOjjy3eX56q4EEcwI1acWw4me0e4WQWkqzwnvqFWqUI7Z1AyhsjlhOXJ1JHVxA23uVCym+J7ut
BCs/0KHxLk+b2j2YurCg3YQIHQpRk3+WuBb3lLU2FSPuTjxlxaSiux3oGZUE8qpshBlWF2czLHOl
WC/LwNJ2JFUf/L//b3ZZSwxaluBQy3pWCuCNcxI/6YB2qym0d/+GVaUN6lEpGaJLgO1XbGTsnaF/
pWxwnDKtB9gWF4A7jjrmjPtfyB2Z1HrTuWKhzh+ECg8RxmY2PjdgqW97mx8SGd/P4oAEUt/lyG3n
VsajqYxD//+reh3viperJGIpGYF6J+KVlOcql1tbAmTv73GkTh8xskEKc2Jyn8irmGUK5zpq3bee
DtBGzIivsOrTZgTEy/GmbDBGoprsN8gs9A4EA9bVvjrPCuI2fxntPDbI9WzmGnSSro//sHkGy7sk
v6BeL/sAur9b1st9Te53tR1vkR6YLjuAfShkfr9NBcyz12fX6Wv2PfGn3jcp3jnGHKqsKlYgW2U7
xl9zAFVt/uFfzHdV59de9rFOEFG0h66lvcyOXsJyd5k3Zy0I2lQKjVl/5yoOGfDl14wKPhx8DYgI
l4lchQ+VxkYKFGC3D/3JNbHrU2LDPB/eSRBs8Hvt/JmfreEwpNdgQ4lv66DT696hc53bOjRIRRx9
7bKDnn+ny0xp8WDcRi4TNAHKa+8ho6aB9SjlBm9D3T4n6ujWVuROEDrNeQp2llNKTcTLb2bWqnJc
UYMxFVv/YNG/KBYIUaghR09HNMP6URvkWEIRS/KuUMaVMGId/osNDwjgRCQsJkTvaPtzNXcX6tIw
+1nWo4KXY0Zb+m4AdV5Xdacz3KGRiNBpEKyD046Jnv6eMap/hUmh8y3Yss8ErMmdlhFCuo6oQUp7
of2+pW/G7q77+yl3wfeaL9Zbhb2EOUvai4FEatrix7mVRsMnSL4TFKbB5pmezUoAxcsYet4iiCzV
nofChC+r1tAlAnjb2gZO2jYheKlyIs5Ml5igz10gpnRHCYi5AT1tjHBElnFkGMZColvSh59RI3Oz
G/aUHsd7vBpE/Pqutt0xk6/6KmjKpVwCrRKlS/rz+7+cGQpVqvF9N3eTs/nSijOR/tjU2dQnvUAm
hRoRLt3rSsPF/qSOaeM6kqP12e2GppGQWYiOUcD9/OxZ/rHNadnKL0ExLWIvdZFnny3MSRjQGBGS
F9aD77kK/FtlfjGep/RBLC0etEsG9+mMftfE4jGbrW5OmM0AGGFjo0QfLF7L6tLYTpvdMeUdL2AE
/EruVb+BttqyvC6/XwZPwF3HIG32SsrPglgZY/bBujVq4fYlTPuIkIjC7LyGKn/MBiYCUrgz0hN5
8UKig/korT94VzLpZxU9jGeqP+VwGO+d1lP2MRV7j7VEome048ROeWUTH+kvzt0WX6sEKEpQVehC
atgA+DsVttT9WPdw8miTRh4Q8LSRV00FG2gf6pxfpkWiZvor8cuauabzBckbAeJRNBGeqi78ctjV
60QYjkn3nwIg58VNxpezWl5MSOcRtbAQ8tXQU6WvIdjXk8/yyvOYy2ZmWw2M48ThybK0A164iMxX
b9tKqK8LDBQlbOQIxtzivMIRhabGqKHA3FtsaT52xQq8/BA2sVKrseqM3fw7BqFLHTrWerLS60c6
K+EUHrNXBsDmblZzJNjS/c+mE2pOibGPw1MleX4QnXl+Xk9/ByeSzNPaGWEfSGR/fe7dgGY0O4Xs
xflc9/4xMQlyBPLm86LAbIyWjgrbGkAsFgNAnzPMsbjNIGHT+a4NMeG1wAJN+06RHPMazwV0nwQ9
uCQE+ecNBmlp30JyGvXunBMJcxICtjm/e7icZW5OFEISvIcwmC+szkg2t9sO81uFkskMoYR95+0P
Kv6saduf19Z9jXsJUl6p4otRBl+JuJP1XIPWf1KzSPRD0i0dm3ZOYLpqjQxkBVjnueaBeLEMk6aJ
gm03YLEOhFUpoJtDmJ2rHfb/Wng01F9ZntTkyEF3j4Kkf690iPRjsVilZ8pODr49YPxDWokn/qkV
bfD4yZ01t4uQpeu6MVtjNkpO00jIgryqgv1g9qx1Z8LezRZjCI7u11lrEYwy99dxaCuB3YnWo/Tl
zLFwsTPyV7RnilcVPWbs4Yny+BroZCQygjb7eJVQYhXzpDmFozpCj1XcNI8ZfGKjejEGVdB3EPbO
wJx2nNhB8FFEeRLt5WbXAVjm0ZoQAU1MaJjPCJlssgTRT13xN7uMMG1omcIKFv9EoqxZH1GhS/xL
iWjlPo/z8y47lOYTdZTk/84+VXz4XvzJmSc268cyxjvTxySLV+jUVRsI1NYKWnN5e2HP4vS+u+02
S+soOAM9qF0DThFZ1Lmsk+N3ENVtPeBJQnZYPFxTtHvJwtvzmnWrbiGMVUUQ4rth01o+6o2YcoVG
n+wiVmxoPliktSo3NPMiuKG2kcqjHQhPv1mSe2G9F+Ji2NwTtKHhtcAI8bAtgQ5kfZJ7z4POLS1w
XLNu2UxavYE2tR/ERF1U8Z09AJcV9U+Fi5X8fOfsq0tdSDCljJLJBsxWVKAmV6HSv/hB8dauMxgB
MVy1Xf4IzOJwPd4Gpfi2YPDjMwQFMa44dp9bo4meDjaDpK8RzJIe8UYNmPHbKRn/eBfBBgLNY34t
vkbQrnEKouKNHXZmLI5rdRmeggKI6NQuep5+Eq9+IkdDOHqS9SW5rvFXE2l/iHJnlkCUyupELz7f
tLftCBMOnMyxpxDpT/LC3Jl8WO0ECXl+Eqq41WlSawV75o7cXt5pC5n4cu6ptxR4zEtbgyS5YJeM
ws8LulU/BCKN9W0+WeQoxk51eE3YhwabMe4oyYTyAybkuNeXcxWXoGTw5cVRaG7DyB6EhvBTR4CX
XGm1UV2L1llz/1kCwfWYY9j4EwJ2jMetUpKNdUweL3begsgqvbGdQ9c/VKy7JXhjX/fernHuMlJ+
o+Xb7BpVTYU/EmSfdIMdMlS8atpqDodCU5oq7itNNe9lFnXmdxIdygLXuV13UBueNlLodU7Ow5nI
UwvyX7CEaNWwBXquY5Y+lu6a2PISsamP8h+ELbNhyxwNfRhMid54Xy4Xn8dbruC4bWws5NFg6Lno
ZvpyExgTHhnTkWcP3rPZKJTtaOHTn/SxCnQ9E+mZPcONOrTrpjNJws3Bj0Wv3j6mUuWd1rk9tcCF
Q9eSC5DTh5qRmucz4EdHkg/n5nXoFJPppAAZy/KW7Dh8dA2gOvYZrsFtvFc5ICSi1LK9fvIB89e4
QggD1gP7ZRw/oktFqb7p0gFDDXdAxofgdYWMhwk15rr9Qo1n6+Fy0TcjKQCnHEY8LA62Kjs4Bp3F
bwH+kBlDdHmetL+D7rHy4DOBsFnHfaDFCzZMEQHofVmOQdACAaiL/7yqCB+zL5c31vv3daIOt63H
/6BMssj1TGekip8q2CKBikfrpgXXmSKulLXBxFKm0ql2FwUAUE7156ENnuB0xSVWmeabdXJ9MYI9
cWX8eC6FHso6F99vTqdX/IDU2SuxawapiJk5twNfxZtX8GmRWG7u5d981QxSbH97sdD+O6aUXV6h
JMYUlzDUA2FZOgDuuCUQxOYWHrW7sxS2TstY94mL8AoWuoW2VzdFBjgoE7ubNlQCfGz+ctmQqm+l
7wuwM/MZldJiZNPdfb46Itpe1kpDyC3L3aIb6nYHYaAU6ND1zel6EcsxVzLCwSU2NRHhRN9wAvXk
VORZh7ttIXsLOWXZALrVj6/M1d4kfV6MGiW5aa3J6gwkt9qAacIDordlEksCG5PIzEasIESmSRLJ
Fuab3935BRC4y54QdkN8fRg80jXH/Y/UsKrGQl97FdQQFh2iwzuBA+RS5It2lUOHPP0VYFrTwf4W
P+TnuYgoaXImna4B1oh8L9Cv5PymGjxh7H0vaq9+k1vfOR3ITZaV8q5/PySIwFMZgGi7BcEDLXDy
S8ZRU9Pmq8p4aUcfyypawKQCGdoOIiGIezxqMJnxdmQ0UWyySjZo52Ts2JEeAXo2wANHcq7tFmUr
Mt19zh8sz21PmQS9NSFRkhoRdEQRAoFBspyVhs1j1ivmzmd1oO+Nm0Wy9bHa7Ylx688fjralUtls
UqjiPwxxRxFqi/cIKzMiRzkSUJhYzRcIBmrFcmHPqCfomfBuApBMEr8dHBKpPLU8JXI+wDM0T0xT
YM6pw703cavQEyFouM8i1GLtShbnbqx2jR4iojBhJL+4oU+ZpP/48HwT4zFh9EBsoQ1qQJ/3e31a
mhB0oERzxm5oeBvkG89OgpJWd3k3IjtC+3kdXeGREt7IFZReiBWt00SiEyY/MD7z0q3WMFRvEuGt
YdIRUinWxXRov2332sVVhOQan1SjWOF1FnDUeRiDc5XT0zzEu+2GarSROkZTcA02kgFZYIylJyNE
9zUbZ7y3UpUnBVjK/Gx83FkZM7YkVJC+a9H/MzFDYQ1oY5sZh+7D7HddEMLYvoaAw+vlwbrU7b65
FumRsXgzaUnS7bBjVKPstA0v50nEAmeGkz0LgJoxXSCcjnRyua2qY5CI4qRVmi9bG/PENriYpSHO
SPEzRub1yq8ilHlEfz4dKwcKngsznKBZ9egKuqymWIgqTdM9hMujaSFPkcADBpYuVnINf5gZy5uG
b7XV1XJrbkB++P6NdryBLT1FLN2MPfkDBtfE3oPzCEDiamRC1Y7Oot/1/yVlkeWBB0HAfNJGSASk
IS3d01VMpXZj67mG5ZQhSrKQ1enhj18y1ZmOQdI0cMvcE8BJruOLA4IALS9yly2BW5I6Rintq6wJ
QOstEz2qZBpuJrBSju6WLjyyTtMmMGoOKMy2d+BI7PHA9xCFZeTwiYFCIN85aR2pQqGHF8ir1rBH
zmYanqa2t/C3Db3JP4uKQovTyj0Z/DXtvpj43d3ktd4hzeUpoRza9/jfj9kzD+XlDlMZ40n4qiIg
9kMK2p00RmF5NyspgjUARw+9MsRCEYdNsWhxbpufcigPdqkyjm1RtpIk8H1Ta5NXD2mXHHz61RVe
33ZKZxQ8iXkiVZpYu7DtDu7psLfg7LVXrirQbbcvvhymlfcSheBywG6qKo8ay/IG7O67eaOcnGCR
XSHeZ8+/c9QJ5HSRBwADUTTeYO2jNBG3GJHSabOfXkchpgM+O87DTRxt3+/ezdaacJKHKczMgcn4
v+/0w+sL6VigFCLsz6DyD0WtGiuf/wMMLmrS8CaJmnwwm1Dl7GQ+cclo39MAAPvDfiPdQCXLn+xF
sAUKPNVjHTBspippNjTGK83P2Y/EnYto0rCxbjodyZJbycekPRJqEYdjq06XWaUp2NBONyRXZZVR
d0JCXeiyNtH1RSCToq3UiFex4eRPE2XXX8X5+dr2WnZYXvHSlMYYOuCStofk3oHaHnvib921Aca4
gQotOk+kFrqWlxFaqZ3qwuc3QuvQn5Tu8JwoGUTmZJXd0Ck+x8g5RTRbG1hJbf/QuJeVnob/EddU
qdUir8d4O9tx3fPtXYdfrlN6y8NyU9A7QeUC0aHmmQolq80jJ+TuA3iSHRcULtOxltw0XTXso5vb
hgo/ziy1RDpsJJ6iGcfFcUn0FALFdLvvk+4CxMvkFNwZkR3f567ooPihxYvpC4TQY4WGfBoWIPEd
sQpAEYsVnwvUBHaKr2cV9h93ChgsQ8HejfmI0XcqyeR/Sf8kTXNk7EfdzIQD55GU0iWpL5fIsOBu
UzmrxDJHNBj1MjlUTf/0PstGHslo66dGCLc/s7/wDdEj8m7PZs1XCSGBgLNpA5FpyVhovJ2SlEhN
xn+qoqg3Z+gkptak8jHhpNkTZThe19DWh5zWzbEsYudURwvd/IB/IAedceEyyZb2gs90HJPBsGxg
FgZk1vqaje4voxGj/FbGOzSh1TrtP0gGZfaSTIsWFjQFHuZr5yUy1caA0uU03HozRIoH4Zc+bWCg
UiNcfyoFSs/ftp7JFGxIKkYKsrrp4YkeJCO+sfKYAogCAJGt4jOT/dAJh71Vikdt5I/L4KsjjzcQ
fo2W7nt4w7mAPGRFM/o8nR7QRSHhizOxAGxETkGVXFdC+amM+XjFImsm/iT8lLdjqvDFoocDgDXT
sNUkDohWwsJvHWbDgoXklNR5AXmENpWdSzqpkX1fJk2rZEb0PyMf0bB+JFrVRrTiIm7bPeRxCp2p
Z/YuzJ47BLWz/c6db01j1Ai5MTAs9l1u7Rs9Sk5ONUkqyqr5FynOCUEPXdR8KgWwfB2qTEq/WqaA
MkFDwmygsBC/kZj6FwuHhsctZVf/T0QfBo5o+x/bUPY3kztJ5BzdfPvs6M8scFwhnHUOuYAmadsc
XvK1sXLxT382EG0UeN9hcu6wGpXzTSTQGdT1aDIAU90ywwCY5bqpidp2T3FusvKUN5fbZDH7kSsA
+HViWZtAD5T2lHmRyfILthVkGDh77w8sCn1viiY4cuEyiFSXIaxDnqDUm5V/2ExT/NVA/gBS9A+E
eRd3Vme3lV2mEuO5csi8NaE491gwl6T5WVfYA3NQoCIe099SCIrAHW+uL88wDnvmEMiaDO9hC/Wf
p6e8NZHMkYiNj/qgI1A8ZGUGg1P1rzueAdAxlFq1SzmNNhConFcxvl8JFwV/SC59EzuYBEihvxqs
FK8tZM9Rg8y6MFrppnhmOawfZIpSwG7JqURh/qBqv+XOlhlO/3zdDM73CzrDHjZEfyOQScwokzS6
fw8Q/iVxtLLQlVZDxQOtUtRpLZCjrTmfmgUPRnLNECm6O7uHbzfgKc7MKwK6SGaJL/tHDgHHkAZ8
sKdhxvCl/DHWicp4F2nW0R0y7ICWeIRU/un48sauiY8sXqiwtVE0rtmJ5EE4vwEixmSCJ3eQb2Zs
uFu+VSDnqsVI9hgF4nwggawPwBtEY8XhT1idi+jlxeul9hROqbZsRq5FXS4dcLd8loiWJwvpkfty
iI3ChLGUTm0PM83IT5ODBfLnzIqvFRRDjQd4Sd21+I1XW1Tq2IOKWu/aiTq5Rl82Yr5wKtmZAR2g
ydMcYBcU3CnXcxMZytbX/9zCuTOuWJNp4h4gXQXCp2L8SfzJMq1oApoQ+iTzDvEoyQDg9XgzUYHd
sF/iG7ge+J81tOg2tk/OVnu1Sd3FHxHU2ynaarQYzVKIcX1fWXI6hUkl0Z9Dzb3JMKYNOEstgOHP
J7wGJZ0TaHozEB0VUbj5vaJaAmJwZuvimtTfEHFaqcy4s28HZGXpBBoRQGiL6rMd61pQisgkta6y
w6B2j2djj5AKaiSQNu6gW1oe86Pdemkl/xJhiYYqGCq91Y3b3V0jJMdS3MIyQmYlzxv168SjmyGC
wQ/ZtMbrWUTzpwmu3a56tMDrtmOSnolmybmMKxrlEFKwZE12RPn1hiHlgdOfIlMXnp+9H++eyLU+
p147HW7B2aTf/XrtUiir+dOKFbMju3Jb2RsfYoS2P1fWsP/HrhFu2yXTXseObkW4CwsPKUJw6iwA
ZDgEJ/t952UyCXMUUmBIkXLUD1sqSZJJAE5agUPSUalH+0EE/IMES+SXVt4zgrovtW0tLtSqSwTq
53l1+DThdElUKZEuKhr5YOXrBuSpWXVnvi1mJ+TGljff8wCY7RKe67h066MdkxE94H664G/pEG2M
nF3P1gdJR8+wRIPL0500Yadk1nl4kwyoRNbDv0FzytTkAxAnxLEjLKM0jTHGjAlqwn5niN1rAQ7f
etJ22fgr0VJv59UQ25qiEizH7oKIRi4d012rFP6k2YdGFZTIuqu/1KLjX9snYZyF0hKVkLnpTuAj
xX1ZtatEWsKgm58SIhiDXIbRRYTulqZiHn6bwJl2xh261bKU3XYOI6bO3+atYS7MGYz/wj/+J1A2
Esb4sYgd8B4MASUpGfYyIjKu4GHCbfqI8fTG939kLO/3j7Y/VGDNyid9wuDIZhWGFSni1rk4hNFY
eWMihbikXo0H95mvpcaWaCK4M+aAY8h/6Sn190Z79mHNHKhfrTk/MzRDjCrKx1fL01jLcz2/sIWd
7n3vTIUu3sNj0ZIeZPTjl3AMgaUN05q9TzQhZegoc/eOEyUk+J+RqwMeX5YtWR9iPH28RQpkYdPH
2l1fwW9TpVA1qhREetHwKGMEAFsdLxGrx2w4VBEm0MjRkaiG8R+YOlY8aIAHVBV+5gv3BW5dcnkJ
jBCU/eysF0kXcamFLXjY+dpXMJBBnXTMZZlurDrCOrqISHLLboAS3mLBu5E+2D5TqfTRbEgFNkV9
Xfz/FBnoUktZc5R3Kbf4WU5DDu4K3jaRKFvbdz81VcuWsDQQgRDO0SdErqLWBD/SKfIzd2bkWDF6
Mabk+FYe5R4kTwUPXfAn4SGOEt1AEu8bZy0YbjoOaOr4vPeZo4wmU6hxV1x05qbP+qqOj7tPswU5
AchexVowcy4mtDWPRv8UsUe1sVIRm3eKISJHY3VRpBGAgBnyzJTZ/q27WKZxjxWNK8Kc0HOB9Hh8
HLxCoOYTIQMLgZN2q8tgdd+IsgDVGQXB0OoVucE9vOtGGUZpwhRK/VLkcTK0F87VvToKeaZV4Bj8
tyiReMCkuSAZSUCLE0YS7a6sEhA3fYWRYJ3NXpjAa31Pp6oU9lY06hVtimwQz3a7WPy46gK6htV8
WK6UIBlJmQxgoE+qGZVLdYXfmC93dvN3WXc8d3ByIth9zo5+znSBokAr3wzc7+x6OoxB3Asg3P4U
OBC5kiP5iNwXvtkUi3g2iG6aRONfXcYeMo+4WlWLIm5dBOn44R7B+Dle9yYgF0b9Djblcv1kpTbB
qkeJQ3cIgZHtbiOJ5AP6dBC4qFAqycqxlfobd3muwGFf62/HMIPQLgeRNcn7SUhavad2nHFmVGNK
LvtNDH9hqgoblWfxu8PU418LJMGmtKr4vwludXoSGW8gk6xmdvRyA9ENzTFhldEi6u9oSWdmMOaj
FuvBzPwSvQLTlQ+rKzPttWGJN3D/Jc52owF7O97NzTDzHEtLSipQAPNYxfOndP0gWxr1xdtaYySt
XZzpfsBzQ2VJuF8fT3VQndGMS4S2FfdYzeG9GPCIeYtWeA+/WpOh7VRtX4UllW855EiW/AjHDMIS
S1V7nToWSf0B8w/t/EpkdsbeTjHeDiAryTwxCuC+/UVYzUa9AMC3AcsYX4R0OxebODH9QcRRAMxd
ELwH1FE2byd5WSFfdtEZwjcTYS9lCckzbUczqGozguW36YJvSufBLv94NOzs2dSOo5CprLncA73L
nGhnFXPbEl5y+1OyhAySeS8pwJRX1MRNqJ2RC7tLPUw+nx0QbnNAZdzaN+jXYXFVfPnT1ArqYKwQ
lTKz68TtgIqazssAK8MSyOyRYkbhx3YuJc8r7BnQ4VGQCQ434W5X866tfJ7qn9aYH8BBJ3Rwl8lp
fZHjd94A0tUS7R5GSqJdyGnorcTGGlIam5KyhNxQOEOo/+5OC5iaJC2et83J/V1/BfhD0Ej1MDNN
hzYdFE59aLXgZls0u6W8SvLYHWE59ns6T5ht9A3AhhsXZiw+CPcvLTr1lE3aI1Ql5btzHRl8GQ1p
R1ILXh+Lb/44YW8YUJtNI4T9UgZlRemnbpMxTxVXbQUrcsM63RBYpDZa7S+ggKX2MF4qe8W3ObX1
crosXoTdCybrlOttKTxtv/CwxbrV9ADML8m9LVPWZL/NvsMbOlwCoF4XLSD9nqMrywK1VBwgcBlZ
kq5dzM89tDVtrJi28iI6sw25k6avIELRNonr4SHuS0FmCKhkMNTzHabMd5FZ/yCvLFyw0NHfbOH4
6Xc0aee7Utui9OMDMJ0g++tIH3SCigWEqsdsHLP40kzBnTgWGXicriBSnD33rr1b/+gltvaI9kZ0
5llTy1pY7jVSlW+b1BT/E0Jc0GL3xAgHcs6QJLja/7drEkJCxj/+Nv/O3eASmeb4KxHCBjS6Iw7+
0O1BJYUzXH8Mu+WtofS3diO1th5lCKSPI7NtgHWYvhCOQ6+YZoOcQV3gtcodjmatvhavH/qTRNNL
H30JctgY1ztFputjgIcpr8DpEWYOjFfg2dG8RRomZcTBAR9tmtT82igHRZZoYim3CAMw3OkiSX5U
rwkeL8tLzLElLLGtLN9oR3h68wpui2T98rmgD82qlXND5Tb5As9LBxMaXRQQ5NJ2IO2bkpLu/SZ0
er+f0nob7ZjZhl/H5+34z2Pr8FI4BUPrsos7oyCL353JQ5fxRVEmMqM6dYvXJ5TwAPMWpdUeg2yF
S/n1qedqlwRLJJ/8MoRSc76qagU0m0El2Y9Z+W3B+8CzMn0RrVES9ZSpUv/Wb5gKIBrhgaEqCg0q
4U7hvuSY011gpk0oOYKVkUv/FROP11TctvItiQYfFXftpnQvd7gRlR4yC4WuQ6xib/fUekR83W1C
OONgB7/kjnmXzekXhmKO+C2VcMqJVFx8L53EbwRUzN+9zdnnux1l0O0VLiDR+fylg+q65hQoUcCi
rlz4Fc/XiHqWkcr4BU25Tx7cUgZ8n3vyj6w3F9cZFdSa4w5PguucGYgMWejIoagEqmRG67YVs2m8
KRw+F+MfbVFRDLhtcGoERoqsr6ovfD2UzxMhQcMphYXoMB/1KDAukmUMKTIsr68p3N510jfJvAjl
ILHpUfH4VqDyLmjuKt6125MsTHwseDWFNOC3K05IAjaRRBBD7d0HcKTmHz9qPxCmR1ayS76mbHj0
oCcQMhG63azmpxhLC4NHRU35y6I4wsbwRsowTPS1ywu1MLNQAg2EupMgTk24j65FvLMvraDzIxIv
ZearhG3jd5iL3sb0i5ifdJtiA4XCEMNC9N26kk6wxOIUjDW8cXcIzU0/0WT85TzdGBgHNgqBrhfx
DrjQY3jXqYD+jn3FkfF894PQyLZD4iPF753Th6YfAKNHe2uDITF7Rv7EcL2g56iJfg7/159NNyF8
Z1yTgiH7mCC5VdjpG11gSQTNk6vqmKufDmGQeyqLgdv5Op8mg3LZunmfv5BNPSO0VagqtJb1w7KY
BhYJIqI+ihuhPosQm1l8fz6oL8CyhHCqIwAhCwkApiiSAvuSFBoLJX8dkgTHdBcs6tP4JYYSWqIQ
r7lsbCYqR6sLCSK/oOWs611pWYK1xYQPV3UmNrpMi/kEyshtn0VsPpnJFndnm5KVCfcl/8ir0fq+
g2DeAgswRImbOwvRQ4Uz2omlUSDxslwC6K48rHYi3NMX3JhjOXUxigz8i3m7BfqeUYk6tuXsj/G0
Rbn1P8N+0GsKwdNpVSLGAP7LSYcS5dbd9UC5dnL7U1sjffyGJvW/z3JK+Ck3k5Ns4LIHt20w3tw8
zEb/PipxBoTKFkGQX+QnOTJOWZE9bU7/uWSJ/VDKDyuwuzzvZ2KhKr+V0CuqIvKmEgCd0Ix+bGy3
VOSiUotLFuKtSxPtGbPIDPIMxQEiZPxt8tmBfR8eEMLIX2Dd2gil1HN1PXgFNOgyjcy/lQqX1bW3
ntZKghDulna+Ly+h7+Q8kKsXtQLPjYIVoVyDL2FjMuGl9847PEEOWB+qlJUVUlTELMNKPaaJRE38
c5hOmNgeST+4P/exdMbP70YM8ekYkWbnguVU0GrMxCoEhUj8Ibx8HfehPEzKuEhggI8f0BkFruuL
pKUp+4X2I2bWMnw15FKQ+VKeP/zFnU4m9oGRSHf5yNcnbwG0aeGZjxfYXdtg70MlWAJa899K1k8l
NIcK1IPdPtdobdbV5bBE24CR2A9Q0UNacX1smiSv4+c3ss07snRLVHDqKSJ/HnkDhv1sx7la1Jov
b0RhheL3wZQexsq2xXxEpYmBXCV2pkTQmeoOFoOBodM0yF8YZpjA3bfxBsdA3p3DBLIhj+rl/WH+
Wqlhx7ZeTZRP15H5NapSB26v1aSqZaUQD3wgAQWNfynuPo+lHKAxb5t+ivaZ6pycxydi4TNPqzb3
3CliLsGXoRqlbFd/nKnodvi88TZXTFoMmo4kM6m0bMrMAZZ8CUyzhypixjRm6ZvYea0qNulzSBWe
bkbTdKcds+6VJWUT8X6SS4xJGGUPBbqH2BeQeZQHAolq/hQsHv0LDKqttIvaNkeRlNreFDdZKlHN
JNs+mjDXLRxcsGf8o0n7XJObI22WT3NVi8BpVBDQ070dJ0ph9Ix4yKN7y5iGnUjxbFlLrhkZck6x
S6fMq1q7W3i+p+MFaTOKtLePZnL4pfLnxu/LMdQkP146y6I1ofsePip4mQ5ybIz7Axti+/z0CFcR
wEiJjtU+Ayh+3mu3FqdjrmmklM0MTYHvbZZXcjrzIZLDoUpVn7g7e9N0ow2Uh9DfHh/82unDVeoU
Vxw4Quy2uL62B33/6RbLIIQX/ZDbATPub5SWZEY2mpZwgHnZPzn3EoMDSokZoc6QlhALmlk4rjt5
LYOCo/NppYIrI+11ZtlJG7wQI4JlckmRumPwrYpcIwtdqfkwp6IHC8gnLEdEK1Lzuip281HaRxCF
V32dNMi18LJa4LdGm9nbxVi++5cJ3cOSOazgg/b8R0a4da5btHR8DKgO/ZQIwfpnXZxA9N0KrOBr
0NOA6hm2191T6Wct9+xR9utb5cP+iGKqsXnSOPl9IMxso6bnq2Z3Tts1ybqz35svlKopIVVVXQmn
XpN4UQh1b1qwp9/cqtlw1yDFGAkBINAGHSJG2sjacjX1WO5jYg09DgsxLGH2kX0XnKuucZ7IdXjF
cxiBwBx6MF7K5rXfTSekJiMVl7BEZbIwcR+KaIjBy8PjiyGqkJz4mljDYnJBUTAMcIQb3gYi93Bf
8LdV6Q+MAU+xgBs4AUSNJCcPCVlcoXXHRYNovfn/HMl1bPM1oDMQYBqaZn6ZIsTgyBLGCYV9VJ5L
2L0r2kqGA6ugkHAObLfEK2O0BrJsiU5UTg9bvWH1cZWo5ygKVlF5sexJZxLYw6vLlcYl6tLnPhTF
gtKtLi/mmSU/SMKQ30hyXfJTI/FxhWVH9XJU0hH4guiBYlYF9E112qvEihBEudoSDew8FiyilASD
qY/pCxBGPPqkfBY5ulfTyqLUYXfuz385L0njBi0/hJuYKHDYnEueBOf+SPV4ftGRVDunMa15Lzes
lTZGwHzc8f32HvYfwx+7+qchEf7Bs4ngD/kHe2XSVQa+CXoDgz2Uku4UyF4VUG0H+RsAby4Ubl5R
GlIr5ibwsH0+3kGDWhCeleDgIizQGi3b0EesU7korwSQXcvZHltHvrl218Ca6m0bOE+jX+QZMR8I
DbhNzgK6hYxEw/DWgPIlQAO+hVdpgfw8q+84U7x7f09fGutFaVJnvpdvb/1LrJktb+7a8tkH9/Q6
FXDcbOCMkw2cgKAba/JwlRppSCcD8Y2LNWq/q6Rouj1zwJBZIk6NQcYchoZo+24+F3Mva4+CVuKz
PL24R821hXQaYrR7TLy161OC6XXCY71Q2kSre0YCywoifF2qgubQR1+V3se8rtkK15h/d/kg28nL
3fyn9F6cNKAa1lA9fX+MQMCh/TZShNoFF3zc3osup7hYMll5zkZA5d2uLLdx1KubEGn0IY5I+PyW
AKlzpfuKqP0lHjOA7nD95AVtflT0W23XBchiSiyR+y26U4jmFwA34RLbnXUGc0kQ8jXHxb0IHeB0
1DOoJujctrC+z+mtPQqMEN0cRqZsXJ0j3KEQKxWDce6lcMs6l9ctyizyMC8a11nfcXgUBY4kppZZ
rLsKYwSzuiM+WtWDswX5ssk1y1eoR0S+1C9lpXdy+s419Itgx2aTnEQ2MFmp8b1qYcJjwyiHY2Hd
yeAneZ76StUMF7+JAbUkTnUda0h3Jv4AQrJ3uf0RX/0/zdAst5khpbzoAPES1xV73DSidHUxMdAm
cL4FFT8uxj5urkTKnORkNr9KWlpfA72ZEAp5Ke0h33FyX1X2YUEtNbv24xbKNVfz/SLLfr2n3Cac
eL+uFDV2LrilHCEYZCs4CZvMceDwntHhjwLbRQHR94iUsu1wC8mk8fiw12WFkDd8kkI5UMsMggQI
swQcegv9FNK3q/P0J/J8qQkWtRt00VXMkK2wa2KjNOiIL+vk68M14Rz1gswOKgWT7prUEYr1WERJ
jpm8DxStxQ3V4TLQ3X3kCU4q6PaBgrkHQGUeLGe6DycSDQI+4EBxGmhPPOOFbjbfuHf3MF0YA+pY
4a8SHke7cMBPeYCsoKtThcuPks3o35mxMbREfwHNgAm5pV2QKup2l0ELbvx8SGCUEd1+oRCHgmE4
iyikrrZDAi4CUNGcr6SysH0EnqljQFJLwsh366QqSl0YZcw11idgDrD2qvLYW8udBK8upMNNxtO6
BNKFXapdnjdDiLL4iqOlTDDpcoMRd9Qfy/9tfCuqTBfs9ycusyd71hOD/HnuJc1i5CA1gtFOzwGX
ZJljSapgrXaCN5iyZCzLsSJ9o61jOPSmlIaEXGty3o5lLzDLOlRsDh/9zeHwDae0cQnVW2TqVQyd
mhEUqLZL0wYHExvmWmvNDOO/wg7bezqJJAvO4DW0a/Yy3RcAoZBI4tv02ChVtOC5liTH2UU9g22J
L+vMxKacf9+f8J/fbwxcDRZ35ZAVs9FqY7V2iAVd0e3e7dsXOXz6LuVfcAFjgCd2YUFAEzbWDJQu
QHrOa1N/hH/SJF+eC0YV9vmBouNDGsDzRDRgjm1G2+78j8AsZJBvOsJNRswxdVq/ye/na/nbQI+x
YkDQ7EO5fkWyZS7zoaeTgngwuwDuT7PMJ8MaLZPCYdlyZWprwST8OqpE5bTly1b5L0veq9rhTF7j
ByIiyi0rqP8XbrWffPg4wrjYbktSSzKlvy4boCDAnKknMf9K22zwpDpdJa0fOZOvVJ3oRRUYV2My
rhSuYPUmTSr/Srkl5o3e++Tr13ffGC94vGpRKYaMBIuZbDL9bLC2IpQGIQQAsELewjI7XiLExlzl
thF4vZh7NnyhFKokpUlr4OTdN8IYGYTpN+CSaPUogJSUiXpoBpn2Nv/kdJRefBU3BSGZhvZSwBRi
C9+PbKA6Wte178YO7YqGvYqvJopjqJAbxasdTUT01u0rJzg8tWw+oQYgyPbAQVIwrxepiQ4ZZvkZ
X5SSSDnb4k5cXmW8IA0HI4qXj/JXBVKLSXKYk88N3JTp+kheU+OiY9/7qlKeSL1NSeeKzaqGfepy
72WXSZjBTZxrqa5lziEKeG386tdHC0y5KM+NA23mSEio94rW4LSRDlRJnoa7p/c7AzHtuo52Gy5p
JcgTew6eAK9nvpUCvZvKa6Slr5tripGFN1rDe3CTwKaY6EVsRdKztYTMGRbJSPfW0HnsOENrXFKC
6wvRXJhCqSDtxz6Kehh51Yxm+Vm625FHyl9HxwxVSc+JMMBD8WsMi4ifc3Yph1R4QOFaP3MbGxQi
cKilmlux0hsgKiWsoU6qLscrOWivVWyOgZJtyPxeLkTuDjKivHHzksW57zL4xuWzY1BFD447cAJI
Q6Y1yRwAxvtYAYmmkdJSEjcTyxz1zjdYsNFop4Y62ntfEu1AmAS5nQcdIHWIiqNiNtTpaLqrPLhc
fKisnbiBalQLa5H6OwRwF4FVwdU10t6J6d89mu60bMtcYwJnm3udXFHESEql2Lnf2y0kg3Sya38x
kxi+ZYQBMjzUnW69RTzbAsKHozeg/maNvKUVOh0rQRBIW5tqPgwxqnQiC0/dvXX9+IW/7YnDszPE
+18tpm+gIVmXbWCevX+o2wnVA6KD0eaiw1QzuHPXKhAIhb9m2czgau6Oy7CmYNcY+40bE0AVW3Wg
MHzgpdU2w9doXMYeyMCvffU7j7CBYH1xGY+x1XkS0M+Tl3LocgD2KECMxEElgXdD0M6ITo4ID3Zp
pYZkiImH5xoIkwoz4c4P2UmT4VWej+0HYbk7uunY0CaFPhxMclDD+Hc75l5TRg8loXiNNML4FAwE
5xo4bZgLFKKWm6lmUS3/ApXtdnwb7N0a9BWwh6OJp0I6KsDdDYoJV4SIHjw9nFIAB094tnxYQoyr
TY/FCY6KWeUn97XAokREgIMu7sOPHFfNlH3ZM+56XrJNnSrV5RIEqcl6gHHusjKDPvb1uI9LpfHD
tNqkYM5EULLNF8LVh9J6ryJdvelpnTrhOezbuVYZ/d0BAfLswFy5yF+Li0Gr0UE90IemIXRTsYch
Ujgj6vZdRmdcMbNSGF/uQdxvfuRqfXYPepaBAsIPhjTsbcWUPEyJJ4atslsOkNzuBwsNOtEs/L7Q
oX7oXFBrRaWT7jte4Uxkc21WvddMwlYqcPthaY9FQ2Y3ByX6FAtGfi6dKua8SFORsJsbMYlUhDBp
cPXNp1zDkHJ6azSk/7Y7MjymmuUMRlbhaSBZ7MhMV7xX38Z5htJqyGEXVRSKVC0qmZfjjTUD/5+j
GI+bBGktxE4WhZVbXSd5xmgydPdzvJbc4balLu1LVzSF5ie2pcsj+N4BD62B9JKS8i8zyH8LVYiR
msrDZ/nNCsBEvW0Rte7ZfMvPrl+Nl+SYQoWVxMX1SHoU5pu8hLoKt1wNzbat2keiDII0qIF9mrWT
1h8wFwTUACoAw/5OCUqP4s7UI/4keNwIrJ5GjTVr//VT9N7Ln5tQE1FtxmJtZZA8ICU2lZp/3FaH
VOcfqrrEFL8qwR7MRcv6/w3EDFA3FX+4kmdAxEwq9oLbqj4s7xhUvLQyHLiavsfXz0GLlSQwre+p
r7sJY5DhXgzKFW8PWK3nVBx1qT+BSR2DPF+Mx9fOKgrkAKB3FrpL4YWXWImUaWCQjSm+j4uQ4+Ih
KidKy/SsH/A03kAUvMuXt+GW6ZDZRSU3L9cvBxlDwmT23ORSfGx1jET6899ue5dgKu7z1PuEuBkT
BVArBRLAplCn9X5s1xTJMrBTvu07AuoYSsG9Dlo24lWtNcdIy5+qI4WHmUuuLFL7RGx/14zXt86g
O8Oau1gX+6cMBHOmSrbFkt50ETAjzcsRjqUBSARSgrgaL4AW8XGBe65HsXgqS6Lf4wDBL7S3yJui
NiQDF+riEgXv784f4h3/dZoj2x/Zk4zUYm6DlJYDm0VMeNpIrONnGXrQTBs6ILoE/zwIKwQhb0nY
mlgtnTdGzAjzVzg5ayew9dPRawiWI3REc4FE7QUcntmsAtDOHF/uvSrdAkXbGy59aqEseNRbq2IL
HX5vBMXLcUCAIASetM72YpnUtr/nHCU3NWxjHVCEdFsp8lLuuu91KNnXgtUb3fejYhturNguLL3M
p/uQSSeMI3I6sqe5hJzmcGYeIxtBpAmSKLW3wmT2NqUxjjNwHNfU/3ZcqeX2TZcKUemk3C10JQPp
Ic+zP707O770wp93qtY9/hn4rH1txaeU64qp2CJ67+u+mzHa1RMyBHWnktDykID8i0GPa5cW/VNT
D6WGJ56hG4TYFQQhW4Tq2NKM9O294QBnX+N0UkPmvjMZ4YIVqc7m/q30s/oqJQI3zAfPnmoG/Rg9
H8DlGua+ooKCT/PlLlA4QK79DnEWr2x6kQrDh3xa4JXIGraA9X9og+8uhmaucMKWsC6Qi8htrhAI
59Bf2d94ON/WVcxybRW08/H/FcFSwrqDJo5njSVSMDkr/urqpZ4AEWqs7P9q2yjqdwM1iOm0RL70
YXuftOgXE/+JGVO1mfEcu4JahrizED3uEQzahxioAX5YDQT7TUc0X+i+gU+cuvWXzgCnNc3QRgrq
AaRMBT6LuiOMWV+TmRWvHPEgmnbKysds7jEZShlvtc68Yy4SQwsPofMQ9DGR7VL1I28lih7ZZJEU
LEttUA4UZPp0zDSlCbN/kVx8DDdrXYeYNQsTHXoPkqg2fvELqw1zdmtNkGgrwqinRcGU+yDdVArH
t0z7nIz8TWB4UKBP+tFp2mjRMCi2fB6h47UgXEiWuwtTr5NSzgEjFWhW/aaCMFqsx2jdDcv2fW7Z
8Wf1EAGpDt9Ng1Vrl7f6oIC0rcCrtZOVNdQ2IUZ/uvYMvKu9SNsE4s13Wt18S5+1XYHc2Oq/A+WN
PEQLQFgn2ciWOiaiB/M7OnP4uOAgnrv9VwyPvAFfUDTw+7Rv5ZNo2mcZE/qrmx7QQtXrwEBzD/FW
eNwUhQd50ISooRsF6tZ+mYEQq8jqHrXVAYyTgOMKr455qZ1ZDfe/QNuLLmHxyX/BSsCl+KGn9jBw
b60W04RB8Rz0wtaGVLJEJzybGGjERVIWZpeDslFMXEAhxVIiHssH0k2yce1gh68vG6QV9EAJ/D0J
hH1S+ZxBG191U4hEmi5rnRlXwM2nG4acITr/Th8HWwJ8HjddbMmxRapB7b6KzU6pA/mc41boRr1G
AxX0ZE5sl4pTJXyQknOZz5KKeOPfAaH/cgoDgyYar0ySjxcsWMguu+ubrXfYNaOEp0tKJxWMo0QU
6b+TGwfPDsfZUjMw2RTDhW7Caen7setpHhd0DWNEuiPuUcWrHncd0YjmETpgbHReHgFS0j2pUcGW
mz6kCH6mjM+tB4N749a1LfEwSngeUTAJkf1f/Dz8X9efMeqWdNag2IDHyjBDDgFG70sV/aq+lq+R
ySCeoAdO2CyYJu7iseLrS/6mbDpgUuUSZ7W6AencE4WwqWcBUrElutnFFe3/WeahootOss0V1HV+
To+c+uWMe3xFsglEK76ZiHm5gPy7nB/RrnvUmcO15ffoX+m+AgiqCSSkp4EpdfM+GqXWd6miq6P5
9A5eKg+7Lm6ZaVQXUac9VHscwtbQVDW8qwxeJkhkMSniDI0GDbJQq5Ku8YQZbe3zYbhIghv+wTk5
YRB1NUSbDxqXSX4bcB0FRL3VYSqQeMA0wYsjTqVl11bKYMXULQGvoxXy+eSquOk/toz2qKOfh+gz
DSvgfxJrqqGSPf5wCZD/a9OXiBUf0RHL0zPb9iirH1zp9tuwN5g6yl0ByzIzpn4dXxcIFfW+b4Df
RqovxZZhsqIOyNxf+u3yMbz8Lw+0/aY7l+mPBgdrHu+dX5pdZXUa+fWvva4oHV8fnpur8mEayrXg
248v5Aa9IRV8cXIkVDFsqhbNsIp00fJzemK+3PMgSLwh6bL3iU7eGVrUw3Vb8KHrlwox/KoKs1cn
KiZOV8QUXaDhM5rhYiSNwqNKsR+UlBxe7XWWSkMyp/PqIk2nx313vvj4AEHRneURB9C4kDSiS5G0
vFQQ3apXpP0owICT1WEPmcdgCqkWGlcNPQzhFDQT5rMZe8bjjw1o8PW5SVXkhw/PiOpyh8OGmjqx
9JFvxZRK5ApWBNl2gdBKNgaS0B00625titC3RI4docTg/CUcJLbsrnFNMtxNCJSHBOIt0U7tTpyj
XOqrmmUdxQuoRCNQqTxmBSCgjEN9IqaTim1wyUqlQ+CA2F0Bc4piW7mSAFo4DGWYYPHYtpVBQq2+
J9XD5f+soVug0Dpn8rdTEBXNNkroZFVs51VFiaLaJqQY5elxYz+RcT3lbNF0rZM0QSgnj49HpcR4
X13oRqxoSp50AFHuzd4yuobmbgyudpertbbhdylHNlQQ2w0NwwNZC0EkANBGnc9upTWo8QivfhHK
YWh6NkcSjlDZTlbEiJOnRMPJIpHTrIYLt9kSrHoe5/kX7zM+WqKQ+cCDrjAddm8gzr1a6iZUs8uQ
XZPVIUJATMQnSqgcT/CjXLZKQpkB+auI1bvRAqIqo072m67gewe/NisXvnut9Vv23ea3Wm1rYs0A
FziuTuqtAv/Ueh9nlDocVQ+MIxjhsP7+UbuI2yMiPrqsqjjIKSjZjBSwzqA/w4IXZWsmkKKZtNQI
/MQL94FocHjvrrxb7sq/xbynEydj7NPdYqY4QmflAKoEYDJCwQNx2B/cv+LkLYEQdQZjr58GSQeL
vdX/+3JcYwmgsh19Axv3GbH0k27RSV5l2rs22fWMtwY5c5MD0/6LDR2+22tNZVXseJKnmrQOTGiL
9bzGu5Pw3bPWibk/rU7LcsVwgn7aMnLLzzuVW74Pt/Bc/BkcMTBA519u5gULZXnCSBiPPkpBOVcB
6h1vR39cfuZFegeN8AxJPivikUwo5IRrQLjc+++yLqyL96wCs4JC1ebIkfJktgCcCbfsteGmztbX
GfdnxgkdoPo+QGhpjRZItOyadLny6UeC2rRiZv90owoaQ1UfSsqeNjghZFfNfWQspQdMsWfyWCzC
FvgHRghUVQq4UP4ZX+00TYRmoa5AWL2vvnzH4DN1MNBDqpDcGSZzmMgWH0l1IJdQFIoMasZRhJgw
RYTbA/94p8kr3hOfD3AjLCBTo9rRj2tQew21k3qf/gb7M8YtLnZcG3Kp7o4kntBc54RKXGdqU3xi
0SiJhQF3HZudYr4ch4xAihSrCru7d/PoHzfa+bOagXD+iFiWbzHnQzKZShLN/kw+rZ6XJySFAMs4
ulxaXITZUu1ob307TskYUfBTAL9vJZpRegVcDypsTWHDg7iDFO4e1sJDcDDceTVpQV8nXcIXDcXc
vzyDzqU6NMu535vYERzF1cQp6Rmiwxu6oiWg1F2fTjQ9czGnqmB/4v8ieesQR5Y1+uWvFojuJjdo
e6mK20C2482XZTI3mDIsGTvh+y8F6Y6aQY0Nqf0yCwnNpgTK5HqEvGgr3mGgZqaD11kCOGDkPHSx
4QdbOlsa5smbD8QpPC1uoNwFfX8QHHwJ/jfdDOehSOW0RLr1iCyOdINAIfduLqU8eMa2RB2ASR38
yN86Axm39G9E/gsXo/Ts+FPE3MlsiEWQZKBRZAa4wI6RfFYr+UF4IRDwdTYymAzX7IDWTJZ8YY71
H62NcBejt2D4WCRNWY2+de4jN8Y7LUMG4NBX+qeHkgMkaewljJHQAGL67MBMLqZj9YMWVOs2dVXj
ZHSNffr+AlTu1dnlhAdbB0nMNSzdiPrSMTAZiXf+n4avoqz/AQuAoFZT1nyoBxn9c/r4Mljrb1rF
yFA1UF7cos4nBSyeJU2dF0AgERcgL4RtQjwqjlxhInqNkf27iA79anca02luXj5r28B/gKe7+roR
oEhUcFNcHxk3rsUU60AFkImdAXaM3zYmvo+E81I3cGxVx/4OE5QmJb8QplFK+L9ol0zckjmgpk0m
qHAMuNzXwFmayyvQ9peoXlEp8g93lEtWWKKzlG9XPfqQhGGewYTqLM/yw0Acmn+utUWbSuVN4oQ9
Jz9ylgCo5rXk8zoKnM+ECkElxDBbyioTaQTyPUfigS68KR0nsVQOb80ZpbCOfh6u2M6p53UiOccR
KC0KqFgtDLizKnVdiyT7d2+WqxkgXfe2u5VV7Q/EPoceodMj3IA/PZiOvTu0HcnAtKaCDOM89Jf9
QwNJasT6HjXCOygAmEQoVYJF77dVUI/+gH6aruWkcYZGN4tvTzoLcd/gKtQn15pLvqf/n7NOF7py
AC3nfJlsF2BkZGdnKbm6dzntmNrk6bNXYuSBEwmSgotPADzh4OW3avi+rh+Ieb+nwS9MfZA0ooJ5
VigWSOUCbOMhpRtXvNXPRZUloRVpXjDbxdhDYX7LURKQMyo6ZgN/TUN9314kMs6JpnVzc3u0wGpA
v8Wonrf/iUszu6xHynmuaT6+bblAi2rSogzXNrqjEPWQ4aAbXlzxE6MIY5qHI1pzEXJV5R6h+Qvm
bTGSDYyP2r8HLGuIPkDUsv+6EESw0ae7NVr79V1UcfEMOWQlPnjkWxgy+kwZm83GufsFXS4KKz46
yt6i6a2qKuIDGMvnMhp5w/xOybgv04El+EntIfcCC9Cxj+6xv4kqIoW41nHvUCxaNrXKzu0QsxJ3
ZkMTYEdV9c8Gi4tIpPJKhGodpGdUxVegwsnCVQ5unRtp5o2YrwanvEBLJHcRNXwqyylKPYll6ERI
KCMRwgV00+iv9JM3t9Q2bDUv9rJg3P11lL4eZVO/n5lYauL+4FD3qPfKAiqG9dRJRbaEJ2yda1lJ
qnfRiVdzFbUrYSHguNFwFlcaNWGyH7n+Hrp7U+TujtS4RGwMKH26EonXKjdsSA/UD6Fchx4RIJL8
jKXeg/KKdakpT/L8eVZfl19p13I6YZD21gd9cZTYwRLPReUXr5nIYrBm3RAwWb/U4U4uYUq0e1WK
u0E4vMCujbC55ecQpn7NMhhat+va+uvLjcLovUJks3cT7gvi7hmuNUp4QLgHM4hKp3BBkuoGSiif
HbAoYvae2p1O9EAYKLpKBdZF4OUTzYl5qcfYiBeckt6FnyiJ0YgA7invxdpl03IBIwmgGdTY7iCZ
nbpu0N8d5eYZpsjtBSIOuORHerwGA/97/y9HFycglqtvQUdH3Ssp+KpDrTlnmCAagZVMTUldDg4Z
yqg8hpGC/u2Uw7h2WJt+5nMU10PA88UGdxitPQlBWXWq7Qrs+PY1/toeTJDyWvXUU8XAtbon8Ajr
VEpFiXbdjtkugutCBR7T0aWAw75tqq/AtvMt6UWG43iTQDzgR2vx7zpbjvqbd02c47NBqmoKeris
AH0DSGgHo/xJOzB+PNcywmaC+OHtb64FLa7caH/qaiRaJKzda84P+Y/y7iZsTzszLNjW253f12/2
RI9e3TU6GnIcj7xij77MhRrY5qUT92L+XgwjQXlhfWtTzpugbjcNr7IWPtgPlt/uu622eredAeIi
i7LgYVhtE1HJ76UU1tRsKSvbsaNVy1HDXuEHOuTXYXn5qxRbXKJ7o2QxAuGHd8sb4V0rkGEx/HFh
I6qvuU59UDqKx6PHbJ4IJIX38N/0jQOWSkdpuNKZ2/zHounXOQ1itSpqroU1XmKSCzWQOjYTi11J
c17N2gRjA4uuiTEnUIAoc9FCSneFWK5GiwHPI1D1Wv6ArbqFIy5K0Kh11EX92Q091AYEzkdU+cI8
DrzAd4YexG9d0Jb3HeWct4LMi85nnpXsy8CLRYEJpoGdvu9eEZ3skweNP3SKRHE4yBuRXaM0COlJ
PKftxDJXnkPvTCsgChbcidOO5+68qd51c4lKZu91xrHhKbTIt1Lotw+JQRbI3HWZz+s9aFj9EY/T
df6P8y5K5jEWJgPswHdqcbSQb/6NzhlzWmN8Nq1nCiF6Re8hGYSfPFf/pm8Da8I0oZWBtqQ8ojCh
Vh/XEVeB5ckEIUgFs/pAkNYOvX17kJCEUgKuhLTTqzCYox6U7JS0qP2cmy8N7Zl3AUWw6YQvHY9O
pJBP/vf8kW2dbXk/cytItRvhedqc9aljoblhzgb7HU/DFHFgGa0qi7iIKWaG9yb+B9OY8Xeb0gtu
aQEEpeaMZNj/7o5pz8rRGaK7XjHNGyyF9t8FZDVebcxezyJN2S3ZF4dZ6jOPoA6GvXsNU7x5GLsY
J2pUrvG0FV3qwWSejtNpYwvEC2fsp7Ehk8v+VjvCuwmmIJl/qk+4aChj4L2v4Tq70u6tFgroitQQ
npVyAuydyrlkC6lEq9+8v+ZjmuVsWOrxrARIOMgkev0evUsIMnTOOUWLI3LbzMM4KGQywooDw9Gd
somOXOyk2DhIsADt7u1v26Lnu1HtqWTMG2XoxrSntK2l/I0AkckashwQVDdOjkZse8UMpeYw6eRz
1lWkkK53uEAcVh6YB4Y+Q5i/uxY+N7bS9mKmJOa7dtjNob09FgYqIv8pDRDWCxaytYtz+UUazqa9
us3/tS/k6lIyF7Izkp+JPqk1oI9ZvY82GwayEbj1KsrIZhRDAFylVCwoEr+lYMfB/zts5e40Sqvy
edwLD1yfVTUD1VPn8K4CfS1ZRDCmBZRYhDVQZGBlwuzd/ZBMrxPTnGddYaE64b/JUNzopb+3SgO2
axF/gwtreovZBGNmblH2/c5t/NrCWP2af58Et+NCKduHpV5QO0Zor/2LNKyCo+MXZOOFipQJNTh/
RFxLCSunsRxGjvd4xioBOJ3Mt45SZ7GQqMNOv7idPd8pROQxuGB6LEvGvKwgvolfjQXk/O9p3Yel
5QPeXwGQ5bnypze2dqF7NWL/yD4ZPcFZMcD9yFe4k+83BzFBFAHdIYwFfvqxLDTWnHCr6oi6QgB+
9oGW3/NvpnfGUkxWmKb+h6Fgs5506VuJcLB5wZPdOGG0iyZU254tzc5761RzbrlLaqp1C2EegEp+
/B447QX4mDvKZj+xSwXGGm6QGoCOUZII5szY/HpB3GW4oBE956JOWD3U/Gr5niNWJoiqgKbfxWpr
mBHWYQ73dLGTk8eekLZqx9E+W783VMO4xqwzKB2qcMPdwyRDT/YHKxR9UEv2/0fmt84rHV239AF6
iyzw5dFeCtILXGxCI197TbjTaJvrVLyqxibdhzqQwHcJo88N966WfeHvz5Taa76zIMrXH6/s2ecU
vV00rxj9Z0LwJEzmpj5PSoVb3deCiHX2Bn1/9Jx5VNKZ7PaXutzLESkmYi9Ac3DWqctt8j/jb+VG
q27Iz8wLgtDQo9475vfzksvEg+HLaaAktub4CIxyDg1k9rRw4seet0XfG6SWHXON7Fsr/+c9RJpj
gAiZJBDaaWMk3QDXzPzsWUQlCx+cE7+oYmNlvkRezQHZz0cWYA+RuUDli10Sry5ZNN6l9D2IBWRV
TCmvsLBxBQfBdzHPy/i520qOPrxNgtS44rkQCj94gVo7+FtL0I5CTVaD6+n4Z5OW88M4u7q2BZap
6EjlSnmPxHZIg7Sd99UA7bc0tUKOO5EgQRe9GjPL3OhwulLH4i3emLnxrcixcHGExewmb+AVUxK/
f2n/g578H16k4NK6b68NryaP99BHuVJ1dgX2rjYEG06ijPnrglbihYZxOYhC7ojVnmnA01MyTQh9
Uwsihbwxf1WTu5sCvi3QMKEXMAGU4kqn6z+DppQsLoMCf1QoDMsqBj7PJ9lRnZocLCIzjbUQzk9v
4a7pUK6G4b5uObLAhOqhlwuUbb49v3BwQiaY0c0UcIBEI41qY2ZiMQrcmU+sqafPloduVk0fVXpi
iFEM3h5bdkl4d/2rYoiM3yfbHuP3pRZdubGTw52cb4+ECDKeMNN/PCSXaTTO+D3jDJ7aJ78sJLS+
5f8WMAsiIW5A+UkGRwBn0UOwkVwR0E3UcxFJbaCY/nLbWQ8NyS/lKKVkL3Glj59uOWVQ+aPAznbG
eA71KZ6ilS2euSw6xi16dXQLzqXmX5BKKp4IJZzq5BCy1CHvcYRrb8ootvDim05+0CgD5eMoaZr7
TLN9HTNz0ubyXBDIdo72B8c2o84rhf5G5gZMNYPjbHw7kAa4oplZFeNOBAcEC8OyiJLQSXw3WiAo
YzHRw4X6PFozN1F8VGJ0xBDzLxq0gcrOC7MTrsqqgOTnsF35Q4tQ2AOeKY0UxSHJou8HpOHQwM5d
hb0uN7Cu8jfjggMFAY8McBLsL3u0Dy3RBG7sffrkvzTWhN/+uHuITpRc9oQ5mnpa3ofdjv7FGfMJ
tFhO3x7VPEMlto7QZvqoNvkE85r43Kz0IT/Cgd3xev1G7hzRbsCiR4dEwZdk+JYQ01wNYO9Nxoce
h6VNCUo31yNj7AFkM3+BwrYz+3K28dsV+NJqZmjTmvk2VRoOCE8pe1vE5y0146vJ0ipW8F2TbXsx
zwHdMLbwOlAzmu0sInhgwj3bos0D5lMa65pgI/T2ZQ7WpzfwyPNrufX3YMjd9Njrnur/SeSP6ymF
2MYag2b2UZsCGziAM3Vaju66j9pKX3/HiDjz0ClSjHRiGxW3Fnuj2/wmM22NaNDMzeuHMltuUNnN
YIL6pYUhXKD2wGh89RWx6CEMBo//4JbnjCJB+rPu8cGdWj5OS9C4zurs9Vjm8nEsrANgJTppL6aS
Nk6n+rhiphcvKmUaMcvfqVbdqD/KULuO633KrAQCsHmG8jKekZlKBcpPDn/qwceZFRYjOMuSIu67
jlcWJStCo7sRUoWf6mKi3htmonuyqvDN8a2lapREO45+lqlkXFHueNK3sZmxTk1Z1RgXE7+80tU2
vo8oTpxFzirZDv7Je383rhD07wW/xf/ucs0Q4N5DQXdmvyLNnKU2xFVwZQ0X9Ww+83KWsK0+emwA
XuK2wlnK7oA5m6OvS2ARKf3skeqkQtWBPnqqqg2Tn1Y2gDJAvIqDKhLe2gbUxehklZ0XgeTG3hv7
ODfDNDt/MXdJbtx6tkBQMHuzEE5xTY3/RTelcGz3nqbpRAI5m7HIy1dGhE3cU+0WBOlmHDuUpOHO
LdGpx7Z49yAnp5ddS2OYAPAjpmppe56qk5yVELaEZfNs2qYkiiYgRBIE4IZkjK53bbKWoxxFmWLS
QPtBa5frSWBPonVmBcgs7pZw8A9qcRKizisWk9VKIyaccAQWZ7tj2hEEAGZ6HNx5vAxF0IugksQx
moA5hSjp452WU7phdXerqDUiDcU2iBJBKBmvSOVHa+69wJv/ofkShnZf/9IIUY/LFVhpRa2CDYNh
4BhPwp4EUS5q9WgMYmDvdRB6URe2FlJcXBBn9/NlFozoh+8D19BDaZT5p7EEIFIiuTe6MPXrjTpQ
+pSguuk7CotbbSbNLwWfpO4N2zp/eXkkF//P91AeHvCV37+ek/NADkPiN2YQb9n9QsvvCxwm1Svq
ftQXAaRZnsqNiHIrW2NOOL/CkFzh8IiMPrHHUfHdu/wGmNEP7T3UuqRcPn/PwEdr7+FoqPQFk//F
OEthRNNYTWnVuzT6h7dMokb5LdDMM4OicWO/Ys33wc0YW7apakDm9USWOAOy//Lv+gMIjPSvzhFj
erKfSBUVXlPYDsq+T2CnFidCYxxxSaAtFjvVHC8Zd2O12+HztnSbJP6BG2SMACYeqU+qr/Nl7quF
oUDv59oh/ru9zroh8A8Di2eUKy4ZZrly2o3xyKW8enygwHEeg/2YpWf9UR7RvHtVlG3wt/XHqqai
kSplYvaPmAdFk0KFJnz2ZihBcfDLlddxHt/qUT5KA+FSYTtmHBhyx+YzzqbcqJVtfVJnrlM7u7CD
SV9nxuVNsNbtzBE7E6lzTqsKBN7C1G6nAu5JaazqPZk+rvvRhcFayZAbUnmm5vytMw85bQPfRUAt
FR/vGBnAQrxlIzqToEwBxZzqUoWs+COcj54XD/CHsguKFkQNrN3e1UdqVNQ0w5eOPii6VBE4dK3N
MUaH55cOSQt5+wD7L76YGI2rSHWqmOVAMkyKgs2ZP+ZVN7RThYKuR4pilDggLLMGYILGnwfoVn1O
r5EjKYPDw9P9hlnTXT78vvtKTfivtwiaOGWwlSSyGmTt6nm4LuY5c8OnFtVilcYA90WOUEMRN9Jl
WeXyXMfHBZ4Q2OtAm4uf1N08OANyCh4JBp/3q7pEhhevqU3LJ8nMAOp5TGkoz4lmhlv1N6qwXj9S
wwt92jaWBFwldN5iIIbh1dH3ExkWcLjAK+NVlQ81//pTsuUN9iigHFB07RrCfsPZiIGfb6Q76XM1
FymEnIeG940XOnWv+oE9pr42aQQy3owdTVwmiLuW7J8UBoFthxejbtOaS3uGG7lqQuxDzyJrI0kX
5CZDR6i2uo5IjeJfiJqdKPiVY48c+288KVZYF/uHdKNRroAQlIU+4CrP2rGyrGAF/LDW1kKIaJUj
RSKDUJaqrqdX+Kf9RoWhW8Yl3FU95D+2DU22iGqWxlQ53RKA1VU1sBtXd4qSRJxf6U5c2isxvODF
M1aGVdyiaba5kTSEa1GbYcWTC1yQp9ZHmRTgP2C2GbesAUrQTBC28o0nORedzWYkElmcj3T8Z5sJ
N9YZpTJDjf+nZ2PQpKM0SEZhvpsFTya8GzoK8NHPwQq7t2m/aH2+VyWDj93WmuNK6o+v40Pti/wB
Oj5zk+1I+i5WOFilziSmd80S8edjfKrrntIo8hCEDL7pyF6WA8+ls5uPHIMjL1luxQnt8jYC6ZS0
xPAw7afSKJ5y55XjlYZBmVMny8iIGPIDiflfOw+rTSbC6WVsof57e2z7M3Zht0XSNkglqT0qSgnu
8xksvNVIv70uCfYlmHruuoN8EvBIdIo7qRKHaOaEz/Cd8bvKqe/0Ef9uZFjv4Bslc4QfXb//WJMu
Js5gQu5Ijp5Q1ssKLUeoVCGrJ8BiSWhqiVNnnyL8elOFCelYwuzvE+EUkSFT/eEPtQJqo+6Ws5Jh
VjOBvNNwG5JQLVHkSzCX9RNaEIlNWlpR4p7tTSemDL03imnzihjZ+kmI6w/ub/bRL/9kvrGy5ds5
RHWtxm9t3IbNb8cKuU4cZp7Z0Xd6CMug0lMIJiakFPVIa75KFTZ+0P4VXAUFnwGDfH59DgmDQBv/
kuqty+sTjpT8LZP0wgAtLI6rTpgwmVQ/DZN1se2QndpJ+oZOVtQO6GfGoU1XcD9Cvuv3Ar6AVTmY
xgxd73gDU0Lusd6XGaNOTjeho0RQu3fYcxcDtwRqDRI8TbqoHFRKkkgGJEPVwfLaMj/PlqmgWK90
Cu3vR1jbsGZS8QkXihLAbitBZgHhpCe/HgibAXTJO+v6smL+o413SrC+4cGbXxKivPIuPmmIDK2S
44PY4dRGCK/zb7K+4AO5heEF3fIhLpt7+PNtMXmSFkQBiR0zYEEDpE05NsacgyaYRrc2T1exSxs8
i4iUU+KHF90iWCtOPBl+BnLJz75NxXNMht5HsFZ6VWNN0lShxPT5vvmoeseQi2IGH1oSGZ15Lzx3
ymZwG45bgN+HpwjS2GxhTthCiTT+O1UfOGnVmFfmT7/77D/LurYmnUhTjy6lH/fXwPOwqNZdZkEb
jI2SBNynjJCZuBX8P7+nQi9ShpYTaAVm6bKMzzi502C+hMFlkdzmfeW1TyHr6MSfN0LKuNfK+HsI
5IQewarxyPo+TPJHHYKLi7jMejbMx9GeDLHpb/8BUAA1sgKvkdE9StpHF9iPjonXqp7BhypzIh06
Xkyq1vU4Yf1+IQuxiOf60KOS1m2Q3mg29OMYdUn1+izBvZmMxyA3vToTWCS6eT4rRhNupG+vr5EN
5qPf9v6QZB/+98dd0T830z6x3YuAlf0DEZNkKs3hfrxp5LB47nIDMjx3LM9LEIC+ThtOO9aQBXYM
MVhdgrycYqsai6SPw20WYouXEdli+2xAURbBSGP9oB874l/eUTy4bZWU+dk/6/Ux5TnN8BgS7yIw
aHGkU6te8ZojAaftYNJrEF7P/9i0o2kYYYNT2kf5AuSnJFzcGOpKKPrLOQKZ3dxPj9IoOdm01FEa
jdQAJr1EWRu8IpBIKTt2Wkzs0ry+20RDu52lpbf/nGUZs5VyrKe6w1dKqGQPemtv+NlE5jgV5WWy
+ZqTwJJgO8LiRBsPs/OG+prosG+VClJU31j05kRN9OfWkwPcpd+hBbboerfsc4p7sg05UHcoJx7V
Co52BhSvufIqe4GpM12LsgEqB6BismPflPE6zOonlg1BaMFNWgJUBBq3UOZ1gi80HsBBDxz3k9Qj
PMuI2N6OCjXf6bHcTpQ0uCkLj4Rq70d5sPaAIjCIgucl51dxCtc3p0KODPe2tX4IW1JBSDeohC8R
9iYMbtL4oqf030Hw89iPWq1oGET71FGvhzEuTBR9fx5bGQhQ2A7VKB4KThOQluVo2cElBginFfqC
V2Q+agSbeuu5wz/udDmw+9TZz56FEA8XnLn3OrOtOuLa1+54yomODJ1UiTEagjCFWSTO6y/rVUl/
BSdsWfS6bxByngXG6aEqZH5EWwMm/NOwS42mXJfZPYImjEkTieIG+ihrfHMiys2ro2t3pGvOk6iM
cQMJn/A89aQGAKlRdXEvnsI7+vfAEruDI/8pxUP8WQPu7o/0x+u7+NGL834/M4znATuKgc/0j5Yo
rE3SgBSVxUUH9En9GtQEEVXL8L6rbl2gWksABc6eBs0ttrGJ2cg6jSCX+fc9tNS3USbNUitYSn9Z
farzf4VDEEmCNrZnyV0rHKdAYsV6aog7/lWXgvO7SCIEpgwz1FwQ02gnG/ZViSGnQGHeLhVY7hJR
5BRf7xKDAizf3jzVbSR/aWC+FN2INz2S9E0CVp3KG528Qo3k+lWmtyl4KTfININR0AcgCWYV2bBm
DM04zVYOfR2NiFfrHAx//gsO5I+2mXne4wGEk9PWmlMcg/bJ5DCinTq/6D22sigOcRiiZ9i4JTGj
HHtDItvtGPtyTIwm9IWdRRcB/Wm2YeFBTX+Zoq6r0sGcjcVB4wQWLPb+8WXZX5oZ+O/EhR6NM1ZG
Og7G00F2y6rh+avgOWKFbQ8POnXCNurUMHfVEXqsNjw+hYleSt9vQKFgKchjfjexaxKV8u4m0h/r
R0z+T6sK72ig7Pf4EAi2F1B6DRSWdOuZkt471lYnWr+mv4JDrSIHfZ2U+c30NF1gduOTG1C8w8ke
F+TaPnK4qLj5rhBzU6TqfT4o4YNbfFKT1Yvdbtl6sl3f2mLzvc2MCmDme8KkGYBVnVn5ZmPhWN9Q
hlzvjgMDE2vDm3yPuM6vqMxrYuV7SGu8Y0Pv6pn0bxY/FsUCf8LO/7X2GaGMSvmJISFRLYPthi+a
nC2pY6MvLDax5qMYZRBn/MpGP3c/yejKFBS6sXd3OedOI24CZgHX08tZgAsdbHcFse0xrSJxmNJv
6jZ57kH1lNSrriblYcZyg0PTfATPdfH3rq8GRkov2rJx/MznAmgJaCS0R9w8F9GHnL7KbrCePr7q
QEATEmgLq6p9QhMnlz0mGmA7wxIYTHzG2kg3K4KxvWvIz4pUH93LPYiTCWcsL//0dKgOOC0R6Erf
uZ/ywFPxMz08aaNqWsZnUOhNLS/ATHFj22y4HmugQDCGRCxLdH5x61mDDz1hDl0Qss7Z3UKus0Kz
NEVR0s8dFt53zBZkpgHhyucVbgK9A4BOhIRCC8ag4pPcVJr5YSNFzqrp/hOCGSo1UScRQ7i2r7Jr
S+dlHqI9v7p/kfgT3fnKwKCYFIm21noMCykKxE9YZ9jz3fmX+7+YQqHgk+bHRBuai0u7BcbbNKSd
PJOvl3VqwcPSnjd/oO2BoOt4FJtrQRP6PXCHQm+9218FwDxRO/QjjgUqCPRVRCI6WP0ztg79xUcg
zZ4pfMMjxkhHYnSaEVDtI3KkFhQ8l1j8V5Uzo4miwTWpHY1DYt8HyLYZzD0opyInQYEkAST0zntK
9Dr9IPd8yvHhkptDzwKH0fF4RfhKVAfXqtbYXtTy8RwcgL1BNbe2mZQEFHuerF42AVmJPRrr9xtR
gyBnN+Z6fZqOdwuhxGMLtox9q2c+1JSYMxRYJt36NUsyDYGlrSgz57p2rf1pN1TFLNc5Z/Y5Di/I
1z5cylpqMWvrxwNImfIG2myaCFE8XWTioF0bWYnU+S80z+nuZsG/+R6qha7+avctEQ6C0NZSHgjd
Tg6KapTYF/gMtkiV5sYGd2JgMtd/oAFfjr6LMOSZg8sqFfyAauJKS9pV3oSmhVEa7TW2l1PPA3Ve
3/Q5laXCUSd9rBxq6kTRSMDu1q17ObkST1++0OZjvyb8PgkR4twNclYNCp/n9R/IpMQKJzS03hlc
Ghu55Y8GvAwV8IADmHkCLWogKIpyxn298UPweEqR97HVSBWTDiirBD++GmnM3f/tBipMPm/ayVbe
PURrVwqAcbyMcWBuqYWZqEhhsK9ldLgxvGsOSFhqxpxZO7UOBh+go17PQMWC2OOeRuVjvZdZai7X
w2riTiUsGWQ4+XU9ChYswxyjT/ttj3UE2GIcJyDsdhTSrtK1XQleqNTpJ1gzG3+Hesu707QO6yEl
R9iPzEZ271zQzlfTFM83eLy4jL7U4XkPSzShEWKEQH5PxLsbPUeraUT5MbtW/r1HytLiZ5wpjNg2
l5rr7nP3tNyVMGu3IL4U+eC2GHPBCNlSjKl36c9WqSs9PpKeiucJgc8Ojj2NT4oTIFQpb6rCJc0E
QZT3UQ5ymVflOdSOiMhD8KN8SIDvPcMkKYOIWwLFgGvxA5qtO37gRMEmOpWmcCUUJNJfas6Jc7ES
XVjEJQ2v268SPrq/dCp4tVwQWVR4qnH3L0Xz+0LxmvSgy84ef38E3Tfj/4oyg5EDdiZvRIM//8vK
JHPj9NP61Ig0pbJqmg+0otvsmV93K0TF8PFPaTPveIV0pSTJf8GDYKolF1iwt3v11f4FQB675feA
DWWrdu8Yqw+TvAYm7rG2CYkmKJRbRW5zUG8hyynWmYHs1YPoMnKmee61zgr1LtptT3io4bLyUHPX
ntlck4obZFcEix7iA1Jnz7z5cKnR6rG5OUl6q7uxv0qtZWUh0/u2fbH4hcDQu5omocePjzozN9NR
od4ps3LvVjc+ffv64aMKy3SvlL7D5V6DSYrTfrnI7JUzkos/5Ry7uAOLp/EDukxn2kGWvyPvKa44
XRsbLEXrzlTGHmt7EqxkVOeUqvBs78rbWnn6ioV1h00bomxwdkISN16Y9y2XAK2kA4gWYao4zFv5
Ad23kPlK2BgJrbGLZyrKFWfL7KVi9hVU6k/4si1TiI6Im8tNbXu4Pi6MPixTeiw6Evjnzz0gT8ab
nDYnDoNW9jKls16En3d9lhMweMVB8KLvhO4/gggwm628KCHi4UZqqf+OCpZufcbB02S0MhRX1zdB
WUMs94IKT9p6MTRygZ/LWGbeSn9FJxtpKgajstQc+V5hahNJ+WwltZApcbbjJ/dmUji7wDWfzM6g
Fg/2yIDoh8Ag6zBMiJEwMYb/X/Q9O8cxW/Qz+NNDrbcLD7AqIPHAaDPQYyAmoXJbY4zbpFWtDuIA
Z3r/JqNVJHCzmixbg1OtcaIHxx6r3NW/PYowudPbXQWlcTWmv35zBph80YbzlHG3qx9RAXSM0aKt
MNgwUAkhD3qLe2IFRw3Yug72i/aOfKU64Ib/0ZotW4loFS4vSrANSA7FkqlwBqJyYe1veOf0Mc76
yCuS5XaLLg6uFM1GvB2k5Jf8DC8/W20mgGr4H6Tm/aoPjv+UL4wcbBCaV2e9fjWifFxzGNO+f/Kw
f6WeYbKrcWsjNnEFS/QD+Pd7QRzQFFbmPopbJEC5YhY0Ue/NzyN6foVKFgA7We3vr47wbJAXtfH+
7+BYbDWurwJeMual0t2mT6suLHxcPER1Iwml5uxmjIGvYxW+IuvkorrH4Two+bNC+voGTwR5ihg8
cmYy163m8dgYSPu/cNnSkR35syE12qMuYl65EoLc7Q/aHXvPOskI5zZB56eC3DQ1Xgopxc8RivlW
m4e/9xzUKkcxxpEaAev68Si1G3IqL+erRuz6TOeO1UCwRspbHXH90K7Cp7t87KM9B+mERq1EaIs/
ntxTGN1YU6A+dvosnTRcJTix2HMKwnrX627OmQPj810MvyZEWEAvGOl4H6Au8ko2aN1rnUeg4OwB
FhBQigD1FhgEDmrY5awfzsCQcR/7M5/Nc7Lqh6dk7akOCzcM/+tmunl3+wqwN3PbCcui7i6UupEc
IUSExBg5FQGGS0HNNSCoIxVGlDvVqr3rDZw0AB60rCzQT00t9wjU09cRvFbGb+DlEgm2SFpnQaPv
S7MxAnu2eo0aiCFVYZq0WpmOhqi2+wlZDOkTnkG3pyAjAFmAebgoqLJHhM0H1orEguiE6K/A5OQp
BRF6NIrd1ZczRP3oF4ClnmxOoazk0hKMV5nsM+idxQ30swGfhU3jyaDTwsXhU+KeUIjM5mFy94/Y
tiAFs4vOs8XKvR0Rz5+XzNZDf8oYEBf4JGDaOBaHK/Uy8+f0AAsCkPJmdXLRpxehtY08pMWCSy2b
Iuj5eo+4ex37wo3KNTB3Ms1lBnyVAFVlUrRPUTzkkC44OjEEKsbDXUeTFWwe8eH95afsy5CdyoY6
kXXj4wlCukb3soDdxmrey1CPMWstP55VCgwALAT1/MbM4Q2Y4FnU5RycTll1DWkmH1xfzmPxLF/6
mfq5Y1F53Mapg2wXSb0yyzGziy3hbBOF/8558RiCwSrIc2T+iDWCKC+AmAzkzMsxeTfNRSdN+L5n
EIRsillgHSKgSgHMaJE4ealUkRtiYdPxG3dy8+M3sJOH7+eI0A5i6+/WSan9JsGkXOLadHUETbKI
kLC1RW+COo2XwPoxGhs51dUb0Jthke2+3qLAe2LknRLLF+CODvM6w01HBlGIAlceGTPVAWRjwwZ9
ySsIMO2tJzITRgRA/wdIiXDrO/F43OPPOuCBRj88bkq2zzTZ0jv6rUSPE/lsc65xQrrgIZb+TjYc
3bU6+k6cKu55yuyHIjA8GlEonVhDMZsY78bDE4Unm65SJEoWwR2/Vd1KKH9pKx1a5/c86koS1ehd
di/vwroPcVdro7BIjxFvJxOLEEZCVxiSlIAnPHAsBXdXOn4/pHqaPHlYqWCQJPl/wyU7nZTNDS0l
HGZYZbzaSfg4W1QmVHVyIgltpd2FMu7JIGP74c971gNLqgsUgM3YeTnY2UbO10v0nUdwnnwmH5sV
4pYnFYff1edPEUFYCryBdDVWe4dgv2wtfOTNx4v+W1jj2ulJtTjyD09rPlUwGOhpNGLV3gWCq2wn
x6Erx87YpYPML3rZsJdvFg3Fvkp1F/EwYlWdGQkWq/47htxNx6FkbkyzoL3DBN72X4B0Gchnt+38
H8cHiI46CfO0Emucs3lj5MN6nWszyYBhU2syu1ujhRIDwdhUVCi5Sy7S0XtBX2QvzGT0oBwJ2G4y
G3tFVzvolTMpVDVtjvdGOirTNXsOV8hiPHiqoM/3nRgc3Vd7SwuaW6WA7Ciwb5Lrx6Lvm0AXrKq4
TFHdjtRqhJRShe6UWS/Lcg2iPbbd/bOwNig31xOPCmVsCNqwGYfxuB54S4LQwy/XKce61YkSCHtX
3rh5Bw9KO411ejrfGYSspLlp1VRIp9njBXUAxAB5NE3umRoKGwb80gHeVN1Yzj7sPlmh2YGQrgMG
pYB4HEqqpdslN/+iqX3oJhuim5ox+SGcTybGMi1NhpAMnnLkgDOfkj8UDlZvNU2KTTIsSwlhu53o
+Mt2XZSwcrAGDhqv/qR/jj+nTODCxBAbweIZALogLNPawts6Q4eTRGErDsaXYwadc/6AhawZhnS/
XNjX/hPpqm7SIzCEHBcLc4m6BDf4oPAE2iNURlu8Ta558/+5iEZtonTRLGaLokxEcz3VLqgjzl3P
GoLfLAvO7e6JQzZNTi++g4Zskha2y0UDUPsoZbw+r/xZYAgnRsQh5K9ndMLh9HpH6gE8yIYtP2vb
x9Ac1KfDCS9LrzNOjs37sSUq+pD126Nj6U7mssoi8fnSRoSbjZrBTxpJtxiCkscy1gLNJ9Ato3QF
d5zSD2KABZS+J/RHY88LQbgySSuJdyboLu61ObCZPuTrOkcxKbXamhbGlRugLB24Ekq444/yf3EF
1XmrWCcfoFf4LU0soWF4OCLx3R5MmTZeHNwvHUnoOKmGgBa312ZJGxbeZ/rrvp+0AvabLRFOJ/3C
48ErSavPKtaJobgNRjT0w+FHtFeB42sZJAsEdQrARVUGIenLmqzqbVs4hZNBxBY8nn6EL0jOpTCt
qMktlz0CSiM3f6Dq2NzrUsH/Y2kXvGdnFPMG7gP1128G+i5QS8lnCXh2Vxjwxsc6RtYw8dem8vWb
TvklIGYDCtHXmdbPh8U7HVIuliBZsM8P9TP+chDhEP/3Tv6fniSffLNvHMbPF8aXDlX0vSg1g13U
Slky0JHz7Y7bgdvXH5UalMJwmFlk7L+bPder5QkrBELzvvFZXzrUEczrDEsuXJpNkOBt5uGWxLqh
Gd7tyvcl15iA3VZ2pg28JUdF+nJBcSjnPEsmjT6iP54KZDNYQJbWK7rWt27rjzUwHxPUXumjhe+x
WVAapVVIZRNQihF9HHcA6KiEi1KwnbFH1+Q1TJqQOikoLi029sfsRyxHzvxqb2eg+GTB/l3cSbu2
24bI4RELtGkbTXUnlsxP2RX8sIbU11oNf7XgN0pWnNzJB8cyJymm7BnBzj6TNFcFQKnyacHSSBZt
X3FNZS4/zcuH599RBgsLoE7noDfxbK+PUo/yn0estKSjWW/GrQjt8mhbkxKiH1nc8lordfnyPbNn
7nRKw70nzf4S1/XaRaXFfvclV4aP0kxDYEbpE/9FqDKIX1653lfKuycSXTRWodbDskmfi8ELGpQ/
t9tqj5/GviX1by+ya8QZ/wAa5cc45SRbiBzgknHwDYYoGA+ux7HnLwV+mPW8eJll1Svua2tgaJok
BU+WHU5lZzeUQwCQHbVDwerH4bJh+MEugY44s//zLZi5LQohM6ha8IX/anlmHhtP4pSl6VVNfXMF
IhvQ3/9p0qA/gDerHJxMRHCEEzdXzCXaBl5IFJLYz+SBuwonJGAiI7ZqiWqTh5XJkJ+y2G8TsWqR
B6WYRmT4wf3qo+TFz0AxvOcrPrt6NPVKEzKi8JSq45jylnM7WFYnEcJBWT9OfT3/DIg6fN2tftIT
TQw0YGOUW/lGDTj4QJJPIW3a0V3gg5eHjGT8QBTTn+C/5NnwA/yG4iCLcVI84WdNguTSgNX0BF36
W0dSbeK2oioakZIQvunWFrUfFB/HAiegIeszL2lzHJUgzRDJZQ4K+rj/rH172IvvqPXcRhBafYU7
iLAMrs9pheCY25iBb/7f/hpiR6h1DKr2LopNNx4AtoubZ1oHMFbqE/KwgVj49WJXAlyBc5M2qEI8
jeNeh32doK7BPirORl2mCjTsNoYCYhIdwhhASz0cJ9rxSJcJSkRlQKbyp4ffTZFHBeNfEkpTWcnm
4KvgvxJQI1Fqa3FCm7ixlovixayUq/arXYFjc/PUXgKA/C+sbrcs2dv8iyeIu+guUiuWVc9qdXt9
XcVKBtYoJjqMtocec/uFiT/sjeYmjH0BtQ9rhFxMupJ0sLTuo9/XRC9hIALij/kpDPCGZCxZqIaZ
JMQChWEciqdPxTliwvD5OWvxgI7XtUq2BteycTbBQDlHxZ81rtPvCJrbjbiNTVNPWNg3n2rnPbKV
FpbVk0e8JtEzlgksqQwlzidBWE6lXg+Rbc8l35ysKj3dIgG7Z7Ocqdz2dvbZ9XQRxCOS0RkNkCCK
EcTICxjo1fYbTFa07DZ5HKkqze1iflJGSJB3W8kILf7U8J0ngPS3cVM7vNkYz2AfdGucloVB4Qoc
XehqDtZWuHrAOUrLZ4cx3x4Up1yrXD1v6Tn2c7HX7pcgc94yaPdI8DBlqmPr7mb3JoBX52Lu8j74
B2IkU7dYynolVdUtk5JMSpeMtGcnONbZxMk9IJSxfHko2mRfsYAIfmrLCBBagGsl4gG+FoyyzBta
FkFDfk9cbbTGhDrsfDcGEewnSGtiKm3CPH9XEn7EM5aO/tdPnvRpS7JUOl0AnQDUc6dT+7fTVbvS
nupJohtjv4bSj3eK2+mKrheK4GGZ19Xr00UvkTRuzPjAkqeitjHNGw7lHk8mNRCW7B6DTCZPq0mu
m0bpZQiWsL7H3+cDZeIhMW+Dr2G+U898gQm+Zc/2E6feJ66l+HO3i1S8uBVPAvOzdvl3W/kzjdpq
rVzaN7bwKHnBjtOeonqwAU4yIO5uSVWSL5rUzUbNGtN1ldZgLSvssqespwUPucsH8+bjjAM20liz
1UsCbn6VOQC69UOu1vQIIVIeZB2HC4hCZjlph4vh3JG2pd6+DSv0sGKerSC5tf4pLAMogVkxN5hG
coqBuzBHptC8v1cfa6UMPht1DDbDQGd28GF2pJtB9i7F4UQwS62wm+gVlV9OG4y92sCNifDApr6X
auQ3/YMREcP8JjPwAz+UNEGAxnkiTfXSqUSapKZzr35+VYxfJ5AujMjMgnRbJI252sbMw21eqWav
4WLGf0gPQhaobZ56QfiiMdwRqW0eEe2E6UW1BRCvZtyBalmB3RL2DQ+7wmy2/D6XzFUxWAL2SL0a
CanrhkyXlThwQMeLuTU/k5dsuF3DQDn3blMfI9BpScdEE54CtlVNqIVutkv1B2/jgBATcXFwrg4k
12UvsTDBemI49o4nJRGqo1++18e08MCUjF3R5azuC2OHmwk1/ori3mfVxZtUlsqAs7PtfWP+cDNJ
NgWskEtc72hGtMfL9o9E+u7P7A8EJO1rkaimv2j+Xj945Y6xL2EMg9LfctMK2SKTCAQ0jCK71C13
9yepnZwsROu2O/fizHwygJE7JkSYAzCN2osJTPHKJdbLMbd/jNrSFdkWWP9csF4D9000Th3M6O7h
eqZnVAwvVfUUbUM0kxvie5uhGG864jWRCU2cV4TLA4U/JXf0iBd8JQW2C2CQdGaclGmoEfsWzcVb
RgETAxW/J/gr2sH+aOFcaby25mQmn2zrjBTkG+lX6fMHM14LstZl4rSw/5ji8xkDu2q4UhAs0Rkq
XThgQ9J1qniGAcD49+BNe9OvFdLeoQ3MN0d7cCaBwMltYF3doga8JFAgul7bPUAjdygmAzZTTaY0
QtUg1LGhjGqtYRrGip7oLzCnM2NJiLg/wM1IoeVjkNzLxHO8NtO+gezetwPREVffZKfhGjewVXBW
I/N0j1/C7jahPdberxSdXbleoSVXejEtf5/cJMpxqw0GgEtGupg5h/9hFcNI67Q0H46ysTbtnPvb
SGdcG5mXZe03358I2YD2kXVLQhgFyL3OBETud+LLR4ibCn4T097H1QCT7kHDNy3HcdjI1lxeOckH
JzgzAqIuqNU+Ijiw1bhHCEDBLzKphlMGtKGjWeWeFEp3cq6+CapSyha3r0t9sQEoYQU3/Sdwb6Ks
HWGS/zMqxoHNypxXSWCSiQbFsu1tDdeIHPdC0uHvcTEwS6+ktSLRGi7TRxCz/nzU/byUlwpKAkCS
JRFmhZrjSRJm7r3cILU3U9rNfqhfjcRAVegH/e8BR3Fvw3ju0OQmojrAQBk7h+3/U52/9UC+hLS8
FQPy1HaeYFvbTG70iZ9ZGUAz/qpZdGEMw+E+ooa4FHT4SP69znAV1h9YKa+/VPWGC93/2IE2Xr43
1zdpukD+U0/rQRWv3//Xea5EzKOgvYAo0i7AnIpwTD0GLED/RGFFmJNk43Pn7fKuTff1eTy971Sy
FCeGK86e0a0No3EjTD7anCO6f+30Klj0vQ+P1/kJGjlSlsUPcDswb9xtk093GZBKm5RPqJrH2e7Z
3ixw6A1FUmYS70mZOkRKAnHvsYlICHsaqsewnlrhN9Lvt8/QQqoegkf3x1aV/L7rMLAHKHvZvvJ6
lO9lky+IDZ+A+rgS5n7NW9JHov87CJ6mVfrlL0RyCP1TOx0JzYETvv4Eeyio95UtR6UwY0WXf35a
7FGPMOUor7wCbxhuxAV/YgcxINm7nJJ/cq4/We/GBir//OCJ9kdsvIPsICRaZH4FlThMGKAgM2rv
+aMMmrwdfmhu8T6OFMSafMtANkn9qVkh61O0usiXyWgHeiddVI+EOl0M84MpAcg6OrqOVwSCasvq
f5jdCdsqcVwBw8ta4Z0gwrdWp7/Pjf7vy3iabyOSGCptp2NNVYTtXDIGu0CTbQf+2uZ2IwOnBa0V
eR/6uN7sIuW8ffxKPCeiVjYVKl6/wTs8gWfSTAiTgaeJIt46Fvy44E04tAlLyHi2x2aOcgRfFFVJ
WMEuZ7u9x+jjdBCf/x4uO/ndAY1dvjz6S/RKNHckPN/mIKEHb7EfutIddfr0xNyru93nZzFSN+mE
ogTfvj2j2OVZ3Qm9mrTG1FaLgMzVeR8baAl7L0oXgyrjpAQ13bb2JzyvdgP8lfk6gfQJ4o5zMSoy
6jVkj6bEGTb/e8tADMmD+L1nErUfNMSjJRyIaSZPNbn9+BdH+P5mXhE2QuThOAaa6fGtuCeJpHK6
aebS1qQ6a802rtutT3z6a8lalue1k1L1N8+EvDkdBew4hXp4XUAEwOi3lbd5nwlcUqOtgNhY5Phj
MjpnakayZ6PXsHB2FU+hlZzIe5JRB3IpIFnUQ32dgcpybvHzb3mrjEK4Bxu8iDGGCnFPxmktEhU3
q1249ceL1NU2sVYwerNaO3Oujo9yTvr0fShI2LlHI9yYaUHBAeCMF2nLbRLrQhEF8Ln75qo2QAPn
AhalJXSc4tInfYnoFBLXlYSyLxhQrPxRznIencFDy0iJPZ93o/HUq/H8iaL9D3Cwn3DZmn6NHxtw
PpryUN0lbDBSJ3Q9egtbCC/y5pA1KpK4ZwbGkAWDg1MaK94MwFrOzrOyqI5ej+MUarChPAzMne+u
2z1moTqhzBr1wsaX4cgxTJYXxuFL73rjUTQa+orSoigoyzfM+iB2w+bATFQZXHpOS58WKN7r5AEx
J77BDrZZQ6spvcnXP2s9abUUOhOua89lnUzXXSK/DG7bYFJ5LNwY6Dyn3P2+nT+lQn0hUeUJrJfh
m6qrAStMgvc16IF1w55vEeHmJIK6DsxEvl6OK85Zj3I1iBqXXdfHRsRgD8i/m+Wav+cLLB2N3xiP
z9jC9e8tCjQc10KMEDvUuNCk8/+nSC8eRQCjpnQdP7Oki+aX2nljtSmgHLpeTagKaDJu4NbSQZwF
PXGIeYP5ZLD8PTxtD0UoZbSLEuXQYoD9IG6SoUQ5400QLAmQRIXxRFKdOffq4J2pWxnVKuu9++v6
/oDxPtWjjWo61mI5X8QY2dpsRjjyjEIdBH6WafU5tOse/Wbz0CJ9mnVk8vXhmTfsyGD72a22DnFl
cp6b302drU867ZwIXmfsStYvWno59X9KyplwnoFGl+yGj2VODqfkMioqVB8nvpGAt+agO+n65YaG
lDl8Dj/L9tkFd9gjZ8RMvAdS/GoIo9tBW/tlajZnGWvBv2xE4ZgXBd102Ng04JEVcg3HNGy1ILy5
h+S3O8faErBwMRePpKgte1KNossCR2OWp3f+wqmK35EUnI6iRO67aSheNdU1Z7y53N+NhQGKzPEE
JuTPlOePZsBwYnDa+Frjy1HepnKnHrzDlwvesYaVZg3nY/LPm63gZtIug+J7gWctz8UEZXuv1P/7
ypZDoERiIxhI+vdvgLknZnsZBwKaJJa/Sv7QNtio5R8HyrucTHJy1OVoIGwiEEWVSAiAhp5rKnr2
lpATRnartuPZkGMXtFH7BBCldmXDUjs70MnnoWtPykUusOQXkR2WKmtnhLf8SCao6AP9Oaq9CZg9
Zz5ftVLFDFwlwISzvwWW5avgQTegrprSnSgmdS0C9nQ3fY3DQAx6BhyfvYGFcxr78OMqW7FvIWhP
vGrIjBicF0CvISohMldhCdAC+UWvo3nLuWoXjRv6Fx+kzCnDxEzpsNR51GA2MIMIp23F+yAMJ76c
aCjkyt27i5XwGmWqEUkzRUYBT0cWg8QmF+/POO3I4UoIRi1Jh3NeuSwGw9nzpKCW1tVUDSNvGAly
bchfJaHwRgYre9ODc9VF/tYf2k2qdOYrBQRGPhLX3EGf4dCm91MOH6FAdJGMI9mfppD1QDMhPaiX
BY9KQYfNZNYPOdDAqOY44FnDjmUvY+rAWoHYFvHSpDreg9wfVthz93HRAMygr+xc7fNPBitf1Jpi
t21gL0H2KkXU/jJvS89AsAs6iPf509Tr0NMPRWdQpnRvYAHUsaB0Pisyokhznp++msQRKN5/osam
WABbSZfyv7Ea5g5YxzQcnfb1yvSbyeAcLUhCeLeIvCbr7s4dbOM4M+gT5t2lZaM/fhBhp+vZiPyh
BpDAAjMxLV7GySSH9H+6IjGyL/UtfFwuzE/uK9mSUr7Jf5ODH13FfMNqPIqFHBmzcJwgegvt+tsl
fSZL4XSedqXsidlZGz19YROX8fgzF2ot1Q4lUKAXXN7ZBrkA+WIQMMNYHEDhYr3YKFWl84WDDlXD
E9dyOpWE5z1mZsbI5x/nwS16QOe4KyBMKmSRvQyUfilPf2nqZ4I2qpwjrQhf6g/ly7joyqKTj+2K
GPKZTCmZqIWU1K3nD1VvRgxnVGeAXa3V3vPT0qmUL5PCI7nLjRmLDVYPItfabWE5Ck1spNL/WEpT
e0rvs1RWjcXWqa3bwTrKJOlmmy9Ug2QK+IxMlU79HO3h/l1xUIcQciIJuOwTGpArXjXwYHrbF/Cn
/dLQiPw+hhS+b+O4aiPO5LX2hFNG8KpNshucUYbOTVXeDc1u9DuLIMLdAhUSmne2w4i3MAo8nIgr
IVfn+/f6v8SoMeHakbrXpkp0DfRJoDAkL2Qm3DilXaAva3fQdfiB1Pf9ROmV0c8NYLfLQcr1pYrS
E5nFKkBjqOJhrtd2CHblQR3kuDiye6RcH7nMf2WOR0JqfT4YkGX3Qsq+s1Xaz6PD5W5WA7SQ4kkU
XQwmvdoIiuqELACppOF5ntjRidTyU5pi7PS36WKhnIazx0IqGT79vhecg8MFgbhSPeo1jpf8PfRy
aHUWgv6HDlQmRd6BfKWnLW6ZDPT1K80HBXMUDd7cpzvWW/RCLXgCbPq77HMjw++ubBLg5qsqC9gM
bP/cs+AOnn4aeGMH/+Sv7+oykVEennHzdG0OHN0YQsN1f4m8HcKoxys6bk4f4SkWNVyUv3IHR1Kb
oYyZCoj6N8sWnCwDiS0gbOM9nZDwFKwvT7fvdHtZ+fog3AtBTE2lTtSzJ5iEDotv7kvt6u3rLcpX
oPqUeM/hcPC+z0R0GU1Nbiunr9pd7q+IRLXCDcbspnO9Mzx3pQfnc3L/riAJrz9Ro+JQ7ojYPuGL
6E5aTTaAvqAMkmvgYeKoHfrdtLimIsT735E3e+HO3d3ZxoWSspqsb23PnZu500ElJryLeGhlJjYL
8Xl4rL5hq0GapIaqOycT9BoyxO1fPOo9Xk4tXOeD+0hWDv3cAS7koqAyudFCaPlOpWle8ZwhMnk9
ksOI1emn/vk0a8sGhJOFCCs/Y9NRrnu+eTl11z2P97iV52BGewaBZp+QC/rKmkyBUvYHqFxX5zQ/
j6UheyVnZo2wg7EFgB8Ac72hBNfLH6OSyMB0sY1tjHWrk66fZap60WNskbFCnpYRz3TN7TS5kyfN
o6AUpQJsJzbS8S/VCBxKZYUrZbYBP4TAV4JXUB6FJzFAMnd1DFaUYRuvwqoIK1cO0/dJGM0mZK/4
WqNNoNWd8JWyM8kDD1g2B0dHWlGIBuc8jfYZyk5h/bkAZeckE8zKCXZQjZosv5MkAEpnHDKUT70P
a8z2OnwUBzgfkwnfgvvmaMPkS1FPYcVZlDhY1rNjfgpYzkdHqqBO1pUhSSY41sVXl/dovKkj4bSO
TJ8iAmvPg6VkERPEraiMjeNa2xc20+M1kOc/gbnS765SxnnZ5Nw/i3/yidR93HOHwW2FBx27T9bH
8h+F7xOSbUGxA5mCJjT7wHMs0OCacUbktLbphmdqxALwGw0l+hhj88jSwYofW7u4BR52qLBWJxsm
RkbAOZdnXAg+BAnWMojA7m9atB6tZesDy6R45FOoxloeT9eTfB80EbEz7qI1vO2iV2CwtN/w+VoB
iBoa81eCkuiYDv+moVJgonDk93rfhzABnc+hYvusc9fDb4zClwxQjXrrGWB8sK1ASqIYfB+56yEP
NOutzW+/Fv6psqj1H/CS+61oDTFTHOqtYwywCRa8W67HtIZJkqbkNwkNN6SvfLKHOqhcR0+Mo7A9
wC+4MxCF3BM6Y2Cboc5D2f9dIT3v6Xp8p8KG8/YfqnlIDuLv4ihT1rIzgFeZdO3RSbFch1cn3UTv
cCplikJicB7c4ApJAEnGp7RRYKbkuuEUKgzEhgc4Kdyo4pByaZyMono8M6ilELJO8EGaXArtuf5d
1zSjpnRaXmjywGtbmvjMOd/BA1pv+Wdd9KwG/ERyBdZic9+U2m2Fb56JPSNpSUz8ZsbKcrzIDpIR
xxnx91hGAmjKrrzwwYFpWYPavrLc1pWTdOScP2325llqzly5aK2XWX1uKn6VG/JevJ2orVYDBWFW
g3TKDTT+WmFdR392HteNlBhFA9nYvXjJauAHfQeCFbiSikuQ0VdZh5349semGNW/Cqcc0Kh9di/e
vaiLuq5fkS8ODl+OkFkre4QuPxlAXQgt6q8bLU7l634Z/0+BomtQYCWAMM2/xDMLJuRrEhrv+tHC
BUBJiU9mTcbYRF40s5dCE3QIV6S3VSopKgh6Tieb7GOEvUHLakksRBJGWG22GqcqMXYuYS2NRu5l
2hwZ11AM+wOQj2f82j2nRPtlB9CHJK7G7YWBAGp+ZbLhCvo9rrDtPuW0NgXGtpiivTlXQrpzjG1S
fnYbeKtwI8VoxxkY/txgAJweLEAAdGVKolRIWi2I9agNzydyPWjTL5Pq7gi3skuKi8I6uxKoI8ZP
Op9Xl2Hx8ZRq3xu9l1/ey7ILZelCVxiI/nd1Q+JhoTWylMQ1nyv3NSWKjVb/BQcFj8Pmc5JNKm5Q
8nksuzPk1lM2uQZkwptSDg5hDvnjpkYfxRoYoV8hW9frAVdaWdXnnrbEdZcBGxZS9vdPwxV+Cvxw
oHGLiVZrokV8ZSXFEv/mgifPYvwateZLwv7Ub3sWVhkHh/hVMw+ZsizYAJbqUM7irPRv2Xjt0iaa
GEgonRXl/u+qXguMSCdPbuqNWZZQxD3UDoEqRhJBskRYZjRiX/WoS7Ffck1c/EX3zIhxkT29shqZ
H2zPooI1ZscoqS90gI53otI3vsW5l+ZYLbDWN3DOLYg02vnAQOpgF6ZvdDe8O/Wa1r668rZisTqn
H+9+k4cHZ7Cx4cB7IkzMU6tyHFC975RsV/QbbKemW0tF6n1ZdfVfdM53TsNHlamtgBazG/Gc6SdS
ka44UX/D3jznWQSEiM0Pa8Ppy7t6dcG5zQCmCKmQCpo0H7oMgxtwfRqumVE4ZBtmPoWH5JJOP1OT
wIQxf6aMQU45RzulR262vJiQWYbPgUD1dxrFRcqDw53Wf3/GEW4ujYxU1LjburDwBgm3snhQGFqj
+/6hEBQnV226HLhY9fgoE7dsK8mpXgvJ5r2wanvpkjJrKmklHEYrGMsjZrl8y6GTqWex/BJFbBvb
9+0ChCkTfz8HIlZKPBAMxV4+Er/9ZyZloJ6pHC2y+0NP6T2Cyq5GGQC9ePrhAIwZ/fRtbf/X9FXN
rvhfxEP5WijoOPeQbEPXvXWM3gwGFaVq70xIcj62q3hqrxrTeCc5BtPi4GVGyVVjPOh8UWZYqrgA
ljoG/c+BRt4VwarxWi63DOAjLWHedH7KswduJuBW991V5LWK/NQPyaz9rrX9IZY1YNsZuhDo7/iV
Yb8V7JlKk3I4/2xNFURRPbsfZIdDPym8IgeRTGBW3qFubjQ3piIEc3iuoHmWqWh4EIpSh4HbPleH
Wiw1TU2rFw/uw7gd6vVQq117S8JODZu16Z3JGl9b+m5z0B0kEfZsd/8JmA5UQgO6TmQTd23yT8Z4
tigw3InGJLuIvcifZQ8P6LhZoh0cSwAcNu55tx4Y/agEZXTht2h7ylWSIX7QNknNwvxwiYS3UeAf
MrA1XUludO//VD0QG/KCI8Cki+e0WXQyrgCRC/YTJcJipmuzs5IW2I8rhHc+AF0V8haJ05bj29A0
TVlQwLTLs3KGD5BvRzrslOZwEtdS3ki+LSpPoD8T/kpvc2vO7CmKVafmHiU/5lmbC/L+trRPHstL
dafs4K86MAB73Qjnf1UimIkiLKhfzIM7wm2PAFm6OfMeKCJ/0UcClkg2XhcMdMvC2MCEyEbQuHEu
SD0wmZCH2yrHKBKWoEyHcf7txtzeU8igb50ibSS00EOBf1kRxuB6VzbCYAyCCOIlCEoHAzb88RmX
ilZ/Til0ZVjxsgjAD2Ht83DiqYc61FeSReZKAbvYHgSCB8l+lpg+33ZfxCeZQ3/aPqYhx2ON2nDp
+sa12CQ6E0LcdhnDozazJqjRJwZcUfIDHoX7ryJfBNQb2n3ENDS9j4NNiN6zELz+i66sBcHPmpvv
njpfM4Eg9xRU4aKQH9kqNicekDnuqSvkUP0RtrZ8entMomipU6MafVxxpj1+VboPmoOAfuEo507Z
HuEMXb3H/9lnfejzQrIoyA+h9yWRGVAV0/70+TY4ZCsV9dKPLOrhTYw8bHtgbRw5ce0n1bxB3AsB
ubdELVKEEwe5DBQK3/lC+3sTiv3zqEmqJ0ueBAw9M9QIr89REG3Q6bfBcBww5vh104RXbd2+NmvI
RU5FxCVfSpa3y1GPsyanj6yO9/MsKIkPFgjrhOLB6MiHmJ4FYkxY0M09PAg+GS+p6a2ltiaaBz93
fUDbEf10vSkDLQ0KxU/rj/3nTmGanouakz4v6zJtVSd3JX6uwuckQ0GgFbUhYoMgLhfJ0fVB+Pq2
g067tgccZ1KvD5Udq2k0mRiQDphoyK3zCFlYQhBYoFEvWi7+wHN9mxQHn3OAaRixSQ5aDl58cf+9
5mBTh6ZyXKUUpkeeb2UTuHMg8larYQmNPEUWQ+XMgKmXVCcewgeNUB3TpxQRH93UPwe5MkDG3CuL
wALbtrpNNo/FbzH6Iy1SmhbghvxXBYIZ6V3ZIaKcWXcm9LyKhonYA376Y4PrYCz/V0frRaEmCcv0
WmsMSl+gB6QfWKmr1ddasZRca0iKe/hOdC5PlbJiSl89KkgwOhEpGXgI2Qu8dHKLvugMtIlKZGBn
/AGqM5RjQxBGX2pVfkuf5qWxBM969oTDZGW3gq/9dCV7fLgp5UqFcVrSyXs/mfRYWo/QmphFsAeK
DQKlkPo7hnMlP7O4WwMkDEprCU5ZpdL9DRUFM6AePW2eUOF52y4Ie5Ja3qFbLAaUFIAREHQmelJF
JowQ23M0CeJNKkUuVLpnFTLIriZVPPCEAKgNaFMRSZBSWfseTSzsbvvazbH6Cqk8ZMlKCA1RkM9k
x7xiEhIak+zkPysmo7TLxD/RLpv2Bi/4coHXDr1Bg3/xCG5Q8Yu6d1oUqNOHtfSk5XfRgfNlZBVo
UDWoE5lV30GNu2VxZibOdQZM5oWQmcYJL3MJs3pFRGM2jtJcDme6uEzrqQpqn7vKzJVj0B0m17yz
NOrmeIkzk+6aiaxIjcLEJm8D/TKp5iyTwOg8m03YQeJ6iSSOKuvf7VCaKyDRnvMulYrNvnEtpAhu
M3coPLGvCOIWpgxNjk7nhYfN0QsmfYjOoD3e4nE7u8fsrosFalSiyDS74l5fMfMIEf/Lz5neIPO0
ED8zoVuJmA1kEPGE+WJEXScg6KyKqCWjZtgNO3jeCvLhINLkDH7O6HbwqYXZJOwZaWkaN+kMLMT0
7ueW+BLqnLH+jl3R/XjOhOsY3+8YOAp53wVtsg4oGqTDnBAOY20BZxYz3MEinSGC/Y9GrjqHnAAS
wE2xVv/Nyk/t5d5ew6ywi4sM7vvK7V7KWqQKWysPnlFp4T2NDoLxHZ7lgSx9ZHjpFEwCPsGRiL/f
4bf+j8SbcxeK9lJ1jJBageLjynq3kuJLuTRXY+kwjdBd11AVTHWm1od12GFX7taiWtt7+HTY4lGm
VMtKiUNkqTW9tFCJ9IiJkh5B2BPq8tKjlL8RZO0vm6fPJIeTTrcQFYsZy/Pltcq3yul+5cHhYgYt
PaR9u0Ok8OWLqbNyVtEo2nxd6WvAXWcFScEoONtiR25CMQS/RMkJ6cUW327RAHWn4VdHZjU1KYq3
i8mJHohJA7rvRn4kLN6zEW7CGfkBEnh8lxqMI2oocEcd5+TOZRv6vbpSDVVlLBC1icMF6k1cguvR
Z79lu4HkeGlvCv1xANc/HnG3Xv0xTkWFTHbI5gN1SUB5WrV3vP0Iuu8b/ybfwxD3eIqEjwYxHp0B
V6YAVOcGTlpWckDPVosJYfS3HX85bxeP944n4CaOrHvKc96JHibQKnJxXhb42b0rOXPwUo5YA7WB
9sASxBub1JNivyBcITfIRQqElCbFzll3/RgGT1v0opfFHF1q4tFKhkhZVVBeIxl9Y3rl5VySgo7s
VHuGHr66YOozTteaP39by3N9+PGWOrZ283zxfWZNm8qLVzkc/6P65yFaoJNrNNZp3R+UbSmXVr14
huqsV71EdHij7cGGNuoI9sQsmnk5NEcG38rUB1fmp1YaDvteoDMGAmFZEmq2ghRDIzfefvDkL8Ih
CLZyAfegdud2jpzPIvQmav2wco0GMr3Log+kHnh/xFKC6JHNwwhWayz2l9yiEfoEQvkfMiCyBzEf
MU2WUZs1eXOnI+ZkQcxl8iH6u4wRMsKs4XI/qB+HqHC+YmHUqWn8HEVB6Jfb3Y5C3nVIbwHNsey5
opKUfFI1t3u/KBYeVb9OvJq1kKuUKxnDkyDEX5IMXxY0/4g4ZVdYK1UzHBYipO3V5zo83UcZNosb
Ga1KG+KjXl5IlZYjzjt5GvZ1u4yLLQ+zwGoegY0e9goXCvE/QnA+qOfntuzSVPNDKBg6pprNjuNR
7KKE6zuLYP2EgQDztEVBs7aCstg9lzSw9lcQ3AeM44T7qoP1JYxJs4MGb1mSAmLtaKJ5O7Ye2QxY
5aWCh46l7gSsMoeo9Dkj6YTcLU0gHGnPImn/eJKILfMCeRwe3xEy3uWxMwTTBfomGdRSiY4bZiFb
gfI9EAeTT25fqMbUSuy/S+xTSyKDpSvQgGhAVIVWkwGfVU8NGcPgYCn1InEeVRwPuJFi8NXglux7
bucLxYQ+GDwfWxcgSZwZVd+yHnanD+1Qu5lOajjv5Np4Y4cRQW1F/edWbetjjBv/XmvcXSjEscmp
yOO+JlCnoOue3iF4mkwfbMPHXrjXOoRYiHSRp4dU1/kqOHNnJeNBRoBNhlLN5ZFlqYq3StoGaRes
aATYLNuitErPRc44+OhE281Gj5iRbYTAV/cOpW23CUoJp66Wt0U+MoM2LySlorkSlVOkCr95z4mf
ASEixVPOckWgR2tdzugiRRYobYOWFyNRfCMZJCr8Swxmiph8SmwKVR3mSQnL2Vkd73XDYl0+2iZZ
SPheoEp3JrXLx+1ry3vtIoTRWkbrj20W+2lRtDjy7MK+/bfUYTNFHXgi49YkZMEMl6+XILmITNSI
aID/4FwD6M8G1RbR8T12bkda6C/TfFJrwNaIEqLadBKpT3qAfAI4OAHK85osrBV3vCiFcUhedgdR
waOrHRkpPrGxKqoKeckscGduaHtZuPjppKqr67oH+6ETh3x5rA64RVTwWGS+H+hCsmZ3EqwPvWQ6
JKVlEw9FQQkD2ZIlJR2iQPFtad/gPQEGrme0BWFfr1Jr/GXsRetYCGglNi7lJHc8a3bJBkPaGkA6
r8G68665y6E8YPSQ5wFeHEFEBaY8pB88gt4kTc6i8vjxhp5edPUoM68e56e9RwU5uDG2zBKn8l+D
9ffooHVPVMQyKZQOE1bH5zkH0Bmh4hwUvEE8dOqAQJyiOAJZ9a1wzcBogrd/IzflWK/UOqTdB4VT
wkzhf7uudiGVc4BGdPBjiUD0bfp7Gaql9XbVk5BI7tqpa7hpxN0GRZVM+QnATQEbp0o/zFGAIPk6
fzpjugTm634LZdYiEm8Qe1ExPmhb/XNzy5pd6yoXWh/n/tFqSzicO/IcLxcxhQAcq7AdX/g76Nhn
z5Z17xsz1WVGofBy6TbDEA+B0l5AqvQe02u9DHxZXNaPxONiyuScUHE3wVH/RDSzWEz25UHaf2GQ
M6J2Y2MLsUJ1AcIu7Euk95nTSm+MEvwA+SqIr5U1LxXjRNHZbgkQ6eeOWwxOYc4BjIbBZPoJZGIJ
XCqB+0aO6tov/Yo7fuAx6oAGYH5nPM/CqZ3X4RZEaiWsSHsdi5d0vvsF9hB/asqC4xAc/8gOS8Ir
DrR6k7QI/0h68OOp+xkDmmM6bxv7SOC03JuvHAiI2ssawNYWW00aZHucTFKJIfwgyI7At5BZ27lK
FJVjPlCOdGr8uxp2faTxwle/7K0VDQxuFf5RKgwoYG6BciJdA70ycjgiZVaTrYk+26ulKDdFwGLn
IIxQpl8nvPQM7f9rNzyb3o1gQ6sdC/m6tQwULfCXS0gGwwV27fMRdKzT/Ps8jb9c5RxpOKmxCS+J
tW0FlIYgDwxBF6xwbtAoz1n+uZYx1JviTDVP7BDBfQ3t/zVgbi3o3pkdMMCkD4m4z3Xui1mmrQKo
1uE4uo1hacbHbjZQtY/WhHtSopMObsEawAW7WIRrksA1W30wlakdmvOPOssr/+WK5490qOg=
`protect end_protected

