

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Kv0N+ODrJQAnD45jVEsSEPytnysm3pvAbJ05V2JaqTdEQNJrijqrY29nJXOyqQOIioMFCyAehxdh
SS8dEy2RvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wl26nrMFXa6fm7UAkMFkRbwMiWczBO907OqYX8JeRapSfb54ShwQXeaNsbVvqp4GNYQWgD8fiWsc
Rg1ZH/ALNgmzzsXH1hqu9qf40O6LpbgjO9M5gvRZkEo/Tsa2oqZnRuXHxvGdfSUWwgm16QfnXWFD
HONMKYo+TnX1BbyoHuA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cF9G3LQheZJrMO7arGfYkxyoON6brspPywtxFKpTvNhoNGqsA1QaxZgfesvqKSR6jIrBuWrdpeSm
PoQl517JxEpEF310dys+9f254GuonHdyipWsWNgWjbTCuw6rYLvLG1y7lYwgHlSqKUNrBaGYERTL
bx0Arf8JZijWzxoSQ9FVJxjXj/PfvGzrh6e0n/oHLpafMxMPZcDI+yx5HuAhNXSr705mAXB8bgRf
GS+N50n6SUyWqcyUqw3kHjqQ2U4vJW+j5ZC3mQaQb3xJkZgzHfCaBKMstoXIjqY6XkB5Su6aeqKF
tsdYwq2h1uyBfljsOFo3IsRsUpNIiryBaM1j5w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fN4hvSzwAQXVTyvBcSPI9qSFGq1b0QWYvne9odu5QkpUwhn44DFKeJSRI90o/blLQLnT5fdJ1IVC
mwqzRlL7DmT25nQgDxB1mM1knf9aPQaDbovHFOWTzAPBPJqGcsU8B7iu5g++kkRlIJA/0D9NUZP/
zdeXDuR/f3RpGDQ9X3WIBcSwde7JdAaZPxu8gycDj+eAg//eJ+Ch+IApwl6KjZF7Lov59CHOoVNR
udrlY4+R4MFUEO48SwDCDlqVGTYZykUVxSqzXifsrNKc0qKvKF4GbqbVHDidoVCoh7f7Jnj0snvM
x3DFGPDnokqNpDBX7xF9L6+GYPELuxQwMV3Yog==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MECPOWJAU4w/UvBGQeSeElgdlWQuUK1on5QTAzUF7zMKC1Dzhpw/yWAmwgERdTOHF4jFwSXDGCYX
dcq7yoSgrYHNe1Z9FD7/4uOTgF7lUDYslV5k/HR/cVW9QWbwl5jLUaoa4U/BsWl+xPk3gCXBhT1o
1qrFxMGkr18FyvER+gYFNuGtJOdwhkp3EWSeT0uUZpww9gD8GQxRUyHQJxyLO7OrJ+p6c8iZL8us
t83ykRj64BZ4A7H8a4gi13wX2JOPHaLBMG6QaY9NxFK4P+cAlJ5tz1UR5CiOSua4Nbo8RZAnEv5U
qSe9Ctk2cb+fZHyT1Jbe89K38c/68dSDrW+q0Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JGQumRp5idVwKA3zzoqht/27epSOGyhvfg4tXP+tPHgo6OfP/FU3H6/X1Nd4Y66ilN9i+iugj0ng
ehLY04ISDe8fLdY/NaZ+qOkmAGDYirT/RxSo79rIeXhylLKnHv9FphaO49Z/wGAPNVJcMj7acDAt
BmSxt3Wb7gOV2zsovZM=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FGXHNsFzSGXjbxp7bvoF47vhF8reHgBm6BrifhO2QcSTwMmIfvC72GA44UQ8v8jHIWHgPlay/nGH
qq6loQoHzagZ/voRdMzWla+HchA2la644cxBm8f8Fq9WGjAfrRKdp+ka7tSEmDbdQiKs1i43XT8z
Q9z55GPf5g5GdS4wXPj3ZM9TkEPcyM6MWas1txHsPj+r/l+N/OJNLRx9g9A23yQcrqoY/ibZoyFW
/7no0S9W9Nh+BPh8OXy4CwqtsvPd0/Zl0/JDLnm5d0hcEAn+3TkTvrZq0NgpjAEEOfrxtp+HqvpD
SE2gPjJVpUBZWou1zkZKYyakXZCQodq+NDtzNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
Lc916Qha2MZzMMf/oLu1x7kg2OP1jh4gJf+1JW1FlwVA7rp+ifm5KzPIy7MNWpd80kkGZvAO4kpP
jINtVWfxYz5FbJsE8/9wOeBDdnH82/eDubGFtM+tmflAlhgagjOM/8zB1Udtx4NoWO9Bn7x+9uhf
ZQPiMp4zIdqIYhtv1wQEpRbc3JI+OLSE2AaUVn0VFGxYhsU2KXR+XWUgnqdL/tgJvgkzZHUZW9oI
+nCybDHpQDgDJF2LLuB/tH4Mx32TYZIPk4i1rAlBbBj8FulkjPL3Bt1J5FG69pWItp3d1lhejER0
6GWYeYffdxyvECSV5Ziwv2AI5eKMPayvNDHRER3ebzZ3xFCbwdiWulgP4LsPxpfzo7Tyt7zr29tt
os/xvzQOjmq3gTx0cD247VkL1jGH8EWEyqV5THSuTY6Ty/dMjs4oI7U6OR2BScw3zr1x9qWsnZZ2
/kpY/5I4W0/c1no/pZ9aqH26NRbTWEPL7vUn2C2JZWXYRgL31SDWbDzQInop5EpEkmG/iJbI28g+
s81aGasIzH8STQiSIl/LyrTMJp99VD7ko5qxaDjrFamIkTFfiaa/bC+cVxdfzDNzlZzbNsHubnTO
/fgdN7M8lQHJJU5a8NXYmfcrBdvsjOfnihcfC/qUVX/YCFF+dgRamrElfIg115NRNm2t1cAn2/IB
emATmC3hLAmPK3Nr09HTfbIj9ox2AzQbNA/v1dC5b8oX3zmsgp0pjL96hWpiw+5HkT6mEzWTTnvH
vtTbMmqNS8h40gnyC0PgBhe5vbdlxBM7pnPgoqo8ZID8TY/PIegJm5GujIpcmQmoUs2byPf2gJ/F
2eSVXZa6A82XbId4vLseD4zpZcnu5k4rbgFCmFL9QZ4p0K4e6bGMdMyRz+zRC0PjjUk3mNjKN4tA
9SxWjXngmjcNaElJOi5YgzF7W8MAXYNebfnQTw/b4K/4+0Co7kTdh+4d/tH7WJT9xK4bSK7GlPJX
7di52C4+K9dqOm3XV6Tzw7DhWSg667fK28Jm93fW+LmGGVL3knittNYQDoJLwNPIIFT/AaCIPW5J
aAxmp+a+7j/55ORV9vGmPLD/iUXK8As73nl6vS5ogI2AtWEyct4KubeNVXb23O6uo+ZnaiLa6ggJ
xx4QGeNn4t1D18qhZLYVuHcnJ/qfewgY5pts9mVFk3UaQLBgWjswHuHgoFFgzXwwUiJqes5CvZi/
hTAjyZj51sasZIU5o35X09DiuON41kSHOYfnxBe/U8dcAFDiLxpELzl0CKQBbqOCl82s1Z6LiO1E
jBniSukRcP2h5oMo43gLRAcZdW8qH/cAqPW0uYh7VPlt6tBdyBKK42sAg4gTFp+HFureG0UcLlPz
GtRo6+ARZgehfL4Xi0IIpHt0FA5KBr+1Hx9VJdsUv+Tdt0yTTafA+Bnyq2Uos8pdBC4PIkR2KTFy
+DV1sMh7WTIPy/bbmwLLfzQCw93EDkZO6V9hqFfihWgVhzp9mqImpC55uNuC32YP0s+gu4aWClps
1rUGZlZDB3PG/FdFpCq0ioMtBdTGOJdn+EelSskGVpotUjg591QHzwo05Z76LQnDXEpHzA3ArXCG
pFKwzIigwRt0MedztnUKj7L451NCkoNGYIs9uqnfzRoj+i+qtFhiggE2MVN0q6PL1aK8hyRlQamy
56OxV/4t3umyMdexumFtaaBiieK8ugFUFW2Hg88d/HfldQmyi+fe6tFRzolvGv57dTcVPRAqfwB3
vDmbmI3t7VWtPcjjkfme5WKpIW5vcRU11MbHnLqlCtoykdCDzif+QVQFhz6tQfbN5bQdnSytCJVN
BvuoC9TIngUJrh6pM603i7f3sWRHVk0g4o5ZZds08uooB+id3/B5LEdcVHPU+94pA1LKzRudkwy7
R5Q+lmepzqPEBzLTiYGnpfxLA7x7DAB4+rbFUGepdnRBMXtKuHQW2ao3VAnf0zxRAUcwjR03Oss2
6vOBHqfkG38fTzkzjul/9JPi6IQLEbAOYBcaShm40piUGSMf31b8m1fC4LQBoEzQFrXthFB5Htc/
b+4CjOqMq13FGYB3loFFZP8DF4VOp11IauXpdCchAy5QW4LoWPYO0SFkzVuRoaLFk6R3d3tOerma
O1C4b9EI6eVF/A3WAIbcfAM1kwwfw9PkSHMs5R9Key/HYkGPfbCZObTJS5BiqFShVUX7HVWVY8zj
stf/3hABDy7XG88ant0evO5KUk7OsGEgkN+a68vd7kB1VqqN8PSCMQ0F3tz9/7eDYQhgzr65DrJn
tLVBc3lUE/M6ZltwChs/ii7oPSK03MEu7kccAP0ldPyjyV+koJE9WCuexo6kxwjfvoAxRDmKYTzY
BAzraMUvLGxudDpHQzHeJftqy7h68iWMk7JfZFfKhqo4kdAtW4vbLlKWZtNWnBMUapNMYr7HE6/l
ivcA66teErbUfD4Bnq4WqiRgznYGnh6nyr2IZfLBN9q3xN1YXouDO37gpljIBab2oditozMMrYjj
J2XhmeHyLL0rt0scmK/NlsbqxEYEaIaT/Y0di+h3pa5clQDnfmp29BT4JyEndKhZB23daP0io1S3
BCIeSZOp0OdiFnvEtBQAfTq4F+/0bGl8ASnycUTj1rRwwe9vW9x0lRQdnMdthXDmVmqa5AYkXy3m
Ry54UW/7iCBzSJeXOp06vqZFP3rnQDVBqc68m/4c5jdkGMDXB6ZSJXJRnxmjFUm27ezyQkOjjOQi
TrHEBZnCFUCgCR2WSY1DXmjvaq8rp2HzGuamJUQakW9n14lXnT3qNGT3R7Ccbmag8Pe3/bizNP52
/BfeYFFwDq+rFSmjZ2BsOuzLmqePzr3PoJ8lOowqCrYtAcEaRFtQ4SXWIumcmDInx1aL7RqkN6hi
4s4xJS9+Cc5qrIvohpw4Kbd75tZnNUcIfaZY5C9a+twJkd8mXwB6x/vM0N3ycahEYGnl4EGcbCuC
QwOU2L63sIa5LY5GuvmzYg6z0bZvW2Vbw0bkeSkGNN/hOX80etHBeOg2maUdAa2bc+woDOBALM8i
GBxU+9CtaFv0iAwdVgWP3QU5W5hkcQJBRrdup1XgtouZ31lU99kBgMRSxEeeo+pNmfPHrnnFbzb9
tcgtRuhPUwgvLDDZ0f3JJ3qayML1NZInICQwkTeCVY9ZM3OlHF4yTZbBhmz8k5rT0rD1N5WleVLN
4nNQYtQDzLBzQ+DSuthrxgURTYsVxRgDww59S8ijt4WfQqRTvBmUHDKVHiBVlkpDcI7UPyMDrwr5
QPwuNIpSxP+cRUk6/DZmyVbe2aJH3AFgl9GEDbqSn6qqC0CpIcmb8oGuWyxzA1XJQpC36dLhxkGx
KesJkHXIj/+tqMhDcwLIQ4VZBEjJVEJDPok09CryQGrG96KU53FGkSf1s8K1UVABBxKbMx3bieVi
DAgVDj+RyyvzTC8GiCqiKX3wDEAB/0KYV3WyqW4m0mt7fMm5tlEsDaZIr6BQmQr4cvcLUy8bw9NK
YWYtF/naa+IvwBBBYH1i3SU4nBuFjC207BjRzr0+ll/rT+mWGV/R8U4VLyA9YAzdl2xm5O/OyjAE
LPoyAEmPdnuG9VlyMIxqTTQ9UC//BRltFpHXUnPvru5ifYbCQlt/+axrj1iPII5D7zoQGCC2Appg
puRHoTCdJEwCFCcTMo/5jVcUP9+VskOdsKVzS0OCgeRzpSHNUIp51yeclji8hW88YNyuxjlcZ53t
jyp3Kjp6Oug9+9DJWUKLeFqoJdUrIUULbL5MtJX7LkVRnvYU/SDUDdrWCAvsHuowWWGa1/S5xtkw
nUVJ1DERnRWGHUscUucauXQrbC5nZfnbTk9POIp196iHgg5e8k1o/2Ee+uPzhvf8SWqg6mPhENRk
uWWLc+r/YS20ayVf5FtYo05QfI8K1lyc/C+TpOXYRZNk8+v0tFz7TiHlEq7Vw498q0hkcr6Ot2ZN
/3D++tcJgQuPN5klx3QVWIqn1iUO+y5a+I5Yv1L+gsJdDg9sNdSElDrq/30KlrdMO3DEGvr1p7Rk
Ni31tXFJEVv0xrYoQE9i+7Rx5+9jREzcRCwUaIYbFlIBz/1zA/LhLWC53p0Voih7U6TJHK/kvyz/
nhhgmSlw9SKyB3c8OBeVtg3O/KKHXlM4evtAaLlI/LyhCp9S48KKdMQqmBaKiWnn1Zjy0bFdOXp4
OlG1WkhRulKAPGWZFBXvO+R7oj6fPw3uhI3dlNQUO08r4Jzbak/v9eT5Cuz+PbyolQn65BJKhP4r
AkjTMO28ZLPAsKDfX7GxXwzHTcdgbFwEng72qT2tcjK1ilcgS+lXK9qC6Y9fs9Sv/EaEGfvVFZXg
TjApfiV405rDF+bwsJwdauEVc5w2kahNJBq7aDf4VGhrIyDCrvUjot+Dw0553UEwkn4ATkv/zbUq
+bb7U9wJM4W6jcNPo/zM1UyxW35HblV9sLioN8ve+4pKgAwOE0kKUsIBXPJ7guvrrGwZDF+xBuxF
rpX3LUNbM8B3FDTV0x1qTAyiFXVGfVHMGgDxPm42eaXtHYwfHCdcwLkIpxI6D3vYjk9yErSFTSDy
3wYFWaUhWu0slyUviLhVFnK+b5vHgyHV/xZll8OaTEIpBndAlqEBNh5CFf7pcCTe04Un+W0I2HI6
LF8WZx/d1+UUGBjuMQ+DuUgkIGamyd1lZEaamVinrBh1bpFW6Lqw6kkVkIVs0fJ6Kl6YDtD9UVTX
fyLpsAb1SI97nefo5HLvEHp5oH3EhsJof22AypdH0Z8u4R7iQbC72RXv8iOKB03ZSQyplIbiBpLC
oNv37j0HoJ891b60/02yeeW9eHIVQesHcyFmCeJZ14pw6sXbB/kkFS7XLne3bSFr3T2MXvOX837g
Pa4zgeny1hpI9+CziUCDXHxM4av7KcuX8+kHenzj10/zYBI2sZ2vupsjr17rY+fBvilC+wsPSgja
OzdS+0J+3Kg6KjQ2jk7WpAPH50N8TPz9WCz7CV8vMn4LBdASi6tysPwuqCxe8S6lPADe3MT/s/BA
wuI7e1nKb2HBljr1GVKe4zfG4qcQttdQSeZBaZIzucAU7+Nt4zhWrJopu6df/VJEAmCBMo5O1q2o
B1+oaFEDu95lnfLgrGUvRHWAXWnrduw50i4JRRYa1a+TmOVSMRxz7E1P/nr27+TNv8S479OnBivW
MfZZx0uCxYpnuSKepG2dAdjl8egDG3211HfKQIR7cP1zDvSuto/CfcxW6+eBNWTG4Iyk0WWu/+Wx
D9neqSw6R4nrCGzMDIxqvJFM+IPzD4vOC3OpQ3QjD/sJiZHAF/FZH617PpAfCiifIetj8AM1Fcgu
icDV29uYUJmGWiGqszrLfsKPrEaCviwC3HttmvfltNz8Sy7taMW1R/fU2B6jshm9xindH7wckr2D
rq1bxMcU434Ij79ETJ8+XtfCfihg+/KdJ1douLJKcx41F41dmFJ4If5Xzp8t+IHX/aEIvaTJV3z/
mXCWUvxSMdxevkxhqG14HEGbBUXR4g9B3Ik/pjuH+C9SYQowraxPIrN1i364qlW7hCQ2i4eKttkB
t+2Im5tyJasjR2rQOfCvbyUQ+PJvXLiHuqLdOhLf4byLwzaeE/XPiL+4wSil9acLAxV6zPJZLVha
PhTMWiEWKh5i3Gk+4oJaT7jQXzegF+2sIwdqjgQfqjRzHYrcj23i6bn+Nl9aVuA7OlvSfRYU8JRX
B5qv/44vblvyDgdKWAGanvvbcrRGKVuhD6X2iQtW6hBUPHKSVPTA+QHOp5+zi7gZdiATKw2O8FyN
0PqO8iJV4etOes3TP58nalCkrm8araKB/JE9hOJHciqLtFHoo/cIKJNQi8TOjg8Us+haUo7gEvob
N8gUKD0tiwftFiRy599AF9+yD5egH8osiQZiQWfFbgk71wPaBq61UfAPrw/AWkIsjKwBa3P5lYc4
ti6SZDxiPgdIwJVrJAqXPDcwyx7LMCF3zOW6WbK2MbiJJwqT43fO2QUM345TZ/rqDQqn78DRxWRN
7rE2kH0/S2HGetrGQFupM4UWVN4ZO/mhA3IJVzudEABcbKzNkeVkGHiRpQzJFMDeGEDaruipawYa
4emxhDgwCfuvR/uqCS4zziM0mV+aDvgCr53vPEZG7BNJCcCQwdlsE7brE7Vru2G8nJA20xfYfvhu
ZL0yD6tz03BzmhXmDprrRUsZsNF8A/+5UMSAcyGDpj9s4MSklaGSZffE4lM/nKLrvbWS6JJ/WJwB
owybIOxtlRoJ7CXgwsiZmnCcrX+SjDnLiHBmp61+GrgnU7drPF+bAXVy4lmgR0J/pErlncc4zfkd
ZVi0K1g86BkMMcFD6GAW1oDgF+aeEq0xS1ywbqK2pvLeNPv8lcr0HNXEp1TVZiLpIWQRwgYlYm3d
bWpobgoQyR4/mA8Nn0j6G18b91WD3nnjLZgxepIW6eAguJiSFZWX/YgiKf5gbInd5KdEuZKqGmKJ
+G8jqZLJhoAQEw59+fmBRE4wVgqga5P7MXz1EUGAqoQRnPf40St8onRHxQxGg2WuNorG6eOFnsbM
G3nZZmH471WWVgbdMfGa9QBccVNDcdE451JwnDsc2aeD/QjhjCD2MvT3FwWh1YPUFcmGom1Kp6to
RGcnsHmZqukw1rhpoNWn1Il6GH5tjTvXjxE7JWGevI8KxxT/2KgT0w3VHfSXBtKSei0dVy6JsJHK
7iByVm1m2xphU9L3zzLo5OUHg7u4VseJ5fitAkNVwTdtuzK2qGEnpFRgR3XnwMl/VrIKEubVilK4
u6tLUuiW8BDEgJ/71mOdmRTnWnA0ORvef5GwGdEi4ubci5KtvXL6HJi9nH2Q8Vo1zzZWDl5hGuaH
7haVrUsmik/YK3a1dVc+ELwHOlluz1v09Bi4vxikkuxL8Y8ZEL90KuYiB2zT7MPB9m0+m+/XPhgO
wIBE4N7jHZ9gGIVOW0tbSft7DO4r94vtxWx0cYVl9WdgKK124vZJOVWRd0+cga0RgL+kAcrubMPX
W055leCypH9pnxk2SwGYSC1OxeyL3AHVIy7gLGSgX1XVczfZ3njLyup3ZvrNwspuwSpB0+axLYK3
Q+Yta9GJivBTtxBgtPjcZq8gEZir89EwYWkKlryyn0ZkJH1Ijhqe/HIHPZF/0P0pktJNqFdu49Jy
I0GQa9bZOTi6+t0MkahUR3Ss+UUMUMIklhwydj+4EEaHBjMV6BQG/6Y8BiLDW5BLdy0/DSWZ/9tn
YWg1ZXjTPLoX0peFJv5T4BGuMNcrlSl5YVM3yIZDcTPePzE2Twym2arPOB9n9Ty1BQXJvYn2EPuv
OBgc0Rwa/YPb4y/pCKMWSiX28QKIBhnMMmtnXBQiz/WyiTWPkikSzPiUhLalN3imuWPqDXkzoLfa
UHG8fZMJ0P9o1oABg1cPLGn+SOTqNrMpGjdWi0Ik16SJO/aa3FyTAe9DIL1AyFpHWafjlStFdrHn
ASdosLosv4dNbOG7j7BYyxiVICTpmOtJ/JCJdoFojyPegIQcVA2iO7rjoEcWZUOlnpuEd8/k3A66
T+KoKMIAGy09YU6QeEbUeEI0IXr7t9Y6/OZLD95e51alx5UYbs5AdZJgimai0rGnwIrfmiv1zCbQ
ysEKJ2wC2GwiB4HwqzrqQIaWVNE7hj4N7j3NEw6Hj6I/X+Qb3JHnDWxUQ+WXYh+J7X1Z2Y2PzUp5
a0i7t9W9sZEZxtTGkNZJj7ICxJfjGVUwc7viaXeQa4aeubs1YIf54vJGS33BLK9vYHZUEzYy3jtR
a8d4gILrmvUAChREzYMMMvRVMuQ+bzAe6TrKZTpfQ+m92AR1NC8vSgTnmj3yQE5qDt8f77T0XG0J
aO7qnPnBMM7aoyqq7wL0mxTFDF2zbk/voMPIOsIpc5rhmtPufWUjtsekTOd8o0Ic8cZvA02vp3z3
iQQi50nSrnAdamvDj1XRI33vPOiFxyxP+dR3j74HDX4H2VFeHSG73npyL1GzHclB5BbskEnpZV9Z
vytcA6VbhQYCOPcs42PeKQLG6ox5+yM47yl/5p6N2VxsUBRTri39B7ubZdxQArVcDvTUeE0aKADr
pOryQivB6n1Pt7HC8IEXdmmFKhE8ZcETJqcrfgqODWqKP5gqZWZznUNeVAIw77PsQbe24IHgDyBb
DT7HMWk99onIVCk3VqgzVTEi+j1RukGbL3T4r9qmG968v/i1VuBnkZi7fkU3kVeRtugNLKopdJKL
ivpqMkjtI1Wy9tBPUrS1xcW6LsgR65DZkMrbKHTnBFn4YBs5OjwHYOifqfNtObVcjEBEFUum0H8H
v7bxNpDcmJDE0gnyfjzMzJwVeGAVdxw9bl/ghKkX6um72zWMt1u3/+mgcb3GMxjDShE6IJ45yNYw
zWUtoM3/MTb8qlW2dWzbyok8ve9DP/GMXeDR8nzBlmy2J4OnLKiB1nHPesP7/vpWMb4IEFK2CFU0
oDFZJ9HTvxFPghhaf4qCCeMf6hbwUBfslW/hHlCcKwBPam7b6/PKB+bFp2lNMYRY58dinsQ6XRxo
s7uc+dAd9tmNsrQjc9P5sKoW3Z0PX/32JYFyLTMW8YXG3++z5tSTbDXrvFiWBeIimtdKG9RmcDtx
V+DXl8sZkAQYQZcmJq8THPRyMElIbpcKZYcJznPRHebS91aDVBk+z8Oq+sM7v6QJ6oeZbWNjKwWU
Mmxbs2XX+Ph2M0QUIgWtcPL8WE9VRA7z3N0IRivchDHewsAw1StiQ6zMxfBxHUglybjMdQ6kWfPG
ca2YPR7fC87elcBULGahoJoVMaljkfVH4lSX6yNnqTnswu762KgYkA7gxhNWVUwmQC0OE90VKVkT
T7sTmCjCBA4rIZT9xX4T2/umZEyo/miyLpXLlt4zK4rzC67z9EhNL/QSizVIwdtbONoay35QgwxL
Uv7MY1bl4F7ZnZ/9PC32ckUfwM9EhuVPdoP5jMuztvYWFB3Zh0jKF17jpB0XaMv+N9RZX264sMr4
RLdrvaCHeeUmAS2uAdADj1G2mU8k9FQ8iw6hfpYJXXEP3bvDTvk1pTFDoGrmsqife/DvckKW1Ayw
PMkD7W428aFJDV6WKft86rXf8YdtqWpG4Qv78GNjSrbmoH71YRIIsgEC6Ftl+1jrh2oybdTSEc4y
NVZEwMwq8G2w6NIw/1O6gSprR1aJ0OPfkAyb+7ybJogoXxVoT2UISvbRZBBYXBM5FaQA8Di3btpe
QryHH5akp80gHwojt/QtaroZL27Ns6eVSyiOzRVEbPJjMGOKgUtQo3IddrRaldiDiN+h2kE7kTNp
KTDACa8M1c+ZNPvTYsKak9WpXLLW5lwyYvRPDIIB3ojZIKYKAy2qnkVY3Y8U9GhGb6uiCDCSsWUq
AFHs5Xf9ETL3wDenQ/qEn5pe8ERCtkFyHuc2KW6cHjhjV2WWldOYjSLSBH49IIc1xlqL8qaqPf2w
K18h16D8UnlUBiLZbeNvKc/GonNXGwxIB5tLmEDH7589V5W4znLAHJHJXuStvQcNKnogqYJe7C99
r/fDolzCq1939GQWFJDcOSe6XVLNZ7I4yQctfNq0v48CBXqmpusP3+7VUCxQccI0RnbzwuvP+qND
LpQjLLyLTHiYdmnTBwQJtiWHyMrpdv31Q4qeCsEePMcMehVWju0qr8pzB3oXUoLMlPrDAfP/imDj
LVmnSgwdvwMOHGShuX+4uxHunWqQ5YqBH/nxJj+T90qxej9yJhPDI4zNHvupkc2KVZDZXQPIzXrt
z/w1YfVMTpVSBB+TcEitk/sFY7v3O1LiyFzOSyvJzqxONU8Rk7zVa6YOkC/MCj4LBjDA+ET2RLkr
6FP0YYhnK6vzOrcFxqw91EAlLi+iVt1jlLuXcLhFRBPqnbnwhUJPOBr5AV2GSfPtUhfMZuH/w+L5
IFARe5WxYDehNQGlFpVqHIPeWCkh1bMx9LvoJ7slOsoog6IDLD3D3i1F6UZGPQFEi3fd/u9tzZv3
rHmE8GZRKkGHVM71zWOv94Lc0h9shq+BDCvYzKjOnFrv2UbLHWlYn7odDqycVlIfi+/IbnHI4uLr
kXGE2fElcWJTe66wxoVW8vcaYI4y1s1auy5EEzcIKFWDaPedZDbNIgN9l5ZDK2PfXFfNgLU+K9gl
2CTWRKJziHgSkqR+NU93x8kqf1rx9Zg5A8NKydXClpDb1Pep/dSRaW7Kvj7t4KOU9TjJeIWYS2Ty
pBRAjkDGC8Areu0HSZU76taBq9AzK6h8sxSPHCOxzO38aExrXIKQi6kmksf52X0tFri3xDjtJe9a
7Do4qTxEH5L3e0Bw6wvYFcaet9rOGh5nXR3SNrd0Hk+IufyWxSQVUTv090VmQ8B1dG9EInUv0xmT
TrYAlkGZBzl4vSz52jhUZTP8QKVQPArInZaQHN+LkplnJYV2ORuquBy+JJIwA3TIdkLJQPrnF+H5
9QXxxFdeZeAKxBLrBF6DKoWRfOWSi7BNov/aZVo0eNEsnUszGWI7mvh1nJltdqyWf5mbSd7gclDV
64tfQyZPaCKQdIt2ujW53rVb4C2MQYfiKYox+b2/4Liru4oa8h1X/pYQs+GFbEXeAHd6CbTCuDEq
BQ0XVDWUWHwSZs66mSUZLpZsyID4FoL/MOCa/ethy0sPJ3DvE3Y04a8FwXbjKl0Ei4hldJ5ScEpk
z/XQUUGuXDCIxVrokQozZ0Nqvov2BdQMPbZZywZS8tcMl5d1+02/dgPfShV3A+ypwZQWm6NCqFOt
+dY5yX9aaxgMAHkM1jX+fiOKVcnlsKlp2bqD2kynn+G6O2mdCIkSS6Dkib9rltUnR71aX8scqTIc
ErcFwG5Gw3uq22/WJvnRJWqNZIih0qzDXSyOVUtiGXKwABWoIv43wLJis8uwf8V2Uf1O+lDnuc8A
kNbYMzLCmRuux1K1K1W88U6g5MGpSMSLo68EglyQvHSUcdbe/8ZXm9l9lDJ/QqX4HWzVq7rNN0pE
7IhfXRCl0FvtF9f7RE2bp7gl0sBq2jXQYVqsU8ftKawKpgbZh3M2BWlJI1ec+yRemr859lE2nKvu
iPk8ii7nzK9DyZ2D7P5x4vHJx09UOV+vYpKOkORz44W1THFzeagK/NpQLTULDabOi3dsGRkoahkl
rBZPCvN/4eXxwyWlS2inPheS9d3QH9vterFYKTMuxgZm/7prEM3G1PcjN69RF+oi7FWms8AA6GHQ
CF2WrvDxSoDcWB5SUmspMTZt1EbBGPGdCLgfatNQPNB4/4+4AhOXdKUl4xbCBkmxnLqhCbxoQ0Ki
Px0qL0eFemlKFgTocJRFpYShmAXnmvCuBVO0VeeJNa5D6F6ciM0n4wpXfdgrfL6S1Cwo4Szd17zO
kGzPcpG1nFiiHfkoZwYNzcCGjdMX+8k0GGd0JQuDK5Kzp/iIROek1eWCutWLw74dtxzGPfDPl/DY
OmuWtHxDfqk3y4vytc+3ttsnpgo+qSdoLxzB7/3jWwRHP3gxl/iXWKHE951XDspCBjOAAlqz4BfN
pzq6AqgTCnMQE0ml/t+mfE7tPr8DeM/j46BwEgkrT2h+SS2UREUIScJLz6LW0QZM1Dr3v7N9rcfq
0cNLVKMOhCDIvsL/SPicfupbnlZ6m5GlN1wqYBXOt8ZRGATv3y9uz/3mPNBeOjPKCsdpYNtHnmu7
GN1DC6cRlRdc1QLZs0eupyRf0RXMcmz6c/K7bpoWcN2jq90oCL8ioHTwvQ/rFf+0V4JhKzjkHLia
DT22V0ZwDu5SkX21nyfPQLekxQeLo+jPoxkWtvFhDLEimVt/Ps+vmOcQkPCOSCgYx3PqAQOMCCfq
AW4YBUlNP8GGGF7QXaSNjFnZrS/AxC4nKyxBnterU6ac53CNAYO7XLkHn8BcjMGECaElaD1DU3iJ
65Nk4YcODeDW7OVghVNaNogoHSrH+o40Ngb0Pn3oz6uCpVQoPnTq8LjTPooTi8gus2JxJ2sVZ7iy
Nf1H9uiPHwfm6qYV6buqBbkATwa69vE1tD/iZ0wt6K5KtSTZDeLVetKEVN7hcnTo4WEhmvE71oPM
xvsACwxAC0BEKY3UycURLtI05CTcrjzHct/63iQ2cl7uerOx5FwAWccH8wf2DZ70Exxq3iZdYCMs
pPocCzUokfOPmH1ukWP4OLe4wJzqItQbMtewUjtrkTnlAPcjzf4y1LboR9Y0i6nDSa6DU+U/sZNd
j+Z4gaM2Yvkj2iD2HK9313J6XnjiQAyXEk8ttCR44iymIN9IyNTheIQWDDJZ5aCkBLzyFEEgwKRl
2lKJ4/1CnvyJapeIzvo1gdViVUZVLkj1S+YfJe5bwaeE5hvObssdiMRrpI0vU7m7bMhX3tsLyYji
vcYRws9Fdx7s6+f7+I/XaYUgZCU/PIiuKpzSqPqx2wnwv3A3hurm1VBw/3p9WDewkrvczB7I/Sn7
LPFUWpFud6qXaww+fvV95mtnbP+oXn6y3nd7WiIUedZ6xAZ0vQ8qP0ZvGqTvwPNPMWGGP3yy1BgM
ZCIf6h/lqvj53AjO7f7AIjRH/K0UdFyg9NuDoSUmOO5KUmWBmSfgfT24FefFyhe4tEGhRNgevdAD
oK/mbUnXrL/1a27VFFkJ1Mfqb5nNd9X8YZ2m9GimknCc4wVbpf3zJqPCKh6syggOL9i5/vCS/lx4
Vh4LdrcQRJDiOMjR9Z7RzcMDMXMyYla07KFjbEqupQjzeLk4taGsvyFKXPfaPaZMKCFpnKUznfyc
G6vIs6KKOcxkgbBOc+VQfntuivXIKR/Q1muZveuYneeyom/c7CRsklNf+FHJHOV5OoJvMhZYj1VJ
B36ZJDNQytjRrq13tXxaIni0JKADJKCnD/uFIGy7Q2eyo9RUJM5Uul4+xyc6fuEERegUjozOuMva
qCl32p//E9nYEikUlyIpPqPa4aRilNZS4cldY+nWRoljmYSMxC8PVl++FkTJU5j31nGi+2bw8wXq
aUPc2l3aqUQVbxNM9a6PgKVEk9YASufCyHHe6vIC952XMGrqVEFH67occG+QzHhBs9tXFhI8IIIq
sgo8YCmWIralwIHpNsiK0iD5HcEB2ZTINYyNLT5IHwUSm/0BncSCkeBvOyujksrUiqOQVdgGbLLf
Mf6rlxSniO3BC8GRZNoKddnJygKM/4iwVdahQMfT/6+Mv16M3MISJdTMLwS0ljTAgHkZYKvcf6om
hcjUj2iwOy+OcVB2W4evAAzS/NPAVtoLeh9RfF+T2aQgfooMcQlpTid8AKC/CXT/IOCFL5+sjjXn
N1oJb70dn4NZe3SdTsbErYJSzVGOvCR9VmwsuyGW1tddgI6UZBYfZZG3s8GaI/ZiNL6SptcNJKWc
MoVl6bbf0/23FgOOIANA66dtVVQcf8PF4ezf7pPhVEWcwwChiyC6dQIASi9zlGHISJyje3XlOMM5
V6JPjfpctLvSbzVnfeI6XQPJUJNXEpp0So3ozEosXNXeM0N8A1+LuuNcbLFVrO6G8a0bElAYmn27
DM3hYtsgnE+W7Q58d67R2Av+msXh41rR9J4EY/YxMzVwICpbPMpN5UrV7UR9xLiyNEFbvc4lGCeJ
b14OLHesR8jnG3u8mjo1G5lGKuqeZpgtcvaIkrwU+S1d+OLf5uLSUv9CPXH9qK6QsQN8klxZRmdt
xRaoI0tJYKpqq9eNGGIDExNEVbNsRnrIdluq8iEPK2aH4Y2Cd/LcAR+uiFF+W7jiweIVdBM/8pbM
aS2/SOZ2d3qNO7/7PGTRj90P532bqnR1sFEkFu4eBAfnNQwBipaPTt96EUKZlZp6TUCHp9OvrgaP
bNSsREKzhLVvjkTV4EOP5PKFKPesHCxn8+ktx9/P5DE8SFeGyJMYzb1e0tuLY7p9gHlaC48g5Xwn
dnvJ/34lvQtJPEEcFJpo7nrW0wPWGjw8mxyVsuYwPt+zwSMPlyEsbkxvrK8h5dJxBxHP3PRgw+dC
Ln2H83Qc3OAROkDmCz8TC8iXEHnrALezJ/qa5S3paJv16/CKYX0/WU7BSQYTdhbpMxeaNphVYx2J
o5uQrAszHrqaybdU+7MDh7eCZo31xYDSXbPhR+IWgb4g6MxH2rRLoX1bSucg4H7FJzFOHqWMjc/A
Mefo7tmATnv+ldSB0psVGK8+AiNrGPpqKn52386Yyv3ILs2UX1R3v6YTiScFcYjo4T+VMRNzDeom
g9f9pGPpz4uu6SVOAQaXMsJ57BlKZunjXFHE0ABAGX+uA65+QcPv7y2FyPlXG4H7AfhhMvXzJlab
Nx4Yq8b44O+dkez1Mzmkhd/ueIGSM3/RuSPRvOLGyOdQDAQXpzMjd2TgOGLFWNf1yUkQliuH+lhV
8poW3752nKeCALpBH9McA4DuQid3m4Yw/wb9aee7fKMILogXq9V5UT94jp2A7Ibw2Who7SGO8kPU
OSkeAdBrujPL6Y/3hr9yGRDPs5naAEG8TMxzdj+MG4ohiPN25wJPXGOanN2wMJr15sGF0QwJ9OgX
RsSgrpE+s7kWY16tF2/uzZKzBtB0jASrG5iELeOGmLQSDJXPZMtNKwX9bxR4o2olH9GR79YuL+rH
Wd6Gr1danKhM9xP9zO80xcCN8o18SDqkYungcAt/ROCbE/SM/vWkfbghrqF3g8+Ab1TJzDiMW00c
cmhHIlnaDhvPHpF4pcEE7+OyQAj8MSwcmusuHTAfe6kpT432afXqvzXu7hVMuMPfNpkFSGU+Vu8+
zgtelacAl3/Equ0q8dT0tCe9s5Oy2bSNglVZIGIwbwoTjcH5GD3/VqlGDWCxj3q7ADkuLQy+HnrO
UmFUz7HODsg3vlsTCYqUSr6RZDu0QaMnGTu6Le6AhgpLX9k/RPuVR2QWjbFeWldMeAOGtCXU5Dfb
HcOfnYGHcGYhJLc8smKccZo+Ml6VhTAaWmHBHxP78okUnFCNzvEpoJ2CvWqcMfuzRGPqxk0LWW6Z
OGUnZDL4FO/S96jEZYGuvS+tZK6FFW+UShDDlZmCwoYEreiNe3YWRfjDgAHmEFoJJ3dbOpouXefJ
GURIQZs56O4Qpa41RYqE5jKnmjVipJkFkadOSXEpBgIFjmWT6/cDtiks3hZVMblX1osEvmr9Y1y9
XuTrPeRGTM89niXswng5q9SNlDnYMxEeTN+Uzyjoo8I7lw3bkDtwScJZwBdteciFXB3xfy6lK1R7
/eXSM9eqorP0TVHjiBg+lZx6KLcVPdkfa3fzhqM+j0+bt8uZmSyQAUmFt6SRad+8W6C1/RV+eaE+
eBOtRBHS2O1LGISOCXrvOumyTAHbcMyMy8JPDgyVcjaGTEH3S5lG/fylJXXyKiOxvJDK7uf27TPs
lMmrtY1fu1RkYMc1KlJegzTxIIPypxg4omxZWa1P3T3VpToUo0jdx8dsrTmpE+ErCQRU6WQ48IQZ
e6bRze0mSBqNSZH7DDQHerxzj+p+tF3OtGIV7CtXxF/ZgG2YajyHDf4hvUERfFx84ChSWRE/qZ4W
LTauaavlR0owFK68ws2C3JqiijxraIHmB+/W5UiU2UcGSr5C6HFIz4SovlBImJSLWTf9U2xtkQBE
gESm81xASCmN7/2GxXLIwzCQdmD5qlmZ2JXJ6ktbTjWKWS4uaf3B9vZb5eYIgf0+pav0oxyxuX9+
5acEXdveVX3QWnsJBhV2Ve/fDwoNHZ1++Cp8Tu+qbymUu0Msl5Dtz2dVDmth6qEkZD3wuzWm8bKJ
RTlpaYjcWYhl5/3PXZvKDNDLfznDiSeRimro6bc05elUG4Z30utCQShynFQT55awtj2UvRnRgvbM
RSoAuBfaNslor3dFh26q9sSSLs9pOYUyOsI092saNt9WdtzstCTILv2P9NT+xRo6/6DeQgbXt7bH
3thie7UGCyFcn3URp1RjNX7WoJSPJwC6I5mlp7XoBwP+IFij8jwL2lc3t+PCzG3KL5sKBWpBT6Vd
+9H1yJ8dG2lZ6BQcPn0va0GX89Qo0bF6zcuh99d4W7ASTHJlSrT8aNgSALvjYt81oVT0zi8iT+rB
XRdghH9vyepsh5obdL0fktC+0+URtmIcdOKXX3Dbt1qUh3RjyuqIwY1c4Z9b/7GbAbsETjVfdsRa
dFS5epySiBNfwy1wEgs7zrvv7ccTgYLwOKgyUAQlfKOcXOUqY1qgNqky6xkefk7haDs6cZ7zf1P8
Ga0RYbACBA7alNo/L92e9q81yR2cxwOCqSMz26jGk6bWl+aYVhWeu0yLFIbP7EWrd6yYokpqmBf7
CtZrc16yO7gXrDpzQA8ZLRcMVE5ld74szwXHLAmZedSEKegdYNUzNBGa/B/ABIQT6T+fXG38SbTk
outofJpBHlifHAEEDUj/YO96luOzZ0B3LDRG7+W5jbIs6XCtZHBEfqF19p+e0mkkPNGcDNoWL7qG
J/u7aIuY3WpRZdk8BkFoA7/UpoVcImkryGdQZYxFEwIm0xNGRdo/YBLkRodQyoveRWwwbXhZDTD9
ieK+IZ+HNBMw1WAAUJdVEnHFSgmEf/kKqsKMzcr8/Rl27mmDx4+1i1fPA8mBvpz76SQu0GliT3/l
aNtu48ZchEZvYvza4/kXruPv/eHl1AOAHCF3AmUHSQAQWAudaAUJhS3bBb8rWP11alA9RqqJSLNE
CHJC6RKwDJ5Dyg7A1BZ1UOIZUOPgohXmZ06+GlZ/9DIRf7j/bQbkATHsSccKBCSTJdDHFn4XMIwL
NpTzt1ZK9ek16oVyvnLqz5zA0x3vAynLae/knGvDSFx/8EcOXR4Hl7IIp1CDZZQ/G/gWVXWgplGG
LBLXxsW4b1m6qJt/FDQRm1B7Ih0alCzbgaTVqI20GuUA2H3jVsKu5FwzVLCzr9ta0msCeMoMdRQc
dts/LKc2O7vhUqhqXIQ6y8DWp3QuXeJqnC/EglhB0xq9klNJTtsOLE9UvxCQnxrp7w32HoFxXQQM
NemnGLrqJnBCXX1im8AtWZeQkhUhNzRVdzDSQpkGeuivg/quAJ4Z2xsUz9ypPAalJ0PZcPSd4tEd
4VWygcTy0nsyi8fR7xoXQiRGYLZJqu1e6vuX/W8wDdXhobtxQdmsuRkftjtKDJpfmldFBkk/1KrB
y1WPhfGS+ki2TqCBGQeCDS1VTsVgAxq5GYR8LSCw9QMEuHS7q24b29llk1+Ym8iBicOx9T9W/ZjC
GddtwP0qHdz+ecco7CRF1OS4WtQNQ0rud29AvD3tEn+DuT+Gg/WQc7niBNnovijlfA9Cz1fak8QP
l8WKnwqYWgOmDtoYLh+ZsbqdfjsJ3vpZhRjBcwoabtcK5f37/FxvE/7YIBoEYQwq5D34GTSkOmka
795ronyqMeRRMKj9wzbquubuOit7GR9/PNOqIWRnybhUUUhxV9XpDW2CXjPJtCYbnu+36ACZQo+S
CrJEDRYtFI1+Bn3gN9zofgVSlIaP60XKERKCLs/8ucEsB2XEA376rDHVwYl9+irTZmg5eH2hRABh
16FXBTHx747TMgGaeXwcUEQBwf1B+NvwrdtyR7rCJf0FSqfcJ90BifMOwTMsrzUrOGVcgb6iP6eU
jpkWtUCfMrZWVWRNmNiL1zRloYhau87QreQyegaALfhI98CFRoCKDtijIf5WZC8GenUDqVkRkpO7
ubkaDMI1I/hSwpOHmELAhhb7GeqsOAglkTXpYJWmlp6yidxRDtwL6ij3gE0ESGGIOGFquDVgqwkO
bB9Kp8vAjl/wbH+w3bVyiJbXfblkfBtgUKMwzp1Z6dM9LCEXobFt2m02MAvZbictYZb+2Ldlri5P
N1E6SUbx7vggowigh1iVX5QHG5Lo6d+zaL3wNwB1jf9eduXO+4snElmmUbeiQrXqne0tNbxBHho1
1Agi/iSbnCjVEtUIQuOjPLHO3c02MjY04GL1ki4/m3xdkVCEMCy2GX2jIsuE3120So3BhYDVeqPy
HLlelgCJPG1iRFywSvOlUFh94hcJggAds5TQ4nc4ZagWW/YXDW1TFfAPpige9PIYmcYNQf97Rsk2
S6iMwzUiWYFh8TvofD/Iys4V2fsmLOud5S79Rfqw3IOUVqUZFp2Q9LnaRPYbZkkj7BwQPoXEiLcu
4m/lPFLrjXWU5ZSYCKEGFVOFkNmnLjqKe9IKJkhk0pWBhUIcAad48e6QOZMXob1oDo7BceZ8u+qm
dxc3pWHoj5DrUVd8IpV/zRHeZFWcPXgETWBXUq79E1JSgIV8C/Ao5tmIFYny1iKceV2vrNE7Qt3Z
MZz6EBa33BOTyKjCbDVT+79CkT2sRh55RiNmYcWxP0+4UlfoiMkNgoSe1JXLjONz2SsNU/aiLaTS
ybuo39c9NuZEv9BKfSz6/fQf6X/szsT5bJF4wiAaspfE2Ya1gGcb56hFXu2OseqHvT1mOK+i34F5
ZfQH1crPkvXknIdnRQo0wnehdOHAVe80YmrCaJRfUFyj/6wS6oTAzDx+lt4xAzy1l+kSSXqwPZM2
HNxrJ2Tv8p/uQmiwu32FtWNG8NuEERDWEh1Ctbu1lP9GTVY4UUW8MVQOedT7p5O/74rRkBio2hKb
qrL1pir1uUQEiE4GWVrpL8otUcUEMh7qdy70ras67At09OHXWKtrOlAKpOAJ4hn5eymJWBgoMGhw
PaovDCZli7TwbnTz9oZuKs4roZbzVvrNwnYO4MVzE9SdZ/4piA8nTcw2OkiJ0tprYWdmxJOj4bQf
49BVVbvJbb5QhYPbHVwaJdB8xQclQWcPExi/pWJ2qNtPWMcyAMYxh+sd7xUeXNYqOR3eQGY5lOq5
vui8FQptrnUgkLP/5QpN6CeQGQVxY+QsmpzH/44Fl6kB4F9P87S1xtDERnQNT/zJdjPJErQ53xWC
99dr4fKNEL7eSvjq6lTECQAOA9btHrIN6I1ImFw//jrBgZRxR0Y2o1tmo2Sco2WDhOVMBP2SY4BM
eSICVsUIM0MNCbnX6UaIFjY5gIMun5JnXKOL9MnfocGqFEs5E6ZjNIlYH3U3yIgEvHPTbGvk8li8
V4GuW7XdTo+auo5ONvjCzuUJQPs3IZDfM0fmsSVeMkQI8mktKv2giUYWC4/Qq8G6ZzzP4G6//185
8ITfwVD6L460JAO6Fmt4ZU9+UhZ1xBNB7dspcQITA9RfyCyUi/ZOUGQKkoU9sHbhHmGFk6zEArG8
d45nhLdzoJo/c2XBAkoUoecZdSrcdfc1rmthThspRv38KoTgC2LYKiHibd5a1Ex+5slvwMagi7vl
Kv2GceQCu3659+6hXqEFeH2C1ppD/ASF73+tz2vRdvHr862DP6hjT+t1d2aoe45pbOgq+im4Ienc
nKYUv/vFkHRoeJjWt97kOvE3ckQ3vEVKSyZZyT8y1vWlIcWxnXfh82uKiTJiUEuKUQvrlly57ucN
KYrJl68VGk11Bd33Tce7bRpqfQAj97ZjQV0cbZfIQTSyUcpPNjtAvGEKEoVBrCI87Eauk2WfCCzw
fKVAeoH1RMKGbqIZNgKrwyM2hNWNHo3cUmYk6or2i6d4ZZAurrTtvzjbVuGjB6EGe8uJYmVfobXa
u304JSM9Us+QxJhSrpbgHFBjyp5Ll+Q6vXVKqeqITLj9sxJL1oLZp0i/sKgc257m0kd2hZPks9sP
eBTwpJIaqTVMEkVMDkNJP1CMG9sw8PiZMBvoVFZDaDvQer2ZrO5MusYKH7zs6v02plADYYT1AiVp
OMKQN6w1blb7QcdY8jV+y9GMezpqIBx8lN5wbP59MRLQT69gNxIwK66wtR0sCNUAq9J0hv0iNQ8I
f70bffpjrrmER0nKoVhXKLj5D/VrWUADRCTUzbM82B+88ShTAIAzkv4ftovwdbiQP3SNnbef0Aqo
63termojVHzueL7RN8oNrokBg+0C9JnfKgCZMIYpTxApmZux7JxdBYLZtHX+13ZNke3JJ9PHzsSI
6QnJNvaWrIADqDuEMOnGi3WPfD3tDBAT8vTL2A15GMDmfV3/3/tMggqevAFWw9RGNRhJpb3/zvSt
LW6qRrGqgXd8rzORgeYoTKlhFy8AeYvkp9pzDrkSizz3N1ewhtFjbGb1w1PnlpOg6igVwhAyaUHX
kQR8/GXr3fB5XSXiDNCVB2RF3/SKAv4AcGRBbCb7fMD8b8FQkIimnl0O2L00jXSm2krm1gevBQUy
6Gb23KGEANuNk7bk6vL+zvgNZR7KE83f+K+qgj1+zLLYeBI79mnRcAUXU2e9m/zwpWjXyAwNPlD6
sY/bXhCD+TcOjJKeTKJpxWOFj5pW7qlTjJnAwYcZ6K6VWrt2KMlHRm+8COectcAwxpGrJ9S8VAKU
/t6VQ1cv2cBLohL81ytEz7PdXB6WxaOjktjxU6Vi7XCXDMhfzlYCJpAWHo31L6IJ4+CZ8KId2tiN
aw49IpT3qzABH09+1+uJ21nMDfkcH3dqaz7tfaust09x63qFVhz1lmaf7t/og4KN0544vNjZxEA1
QEDCsC5zwVcqtmnasSwRW+MO2Y9aI07Cti37kjY+SXeCJAcOAh67KMgs/C/37MWxW/tKwt7egLtj
IpHPcsAVSZCHpvmM9g6riZVQT3RI7HMd3magRKgxSYOIahIJuG+W38+Ql5DCQI7eWutRw1zqKnO5
iSy1uBnVECCYFM1BlpBxHx/MWkQ/Pw7eZFv8dWYxKv66WTZIIjnHBUUw6uOWenOJ+2pWiRdDwL1c
JWtQpkrbNcnfiPxe3QH3yZbplk/U5tQdAChyHvE00zVqH66RmH6SgInncj5kU9gsxRxoTiK7s/MV
0z56rf9h6xNDLfNJvTfgky/KGt2KyxEfvSZS0u0Cs9vpNp099bQqcGKOBjmQm8BEfL8oMYtP7eRj
oiuWzKaRs/MJNQ7uSzXn5D4VrR6WF086jW+ybt16hiILcsO55IVT1P7lCQ5NnZX2ZBvwHpDBDgzf
LArY3X9Y+dYV6cNp4akj1JdYu0jbkmli6B52krcrBD8k2cmVpFFhnVuz2NsEjJ+t0cXYtLnpVHqV
YuUg9sgplDei7dTQQe7/cFS1knHDoTJScBitq50UAJrOX91sCveOxkXigV0jtfEw3ngLyfWbbimr
T/U+v+lwmtayMrcisicWVmi58XPT3hhp34xi+8RLCk5b3i4CCQgETRGl677FTrHTRwQBtRFf6wAX
phPA1un8+5IFmndYJK35KFDdclQ0fAeIYynkJ4f5WDOq/4hC6X6bJZkoQN1qnGZoyrCTOHBBVQdX
e2JBVQjDZx+FIR6+QzN7rTMLGCyYGbDvIf1mYCJMlWsn02wRW24GLGHIKCYmJ2US0iA/7jazkMu6
DCwrNx+z4Q3JckYcOYk7hB9HTrYfqod1Ut8aJxamq70s4JQl9mkPAcrNeuzcr44EVkvswA3TfznM
U5nsb8w/uKcC4v+sjsD2KGEP1fmPMR7VYbeyaMohD5NkIgw0S/fuIdBJItCti1wZfeySPQZgtAJ7
8LhFZS73lTT1WXWuZY/qsDtOHpAuyD0hD2JckHfYOsjwthlKB5UtvMqCWw70GCZKZDgfrR1N+Ydq
LyEJg/GdGeKOg9gcBwtGTcjc8z8EMMpSIhAQDG/jvmtbyfUYzkwFFX5ra/X1RzbUvSTBZc9TOf23
9S0VS5zPb0Lcth1EbNtLvWGtuZ9tICSiFipyV3L2a2wcwXLkYepxIeOla1udljNFHMTGw58zFgCi
Nhi709UKViJ92FL4b3JRMybju8In/jvVu9HMZdFRWFuTsdt5+L7Xb1rjT3tKzTHdQRmpSuc6p16x
x2ZJul26txZXIiRagQ92n2XWbun2iAT3f6PxywKDOfr3e37lZL+WuEBFPjCdC+KEUb/aoX4Fgo2k
YwkmM6aG8WLQBI+T4lIFwwoneqvNY3G+xr2DbNP4cJWipIKyW6vNaioU7IvfabeLRYa2dwBH4i2+
W/vye1gbG0nBnnT5lSuVv3faNXRdoa2r9XW6Gu92rnjx3ueDhshjDhvCbL3Z2zlKK29qLZcrCb2v
Teygf2gFoDNMo6u8kXkz3tyuZX+PQ0Q0v6TGKOGQXY+JP6dsuCIHWqVjc3iOXTwURZVZsFO8MVqH
0soC9l+pcmqLuIGScBgSbWjTJ6Fy1P89yGvcLQYBE/tSj0LeY8qGRUPR0KzwmCkce6TJ5LlCcmcb
83jW5QM0UsgLtu7H1GLsAdpYpg+S1Jcj+dgYvLyDkuJfTlRQF1IW9mUwFelkge8v8W4D0nD54/CR
LyqqCk2zVzsabwLxNhxxExiVph58FQ7h4mtNe3Js/CSGMikshpt4B5nGVAmSz8PgVUP1itPQZ6Fl
vJGEip4JrBDFTbeP6vjpQPcvRkLKifqRhWSMZMwiXilMY9RxGK+n+ed2SrFqRSF1Pe3N4Ug7FzyB
PzHmnwAgU03jz/YQInTAJ6IT4G69oOhr6XTSJhC7VlPxEHUVStpqhECAt0Jgg+3gysEKd9UHHmON
Z/yHpwOJuETL/YP403uP5gyja2gVOru5X+CZ+bNpw401bqlH8c9yxIAGUpa/IgBwJYi9omg2ohoI
FRF0oDjbqDXvv4S97GwOjsOOS3iEQ1t3C1Q4c4f0Hcnwy0Xx9SznycHJ5pkmTiKDqwnJLyMVxMTd
wx5Br2/ZM1v59/MxbQTSmBWHDQJQ1d7gFU/J9yOexFSY/Dyo1lr31qvUlt+RU0Loq27bIPAsVzi+
hSP36K6YjQTlYGaCduoS+CWtKSxqpOqXBOe36dL1kVc5hiiSCca+S+8wqU1MRlRfxanofhWk9Qh5
wHgcNAs8kkY5lewof/HeZNG3jj1HaDKFp7hhvq/Rdd+d1D/cFYmFhBgfpKzQp77km3CKx5vtyC4t
VMNyOJ4d4d9CZBEzFGrULcnj1gR6DSBT3dtBsegpQrb/UY3XS6JWyqPRu0KQDgOinpk8ox0uJ0VX
f9xHk+Y+uK0uceWEmEcYoWfjmoQc5zfPDBuf6kXEqVTsOr6S+p/P0R8V/an+FJQu3wpb7EZYJs61
SXOZtK0VQfwJWXFz2XSRa6gF9k/zc5M+MbC1N0KUo8w4gO6lCed69eq4EIqYE+3+TmG8eZDYwJLO
eN5/RhBDxLQsNfJeRYKdOhR96ohFNWC6SSHy93aIEpsdYjXVb56wMag6uxM7WH0J5Z7G5u9//vLh
e22l01G7t+cuIgFnXRDNC0o7lBl52eHvHpcNs+pLLbWtID+XHb8xPZUuBdt7ngFsO1tR2plHncom
vsMUvPHmMSsV0HjID8U5Dm3YkS+igPhFku/XV3fJq+xgXCxu6SAHLfk1JkHPdYfzwJOYifSOV1RI
pGHsBb9LoB8KIFVy5hKepU340txKYLs7Hq+ZNklwAbsHGGdjwt5twzhYeAVOC6hbY3tz0zDHt1J+
59JIkg3QI2EI5tjb3SvcA+J6AwuZdUURfUcZRw6SJZUkf4hzTpynA7VlfJpHqx1WEZHDGBa17T3i
UTU6WNCxHUoyJTuU+ByfA4NLnLT4KYoIzwkkKOn1Vf6G2k+0E9a5asAJM7fKGAnphiYP/bm4BIYe
LEmVEzk8HIjEyjkfw2ej9nA0ljEsl1UBI3s0hCa61pbhC0T/lW5rHYMyuu0hHd1EgKi+vPUmO+w9
0sdffPJc07M+S0BksTTEOXNLnBg1y2a8XHIPv7b7f1IkuLbz16iCjlP5hN8Ub5FRSjO3EtM1YY4o
y6mVi4jVQXTHhU2uzeYpfZi1V0ARYR1a4nHjRvFKHxs+lZvNM7uOsJ4aQ+jjoHEyf1DT0yyqXhCJ
dfi23EGrXT/EXEfFWGSAf13OveSB//9HtujZoBvEVGkCegiaIQ3op2lI/P2bEujpeS9bBc2hdlyU
2kQdab6OI7AyrbTKkKotXctgtKgQOMcBJ4jtEXV/LEQixP6ow0xMun2Q+LVSkE19XOTK+p/iXSer
NbjMo70L2uP+76i8jPXF0+mzPhBuPii3kCoiFjaD/ADiUIP9F/SaFCzy7IneIJ2r/xHZz4CXsjMH
8UUnysWMsTU/g96m+bokLJeebvKjlRbZWSYTSK3Ra3L9SStqvmmoeVmHqNh7SlQlJ4E3hr9PZkap
NclLR/1WXAh6b7khqlpyHYJI0EpyvZuwa5U1RQVHB2F/zCBpMrD9oSW7uCyBH+wEHCc2Maf1BaZ2
MuNn7AFfDwFvz0Z9tlmAJAnr3OG8verMFBAgMtRTvtCFltocN33dmmoqP0tldoqyUaHF1ndALqoG
dJKBDOSvgsgndGnHo/bH2XgsWblAJp54TUyD+lDhVH3+myyeUI/CZn+aJB+bWswUr3hRx6ZlBLAJ
XPM5E0iNdbDTQx6gF3UsAOg3JpND0LYe+y6uLonzpvJO8443XcCi5bnOV/jfqu6l73O/L7qj1ueL
g1JJeIIvO2hr29UjtM/mK0W4LAznQyI8V/MCzcIW7pktCq+kvg3WwSLq+uvnnpO8r9or0WZRWQOt
+nppO+kmHnx0wqOv5PTW+GuZ8bLaoL84Fq31ZNChO/R4xVldaBU9yA3fMj8S7dH2JQ9Fo6Cgfj9h
xCXHgMCsJkyUVLeFrjywGjvu633f7LrzVUE7xSaARwmHRnOymq8tmbyIsq9EEcKKAThYzwMwhgMh
qWcFbcTJEv6c5V9MmERwR1oveiPVdvG6+FfvwiWZqD64k4+jPB3iqC+yQ5e7DrO8mO8q7euDFdyn
4ATEGS6k+om1zEjRb/vsInD+duQ9ykp00YY4j7GSWdzO2pCDO0oLqr2USdva8ZFdNPh+xt8uahL6
UWE+S3FMGkaZhycuhwq//3vUsKvr8L70fyAg2jbJz2da1oYjazRQJZmUDw4SH3ccLF7AgPP289v4
CV1sU7I1sVDFssd32rK+Z+FiGM28R9rlt5i6LD6KHNeZ0aum3fWcwnlZJl/WwI69g/TIi0EZqUGZ
vkxxAd4ADSUhPHcIuthf96tCxP4RoWSJt0THrz1tj2TnlSJ/wo369tYSfQbtCtFhxiwPewIWyP7C
2rCjlTHRbAgSNWdgBxmc/PqK8QJM5RokvAHT1icpxdpaHihEo4xFVjY8HVolQdNxZO+Oe2IWjfL8
z2kwPifdDwhD9Nxw+DC3duLYjjo5j8zpszILZd3jB6fdfYvjKJXUspC+UIuJpz+uCxf4ZbXi0GEX
41xmtHLWWTL9bJPfqehVtzYHyVc+rtiFkBJDAcSfEG4nRZU4KsQY99UCjBiS/GyayfQXV7rCY37t
C5nmmjQNboWke/abPytgwlpxItWygrhb1EL9gpG6pnpBFQtpdncN2eUytPcO0VRKjOPZe9paN5DI
HKx8FyFJLUyGK8MI2aFZw1qzB/KYC0pKs/Nw6ZYkP3V3djU1mKFaKLhD2GFCnoy+UwLOHONFho8T
BZ9jywqXowfVad9KJDA5BI8YYWH+rflpxyV4FptFaS9ilbm0QeCR1SAk3KuZh2O7pL1dcr9cZinp
ERflvwblwx2XhfJRlDK31N2kVG/mzao7fAD28o+t45JlMyGNVibs8IG/vXzkbiefQCumqEpl0XCv
bzkfVEtEdCI//UOTdsMxcmNeLi3JVbO3R0Q7uvniYaHVsXYv7aPVc0ChJsk4Hmgt3hPZz9FtN6nr
8JtATnCYbPB+9R4SnEVyU/xCvpW0WgRuvRLnRUqsRzb3U5taogap7541dGbeNn/EL4N7hX9QvsGS
wpreBHpsZDIXAXcPUDKdud7xnNB4wJgkOL6MxPBSJLAvODP8TFrbQB8V0Krsh/tIDUcxYEkfa+6r
kP+mAYVou0C7rhueMTBCgpbA+5yFXnlj77FnOOmyRyxPumVM0Ui8j3iLpek6XiPw9P16PzsKE243
HOV2XtVLu+P7h6urMrHaYO8mJYwdQazv08f0vwIqhsydTLRbT1zEDQS+LmEZ9ppojjr714D4V3OD
b29sIelnRASnlUPYCKBTI0ckO82GVIIf3NZgWrk3wBZc6eXMgPm35hI+/7xkn1jZPmy4HnIQzh2N
TN7UQA78MtwdgVqM7snNuvOm7B2r7SxkeL8VteGQxyKIMRPI6YEyGHbeuJxRJovc1FzxOmAD7vyM
fYejaPCVJcAIi1buPGPyo8T2o4dWrOxNJzvOpw7A8J4zkDoTh0Tx3P770l0tx5wAs9v+8kNdJQt+
LzeV7K6w7zcNlAeacjDMK+Snw6YRhGgPrmU4TsVq1M0ORi25rt5NOxncuDJ8tX/k0k3/KQsuWhqo
SL2v2qZvylXkoPMqzTpDJdzlNRcmKv5WqMrd1DaskAF4E+zCeZGGhYdVjfEBm4ZjVt7aQOkHhA8X
4qbaIRggXJDWE3flUrdrk7G443rZ+YWM0qR6H6GgUKvVf5ezGVYRMW8mx1VB2LHUzEfTiPFcAwTs
1v9FkTcrb2+TlGM7m7HvmZlxnsRPJmgHtZ6Uabtz2rFEnmv3VIHjEn9JbQrb76sL511UT2HT0i/M
i4KJCxwxYqRPJVtHTqrm7SYbpD7R7+Q8fUeMIKzVfD0mmTrgP9nTk2rO+TXL+WuGikkXhpfTPd7Z
AIr3/goB1HPQXL7Lea5vvJqt1o1H2XNmerfh9KfA2zgjBr7m4Ch+oB0ePtXMyMksX0ykTDkea7qz
Umxo0autxGrYMyOLR8PUOWyxi6AnfAXJnS/iVmV+DNKWh8SSkuTixVlThFHgREhCDuilvjtoqhVp
YalPKy4ecKLbVus7MkMkIHmL+49+X0OBDL/CC1ONPPX1OGBHxGR3CjgwXigvFnIQGkGVtCAF7dDw
eY8VMKdS6QcoDxB68+GIiZrVu7ZQ+MaCFUN6BNe52vQrIjCo12bApue3nLpNs+Y8oyfRew6k3Yld
zVULecLH5Lp94B/KwKTtNxjjeIZsvI6Q3H/n6cYHbuRpDAESPTcTJda+QMLfZMOG6tub9G/3cTfN
Q83Qj09j5tkHwZPDjPeSTn4cDybD5zg6uPZP0fnQLxNgyS7/he0GB/EXVHl/Z4akoG+9OxV/w76z
5C0njwkSDA==
`protect end_protected

