

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DKaw2YF5X/sI0l9aLdTgbK/M5GUdtEMTnIFmxvSMohXCNpaRunL9ipaA59Dc71YrenIGtec5QT4M
zCoGKmFbyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QRHRuF+/6jbJdc98CuDuU1RSPkw4Mrd2rWInSv90clZq9I1OTAA5/xdv3Hk99Vg2prXDV3YjNqoB
pcpnTJxql+YZ6VAzN0qCk+oUeO1cCu3qiinofcBjVXCdgYxomUKUeE7FJeYz3Js2G/kJGoeHFW9U
+zAl6jadwyF9Jbvv+i4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lb7wQIOJLuT7MorOQ8eHbXO7nLYJ4w6DRb/CRc0KXgD29tV/pKu8nH2e+iVICJbGwJJtQ3k8P1j/
LscOU8Hk23tTbvsi/KP4jYIAhUNpSlUfm6H0KJ2yht05tm7/nGOSq+YwUD5ni46LH6TZmw9wRjLo
RAHSpBohLboc3y/hVTXta9kQmKPnqAmdZWZqkVyyS5o93+63/fdqbFaxxtwx1mXeZDQ2+2zbTCKf
tbrO065IQsNhLqpQ6GmWS0y4Yk762FiY/PW8xLoCZ1V1Fh8ocFk7LKyATUlQjo3T4vsNks0JLfh6
k4wW0gpjLf86zBHim396ye0D0jCoECOhPpGtaQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZXacKhqAwgw8zLrWO0Oej9oQ1uNqsfSW24Ju9AdSqiO9hJgeX3QSs/Auka01BXmxZF02hREfAK/G
6uXtwOuytUDW3C0vu69znjuzfKa65iqAvitXfuV2wV2SBDUohxstI576S9cHfGPfoJ7tVzjIg2t8
+fXxMYGWVW/hL5Dt3LeBc+ul5BEG9/vwugVmMP2uMG9nGEtDEQeLb7bWAsdsP6jyz5L4K49swiWc
6TrDCW/53r7o1y18s7qcumMrH+8e09lZWlV7gV/qSGCmNFjNoXkvbq7X5+RT29nF6kaEY/1Y1wcM
sqDv/0rI3Yh5PZatD+o2YnHnz7Es16C87EBZrw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pkb010SLYsAhKXcWm+QlAA9Be33Kx3pWG3KQ8c4OXZxiNI+ziOzdNGDZkUALVJhYeeODAczIsICK
xPobg5BZJdmnFjXMkYzJiVNc7H8OtQ+xwCOlZfGQy0nG30bs3aCt+0ciZZz0ed8EJ3QfOUNUrA8S
ACDctQvzk535zqal7JGqVOcbax0rksASegZXl9TYHMAWSFXsQNDtHG7HCq8QaEGySiiJnEz1Zygi
CXmAaOXrSZ/75eRU/jV0Zmfl2uX9M3RD4WyT2L0mtTPVI1Jo5riNKDciMqi09G5yCgGBizlVK0Le
ynsKW0Fvo5j+TrmGuES2+DcsvwzxQUmrQ9n9YA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
saU9xQVocYCNVhmm+/jaIKt7f7lGDiBCwD7GUeN8jk+fV3dDx7VH8BXnwqh3bO2UtgQTq4TYazR5
PsEJU9lk5Y+2uIztywixaUOcY0t6PGvi6DZ5S1UapcNaqz1GzVDJNMdFrGWeodfXgyVpIeng6Jtk
EKceFNW0p1SgbLjlCjU=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pbTosJ4LwLIDFDsIbDQWyryoCwFpua23V6z9HaJa95eQ/VgCaYwQRc0pJmp/UgRFI8GxRIcCfLjR
nDQiDTQUzYsgXuFi39wSqyum1ybk+zJc/c0tfa3zo7fAh7WEKBR6EfegxJoOfQ6umn8yMUOq35ku
5cQGVgAH0mV2j7kgcszzSTcMNu1shLKlPJejpCdXAsAct77F4/JiYgr35R62Nw5TiOPHxLGWKlD0
S4rOzGqDzYI4jb5eYbnrBMtpHWXse9ybFZPj47SvpsioKcFIHeUE7GrNOvNDQPdNPahScNll6gSb
fa6tuXH+3Q3DQNGg7RW23POGEp2w+WE6Kef4qQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
gX/gXFWLvKIaWicHHwOVelTJNYGD6JUfgY9YEz9DRRjJWsrfB36akg730sAcPvv15V8OrATXjDGK
0qBSXGFkEQ7WV3eJZxe49/yc7CyWnJe6wmD5YDa9BPFHQ5sGt19ie5Ey/zpikFtjTIU83geZieS/
yFl6nqEUo36sZ9NDaeG5Wh2ID8ka/LIam960u+LZ7E7kfZPuCdAdBSNpwls0X+BUY7Bgbvc6+W0u
Q3HZ+I95C4X+TU3ow9Hq0PC1EOc64K+V6vjKps+2IbDO5gMcGCrq65KQ7F2g5G27IGbzT4/OWmD6
VTYBmkFhLiW4zRn6z9aOIVDaxWhrG/0kZ8u/N2kqkIT1nrhDmTjSx0BtMDgs/oe+FJK8zQ+hPjZj
wYNrETrSeS8Wg9Ont7OAznUB9novBq+cIw9Np/aq3fA0aqSia9KIX4FKZUuv76TaJhGGX6X17mea
VaYNUU80/2h3UDzZGyxYWpaNHOBCqkGahDfJkL4J5MnUD12QImPEJ37aFyvGwB0GvTzyW+jXJv54
VRZsemBbYWehfFM7nbijZS4FI/bxC2bRBnFJlwISECJ5aZ1ok9z6/gk8QkCjcn7Aj5HBVUkh6RB2
f/p5eszFTU/6UDTIz98hJ+xrPXOsqlG1hIDzy/N+sKYNFPP8xVpywsGI3WmsbfoB6ysgtnQEj06f
HWVNA13WViLIuIg+4+1rwpz5+VYoeYYIYKTcLTUrYn1E/7OAMF3dGx9OBaDNH+4SUXhL0IbBQWb2
hqSC8biFSLluW1pggYFaFjoFDsGY80Qfkd+HgknuSi198JxCsgbhdJhQfR4dghwsg/TpiC5DErLo
T5FPqCe7orhaksuoRcu2xzWUfqOpmFE+9gRj2FwCSTZ8N6n/i8e6k0u4TsXmLnhjAGchpiahbe3j
WUhQ3vu/WhLxWZ0W5GYdfJ1rVv9gTEOUJWK2s/Klym091WbIkt5sxAo+FuJnNcomVUI622AQnWvM
75WiXP+QODoMGN8YQUyn4jl63NQAVmyHmrPNHrokKAbLrJRBOaBRHr2cb3hhekQpC1wyIvf1cjk3
+zTV5ngGgV4PeFQYPpQJ2P4u0YJ7MCYTqu9s1UaekDmCbWtWA4L0/0V8i9vQoVfSPAjH0omFB9/z
5cbEACXEcsI/cZju9AU2NwfvvVcEWXoyZ6vhe2Ffcv4bewkEJzomHQaLiwjVjpscHgKj3EgUCO+Q
360pIMEwRQQCiFLmV//EbxVHre+24OHDZObs84XV6EIqi4In2M/iafTf/J2xfYyhtmhhBDtpqwyM
SyWN1Pr2NUdmKLQbRswKx1MeLQngLBoRpY3FP1PQrBA9KxESOVpElsoM3JbxAnfxz2S3M8/YLAOD
0xCEz9rTj+Xw1LEMcNUl91ZByfDFJ+wNk7SInEqLW9gRgdoXM5Rm9g6WDOwyXFVpPZ3vtyugqQLq
F84aWXWplQiovqeShpgxc7I/nH9MSR0gf5kB3kLPHNPwMRtK9g1pffx1VCHpqRj1FMinr+wPzuao
2ZR4xGIBKNqwdoNkH6MKCi7R4wFohiYbaZbAGMiJduZrjrxxIWKvxUHYNcpINKNNG7QY1EIn6Kcy
pZ7U/G8V3gdBfW99+xmOicEFnbSchwdTOQ/23vGmYB3PSmMzNCmkfflPXIaJlGp8F+hAXqBXxW+p
nfWEtGJpZRbUhly78g1VukVWIN67yBG86RF9gI2zS7TIt5kIZZVNMCEQuEx/eoLOaQvHpNL3gSUW
GFvEpyNWnYxPRS1a7drBZzjCykm1ZQ5yrtWSWFWXFQktv8FTlgRhxne8pID4x3gegco+mJAhgWO6
Nq+M2YU+irw4uGVHdZ788CDl9V09zEpofeFNaBf/Sgc3L5wP1Tp8mIuCrrPgJHEXx+1rFO8kVzSw
bJykdw97H+HKtaeJeZdoPJloLM672rJUHsW8AH1IZ2xViW2y907KdesI0uLDsajzKqdswSxmskAN
XiEd2sgZs8gyOpd5md97JNt135XT2iIOaDptL/7P3UdjwFiexrTxs59IvoFpMas76Pejv0P8Ye+Z
Gd4SHr93qfEHKStBZwiqxP4+THuHYhnzbnO/IRuh3dfgrHtgawc/qD0PkXk8Ru/sYJPiwmgcbh1Y
e5s+1vj91gnHUUupatr/XINeGSK8kEOyn/MRx4rzvJkOPvB9FI1reQgjM508HV0wjnRkUvnrSme2
UAAWQK0sHN+hO6PoqLdWogvV5nqmbwVW1/dJqPrR7G8g84l2arnRKKnDwCb5S9kZdejsRVzKxkvb
Gv7sOa0KZO1Uli6rJtCgK3K4XF1K9LdoDgpR+L+OFFQRCPnH4dV4Mk8q9HBMqLVR0gXWOthOUcpj
zXmAVldnJWwod78C4lmKUg7LYog68C1Lr2rswsarcXEiUuOxEzzPPo8aO1DtTTosBJfq9vCL98AS
HlrAYlw2ZKr9kMB/XJFP5PLuWJNFR550XJTUVNIMnRS/lzY/Zj6PR7twURCTQ7831nK/bqzHA6K1
AeKuKADLciCQk/jctFmkG7Yx/FeEoY/UHAzk+5NQY7Lx+E6Y6bYfYpQXqc/udUP6fuhTBZArUgj9
WFR2R5zZ8/F9p0kqKkJY/alu25iNOVUaRuS6S5Ra7CFeeuAuxuEiravTyUssZd4ZoBk5DWH62mce
cHKBOSW0mdAlJdWjI22Ty3FwzTPYEg0sxOIdxhV+V3p8jD85t0LSnr0QlESb+LrzD1I6yinnrTGg
mvi22UoF6ZWsRLnSgx3LPhrieQUuen5TcfN3APl9Q1tiNbtLNJYV0rvyXBxXR02tTzQZSjq1ImVy
w4w1lBZe0QtoGlIJjWcRnstKlikTtM2xWHU0JX8ErGpOi2i2BEkxs9Ls2tlDs6fjsThMU7J7PD0Q
P0fJUvpfUQjkj5w7ou2Zub0jk6RYeTh01DxJCrDxS+l7f85BsdLbyBWfeh/eOUgxBJHeg+4fnxd1
o/D2Xn4J6MsEO2DpcT5n7P/VYKkkqVc1sJ6xnp8N7NW5q5/qWGt4av+xAO4s7ELU8kCY8wcYOsF7
sT4UWIeVmMh0zf5StIqJdEEWk3Hj/I1l3e1F4kdTSKugmCALg6CTMaAPjAHksPQW349ZcyqWXXyR
whh9Bk4Sos6xCb5dwx+b7uQnmTP/zlIr0jQWxwBx2NNJPYfEI6yrgsHP4J1BUMIOl7a/+sPITXY4
IdNg1bMkieAfsRHMyQisJ9ig0Q9W3Lz7llScu9Y3uqs/oVQrJyf4Sp5wbSf2q6jNW2rZ/Khu4KnA
+ibuKkgCQPdDVH2nH+k/Fh1fHTql+DI13MPXZBOrjf49RUXIxOHzesRJ+aAewhjB3LshXgz9ZBOh
dHnYuYw1h+o5Ukixs6ov5pHTU2PCEjV+ELwLV9m8CVa7QewsPXg7V9BUokZvV3RLgsSAcpmEhbut
rNkkzXQ2KdY6P6rqOxXProU4cSTU06XJvZs8uunSbG6pLBouErN2IBbT0B4Zf89y+b2VKXuS56Sp
hKNLAlnvR8CyDpN7N/r3pjNiEVEq3qA37SLeWKW/pDgDAxQ+LuD4ih8HSqBBRoqHV0venY6LhBxa
U2/yZo4Tzm68H8vxBRbAt/54mTHFWwANYQ7P01ypO7P2PNyjYi28FbtToTUBLXZo7N/iSo/tNX2G
yVF0LaLD85062BTqBkEgCvVaT87LbiDtq1c2ZtEVfaK59/kHR2YpZD/Dsp/126YDQ9cxni7Kdbgj
2MyRiONtgexAvsPnkiUZrTmbRjUrPKqeZX6162imvUynkB15GTMBrbT7CDxhO3+K1V0EXIp057gn
2+CRZyNs6wdM0BEX5hsWpm6OQ/96ZeuSLznAq2T70ex4kiONDkTMEc2G9kVnBAhwFAmyW8yq95w3
nl0msWCRJywd8G8wtYyaWQnHMmNUnJSjgiEJgdCCXf4NGeNqXI4UFTUi9SyJNqGDVC+mqpSRDFWz
FHdORAQgTtZv6khdLkFkdqli6je9qx5YfAjVkwF/MQzW1YF6RbMYEvAC7zcaeGWGNy92GkjKWTuT
dVjK9CX74D3GJ2C3Q9HvlauhpJjX6Bhk2ySwfS5SEfSC0XJ9/UOfGsUixqVd+aShETqMFqECZ7y2
zic3r57MDnfeXfwoKQsnViIIWGPH0LOXdnjx/F9ZXTsBLsd29nWkaeiiyypo0WAkzvjW8ARJmTtt
2Ww4QqQRGVP5+prXmjupEjc/e13N4dtAUqmqx2g2RjnaJwlbOnYI9eTwCiXIUP6FVOKcI7RUBpP0
jQD+3zYbeDTp7QHZt7frMWP7XyiOqr6NLrHC4VM1tkMzkTfurYuqmvFWFvg3xGj3PXBlXPsO+7Lq
R45Z8KSOGoOV/7Nt56P9AqN5rL9ruvcEtnc8mZekXJ2mwhPSYjrkrsGh2pOLp5Xt+1fncuRk+7VS
D9FEAw/8CDa7qNnbTyv3ZZWDfk1U1Sr+I0g8WxwbNO+mcyay2XYOQ9YeVnVaN6SUWAxVOON4hu/L
s6T1aHIc+3ZKRVw1xgtgy3DbZsn1yytm6xfv4ojMi0ztHi92f9OGbME775eDlNiebsYuHdk9Za55
wC2QsvmLX8f0G1O/XZr5aw8ejJ0Gg4xfD7T1ZdOc0l9bLx5R7kt9aSmfTXaJV7Wt0uECAO8yzHyO
rUB4PiS3E3KJEIHHe3zKPo7t21HK6iBsUSVtJQriuDD4I+87WsnN52HjGoml3T0r2BWI7aFXhZZ9
8eaXZn4Y1Ny2EMhKF09CIEhYIi9H8QxRJmn0mMv7O7ZeBCJcbF4R6/xcE1KyQdwqX54MVJLOe6RL
BZNCMspNumysvAyXx2iNjfHXbkpLH8H9luMf8IbsWFM4EyJpyN9j4HCK6cipcTxBrg5Ez1af4Af1
bfaT8Xj3PstzG3+svq/ToZX360tfqNVnIUGdonNdoTKhOQpuGsMVTsNBmVCr0AsDOvyF2eLa/E8h
FOFovoXR9MPBtXrqIIJXOH3917+fHVHPjAD5Xh/4synenNB98nwf5A2J7bnPdJV0vfbOz7FNCnlt
5oXgcegZaAAMKH3J/XaPEKIeAN4WYFKjNuVL0ZIuxC41GVhYzRti0SwwkKzbhliUVNxM+31OhjKE
QKDzASR9uZibAW0+I6PvGQ5tu2rg1QUxfwi912ojoEmOxltefbZF8wwc2QmntxX19iy9lLeepJLa
BycDdHhkJt62rnlr2cjVE7QOtLilz9mQPe75s6rNOKeqDlfBuLIhl8On27FgCJk3O8BQeiuY3QmK
Y44w2VpYGzvX7PuW4RB0v8zuKBJpb0j5w2kvmDVI8vCqxvrur3lDrncZbhziAdioNGtpsbWJmPQI
LYJI9M+aeqsN3ASHqnaVk4neVojNJqOKK0WFUz7Y2NoTEzftw5yajxLJ7GDyp0vc/uhrAODG11wY
elcWjW/vO76tEsI1nLjzDG/NzuuNu92gg0KTNh0DLLfyCV3xOXUkkvb3VOIgPf+XNyU+I9XqoNvq
ZIbxqeId71IGfm35NFDYtimNeHDiVNi9w1UUOqhL6KxkaBriEdisNd3ckPFxxRlxTfaRqnEe6gl4
hgS2lTZEobeu/3RvvpRm1iQoApjX8amtJmQ41+axzaIHrBTzNNe/nRV4Ck1AYJuBHOfnyoUO2UQq
aOxV3xI0FTN7HmKQdOeV91oDKp7jWnriasgehfhxXED1Qx1S29enR0xfJCAljoRs0IBVOBmWG4bz
wixohV9CtiitJS10xXNXzTiRKffu/wB/NbhkOmdFErhvHYlXup5KuF/feRsbCJiv72gPUsFdI8Cl
BMtsxy4BAq2K5EzRdc95fu69F/UP54glMsCy9hq5FrEqxlozlRYlR0OKLxYwnAiFdF9M6PG2fS82
w3hODwCJrT6MKX157dstly4NK9WGBGuxQrQ/Bxhdig/nUZZbN9d9gtFgYRhBdFAaiA6UXOvj+PHV
Ml8YgcYJmqtxsS5lSITPoiATllwxOjyKcW5ER670iEAJFFr7ipyA+CHEmSc1KOFAGhneG8CGsHqI
EZmyADsmkGaJzw6RY+8kp2GfTylNvSWtExopwXZyU5k6P8g0GvJcYqZGpnVprHmWSsjaWCx0MVr/
xuYeFE99h/76G3bS8wYEsFfNNfi6nggY37ox9SwLZ5pB9i/iRm5fAfMbjw5IGa/LkNMJHYFm7FPK
4XrGaDLRhBiB7ScrGV+TkTj7MxJKjmqdyRJ/Ato1tN8eEoEM5sweGjqngrqfgX6GtkppIfn3AyFN
Y7pbxUinfC82xZ/VhuSuhFpX2WVyiJsihnrptPp/EBpv/TZQ+4ymKiItupX+karJoFkb3EC0AQ+X
CogFcaZLvsaRkkAbNQYA26wWUqgRVtOilRwzZULzDq8C6xKN1FSRguxcDxhtFsHd2MYpQxJPDDtn
9A+1I8agMkkg/2seO14c0N6hBXDsv5dB4gUon9RBhqSpoIcUE/bPEKjLn6xrpua/sylcxEblQncM
ZWWx/W4gjDYzJS4tINgBWu1Ua5IxRfh6kubRhB5rIk67ccM5L6qmlEQe9aGxqtgqYcjwOco1wkEh
wVSd7ILt0rMcko/g8OJzaV+8fw1VGBzpY/fEdwyzy4scYoRvX4S9TByf8cQ/y3TheNjKsR+QSs0L
f8pS1Ac7oS47DGln2SYXL+KyALzfnHqohlCwWlZEaIKXcap/p4QU6zpvz+WqXUZ+PcbI/BUkh55G
s/BtnGDn5708+KMSGyjGM7o/9dxmp2Dfqya2GgtSZK2w8kDNF9HA5J5oCCHDTDNuuPveIrFyEmju
3tEorXpT1ijAPPu2H6N5D3MAB/WtdoJ9Biy0DJePkJP/54TNivgVykw6H3A/H0WMShhyz50tThxq
q4BgzHk6uac1B4V67AuknZCk6k9ky8Jcc8vnGPADEdL5m1Syy6ZteiJcJ1ecRBLMAzYzHWlVSfDO
UQrt5N3/wfqOAZC4VUGmSGbeJcX8CI4DTI3msGhs5EaRWevtQaVk4w18s15bUlpzaptvqjLpcGJC
2o3Lk2PVsWl8Yznwce4DoxXIcaWJuy170w2zXo1/V7iXsFw8LZwXMyaTSqTCwHiw5z10UABCAz6K
d55DMO8nf7tuE2wTXxpvo93SCbRMWaE1pliW/DQWb7j01tHXUfYl5aZl6Mn4tZdbfIxZzBy4iw3m
yp3R1SmjcI2yeNmDIAIQF9qsoU8+hXLcnpUW8hEvlMcPzrOnJ5d502otRhxvl6jn1yu5FSMa498z
N+GS3t0A6HlonR8JcS2RLAZwu4Y9C0sRDKOkX6iEwKIWY4imfS0FCNemtPE+29qsrirBWEn5nqG7
NOCjsFL8riNB0GQgBn3+zuIbOJE8lDkIUVdh10TaFraDn0wJRg8jddtpPghBLSq1o+4gGVCSVu62
15XMq0jhEBMP/nC3kZCAV9FuSKDAX9BALcRdYcxHKg29e0TN9tTDmUDycCEaSW4kUulxC2ou9Oy6
7oKjOBfz37GTqhOFwvGyEtM28xz/sym775WvSJXkANjPrSnzuNF+ENeVTaccpmFFU4KKfKby+GwL
dL4za1LRCG2LDl7LEmP7F8v8nr9S4i2FW32dImjyZr1uqcEC3LkYVm2xHV1X111UQbTPEP8iPTf8
jWmeBFsSmrkJ4uxvV4U5L4Siy8ElTLNkETrtqK8AYtdkxOGUs5wTbbhojtdd1ythn8/0KjpnMVMw
dS5EDkodcbDZ0NDllp/PG3Jf7fL2TqKux/ASxd7vHDiGeDvk/w7364P/JtwLr73V/JzflseNOTOl
Ubmy5eqf/2Pbyh4r3opguEMUrD9U7pP12p9gMs8fVS0BCWvqDRcVvE3pPK0laedDk1E7b3PMrRno
x8gDSd/vCbIGP+8L5M0uPZ3IFDt1bULEWmEKjyV3YoqZ/RSTq2Ca2KW7rMPxcN0R+aJXstoJnRpc
8NaghIqAD+TyEFzRV89B0dz+Lamlqx22i5IPpFskj3tlX0B+bPvzvKXUuWw0Tww7wHI449r+GQrx
3DB9p/ESiGsKibAoAIu3lvTUZm6j6j5ubBhurSIpm4Hehr+w6W1ptQMBzlA6/4Af4PaOcL/Q2Rgv
AJgmyLXvNBwedHWpPv43o4AMWNq9pjtPXW8ylNEYpq7zejGfxWxjXY0hzwLavug0FW2ZZtAh/9md
Tzc9OHzYiysfLfN5OcGjYm6yAOpmsR9BzARVnACeJdpR5GxV/3PryXEL1YtlCIsEeMDdH4W00hIA
2ZGitv3e+LmiZsDdWpsuUirxNjY+Vnyarm5vtTjNwBO7r83bhvca6sca869+jvowXtOk3edNMJA1
NLZjCdA1LJm957UCDm7HDQhNIq8/GFVcGcgeBRHWHzetsYWdg+TKPSnx8M2X6LruF/4RssLAj2Es
WS8viEwGwFtohOJJTGYFirbrz7rIX/03o8c4PzhhKVT+fX/lTx0crI318qyQ1j4iSbMdVyw5yoBN
JJ8WVxfu95sLXn9bA+u0HAAqqCE/MRCH0IZs+k3VcrBuh95hZjEJGHW2aGqJ6KM1DBke5PBN/636
oIdcusCBmz7v6bkAFtW7UlRtLkjx5GgpxJkh2pXoWWWuWoHtN+CQUqHA6X6nbTqP6zdV2NhfsKr7
lXxVeuwRgbpO1R1MxYIZm/+Ihy7OSP6k2HgGuG64+87/JAoDTaj96vtvmhr3DMtFpRvIQ61UT2jb
5QF2QAdQdPCnI1J4PD1a+fT4cbS8zwrz57vCAQbBQnWuGyAOgLA+15//M5ph7Y+QxjNdTExW9vtC
IvEasqmXxlxiWyb5BxKamvL1yFw6t7xEffOoZgVsm09lXkI3c19yJZHsfB+psZxeiU+c/wImmXtN
ulfjPICQNcuc4CkNWwTZRczncTWdiZXY6+H9wCHeASjgRO2jIMBpn/17Y7PQ0+Ce3Mbm9PPYo+1c
ROTie9rn0z3+j1NbqwTT1kzv1//xH4T7xvMhNhDrf6CMkGdk6IqXrY5Y6go5ZPn4Rb+CNl6wAHDC
6k40wuxeA7Pup15HrmJw3c579SXFaM31x20nuf11wqs3IXw2k5JajIupGIxx9Y4lNnA16YiY/1Uv
myXAEUCyYBi+H3tJSCOqo2xf/uO/rKUCBgWtTDXJjjTSAyq/ikfr2Ve5P4DZpc8p796OkxsIzZTA
VgpwUY07SRtAsK5+WCsBqQ9KV0xK0BPXJ3AKVTgpRAnFHZpLkeycvRXm/XfK3lHX7bo1rgw1VwqY
zYaV5Ut6JldGyZqCbYIjnIA4hZ0RZW5nEUyFma07LNe01TkbYqndUxeqbXDI4hAs/FOSTxQbiw10
S7tcE5dcF2RtwTdNY2kHshIWlwBeGYpS7SMs0ZXbPEZlM3sdSGy/ww3cVOiO08NNGG+n1BwyT1hC
9WWu7u06kNLIdG+YG+aWHjuvbZGWV0RAzY1Dnai78a/0yxj62llkW4RJgcXOBvg9WmMXdUjZN0/4
/+vhcNJcLQpBf5o/4YmCnOrPsVQcQC7G/IU+s0STS2DTEIyE69aJGPu3le3tiA0buC63xAy4sPfO
HK5epefSYuStiOxy6HVuxfG+DXvCKzAcjjjlcEErt4aSUO8qgoQm2hSSlnarLYe3gFbyURJlT5ru
xaFnJjL4rQnO36VlIw41ind76vqowWeKM8TCjoLG0PKVnFDU1wyChBlEm0Al0wxVqMP6EEEruLC/
jL+FAkkE4bTSBnGHuIIKcanUMarnqwn27RoZsOmR9muVPRXWUfJtIFGFPgCvscYkGiw21brjqLFx
YcfUhXVjnKzPIISTXlaV5rI4f6p2L8Qs7zyzAVD/VyKpB9h+KTv3zwjZ9pxKnPMXe8RsR4Mi/qaX
2fxgjJE1b7epW00BA1AUL9/bXJKvVtFQeuSVPDJUqeQntT2lB195MovrKpe1TTRU44E4/CllyBRc
igdXlhqxy0DFyvZ0PVaYnUkakvlLm9qIS69GM7Ud0K1UugznkLn2//Ta9p+Op/6Wdk6s3Ldf1aoL
FLRt0/+SNrGQ21IHpZcFKZM/KXQUNo87RKCesTVsdQNxIpuLjmAcxByviaeX10tGclc/x57QPNG7
w6jD3cZsurljeL2Fg0h/19hC2mR3fuBx+/D2pU8NzxsIJY9NyjzvbjHhVXyPEJBtt25pPL66xl/K
nNp3RyndfC39iheok/95XmyzNUiXCy/OITXDj1jCK+nHYW7AQ8z+ZCzmxJDIqyQYCQBxWBcX44a1
58UTjHlOi7eMGd74XU1FdfQ2lbw9V/jb6tO7tx+XhWDc2JcpXlGp5V0Fh4YWmVoGhKkvo2n1WRJY
Hlv1PMtF9l7d62GLFRrWM5eB/djdDSxMpDyHCXevG2qlAYnlcsSwW37e+DtpX07+V4ghbHbMEhV/
pjwirBv9qZT2xlC0O+1xDUHMV23+VcaqOPYxQG1pj7RMqBqkiK6zgxog5XYv4wRQPRH1A6m2zvVw
TVPI52q+D5i2ptZwxoeAjzUufeUo5kCIbtqOitmyUHiB5Oz7qp1wYdr7TRUzlhiHgN2j6/qpW54F
6xYgkA9mKX+X4/zlekfEpq3tuVTSrVexJHJmyr35i4oVd9RuokD+Gd0XdQM3TuNC8NxDXx/2lARi
5HUOaSvgvKT/UDwMtaWeYHHJReY5FXVaQaw7Io4GER7HZSpctdW6ku6/TKYp7w8+RF3NbX9fMHna
eFpyTvBZ/wL4/JJoWg4YIMtplvrcHfyWMXOZI8EOC/9UXYNCiT2Bwk+jTW7Srqt5a2jyI+FZvEx4
e7U1rutjEFWYsP4HwtyHYQt0XOb349AhvfZSlTKpFnbR84SqW0IAfzy+b9KZOoFXqJDh8INdDGL4
5TxASfGJPTFXgc7DY7vKTShO4TpNUSn1SYM09eRM3nWxHDmVGfAEcgyZ+dtL7tt0mGI+U8UA/9UP
KuPYgF65h6/RWwDdqPD6QVfBd3ZPCW6aGp9AMdJuWad2HSWQdeAMIp/vMc1CIPp11GjvDhZV/COD
mOTRf0ghg2OUipc16AI0HrkhR9Zpn1nCNYmSG1PQSZfCUbQTuQ3VYO8EMRDvs3Hmi8+lQ8X7xjlX
fgwIB60McOJSl0RlIdBGIjD6zd/TE7NAOX/jdGXX+Cpq8PbwzTplB9UIG1kSVEuezuyBrMy+xr8g
kwfBY41Sf9INO6tedI2CPpNClsxw9sPaSwRF0JLwGUByUtX8ZpdmvSG4GYKji6JOYkHFWNpU4VHj
5GUVqci/bfJVeG6EcXO/ChQuu4y6bkNg8N3rCmyhYjUmDssrD0jcM55+MeXJh6uyrxM27NCXNWzB
xVFks5H3KeQEC7166K1tJ5Vbe+gcrTZ5HyhPO8m/88dFsDfU8SrLai/SSZyY4nsT5bKgdzBp38Uy
wBmXy0qqLhzbTk5jxhkKJuVBoK3rjvoqL7ukhmdA+xUDmUJz8OR+gk27RE0idAcXv4xd6SndyEdM
HzLgidVqVlpBXuSQ7UZA1CGBMK/QNpgfsfE8xpifIoryjFvxfpZzrHwVkjnFYq7ivD41aJLy9hzY
l99BO8p3q2ByoSZkhvrW2BlYwGkcvEqnlNe0v5SYZpsodVus9kmZvddV9rSqt0JNNTHKJioKnDvP
1Gyf1rHM5LJiQeMRWJ5tj+7N9djSIwgwi33UnVe3JbVlARHN4Zbx1mOAgdAxRl4H+EeTMGivygyk
VmqTeB3I0sGqv91UJlPtDhrLeIha3qYKwePBXjcq5tJ/LOFXQfrzX/FmsQm6CEpVC+k2iYkqVE0e
pO3WRzgle5J5aa2dDNaJIrCMlnXQQsJ+wGV+S32EtpZGNzekCcTHqet2Syk0o97JQ7FfsHgUBJgn
/i5aSD2r7XIRGDa8rJCPppYLVAkZ8qBHQmKAxtHcF4X06U2l7imrY7O9aVS7qu/IOaiWbGQbgMCx
LfaWRwh/Nw/z1zlNzEuKlnC19WdASRI1BAivitcfD48Oqjv9dM1VbLORLmKjffqtUoMTwa5aTvf3
Hu5hkCDcSm0yHwgrWk/bIt1C/OXzbMqmqLp8wNmq+N7mYalLNv0pmJA8RA/kwR/4DEbWLo8T1neQ
4eI4twTwY30B1mU4jmBGoMcWaQC5bS0WPYLpjpFzD1AlHWr5SHKQTvorLL8QC7PdriFfCixvwPNa
iR/C/PHqOL15vo8u4YngBI4KPjKJebeRcbf/SMAUgzIOxqKBqk2EWJT8MvtXohUvIlbN19NKvpfp
uggPj9ebjxwrGUC1NyUWGEbcbaxoxjy8jbUWFdlB2F+URWP7J/O2iDAaUTsaoM3Z2xqnEDxpY3se
3+8t1BmwPvpknlLrWaqp4fYTBADVdSjjXJZ+vbvHtvpSC771pStrX9m0oERFk+ef6CUD6qSfl/Ul
QHcdd0Gw2HQB9f6a/CCscpb9NGe9AUK75SYAJgVA5l0Ms6pUlI8wop7kZOcA72YACo85h9gZov2+
OKZE6fHfaIF7QSR2EieQhq/ww7KqVdUaG1wQD+PO4UtW2Ehfj/v1Oz/5gfUfLc93TSwNHynsmgP/
Kr6Sewb/6CUrzmkAhxoU2N+TC3P/qf+7hNi+R3yCvxoMqpADQ+Bs9/6fs+sTSX/5ZFP7E1XiYwSF
fH3LAnvhDke2RrGTnuKnpcggtutfpEO5SfT//Zp8tl6g2Jin2EQENSmB2lOwXkKVMgbaSD3SQBj0
cbRymTzdc7P2TSTPFnT4dHj9Yac8Y39tFBhslbxBaB30PQhexkZ/m9Qo+sFth0AqGz/dkm89F0Z/
tTgExCiQn93VlgAw861iAB3l2TfmU8N9svNaYCYL0gFqupGwmH5TFu8nQPpZEtJ6zBuTVPCkALl/
3swO1kln+t3slC3i475SdmM6qfyH1HvPI6gF8JcjYIDnBrkPzb3cUyWm0iPVrFs0PhooGRI7POpa
lgEsSR4rFCydZyHlkgZX1nL9/jb8qyKXxKf2inVYkp4xrPbRodFteR/QYcy+f3AsGn3G4Ra99ifG
RFrlFcc58VMbYLQNl4S8p7vgfgdYKdMO5X6uMc6HzGSbKnL8CmtFLmz0kAmee4mmFbvxQJ2OJ4Vd
CBLRT11XtPY2PmsALz8elFZMizDKANqnQtJ8AH2bc+T2Okl/eILFQqOM4kNqHfvRMIzf6jcTeNnw
5+izaZSPS4VacQVjxYRpnw0J65ieSfh8NedKb9ugO44d5Ij/z12OOcT7JqOohZwRv87Xs7ZA5GbF
EhZv/HoKztI8kx+MX2jnhwJfDbpB7suhei7Bbi54qgj7veqWJDiUBe28Ql+HaZO9i0aHFARwT5l8
pdAlpi2euDU1BYaDm4OpAK2NRakZHwLz4F691N+L4PJIG/htBY2+86r3nFPeoRLqRx7/u8szgIKF
l+9fLLvStcn8dTH619GxwCL1YYtP8kOrhXh3MkV9fk6ZuurMwpd4uFkTeQuS4kGQHX2XpLmpGIz6
xjQhSBpH7n0ILaMyP0I4oqUKxqWPmW5WCg+xPbOms7GyWkkAyvXZzJAqIVgggArNQf1G8+kbFueV
/s8+riSIQR31hPUgPEJm/1QSmT7tMGqnPj91JDs6p8zyyz+tmTZcwRjpMDa1pjkTSqXjNjWX/fk1
/TtokJnYP2QiW/Wusp2T/djs6WYlkxM1mx6TPqTUzJ588eNo+FifksZpb4cT0DFOeAeg8TYGVWjD
0NpzV7WJNfYUcyN9z4jvWxqEFeMWT2D4IkCAbPO1kvKrghjtCI0qu3RJsC+luSoO+65kMaLIZKMO
U0zj05nGOuttnc+GsBGTVSvTtJ7hRIn24gFqUlWGbuvIZ8ZOLiPDRfAnoE9OQMndXjyyfKL4mrPM
u5VNhdbBXOASULXX/dgvOqn6NF83Y4EpNbt5xLj/TgdVJqnFnupRx0YTSv19LfKUB1+QgWdSrMCT
LpYnWs72zl6WGwMWxlfutRk4xf0xZ24kxcvvxCpmayDBZUhf4P0Pn/SGkqCCp1MOjp4JRhbxB4Cw
o8dRZ/MbW468P/cRARE6HFJsCf+14yeh5MKJKBw3vUB1LdSAqbn9hN1wCGkdk4WGgdpTXvaD15g4
UnTngzjsT9ZVyeuW1bkLtK9nHXW6O4n0WSOxYM0J5Id+ewXSjBkyNrOfBsJQIKNuhyuYz9OhMhFS
+u3V4pfUZf344CtvAJoNZx5itOgKCDVvQOy49ewoNcxDtEraBAijR+RvUKP/InFWTje1PGaH1I/7
Bvx5x1FRst6/JKbHOE7GehyMVei7KKUrATWAPEagLWi/FFCVVvx5CyDCPhQCF5aF+XWclIycW+Rg
cUWVCxr+EC7n16J6Qio4BgL8WqoSZbi6vkzGRIVkCLuhJaMb+/Ntxnuk6QrHTFejtZcRVC6ZHde3
hnyaqeQ3RiyGGrABfjPqkAjt27IiaPK+WV0XHhwDFKAlAaTWzxS1ugy1wxfj+tx95fbL6UIH68O7
Rv5THxBwaUI8VwB3xbNHpZBi/kOzpqASgPoRf6Pv8MOlHoOizuS3URKC5V5ApSUYhqpm0CFF60yF
D/e3p4bh+5dHAa2l0BGIi62gYqsd2U87lzcOnkL9KbpW5bdbiiMVe2clZ5aenWXGv6+VP/9zuhk8
IrD4m/gBEkb94mR4BBnh7pUwocLvQ69x00xXgoEve/85Hs5KxLe1MluWuM557ImLIBTxZf5kXfNk
ppRkHQCmNhQB0oE9P1mfDmHC61iNeEkwpD3r+Yl9UJkCp/q+i95KlMw0JplPGYm9O84knD9EsJAL
V4hKesHM6SL9YHLrSSxIg3Z37bJxLf+xdroL6AjT2WCURZ7n7MM0rTmFHzvydCrNlhotA89MA5Ed
DCQ06U45GIR+ZDCk1XrJr5MM7FWpFb1Jk/p5dFLimQ5yqrSLfQ9Ix2kKJJ1vwnZ8s1FqF9HJOo7c
oep2FNj4dozDGtcLeQvhlFw9f2CyGGCIL+OpaysXkIicoVbmaZwnQcuXiKVtkL59SBL+rVc+3cr3
xLeWHXIarZVkkbOiYsXFrpOJd4l/Q5E6RrevOo0CafI84GEzFRJD/ILlekr9cdQTRld9HJ8lIk3k
5EZ+WSLxDnn1yr+DxY38dNePp4eg4cHoz9x1QbB4dJnmN9LCVveN7XPgP11AKSukcD1jvsi24wZ8
mL4guBTEdZ5lTjjZAKo2e2A5emEMbOpuF/xrqS7I4hHCpc4r2MSpsH/FlslQKSYHMrt0/2qcDpRe
2ypvoUlDOtVYL+yfo8uacCAc7ciUpvDYDhH8DxEBFW7NVwpLN8E5ZvpDQHwtko+hE5JAxSvgJrwb
4oJHiiLNv7WwdpTpy7uT2yMYKA/W3iKAtQLz58wKOu+ykXYeEcdHwWhUefNvVP5R8m8HJpoL/yQg
P6CMKiZbaP10ZA9B1b9MfFbuTKZ5+pa2WKrr0JiBoSI5zUXRl+neB897eszRxIB7FNDJnZmkwIQq
2yE3eWAahrNzRwi2l6U7cZpTcG5UFMFWFt2uOxpL/bZA6PtTjfpNrHXkGNbRTLa+tsWwj0Pn4uoM
VGzB2WZ08YTK7eHlOtQpDITBrBunqa+BfXqwRnzve72Q7S+yMJAzch0+1kQql8DBIxyx36LLsTXK
Xh4jaHoLKFYFqcZXLJLRMdDOr0aoS0/0VTM2LpmMMhHolhT8ZV5XcIWZlrsumFGWqxz/Tg5VbCOF
Ae6LcsI3tK33ZXKTj//mSjL8WWEdiaC/EWr73MU9SqF81ndaUJvZsvbf3voLg87txATNzjYoD+o2
1fJxev/xNyKQhcYXSSvRjwY0CG+zCEFkNNvnOsjE35Nb+kxiL2BhlFT4CRKtPRiK6Rwt4wjRQk5y
imcego4XYOXSL7jA2HqUhllrykQMEZOQ47Ut20O7snpHoUT09SoXrhCLCnjmkJTnlo0EhRk2En+4
lVzIMiplB8ole+6IIQdNWt7TPewCgx5ggtswnkg5wMUnud/ohhUdkwa4JaeP2TclqGu+X1s5RI4s
4mpoYFGsw7yXRZKdPz0pR8X2bGFlbVYDadwPW06gFpYfyWi+RvigX+DsGzRRCGedpAipSqRJYBWY
qApq9gpqTZFGthDRTi6/k4uMxGkTTy+I2uzx78PAV4UrgtxVfMbRJ9Ea7X10EXHEzr53rGWW0al1
K8bt52wLiZm5lnUqLFh16TXpQQXJOhpn9k/oZ6UCd74cylBMhNiaPqJYpdu5HimcZTJNaCJzjVMo
PJbA0hXPR4hSyowpEapaLD0cpxSNiv3s7YqGQdCmICLmSOBjqqreDAwt38MeO7j3HkUPcJW6WvZi
A+jekBGW80uETbyBiR72ZKXbyY/5HI+9QBca8mX/hYCZyUytoJUkp5rrRSbKMHSvoVfYG4A18wqU
7k3w4yh6aqE18lgUq9FfDwBZBtRQ90R8rku14Iw9WvblnaMhIz3Jtyumboo+NX7dyget7BfE76j0
jl/SW2HuBWbeVJfkpEe1qFCPovNndCB/vFnIsR323xba6TLr51PyutbqNcJ0FVj/+42KqSB3Qn5p
0gL47wL+O4i4x1mhCqTCx7eX2zhPPNATAuwb+x4w9Q+Oy0Xi6mfSbe4ubIIDZie5e/XJARYKep/D
4W9DpQ8iJmVwM9sisr8J8jig2QqOiw6U0Afnm68WUx3us+qUQbGQelNnL8nKVrgJLyRdBkozjwzm
NEXBKy9I/xQ2JEb1B+juwxQT+bOIFU7dDz51ogQkPoRSaTvSnllF3AHwftb7M+pTnctBbBZnfeZi
RnbXjKm4TdYQ2e4qkNieS/TZ361WmjNHIoDAycv/1FY0pLM1gzgKxeNvPcp8jgUU2n1KOEdYCkVZ
eRex9lHYsjOpLFnWnd7CvMoknriFduhZIgSq2FKsUiwQ+Qic+1ZZZW+7GJsecz0m2SdzDL9lVGgP
Rs/q9WXyUp/zQYj2gYLU3AfpKpA0C9BvZWBm9orgx+tjOGbDnWypQRdTm3pSHUN7dcVJ6TobwWVW
K+bx0j7ll9aVCN/WR5DLH3dVTtbvCFIGw1UGor1Zv2pE6A/asePY8+1aL3ka4QxrH+wsiwG+iRxd
kqqyA+DT1DfpB3Gu1SZucRAFdY87NFnZ13/q2GApHuE8wppxqX8Cl7y/mFr/4xhfa7lwe4UkkayF
day8f5Av8mLP9UV7C0bb3qVk1AqzOabszKK6e64DI9fnLk7b1uwYuQx72RI5QJ6o0WtmHYlbe5mu
ZX8QclFX7M5aoh9qup+hsjUD2DSAUCQgDG3I375ad9qq1r8++ggY1W/+ZRhjoxZqX1flOFlP2AE2
oeHdMDojow0kL97eAVvLqmXaWcwE+xrmaZt4q9XxvqCQNqJCnV54NVUDfD7a7apl3Uodp6WdcmQk
K51/0WvszFkIyN6JFwgxHkBoJu41C7nWhycQ/swncrjmEuJeifHi/vatzbDiZd6j6TQmFecn3ntj
R7Q/A5ngmVld/GCMdi+b1RjxJDicf1iy1ekIRsq9mQ3yK5+m/KUpym0Ht1/oo7b86GMEzphk1nam
CLarG3jTmYFZiZBMaljtmsnOFmRTwtQMeNAv7C7gHRqK/Fnmr4bvIuQF7XbHUOSHcbSGwY3S7Ei4
sqwLpgZutBgWsgRrWb3sLH1vhyDO+RQo9uK2s9ZG6sPWFVuxqigq0JZo1MO7TGJdPj8TXSUKowqC
sAhhSa9uBbpuIvLozOxuN9odCufjLXCNPedU4MBiJAbpIjszmnFHiOtOTjs4k+FGeCIK640givGd
RK4T7VeO48bPgsWo8nZheN4rVAdpK3MkYsJwR1zuT7EqpoarmdkQARHpI3kRpd4MkVOSsmSu8dkR
2y3aDFSTXRTX4JyfbGRKzvm8c2sYOkSf6CvP6bIKCu9g5rh+b3EyI7Iwvf6X0z8RyD9kOx8grOFH
TmMX6HRCatebHl9RW/zG2QT/2uWt4VaG2A78v3+pCE44D0DLx2kkgzTXzpsRywiD7Te1G9E4VPH/
aDLHVV4rDRFoIPwrc0uF0ojTKsuqUxGNNPH+KMjnDaZ8u35QAE6jFlqRV7TxLlETwBtTrTrVeKp2
LeYaobErAq9rMD4cOY3/kq6IJqapeIDRrsHwVv/47FhBCd6jtTiJfHYe8jO3QSFD+nEvCsiIAEqE
wbsI9e//GjYNwgLa5JseCVij9GZLzfHO7tySyzpQvNI+Yt1tnnBEGknX+MsVOk7cM4mFobxqgDtT
bW74lf5tJhN3gcmbE38v1FpNEZCojC2rJOMpyWVau7+gLpLNT32bYuWHuoJp30onepvDtQs5ff3r
BA3PtxONGCoF7E6kQeJu1kh60kYAcUMhqF691sMayQNNYJYCU8lLs4hmb8b8JIeJtnVO+zapMNU+
NbjbLSHsJ286BjmHABcqBf5/snKF/8NGzQh+/KKzdUUL0S2VzZGkqoDey21KGOiqEwg/e/czUuxi
Bnne6fTyHNCaFKzthf9Eryff3M6wVsc2OQxgMabDRPhuu0Ylwy13vMIXcC++vawaSFQE54v5GSGj
odXMZPWQOeQmQkm/9kXmNdJ8BJ1gqvi+k4KN/o2AQiDLH1GcFZhkeVFuQ5P4asyhJWbf/W+36y4+
EZHKwOmEGZE+5R2n5sXTvrlRtPZqaU0PJ0dkJYcGsQoPmB+8Bwn92uJkcst+Zs3LzLZgUvNPM66B
ueGJv7Gxx5jfEaIntj77aGFmpZLq7PT6pjaiuyNGmL777bdlk18bEvwaRgUna1ybHJCxy6B2kB6R
i2x9mI6dG5jnaxeYxKFpwKV2V0xRw7PiPtMVxqMyvHT+lC/4geWieubAxUn1SGc06dYahnKarpO7
9zHVQTz2eFJGf8zK/hdwNOJd4pBNx13yI/OBWigkHVLmWPWm9mx/idvwqrLRhquRoO2z2QFKgDG2
ifntI6xJq/eYEtUx3fwZng735t5YB0yIVEtGlj15mBJXXGWrzqtxDWhbVofXQzyQZa9bBmqhq4O8
WVEHjwU5isJPg9Z7mnLfLCYNhYhbOUoz/+lmiAXRw53t0mazRboW2QiZyKyZCkC+n4Ps+dCw+KIj
JJb269rTWh39xDTb+2tstQiLSZ0h0ot1qyB9ZacYdNWFK8LvMgwvVHe4agkhgyrcYGiAQhhd0Xrj
rHl2LyrRrbrLGd47/RzbiqWZJiwHoTRyUyvfO2hLIK3r4TRZfhWzdIh0/EvltGjJP36sWySOpApX
BM1wiQSJsT0rB6GW6pojlHhE3COh3hFnlZ0T81m+Zm348r86xfgox5NRtSiB2AdCQ90maATzAA2p
6fnnoMCz0C2fdcqC3rRy+uDAY1jpooUeh+Ziguj0HF42+vwxkDlobE4cjgvNNMNwZ1EJGTtdIhuh
/Uj8hW0rPVctHsq+vVWFyBpLT9ulRT4MSXkJgIkVkJvcrteE4sg3sABCzxM5EzQtKezJX9Pf4y+T
NmSRNcCebKLSJqqBgVYDnFtzOkDy0VaOYDSxsa9TDU3GjfyRxLDRfeLijVbiBviMqIS4zZl6srgQ
QIvjMxSITiGPIpZvThyT1Bc29kRy1E7qX7YrF6TFRjOm8q2bm5W3bF8nKlTfCVZXjJBex4uOTLW0
TwXx14CMBw3kr/03966zSG0g19RTLBw9U0orlj8VG65XGKSkwp84TMUp833LCDpqeot8Yli92kbR
lkW8f5oPK+u/1VT4KUn/3Jz8JVpQ1kGnoemImj7vBY0F5dvg82Gx/ZyQ9quaEPVwwzHUGGxfjngK
TaHKW1efUEfOSomlszklAmaHNNAQep1ngVFANfsmTFB6GLqIllQwKYonw3QY0VmdsP5skJsEpZZ4
Lcj9zIrhFpjo2EecvGULK5V7OY32323eM/DT/CcuDluQw0iBEWD8BxdFFrvxCKNi+NYz21u5HfT+
XFqtzl3XurUbrqV1zb0bqX00ZtSBO+FUyS7+00iAg8awczCe0lUk7VQeHALOv07uLBrzol+38aI4
Im6XGhPF2kozIZ6SHdkCujW1juGCLtKuNIPUKI7NlUlqxqrBHcGibJFUCW/GHOqXoDhr2ovGWJZ+
nCSvnl4QsFLy0ShzgcGa+C2GupaLPRQkYMe7VzTnP4iorrGAOVQR4XoMvpQ5krUdSi87hcm0jRAu
Ck06RcaiC3lO09MiGtJw+p4O0xMPSj2C3nxeZFx7DAJQNnGNBE+5lhDeibVU1NLswxxxbggSQruj
YYPdbrry2r8Rnh0RPlRx1iMK2qVghJUCVqu8cs14VdyprGddZG3/8i5YNqOAWd3ABqvVrNJGe6NQ
93qAMhwR7vBA3eDn76j2qerhkHgwSrFPNfKxG5U3OPEC0La01SkDe9HA9rbUEPAaX2i+V6HhPm9p
qSOLzor+UuL0ZCq8bkP4Ld38AnQB8p4wvxJ1MgeRp6zFzDyM7BLVPuXHhShwyvcD4bBWxapHNwHM
+QsWmnbYz0libprm5WytIKuNoz0BE/w44vR61J23XdSiAWnEHCKLJ+hF15RmyeZiOnqPf0KDLK6v
1J2qqxyMeBYhzOfY+rtHM52i+E9h3LNCNE5SzK/anzX1jA7RxfDgcLuEYoYdrSg5b7ACfjVF/Asl
L5qyZdWoOJHBqoMUsByT3j/9SOpGCYJbI2wxcaJgsjXG8dzRwHgE5CO/0BzfXDcJD+7IgLLsHP40
AumzndfSmaXqOxPyH7wUpUJtABgDRFMRaw1j1ChUg8WVsZwKwDC1pcpcNx24pTp+TNxRjlRXvB2u
cLlar64JA6aUUIV6x74AK+j59ZUhULQtmCXsGfD63Fcr6Y5UfFoSEgz/4Ft+nKTc0gTO2+WE388J
9YeAqof9L3Tt7Zh3a4dZKmGPlA35brvVJkDX4uCmi+THuSD1R8+FrLu9MsSuOvTSMCXTUkU+9YSe
Gx0FYtT3F6bAc0YdQZ9VgGSfUcNRqZliOwZK9yU7c+xagmvcb3wuL77DmUbmHMjJRrZ7+1wEnlXb
N8QLEPPIj+uHpbKpIqRweXkF+8g9liMtN5Z9Dds8szFQpqUuR9H9i03ES/1CEjgCzcl7FcHSGGlB
2OquOGSgi4FG6AwNV9aK8V1vXUbcYUDtr8R1yedfIeIY8rMouEA/PZIFW6XN9FZkRQrbbdpftQ66
aolqvPSnRWl6yZIpVc48tbwc6k8zmdzmZljRTOJu+oW+mHbPyGcx4ktmFipo6wu0GaLMhnPQ3/fZ
/JqY82i7pgQEMU6PAIdMGl0DHV9t8Kzps8QnB+IsrIhqChGibP6kBh/4DHcDtkNKl0z5739sfSgb
IBzwgE6uO0EMrM2ezMSu6OuFlOxmUF4zOe0uMZW9tNQ+Gj0CKrkpOGyXE8QstnjeaI86UwnBuKB7
vEsN8Vl8GB0YKUlCw+BbJQnX/BH4yOj7kOKXA5rTcFokfENkQgssU0Qbjn4Cy47vYmrIK7u5d0p8
Wxr3SoW968I7YUgEK7AKisvM61sNUVfsP9KoT12KIf0Dw0oQPVNgbV8KxS2Qcwjol0oXYTSt4ZI0
I9/JfUAyNxQ851RSnYxaqD7CCDyMelq4SRS4jaAG9ZNFxJaLWmxmbXkkEnVZdEPbjUq+f2DyE/09
9PSG7820V7LcqK57PiipK9K4ySEyZTD0RanlYKDZjhhmFTTUc6BuvDDaLPvyUnOmUnoOgqRMJ4jC
aqDOgsoMNQFqnCjFmq2YxOD5VzrFwK14qH3cb8xuxFkYeMoNrpX0dYT8osuO+A4AtFX1IvZzYVRg
+iGOnbbaHbKPKmXhJOoiHpJYw2jLUlWKp67vzaZitZzylRPBZz6d+ywh4TCo7AvQ+JyJD1ADev+v
3foiELsjc78kilDdV67xrxQpJjHka676z+W+F2ZSo/R9Ue7YaFkwBuQ3g/b8/YaVgRUvqY+ffrRk
97GKxilYLaol+z+NYpvhT8fzlSnocV+eHNzY43SvYuVC4i3cpeyuFf5odpIiuaeQt1WLW9j3HohQ
pe69duNMRYl8IoIltTW5em9bZekyDOQ6bntquVWF/lTi0KpmFEnCn3LB90jOCVAWLlmUB/24kuQn
x0y82eNFJ+ulr3QF+XPo645B7fT6/33po+RMlM72JU73ESqkDDQuOkJniAW+t3Q+ctrnf8krm15s
AtZLis5bUDIw24lltSoVTusmwhQmQYc1oXITU5Zxysegq5cibgxR71pf95oCxbMw3Yv0tqXK/Ltb
2ehYRcsu2iD7q7U9ulpzKCWlDDuqbJMCGsjIRK9iaL9YcjGLEKVdkcUXAL2a1UtFx3ZfKFhpMh6w
Iw5YP2X4q7W+F9C1zxk0yBcwPG864FPi/8pRDK3ak/9tN9OFrPuShcl7rq1/dN7EMPWoAkF6yyc/
SqNGEVz85XlEtAav2OxM/07ecfnd/rbyfet/uONUBDAXHmHvcBjQnjPH3qoZg/WrBa6QswehAPZ8
bZ2lBZm/5ahri5Jvlv7tcC+8t2SQn6QL+dDACAHkBCywj/ItC9eWzDLxGX3qBCp57OGwwCnIkFVO
y37aXXyAougTi3kb5Gof6W+Ng6Ywchz9zCax5iWqSnKsPPDKEZTqQH0kE8iYxyq+CVeOL4O3EZ5u
TiX0DGUyPfbTApzeyWKU8kUOrGLWmifqnwlFta0BLKFvEyZ9Lv8Z23eZihtYhI1f8ByiQJBo3Gr9
t98IMfGaFs3pxaRMOA5RgpgHD0g5CZamH70/3GZyr8X21v170VHRC8sr4tTPurGXDPU2OlPGM1i9
pk0OMydvaZKZ+ZD4fj/bK2OYlexzaNkFWs8lqpTY/PZOH1J1AZ2T/HuGxGlHWykQ81L/HpR2hiuQ
B2z6Cy91qxSHSW7yDnrHIwaw8DaKN5hf5rJnTf4c+aIkSU78+SYIIPPRMerRZNOePxCWxxcgxAeQ
87ZmyzdBeIreo4WFe7tm2W6nYJpOkvI/arW6dynQAOrkyLtBCu9nhyssIc1/cegLjQBykem3Y5np
mNxGWezdDCmoq+2VRwjwQdKG27m0idv0LMKfaprOOMG9teUDTdCR5O27GQa5r9TFvhoLo1oQDlNT
O5NglpvjsdQILUuZOmNWNLitqVSPGBETKyHo/FCBlYRdABWrKWS1183wLk7oJSdmg1HQobd1ZsTH
7X6+5W5wG5VoquknlOCmgTh+ksvbXJUEiOtynYz1S3LkGadnI7SiO5AWZ+uwcxXECaStpZwUdFst
oXsNXGJysw6is3UrBky0Na0WKGKGTiu4ftdM7by1RFwv88E7dpCVMSK3zwGKfITIgfPPoUed4sde
1MB1qyvQY21UgybGuQn7LvmRLMbdpIAd6YpaFs8daR/uub6NSRpNfVI1ao0zTL9EL/bIUlhoUb4l
U6pOlhh5gXhOVbaa0NCuJ0cBUnmCPhs7ZC01U+2WZUSm+jT59/1DcNWN3kwj1I3xFZO8aTr+rUBO
yUYG5aOH774d8jMmnGy6rCAwVhgyBgX4xybnEa6oL3I3fc7dUnLcaAIsRXi6+8UIahsrUJHMB70+
eQiafZ02zAi9Mf8yXZ6n/Yj8OT3RelbjW43RnAGixD71KZluXUu3lXeKo39NnRIQEmSU/NGhXT50
AM54uOfxozQGKHbPMiKufMF8Z6eC66iWkxzXm7xMluS7qS93uf6bErXr5zct/nvfBOzF3bBagk0A
Z6L+cknorOKZNxFhBYEmDhdYqbngUQtiztQERekX6mVTR6X22YBCyhbg7ejJqNwTGsrNzEFW5pPc
jhmmNXMqCr3XFgtHWpt90kOvEN+vGOvl8TmLKA81LWsPox/YSzX3UEIkkwYBOQqbHCee5d0IhReU
5TGYTOcg5Z2SHKY/GKtq3EBSmsfS5dvBcAW62/ioO1y7nQY1aq3xTS03FKIgtLbP/uoH8G6nt+A0
ANUZf1fanG48Sh9Gt47vGef5REZy5eanY0hu8LKu6oDRS0lmuktP7Pk7ar+BSCh1BKV7x1uyfl0A
hKBsL9Ta8n/osnl95OutKr80ovsitoNC7kHM49oz3TZoRyGy9DQ4odkXyGpynXpyQN2RmtsYR/Zj
xYm+QutPyAfLR6ULRmzoqHuQe7EuCORzzuqQIl7cPW7H/4ORI7c39Yzj1WcxWSXEDKl+cQuKp0xr
m9NyGo0KZ8MevH/qVZ2CYpAq3T/TTcmYeZdvziT67bDpsuocb4aQacE4xD0Y8Fwtm9T69t3ESAt8
WD/2m81QRka0Xx5qieDeDphBmJApuIcpJvcLHn0lSF7xIrfT1oAxwp+HFR7XKE+X8Mvu2oovYg4o
ZeQJrBUpEV3+zOl2/S/ohlK9RVWSzwcdAsiOsT9bNP2/Rmzw4RTQrhWqhfDytE/UrTrPCmFpNv/e
5W9tFkoRKQFuK59jrj3tJVWDUvxBN3vxkAhSKS9Zxojtds8mxjH3ldp8QjASzHtirkDq1SuojFIj
9B/nhlRXZrDtd3shONLE+0LKfrfTML9SZcj1Fe7yx1+3LwRbruU4QPNQwuSRIVyn6iVHqWxRpD0v
VvnTt76PkXf+0ShD+q0wnSDTQA/X2xfMAR/PuLnQHLSzmv7ck3jSOky8yV1jRJElZ4CHypEavj51
7oh0B054Oiz9X6HuTjhnkMLOaVWcIe8/CsbbUIfHQTNLZ7iySgg+L6e5cXzQ571m5M2FR/+N9khD
oZWLF+nTlKQ55mSQvH1LrM+tFqtDXNhnbk2bIT8haWEnPIya4KOOyUW7hyrv+IOkTmLFDc1mFqz5
9ZtIbmWjoaRAoA9cQwfhwoN80wkJissxajsUSrLSsWFjMTsVWaY85Hnoc/fMw/Juaiqz0x6iPaTY
XUnM3COD2Q2DxdaUQc5PM2EJwSZfyOaHge0WAgWmVmAIdwT/evnPq7BFmes6mtyupAnod+kuMTNd
CqY2icfHfYDqHnxjQDetHijcJrwvvj9mEinYkl16gd10QG8FKdSm+FhpGOpYn4dfuRyogPM7Zifa
/B5CDqoH39yD4Uh5eXlI/e2+v+iDhslOY39AhY1HRLar6gdll+2cLwcuq1B+WHG7UhHkJvfoVXlq
Ej0aPMEOP9lwwA0d+LTexVcX3mzHim6IgPFrZcajl9mpwWVk6mPjufCZho+vQspAOaQq3IDjZjKO
V5WNBQEKWhUZsgsJoG3TropHlxv7jXmqNuNyGop5vSCNpMYo2O4vRI517NTFfMN2RkOnRm3zXQMj
IZ/R1Fhp3skuN4LduRKUGf/eXJYeDtNh/KHitqZrHsHlO3DgqaJtKBLe6gkBM1Op1fxkudLvSlYu
IClp0OEq+cibX4pyvEAFvXkOEBPC7qSxOgTjJKUbaUfEiZEir6SneukH0S6qWtesbjBxon+Cegt3
4Wx2hZG+FyfoANASnKHVQt6dPf3iWYNxCQUmM2Wimdn+2LOrYl3843ORcXF81V6YpFAuSKVgDUpF
ZWbYkFc349/3fEH8obrfr9DXvP/1b4NKZac2+xGLqHqLvEkwQcniMxnEeFu5K76S/NCGBdvNGQ4+
0X1NlAhaTipNgboq0MWt1j5xdt4M6bKY4IS3CS6osEf+8412o6CQjT+40G/eDwZSx4Ni1zLO2ucb
vumikFP60NvinqJD5qyuASeZnqME4r9g0LfhWkvHge0pMIW/JHc0oIsD3LTceSRjWRv8nu3q/JEX
uiyaZMY6A+EzM/Lz0L909wRmkHWhkBpbr6ruKiEB9UKLUoe7a754h/VWY2CMhFFti2rZims+Om4Z
ODr6zsrHCjJBGOLRE/6dYkneoeAYwVyyVe5WLAL4T87iPQROthuKlaEGhpkT5qfo0vGcSDas/ZuL
WK45B4DGFyfEYzGzdKIQISLf6c3fRGuKh7HEPIyIodXswAn9SzwxMaocaKrLZ+ql6ChRO5STCc3s
RL5u3ajutgoVArb2EPrpkmcFwnryZzEE7pKqWmVKada6y42JHd3yusnGmCrLONxOCno2rdr4y+4N
LhKHs9nEryUx2z2m73HajJEArNFSMwrt+B1kVB+Qh32Zeu95lajBqvNrZ1Z+1bjOL0PucssmhqdL
GBLCiJlDJSC9lYGbrXpSbx/e+b1VstZO6/E7hONI4S9yQjAzH2f9qoJt5Nfgq3oQWYQ2nKX+6Rly
/HzpBy+HVnYXTKqMbrOK/CWQk6vuCldsdi9kJFGTDeKkkrtWvNf1ddVn6vGvAZoP5CF0MCjdFoKa
01krWmyiQj4Lnl4g8VfzJimjTVtlN06nMDVSiIy83xZJXYStWAUeIHh4F3Q01iFLsPH4fhtZd/Z4
aUNK1NFqCoD1amZYrGM+GlQQxLxfKv60Rg4paOccKQHz7loDpYR8HwbRE9Y65zJnz21ncpVzsHaA
eeJ+tl+aOHQUA4rwvqFUeIuYSeu+IvE7Zyz9gCo3OPo6AyZT/+hohOskA8vzPM5YI+0ROr7ChK8d
g3koe7RHCv+UY4fgZxXxth0m95DDCaaEeh1KDP08SMNP/Cq7FcKGAZXadOTvB2AG4syW7h9+Rikl
4/lavdR6LkxuUHWdJa/CNh7D7hKy+Tzn5MEhR0d+tZtdUESefqt3ENDGR/cgwrANKGXJIUYejJPE
ye1pCqlZSEhzXnIEVJkRR2ges6Vc9h2IKEs9W3LeoHety7RxUpCpCCAeOKn1NCiPhQ1+mSeW+ZQB
Cr4nBDPWi6d8pSGIvi7DalnK+J/5busYN+WODbayNipxN+2l+GTDHqvCPWAp5OGg5+9yzGEb1nEh
lEbYyMrAxiK4fBSEjXDRjAUklzJXNC0PJLrSCRpJ/mdWiz6cYJWkSBROC+Yk8qTSQcdQYg8/j6MU
L6aibWe9tQPDqG05imqcNVxnkx3FOmfggJUZV/mMbL8Q838qgcPrCILI/kK6ay81o7joU+mgdsV7
J2u26A6nSy3wUq6wWLq6oBb75BU2D1LMU396yYl2lyqgSpH8WnTt3QUpKkjZwmRVOhzWvYINc7re
LjABHhDD8mlIPYimnm4wTS/74B4ER/FyNSQwvm3PM736ipfrR0qRWUCztEYm6cqlWEACAem5q3aL
QiOmDLjjfXobDRmLszRKF6OnSvhtUnoI7XY2wosPBkJdmgjxrHZ1SXWcE3ssKn5CCABBYid6Z4u4
VNqHn+al4kTUJg9PVW9wSfjBDjllwQgtL4KobZzoyK0TtPpzr1xN/MunKc14ITUjdyN6b1mbFFLU
BC61bAkUrFrM2DAIHx7BYnQKzpGFIcGTlY28oHz/QDT4anslKrk0pr5kcvAD6Z+yWd98efGwJ4bO
g2NIxriuKeMBgaiU1X99Y2B+hGNyO6t8ylEgMN6RBMWnyRiv8re5FYjMAbPeqKdwWVXeGQ4LEAN0
npPzx+ZXWeYp7vN3SkDq206Is1zAHFFjt0DeH4UsNcGhKPD2U7iS69N0E5krfTREW+bcChoHqyNT
HkzLSxDfM98DFEfScT6Igl/SXE86ALLpQV+dGkAePw3XeiDIfMMmYJEV0HaDrLuqD4W6hRfx81uO
6BwhMnzq58s6WwoMQB7V3Qc8ImhYXECczKxA5O+phJ4xrIaWk1Ps+/Em6Hs5iSXbN7GEBlobO30u
eBbziV4GJJDNqu+cHOD6+XmdxLPDJeDUFRY42bKUZQeDvrXcJeCYwTibZxxKCp/U8phnfUchhUYY
XDags8ol2Tp7LpagjQZrFSG7SZwYUZToO5i+Wl7QcpVAXyn5wEBt43Ozz5kJCLhTf9ClC3LuZWTJ
3mU2jgFOSN67yjUuEXBpSDFjm2KAYhUMG0aQqa2KHVr1xvhReWf6athi5Uak7U0qkREI+rwdVdfv
iHP3YBNW/kljJobCXbf9hoXb90k7fkuYMHXeYuiygB0fhMc+MjOHDThNsXwVQ3/Li4QLt5IBOYlh
9MhmXleQGXU57YgrTiRznxUMWYsETf9d8n/gcfW7gCr0TLhOJXl8ImCp2AF8VOmyYahpMM13yC4R
dYev2PvuKe7AIyM8V5UCPszUfS1PBu+ZcqxEFfvFEYVGe/QwoizMo7ROVSYmwx2SqhIRROnUT5kM
8MNmaw7biO9OVYRuwu/JCkHeicvPi005PHwTzWSNmgXQVxP1gbliAaqjANdj7L89fDg/Z2R4nSRC
5KJ2cSN22xr6sWui1L2VU8Jz12vu2BHbxw+kpmVqEKz3jZLXraaatp1C0QEywbrloP8nq9m8Kc4o
B0KpU6xbmo+NUUiIFyV3yCHAk8aiq0gL9mckfMmlVtdbPp5BTXI9bdcdenGbBlwfiToYFnJQwBYl
0+Zd78iUT6DE2VAtZI8S1EnEwxYHEuw1l6dR04QFrc6fBAml6zepYozP+iUtXDng20kiJf4Wydob
blot3Oi2dqIJmQPqHYro3AAgbj7J4N75FW8ixNlN3bGP+C9jGrpLbrAGnfzZTsm8uYClxC3iqb8h
GVN1BaPOR4Sejcud5JnlZlehkuaS95W28AkzoPauwINSM4LN1uPNoEIRzAwWV81ktLSLstbNTo/F
7q48wdCKF+X5GAh+Xne4mvrNJ/Rx/szpotNXUQ1TMjFJlxalWtHnx8FySfusnA4+zCC2R3+zvbKn
nFCRad0O3Vvpm2YFOETN+HEoRjD21cRWseVo7AavQ4Eb+ZevJXW0QTULr0hqK+1pmdghFWhflFbZ
6X8+i7pi6hUGcsjRw2tIiPSkGP+PPyeY9Ma4akJpYVFU6yCASr010NwuAatpCe2rQ8B4LqCcWPYr
j6SvsGYfzUex/fFMDLJwpWp0qy9KpOnnCy0WGqLSrGErCX362OyGvhezmF6GfDsXSkhd85Aq4Mu5
OSIXTgCmH0ow7AGo7krG2FMLPbWNqpr1hes3ZLGQHE6ytRxqj0pDf10JMZQlfwVJUSwKaS5qbrmH
thlga6Kqn0ahx54CtxbNqKjiTzddynsa12zd87L1/pYCzM8x0eQT+HGNbS9r+knE8yxumDGFmbWg
Sjs8UP5N4Br1GdoC8Q4mFYgZMnlO7eHqVldO3CxJzB8tOQcj139pCMgMkdWXqN3AHP+gP8IafotY
BaBXuLMVYiXsciI7Mk294wf8jMHCzaIyjLHK2P00pDuSCf5xdby0RBB/TVoQKX8FKwMRzJv3QYpV
roINjW5SvIc+Q+4BmzxHo2I2+4D3mEyKq7CAAwsT18o1d1CvTRaY4PNa8ke0k5kAeawxkdRaTVyP
z+KTdPivPaoPJ/je/WUd4/rBeZa9pe/IoMlcsetBWcloKSL2mbbqGgkVWu5gnBDxL1UUoJPOeA6N
blgzyr1lFw/7z3ZD8X6RwYaidQv4FUdaD+aa17UhHoIgLwB0yONIthwoA3gUa6M50ehTRaAodRXZ
T3dhHAZrGLgnW5OnP8fK4dxbN/K88UxFnsnnX8/a9OHkfqPvnHU7DcyiXthIXxdq7vpW/vbpUk74
783W6RrzgdBnSuFtZ67VF/u6s6ItP3b2X7rTiOhYglxQJjRDqUZH+DUZTC2GzJos2NZWFDjmzjXw
YOHsg3a3CToirVjttY2iNbzPhOh7jDCwsCPex/IZizRe61Vi1TZJL3PDEKp8fwXKXzlLm8ptO6wA
p5+QLF5ZPWQLM74wfUu3TxgBkgSeKi49z+b6QXQyvMkKpTzUVB1oGwhIx2MJSWmgHavuKCih1DFQ
ftn3yPQyqIq+60pyZxqalw0HRkGWVW7IeHMbQ2R4jp6vzaeu5BYsBs4IHu2vkiBPA/bjI9E1nQTi
updGJqhpvF+s8fMyzqmr/KGRy4o/0S1w2RmhcxPZ77kRHv1rPpK47mDA4ovPzxYdl9AGMhlUkG91
dy2eXqmCGpIFVofzUDwoED17vb0ayqALq3eI3rHexJSPLYqyg9HOn1VFvONQHa/4q/lLvNcLO9IR
UBhPn2BiFZdEk9PaRXClhSc0AAWvVhthlPG/XEDyrh/b9mSE0yBs1fpRf3mpyF/sAOenAUL/+IAk
eydZIGseMicNoD5evAW0ie8zqYcaumFCEBvEkpWZF75Vu+s8uQPX9YsTSG9xiLSmMPkA+Ez7b4yC
OCm2L1DXwxYBQ9pjRLxzSu9imAjOgTztA61C2r03/XuabK+BSpslwUvn/NUKVFeCn39/1pT3+C5V
jgLp7lK+29KEVuYrhb8g8J78i1y4OP4bSXg2BxgzxwjJb3Z0p9Cy6tcrEGTKGTIfDLy6LKUB1zX4
sFw3loqft2a9tanFuKznHtc+tMKx9qF7/Zh8pyuY7bO2uwok8cyV/WfL7x5jIcrZDumZGVA1vJs4
KY4MimELUDqONFMt8LTh1KV6oDbjKtbPf4eYe+y/kre+lezzTuACGgjglyZpHjkoMPf8Fkm8e4Mf
9sac5+dKPqIoBF/fZRxwQZRsFOk/pmu11ROQUrgbRx/6OKhuAJZ/N9PUza/rD4wTcpo+LfJ8dYz5
n2X+nkKXtVHiudfuJGyeE/gRAz2HjOrG2hwcV8IMGJw94Z2WvnefxxyMlOslANSUW2loNfrjb+30
Yvj18FWM/0WlQXsdXbEPT4fzLxqTX8NJNwFhqHTVpLE1TVpWucN3nL5UNKhYfQBDBAXp/MW5a7NJ
p7DR07YKWxIXz4P6xARcbyjrug3xiMBqw2hANo2brtehjhnMHlkfV8HQlXarpGw0XVZt681PChMh
J/3Hq9IcxYH80yHWn3MsBAchmUFCTr9SXsfrYYm/dkY7/C5QfQGnWtMigPBKR4yjR3OA81h/73E2
Lll4Q6uxfBYZ+cf8efYpIvyOQnDt57Gfn+YRSltfUygbBPmW3AL9z8mp34QhdqRKAGzjLHpKCU/z
fHmbaMqZigrrJW0GGnuI3JEE9xUtehUv1aPXWmymUDz+Eqgur0GxZBedQDy5DeAO0uvEQ6uhkLti
RXgfUw44+t4prLOCNCKb/ismwx6HME1trBGlYRGY+7QUrQq4e/BiAJrg7e9AtJfmkdolQJlfGXe/
QTxuZQVboT7t9M0EAYo9u3BHuBmHoIphoPJ/sPZnjVBc6wOgCqPyFVlWD6SR9AgFYbHI6FQ0wYCs
t4Cu0Vs+eS3xV92QNxiDuMwyiAvUcsqgw8Iz2ZpaWf3t7vt6mjIYhnCgQyQ/c1PC8pmi1PPU4MDO
OYNjLFNLoQMrjFAkzPylcaeyM7LEt18ifvHld1n0aDAJf3XI9UwQ7Smc5dGNCxmwmME09t7bDau/
PKVouylPJhtEW/uFI1qOXKKdGuz34y9Zx8dnrEfoVuo5iLH8QwqOKj7+gR7aWjgqeDJCnp3k7Q41
LURkQV6VMlWXI9mDGuUmghafITb1spsf1qSrYjZgK4P2BtmiNkhWrJ5QsmVa6/ZIzWWrp/17qGW2
kPNhKgTLwSHiwRe23BF7djXhxyTfg8D4O5RPne4B5pIUeMq0H/kvzAH+mV3LXHwBlUicMUB1jIsa
qApXYzGRV95T2nM3Mv/NXLYJdcyvtUTi3xIaL+bQqzKbOkMjQooxgP9onR/keWhp6q2uS3UCagTN
xXTlZIa8QTtsEQDapTcaWuU9sGYkCMUCFnPA3Yj98HbxhooG9rSAgMPN/Dr20MnCWPeTy1P/GddM
OSHVZlnvtCK3JAQEm/HUXr4y+iBcoxD0iQT2OL2ofCtfg6foShCn6jx363teL4ODVfe2iJAdZj2w
erEtjwDvteifjv7hts2MzNjUWjIZVOUGhg5rRuhR+fvhdSRaCpVhs/z3EwGRxVk1TepBg6YIU1k2
LKuSAJ7k2amhgOJMFJFH3tXQ+wlI8GLZbZowYtzdS1/egAj36ULSKwtlq82F/EKKY2Kt44tEeVz5
dh6CRNc4Zz10OYwNbOSIhHyHwGSzyDgwmawdyy/QK38pYMPIf/577lsh9ea9Ie3qSXFDyrduvI+F
q3OQDM/ZiORxmJBBHgw/+pex1GsxG6z5vBc6sUXhhgfo7AHQDq/bP8NsIuRgNyOkEq+ni3qjq4pC
OKOcjUTuC4aQLVfznIhFgTGDT1+ybiFo5/f2Q21tGH6+HCO92fOzMO1QRlJXipGYIS+TaGQ/hV1Q
XwfGbDQS6vo5f+qARbRKCfprOegoUl82TmaUO/YCf1cGNrnxyWwdzRQ8iU55HCa8OSRpAgQVj/0c
4iEVjc4AIrRoSsIb0iXlXF8zA8VciHO6/iT0PCbxETbNSQ0T4qrOdtJDSDmjr9NdFQsfNcoBr4BY
lX+//WTCAgXf9ShgzpwzKvPhV4Ast4XINVM3r7XR+ye0FLDbHfl5gQZ7J1u44dMAigppZYBC1i/4
SpcVqmjyo3sIZPgcnmPBx20k7iyA3+oFFX9O0Vzz6owAOiw8Au50SKnTgvV/afnivPyiLl4fHGKC
kl3Lf30F0DmqD4fCfBoIJnA9ODk9t1oYRJej1lD4YSKpQyKzBZCxgoKnoRl13VT1f0BhLS+u4ZYA
M5kuNaNwRnPUINCS0MbJEJlNoDCj6o5RJNENJoIOQBl4TTCDl1H9LaItIGVYBGt6qdLjgzXMbNzw
UTzHq1dfulTH/xxHUmjokGp/+XO4oCa894xpfWEYEx1Mio1Ld05F/6Riodsmy9WX4UaQHwiTkZbJ
8DXAPHFZjX/PJ75P8DWlBfXu7y7tO52qqnn0gZQqwY8hAtSYXvDoWFIs0WFLcsd9sFbE9e62279F
8GPXqVwFlo4Cs4SK6aF2rljUoS/5AMNzWfPEokOyfObcPeOAi8Q9ZOVIErwSV8ZLWKQ4qPe5/srt
ls+52lO2CmSR3EDghcWhJRkt1ARuzb9b944n2zXALjcDcnXlfJU7FjSCQ3wM28Mtdn9VQdZT72qR
oKfV1bwuJkufs6mM/SVHY8hUzi108XRo8KzOspWVyUuiqcZIyh1FrzZFX1AzqJfnZpDh6T83Rr1N
fJ2vFp1TGb1EXGFNCh/J3Ft8IIeZ+8MNm4271nTLANLfJDkGKk5w88UzqQdYMIetOtT/lMyOgosw
8zuOdY6tC/G2UW3MfrAJWeH1VLP2L6/FREEddne9s0PhNdZUm4qeJ9k/r9aUN4DurVSdAhZM2D9i
Wnw2LhSNe4HTAqI5qzJdDcVSqTbFQ8Fqojan6tXjEkWGOkBnX/n9nLlHoauvX2gc7jOpNed1y9AV
M6yRYE+dkfpPHbvJix+HLOwzTMVPnQShTK7VLhhORe1er/lEKKKlGf+3F3KaqMSbxGFk0zz2x+IX
Zo/qINO3koTmwwiHd1fV3vaBbuFRl6XoujddHfQMbkQj0Zzg5t1GMMWUFh6j/RFtmgnQC46uRe4q
XozjzlLls2WtlAaiKyuFU6osfZZLiEDQ0MU4N6RpjmHSWvh8cixPMb2YyYZoviBPSIXWtjOTPrx3
cY4/7YCDyq/FgY+UApEuq8FRs68z5gBIKDlCrbgz7VjwU8ybAVL02VzsDMNoBU48imJ4u3Sn1E/e
jn4zrt0J94+LZam71oEK21x956X34Uc8V3PdJB3I0KYY/fBxp1d9nWvRH3sEqVv5kl1BiAuT5eLY
N3dxfiwmC6LjlXlmm/pgOBHcTr+6aFdwuObMHVEA0GhJzSb26ov5+79XX+/SAHrlehfnX9KzDtQ4
N1ti4+BmU+nfUDhi19IcTuSyczjQqs2UiEDPNloExwh4cQDl/kPjJ2MALuLQ5fcmKqUpTPOgigJg
/vW1ZeNSpvM1F7w9LvHhUFPL6TYyaixaVutJbMl/s3l5AUBShjNLiyOC+rwRBBz6YcGKMvswzaQX
F+J51AL6sDLWfMhMBFoWHdUmqfffiNnRudz2ynh57aWgSEpcIfdeKq469jrQ9SAgdm2B+J3Ioq94
0f2CsvQbmMSuQJxfyPi7R9pIH68lIwqMh+gYK112kINuqJ/rPD1Ea8ITv58oHoFSbbb7vyXx4fCy
J/r33m20H30XcE6nvX3JM1G/x7PTLoCf1YNa1y/6TOaD0ZpJAU445V0sFVLzYSfikrbQhpkaRI2f
H/jkt57OKjQ89gjOxBTUYBYU6IJRI03v6ndXne6OgRsRghuN40JoFd3b6T8YjIXw9F0y0j2CAu51
EXhMhyif3TDcLKfhjkBMs9K7+Mk98l0ZTh+ozXi4Df9vy/HPqHkMPIFTF4dM88r5V3GDgZEAlDZg
VfssugIW5si8gyJ1JcT95SsVDGfGC3WiiLSVKmJIcKmlti/tRDbPQAXdouKUcFUX6TdqonTte2aj
pgVxMjNmEWDt0KVuYxu6e0hzZlRLcMZDqAAoS1W5FNM7sBiBHtmaWmqJf8kR47er/aNZwt5fnC72
boz5F1dwSrHgurCduDKYKTtV4h0j2o2fmj7uquMnm4368hk+NeuALdOL3SJbbQDd5nJbd8jVoktp
qx3SJw75ydFahKlxIKLkhIJrGZKdwPybv0mWcMIPvBXCGxLhSJzbToahuG/4kyO697FqqlUWnyE0
EdBkcqLERaHO++PZsfnPTz/pVbsHttmiTmPa42ZmwvhNtTZhsqFVBjOz9HzhnO+MF+1C5Ob9Qca7
0N97/Yse00Q41pRmqnj90xlf5F2XRWdEfCYlI3l4XbWaF+Dlvus3838mN2mnEjJLrT4ab3D69KxJ
cUXnu84AYonPeibvehmFGtR8/oXGT/ZyVRz8ZjS4HG8egCFwe8bfzUptALeMhgeoFv2idlqhl1x5
OzYbOEO268ESCYEziDLWBJ0Nr7W2OT7PQyLIkyyqWdNl74ewZezVk7XBPECE4j5xMp5cDVeSSOun
L+munZ6llfVATCLfs96khOpHkTP3TeHydJPD2eRlrjp2DB+kZeOt5xHA7sVmavSt0uJcTjxHm7wM
dBgnLQS+iDLsrctjc4r8G79iXqwcectxQCkNNRaCUsnSU9Jmz746MBW5hxVlW/aoNZTMKm6XzuVa
O9r3At0pRpJXT9P1poryhMUGdshevpWMiMaJHNPu5Tdr4G9++KQ0PuGQH3wQ5mHZeDP9/cFXvFgZ
9Edyz9cCgNOMKuXljCFWpfSfR/7jTYzt/UifPhfusDpE1mIu+UIcg6IlQh0nOsaUvUu48Am07eSM
xncDFLTQZyeG68tudft1sjkc7oPMR3dYYd9ZcOyuWk8eLxpPl5aqC7JS0ATVvx85uZ0U+nDoDAYT
GjatDy6gAjMT6uz0G6Fh0aUKzOzPeu6s0hkf0c+bC4EYmpOdh9TBWpQ6icEIkbfvYRgnI0zHJh0/
H2mYGSSWlr9spD3WJVeWjZ3yb4Y84wARZcPJAs35SRIZSE7Gczsr/MiD6heiFVZgW9CYBpwuP7gU
ClanuQLbyeqGdHnFwRZCa3PJ2iKKbXuGsrA+nPTgILmvfoxoQFYysRlb0bGn57wZ5Xr2SobORv+s
JXQukklJ3OP6JWm7LVX86i9wShe1ZFys2e78XyDI590vCyJ1hxyh2yrjkjC8afZMgDb+5/e8Lhaq
FjmHBeaHZQW6gRcIwlO5TQR65ZMZ8l4WONLQTgcISyJEr7w2/OULHK9ypDWJDwFSKIL+0qjzz7CU
IkF3aiN1vzYvZTcZrcJrkFhMzhDW4/v158dfSwPx+eAwH1MqJcl82yb0bG0ehvNBQHT8ksceLc23
AkrRMrOocetbbGva1ePnAUd777ThO0iRfb+ipvbS6vKmx5Va7fh8F4Jg2gwHhLjzL4LxiVUoUTsa
+ytLSed356ZJ0Os8D/tRaQ/wik2U6uze7VxC796kG6S42/cHb+uOIVGz+q2zV46H3h/3vqCdAYl3
n4fOoXnSpl75LWTD1kihWfBOFWY5PlStBH4M2Zdf8Q0DpuELUjVy5+Thx9yIikDKjU667JgXO5gd
0xUodeAvtct2TH1MeKAiFOF4e9jTSFzGq0KXGYgB4lWqmiDtcJMuXkUce0FFi6bf66CyDlJNGBcx
mNrU6J5bvqGm1BGAV0ItCM2X1JNh+hlps4nPvToAH9NfkNLCo/6dJiEewSwCyGppEAB+C4OulK0H
39ubZBDK7AjEH5DXdUSgCQiDOQ726tuCrUFRS5IapeHPGFmCP6XIWaGvAZulPkR5D1MssvuJczTa
fsLVJZpJURbY+5Wd9wPUbD/my5N26IRV4ZisUXXNK2I/rHYInqs2i9qINLSsI/SQLQ8pS8jS3UQh
AtiydNlm2ukWf9YL6DKhQxXXjqqmfBR1z1z/c8CqH1HRhl3t4jZwiiE4ITkIQ8Jd+JqQcNC89mO7
gGBOi7qpkcHRTBnbZTLWLZwp96sJEySDjrWrYElAzR9BqBh2h64dNTYG6BnFNA5sz6Pog/maL1+k
SYEkk2jDrjkOXHGfVR8KCb7mrOz5cz9fW5yHvzQM7nkRs49FJKi9KOZL5eLbcCkTM9wRLrUuqFTH
xsXmViIfiQnQ9TjTcahTfHi7jr7nbBNifBUWOP76iCUhQ5LWLTUZEegurtA5R9YnfWoTIthLAgpM
4uxAB9qKLb0bTMcGzkFk8g5/PBoigjqJxK5wdlGxa19683yF69mZmFuTF4zpByQcXLh9/Ipy52ec
UfKLVBYfHXgW4lTLBjjR+cSHcU3hpv3U1pwE64J51Wc5OIkzrNTWpH22O8pBF1aonJo8g3sKYJ+G
FcaDvWJyL1by+J07+OR8/dG8+FH32WCA77etF2CCR4X1F/pNPeZndV0eSJWWJUclC9bzBNdq1HSo
sjq7kn9VXYsmVwgl17AgLr6vrKaJp1p5ahtBCOOZquchYy2eY/acgM+KxoTMcnWi6DD4BTnr9tot
dd85RMdc8ywELWoSUpv+hgiyeT797OEgNhHE/f5wBIIfIMwWZNvWJpAUay6h0/AwD6ZvBw4yrJAr
uHIqSQeLWkXKZuhMBEbMKAshpofFvVPayymFbzz37JV4719CDj/6nT8SXmk9Lgh/3pn4BT8uT8jv
KL8kbkXFfYqoGFYxt3xnNtw41IEfet6l35YaVro+VjZEQAvTXLZ/gwVw5FcoNzOt0/ZDs5LF6BYk
rDzQieKBdzpCiDLIVNpytlB/ciSVZxlWW31LFZ+fsNbhsNPDYUBS1wsxTb3P36Axs3p5DWv6Czhr
zF6MwX/RzcBVz7yy7u9kiO3ZS2GyNe/GjGZPiS6Akt4AqnHUvlCAfllQmpneyL0nKzy76xC1NGwv
rsmFxxbuetWts3/n46MEgYzYSQSMGor4ANlDVIOCi2Ih0L0bbvUPUlbvoO9J80EErTbsQpuyV8HH
36I3vj7EDkXalf0pVwfoCe9UCFSgc41lTO+7KDMYabUxfl6r0OX0f3BVR4bkMHgWfy996DMnJpdQ
FhdvNxzLTBVKeMDv+ha+KugeHX05vMHOsCYB7kbvYhYxZSkmkidCGUXb3JDmnkX8AUJ50MtehQbs
CwWEr3D6jYdbGOPFELGITaCiyNAfpDJW4QmTHsBANDHorcU8gsbP5e1J13y67PcmI3K6BxqqYkN0
BcZ6FLBnaGRRz7HE2FFNbit/xVO4JGz6q7zdyhmTSDAIPbvVv2mYGR/zT0ROK28jrpCJ2v7FdZ1R
qYgJUsb18xssCwdXnypdcqRyesk+CJAo4fbg+/xjn3VPwIt01N0LUtFoDCRFBW5SNhaEgTVFGght
R5HN9bxx3BUfQ8TfmKsijqHIV0e52qqhQgU9BfyHLimmAqXhrygRR2c5knqkZSkQQYIqIWhc9Fy4
DEDAJd6E8JhDlIqmJFJnC59IYBQPe544P9cLcc9b4yI4HW7ZiCLVq6PLYwRb1lWBBr+X6F41lX0N
GknftttlG71y/IiMKMCdokfpO5hwHDns3zB06SAJ9DzCv3DlP759N/+8T3IrcWNRdwu//7DR9k5T
p/+YBJRj6l1aK08o6whS4hmjPGQ6dguI5MjJ26h5ddqZH8b6AmW3cgIACgjYzeytHDAsb2IIStfb
kHkQ/ETzo2QTXkZcwF+KXVIhuNmaIuTSmDd2Nk32wAHpzMTmLVfyZOZdURqenfcVEW9v907cWgkA
YNCzKtbrs7Rtzzwn6R8LmdtI67fYVAwb6RrX8B87/J+189dxW+QnjG/eYnWHqP40UWjDSOL5rhg4
C9Np8KQfWvOOtVCFsIivJXKGgDKQFMLqLkMn9lNSBQe1sFAcDXgdOJrzGnyjLw31UGstaeorN3BR
TmMCaj8fqXZkCu5kjH7u70aMeSsoq8VGKrSra66nV2//JUSykdU37u9pWfBSTABrk/+NsXzv6DhP
J4k96PfptILTYl4j+RsJQqgxdib9lrEnEuNBrDhq0wXzBlv/j1U5is+w6P5Z9bxPSALJbj2ehKju
8JTjAtUiAaXnU/UST0dzyUDVGZQdm2U4MGCPWK5t5cuNQegu7KQT2Hhdb+7tx9mFHaOmXqQ27FRO
ELLCtVMxTakBZUhmoi17thrSBr6YC4y4cWZ2wMGjk4GPVFDKQw7quUYkLEgnm+nhJDTblSDnWv9E
KIU1EhtSIKV6iy8g0R1vI04BMc/5p2yRmA1hyCj5zXi5Ti4hScsZubRhO0C9iauz5b7Mh6P3ES72
0TaWdcMcTNC2Tn50amXaj7kqTHJdgPp0ktrVp7gKfExAYOXev+obopKIDwYmijzo8N+yaTq0+GQa
F++mey10YAZnwvrBrO0JsU8ORVz3tN7puvOYzZucL9ZyoF8uNQmEUAtJbPH05w0Pw+oy7eLJCSoU
dtW4b3bof6rzuUtFzpUP+NrjtHkn8UvMg1BFx2uciYMm2axaoN4/avGzWeMj2FrmvwFjzO2OrKDZ
MWTfERp+6B838Ze3/ot9OEmc7Ik2t5arLfLf8MyyT2evZ3NpCPn/cA4qes+0zc6EODshwpUijnQX
lz6JJsmFSxd7/ANTFJHxc6Zs8rH0XnxlMKYkeVkK4UdAbQAGnWBfFaYOUzKSW9I3BaGhm9y47t2m
z1U5A3p+BR5uIfILCFh+IRh+aFb4HbxpA+ZpQXv6dSKjPKcs0OjgMPiyG5fjoUYsOmsbtKu4Uai9
r/Mkd5nBTE66Lc2ypCnpdEGSSuokvqU73gsyYAmuHmsur+vGrMtHjFes0ElIJh+wB7+2iQZ0yWSj
7Zr9EQ5y3D11I8+UMoiBRXhs1rZVIGL530Z1fvUZeJ+KqcVQOLWhqYwi4w9+94Go5htLXWwUe/LU
/twDXqdxasxzAhkb3LW0pxj87kFEz7DshukGf2EgFlV2UVMRXuTiRP1Yzp/N68jvqyXijVMAC3zl
XhHlbbHJAh5QZxO6I0peKGCJbi8Ey5IcFRNM5skM5S8le79ITsJicgTCWq8wySuCp6Zq3QxnXtpb
6RzMJuHn0Icu8+/VGN/7L7lgAv/bmseE1LvYB995t14UdC6XaL3kuG7ZoXmdveIdipyIzSh3ddgz
6d1FA6qfzzArCRCn7oK3gQAEA6gOfIL7zXEVjRIJ3rW/3MrCQgvPyKaeSClMBoo4fPlC9YhSpkIl
BjsQimwJkAoUC1j7Aje6jHfpASocnNAIpXOEYjY7ND2Z9XPx58IcgjCd3v+QvCKAEGyONVlJWZTB
cUJHq+uHJJbBMxBTdocktXLsTnpVkRzNziGlV/Ys6Hd1MH7IlP06NV1OxTjC8C5FXT87vWJ13jAU
NZl24+DQ/pHmv99K1g8h7Lw42EaWpCvjMe5d3qFYHpfHuU238latkPRQgfF04n8CMCbsr7rzlRhI
8NPnUy6Tg8g6qKyo8NdYcEWZOCRhS1N49RTyzgXNBoahj039jwk9k/UFyG7CEjY0dtN3nHUrQwcb
r8ZSf9s8LTFFug6TN5aPXEUA+UaQXtna0nKN/B9VH+97BMUmCCOjzgM+1KS59wzvMadJCFewhIXY
rgq1dC4wq8GuCK/YD6zNwIOVO3YMBacuuqlhlNwckEl1HbHa5th++0A/spjnzA615TWzs1iw/k3O
r7LSpjOK9fccbtoIUa2z2+gH8Suj3niGf5FYSI1ePmXlw7TLqfquqjxqxtfwLsS0XyARCkyl6b+I
zdGx5jkl0sTsbRFqo4X6XtUyn12wxKOH9qCa4vQFWtEm1qx/Tk5P938RIUqQrCI656pQuO+uvUBU
9sE7ZtBz4w2rpWaGiq0q358S2UzliPgXWZ2D6JzOjEaHVGXgUu7bkuQ6BpDLF/6BrvIsx64gRqBx
6Xddz5HWIgyjitDzCwc6DGgaGUUgfAW62LlMHCH+fjZnQPun3ZCsXht67+PGkqwYm0zS5BKvyeZM
l2vK1D75FBdErDhglaYGI2E4bWc+lrDfqurHtcUAc9JYBbMJ1CggPuy2KGSlzijUXWyXwecnDob+
YP26PPLYD3FPgkdtVowoG8thxtg0y1Jtd4GWslaYjhttalDRrP853bNQsj7kor+DXxOhF2wT7JFs
Pi1c9ZJTXgPkMMtn3sekfIKt6Yi3p2vfcJpc/z15yvd+nIChd0uFtdKOFKJ5lECYPKMzktu66kSJ
t+VAaMrIYrMxSIdwThztKmdJG3+xeEYTR+mhuOJC3GdlLLzIf8uLeHoLe10jCaIHmxk9Nic56ozi
XV0v+ogH7vAK21ohf4Uukv/uOrJvSJiRu/ylbrd7/nBipeVZjUsGSRCqC7ilfqYQaCI4m5+9ua4q
gYYvDhm9ngnZbKxliNop41e1vZ/XM4SaPP4uUcOnfbqEnn6M3yBiBmy1/8UvgcAqt4iBImE1V0Ql
2W5eTxr2RCuQHqyNiM3uu8TSzhtweMHkQpLvKZSAh4s31snlXwy4Qin5oAyOeTPOgEepz6HQJTZu
GZcF/pk9YX4nWxDTVjmVxQA5A4/PgznqisOmsex+JoEco2xytu8gA+O0trJNN0vM6y5vhRFp/ISF
xn/wJwGdq1g1eMMmHkcjeDElYnJcF5tI5ILeQMgv3TXudMSqs8uv8NGuV/KsWejDVj5kt0KLeW1T
Jbq9NFmZxvDVk9TnMtxdOCJApkBvJrOY5J+4m0L4zhXyZ14sFgsrBxIasR2jGwH3blsdeSCyvywA
QQZBY36lHRrQXDLwP6BCLl0d+d1iwl9nNgCxvoxOZkb7ZNCQaKhc3LadTYQPArnT7dLDLSLV1z5t
0eKX0aKtbLi7AgccyvLE0SvxQ9dAy7fV9Fm/vdjXh/ZxObCiRC69VVHjjU3K29lLXheBnw4wZlOl
JJx7y2fh9/ArbGKHDUvC8NCDuoYh2UTOhwcZYA9f+b9z5+VW4WFJjPNiXQerpcBGaY8iIbvtRJHJ
znE1kaQIJPOE9RLTeKHj1n+tJkMK9dpIo4PlJK4E7kJ4Tln0q87W22G06HW6zN+6r9hdFNO36rS+
DthU1vI06+eyJ/Ogbw2R/CMkU2yR/VFDBSs6vwD/7DlygN4TiuYg9E+orMCKkSqQwh8gzXhKkxms
kD/5UGvmAWvCe6uKkTpJlgynAsZuLM2iqYzF3uSyJikBkDzn8DNQcO6TXtojuD7R3oPdq6mlcTzK
gQHrLQmK5jZeR6+DPJCTe7WN4Wch2KOBNIkPWVPCJ7dHLzsRLUugU7SRNhTCTPpmLHT7ll58giKC
Xo/2IfZwvctSwHJtctudT1/UjTmevuTLMRq9ALvkmWmPE1qdR8WH/C6QgPKrCmFXtAbSoFr/czXF
ucph7hdqvi/KtiiDz24AmxlivOBnrTdRsjApTgJ9ixtdTZ6aZ4NtJuD82er/fftMJlXJesApFJbS
FdenD9CUkd39r8yOdiyq3bc2ExjFdjcY1oeL94GAr1Q+yp2H44IRpYLe4YaSYRr9sKExFN88wnUX
eSvEKxYDvNtxCUT26JsNa3IjueHHo1GMeFvih02k6PbgaJHRN1LxPviuPk36hyss/X6I6u9vkcAN
uz2sZuHS2aOOm2B77OfPQMucPLsCqyI1b/jgHwlakTBgmXGkRluWuqf14QF5pAXLh7/d/x9U1rH7
/wD1xeh4sFIDLtsfWSRgioEscUYiR0E7CctTmcxsBKcmjTUdwk2xzdZh6SiFhbTKF1f5JbPR7ffo
AsMEdFTy+jJop91NZWy+5KK/scIdsJOuXEa42Hb3lz/xU4W+M+2SnBYokbqd9x+UHXxUyxkwblo4
MmpgVx2a3RO5Kz13TmzSCTnkuCf/T3f4TGePQf/ctLIUb4tvh2bcxJZql2eysvcyLHXhWoyOoeig
c+WpDSlO/XK8LwDFGekLbq3ePalRgiOtydixQh0GXUu3Y3Z2HuCgK9hYv8zl+/kXaCq0geXT2aDt
od4X57GBv6HUsvQmXu4VUqn027JeBhQRxJwfsjZeQIEsYj3ZBskAhZ1w4gaU9Obtlb/q/dTZbuzh
yDDVpGiSKNJwZr4z5/oBBI+EZK2RM64yUfJ92QjxGiDhPpHrv1Se+dQDXQRE1PAHXsAZf8Z/2xcl
0k8oPSUBxS7Q0XMk1+awleK2eoEv9AEbnt8XvPx9Fhm+q9q+kVA0hLETxmt6JbxcOAQBwsAMig8G
vRP3K5T3U/tdRE+6UUZUFAZ8/jdGbklMQ1G07fG6tK5tJD1ZNIr0xBsHORHV2vmqSSWd8nW60Onk
UZLrLygW+gg0hZK1sJx62zXFvLF32WIeCrp732kK55d0fIb2NwvfTfzY9vp0OZ+7Uscc7gZAoL2N
OvrOvzAqXlIytuP1Z8q8oIdoWefjvbhwHiMHwSCiIPvhMzvPSm8Kkmzwznz8RzlhOpSN6YOe2Uqb
FcwtLcQCPoVrSW8wwXLqXKJmzPisOHMDem7EqoN/DYUxV4TXIPrfgyF5eE7WzM+9m8Dhh0fTsBo2
i1b+avA48YER592zU64njmPXlieufmKEwLnk2PFoiycHAvYQp6boDednxE2NyBSQyzf27Nbzue0U
0CZMYqLcutSoeUp6yP4L+M5buRt3HQJ+V0zl2hUfoiSGRZVbXTOV6j0uviPKM905rwK7dLGP/R2z
YwCi32aXDsoBx7LycYdzAIhdAqrYV1bxd+3mH4tOCkRAeHeWAX1vtcKFKkHcumlqbp8d5alxt4YS
mBetpx3LBZHn+zJn3PdvxZX9obeDfDwKOB76gmQoa2UAUjVuHmk5ORr47CuoQ2uvYdwQG+iz8zdk
QyshiLE136sODpdVVzMJph0hujs/xFeZ0rSIT1qN0vCB6HOFxpuCgf4oDs0YYjuL6UUChZs5oaRz
/ufoosAdsrfnYfLGehulaegwS7puhR9uvpirFhf818aPKouvwR4o8v7097BvwGfxTldzi7g8axZf
NvnSKOPwXBCZiIb8hBDggUoWT6fM1W/HVSHO8F5rKAW4NNfVcVVkaUD0/y3+MurSLvzf+RTTIhKM
ddYjFAuG4WeJzcHJiBJee4Kt5qPysgJ/1vEZ3lGQ5YuZKHDqEgJdLZtmwKaP9HFK5wdlppv8fsns
lA9V7RWnbR31IdiGBW6A8y6hwUhZDuVu4djCF97ATadP8CNYNtX08zSKgAavKGE++yQdFQFnMhqx
Rgx9EYMx6Qe0sQlEYENXPrC1iZ2nevk9T/OTlliJ4uG473rRE2gVL/bnrybIfLy8QOJh57Z8hNyR
ydKYWAZJa/534EPFrWUOmxhglvwCoBkHbea0fEGY9bx8zDpaIf++DT84WNCIwbGZ/Ai6YSR/jgar
2NIxAKfV9UPIdEASwWHQSMLdzPtMiaiO1iZbVW7JWUfyavut896Iu+U5Ee+zVwGrRetsyZM5xn47
JULP9m+Xe9VwueTog/ap1hxxQcfa9jIGyO17TGb08R/8x2iK/Y2B4dUD/xnmTw5k2DXt+4a3oxcd
RySu2m+RlqBhd2juNjUtqEiux2J+dlTgDtEAPAU8IdgCE+U0uy/hDCaUuvhSSM9Sp//NGHrVrpar
QuT+2Z6lyrDzig2mLdmPlicgLbNMHLoYTZdj2t2ltXxiHx/bBH3MWlimImya4pPqcr80/MZNZPBk
P+Oj+kTPkSp0YArLOyd+WX3JyQ5D8FSYtu5sQauQAjkoq0sgDm5QVfMghMX/ohvVKAI9/JQ5fCk5
uMY5RAOV6VSNQHmvLBDvf6jlgrkUhausG457Ush1nMD9NVGKDnW4rqKgRbgMM5z++iPoudnQD9wi
Qg3eVTc5Aj/FxoTM4G2S4lhAAjkcnayRBdpNqTHiKyhd9TVK80XBd9MxWQirJDdLAnpH7TQ7Cdsr
9fmcJAD5Mqqq0BU5mLXLyrN5EBbOTfqpkcyvzMVHSGi3qxtdZrnxtfUiuZ3BjmjxQv/OgLW7jEjl
d01dRGsTZZJ/WUhmpALSOoJk5wW0YOumgpUtbpov4fCx4nRE9d/3Ix5s8OlAUDQzzEj+2f4NfvAx
Cm+i6HbmVMrsKE5XaUUIAt6Tc5Qj23SWaKEeO/kwnNXLeN0b7nITQQyq0SC3jnc9I7yy/aUz+pdo
Cf6dOj6mNcU5fgltVIqG4N/qnkBis1dfPwUX7xRGkSD0aMta6QeySXjo2IffL4Gm5MYcSWb37Da2
LQMc+uOLdLW9gi480ILcYvarcqcsfo50qgEr1Q1vgdffMkDS2KFqdlqha/yQJVME435S2uWEvXsz
rpRZ1axkp0zyopCr9WJbj7N6UyXAh5SVuQgmRhBfMtTUFiy8brp5IeOXxM3x4qgTTjSwSPHfPq+i
4AQ39CAekwMtGkjMnkUUURgM2AFb0HGupGMLOz6xfozJ9HuGBq7xDuT5jtzLDM7bI04+tvQxYNY9
zA3svOjmVJ6TE1pyXy/yNrRxI6duZQZaUM8ez0A3GfjFeJFzrvNyov4JQybysLkEgfGVLe+DbckL
MCu7CdxFUgc8l2T3zL1Vr/2OsnSGiQuy3z7HIm6Vnojgimmg70rC715Gic7D7KACLCOkD3yJ6wm0
/F8uPeEB8xAims8xXftFDNTVLD0fnlyJ2jeF8HnhftzIbm1l0ZOyYfTSYFigkBX5wry8g5NgTVmU
dv8LrryPer+1xYjNzWv2HB0Z0M9TRPvxZQZ8VsxGVvBvIzkBZSyMg3EGVeDdJg4T/1Rw2MQLreNY
FkG/xhVsKwzEUxUyvHR/7WZ8XYK2fs1252CLedzAN47tYhRRXZAPXSiroO3G6eQvztU6Uh/KzhLg
/ZSyukisZ13D1qLhmbXc6IE83nMo0MALpfmXPCvVV5WHhk+NcTnQz5g2/ozjQCSPqs0Auw83yrVm
R5+X7Yc3J8eeqW+aJQddqdj9VwkgdYOEIBiqhzaiPxb9Bae/DDwkj9GCE5O3o0Vx/CARJBmiqTDG
Hd1HmRieX9b6xD5eHNhplfS+VDKTSX/niiv42vEdVIbwzha+8Ytx67QDskSV8GdC8eb0qOZ9Bo01
KkFw2xE9dqTvo0VofkXnM7IE4BkwkC+7YB11ScwUEVR1O0pl1VtGxNJhx8fVOGIPfY6Ly+tvvWu4
hc9+DC0/JXqif9TVnc6xROwj6e3cuiukf6aszWiwgpoumBAHm/mQMJp69vULb/NqKgzYfqB4j0VQ
pTlVm0Jz2IJkZfmFwO4o/t9WA9EoIj+GVPVN7/7srrt6VchLCBf/VJ/3akg4bhYwR9L0NKVmgoKJ
9EuN/xkRswHXVIKwURFW/bHWfWPG5MUwVsoPEdCqsR/LBMUKk9+Qar6/hV1ZxettqZigxMogE3Jn
1JgwrFEy9gr7M4cqhzFrGsiaQbUQNyppfGTRMhzZpuv+XQw3s9acH+Rw3+ZMpAC5HHvTHk2p7M6O
Ta1J0gwPFAvO4AKVIkhvZYcv8OuRIHMP1E46DpJWMspt4NHjsty033NPXxpvneaGITvXiEf/ekub
e7Gk631C4yucy1PQpWyQMmMYyKRWJnF8zM8xiT9tzPEb4T4aUS3c+ZoHmto13ZZaVytHKor+GtGJ
unMQPldeJ2Jdu9Y1CCiDKQWJ14Ycc6ECSeSUKOu3PZoTT9y+HteHp0O6BQhtswcJt4RbLiEgOkW7
Y05UWZSNeRa753z2yaIZ8P9kGDZ10ReK9c36/T9gsHXVOvE7xFkgNjDZHH9iAorfHzs5ybihyg+v
GC9JciWaRDiKOP9cjEuogUfOGa4QhDt4XD0teabpTWb45LA56i7tbKqAzgVQp0cXvSw408hrwYu7
JxVvNcJlt9D3W2DP8qZ21FIP9F88uaYdKtzRn8UKCUFo/PsFVnfKGPfbdY+5TQex1/46iot5o5uQ
Ueg7JWVkL/pEL6U7VlBKQ8GeaxdQ995p9tuv+kTPLBmHjCF4ynHrpwmdw1oQ7VruBtr8Czb5Gu/q
f+XKdcw6PAKWAaWPxprEq+MGcHnKSa8yifWoeDWmcogHNauqkVm3Iujwpv5I38l4ouRMFg2ksU/x
75K2FyddjFD41STxhT1GPUXhQdHcJ4EFOVu+VJFVX4CMg/FnXI2KI0/H/a7WBvcA4gMl1iJM9XxV
KXvKza/3QF0brcR+M41QGbuqaZ/esUHOt/nMKMK8N/upkOZqUJsgzZX9TI8qGZDkkC5gBXhOPQYU
213Fwf7hzeXobvuJ1EbchRW5PVXiL3wjB4gnEE1NJa+DfRSkwyZXENpAKcshNXkV7Iq3nFb6e1Mh
Avvg7mEmaF8E+REXEVJdlU6P1SYN/crc6UvryffZoG+juvXXKX67bht/saVD5kEmmYQi9FpQ7lej
JbLXvfMpGj/xTG688lYhdT+qaTycGRmXE72lGzINKKNKEv7J6bm4OXIVuVoTeFVK+CJ4ARGcqxuR
6z69BICBqzF98SD08ajpX5lfCItjcVXic+3EwPRiwdnl19m8vMqLkWa3l4qbxoePnCiNr/jT+BMc
1fjkk1FA9ZDHTA8kuUCYxx3Ag4VTiSaHQXMLDhU3UBjeNwYfFglfa1sea8o4qFHh3AJef1kY/vX6
lUx2Ufdh18h245DLpg5YoKxJ+wdAxJ6wz2IRU1Tle0pCeORw2sSu9i9OGN52LdS4Tegu1ne77YpH
d3a7nvkIHH9DCgIqwYp0R3AVB0kzjQrgN4JBlqMGVSqsGHT6P6pmY9V6rHpgjtN/qnoBgluRtQno
/S7Dd/tsK/d5SdFm4hj0Vtw/f3DvLeWEABycXXe9MN7T0Bkf59uJTLRskls+umZj/ShN6HXWH0+L
iHH662fApaNJ897EH8Kqxh30y9XFg4oGX4lCHH7AO3xhpSDoy7v8P5EPqJxpEoaCCnAnXlDNjg2d
vAOq6XfZ4y1RDKauLsg8NiUzalaWRP5LBCt4/fVzITvhh4bWOWZPjh8j9rqGs229pNCfACGcGcNL
U33SxeDbdMttw+jExzpjJvYDnr2X3/qUlWiJoSPbKsoRQs++huMYbb89uDSCJaxOrFWuRdtASyJI
d0n/9BDdZZ14+lBpDldLdnt6Di95QIbJAO5bp34PGgH12etomcVF5pxslsLXR0vlON0l3mR7xvcp
JDgsPhadL1RDa6co+fn4jmrlP1iysR73RqHO1hVlheILHli+OOjuYbaXIfNR53iAA0w73q0qE2H2
vC9CZt41wy5buK+0kdeoE2ezoARj/xSnH6eU9TxC/NWV3pH1xXBBT3qqHRtveI2k4gZsK8gJLFDB
RKLCoRzFjO/LIdtq5XAdNR2bjGvGbeIW7LkTfu10DRs+MHrxuzXmAaABgf5JNOIwR0oJ/OmexdVB
lu63lhcnIZtgzYWi2DtW/NC0m9UsXD+s6MPAnY88PDLgK81CB38IekelgLXvEoNIhbe4qMTDQYr/
HlEKn0+/WtmI9gKtq5OZF3L8AaFSsGu1Sa3K72bFc/Pbv9EK/xlo6Emw2GlTp7a0HFvFt1YMNnx+
GOONWtWihgYquoSKKWnamRXPzXQqIpLCURIf6rnsdUf34gX9xobNNWvgfolMulbgiaQEcXQx7teV
AU1rHgNMikTMtH2iGMB5KLooOM/F73NIMu/A2ipwOItU2csFU0JP9iSnWL2VrHnkP4UxElRrkaAk
U5BglhNd1lpV89QkCCA/deRb+92Q/GXnuE5SHNR0VPbR9MApteHjHFnMKGrQnQbhl+ZCx04c0i9S
7n7YsK7opqEkYBR1qlWbFpYn7yPw/jX8yy1/tgKdYZsCe+OZak72Y2GWmdJqzXTbzAlKNR1x8f9w
IHQLApAWk+6EQ2w3E47Ees/QWaDz29coYu6tVK1oRG+XNnJQ188mUqv5393a9aVHdBjIsiJdjid8
3JDwvuZ8IYYTA/Q245R+HGGgV3oZh+I/BA0MOfQiUSwNDYMBwOOWPVQYWxecI3v4FWxNymVuicaP
uygtlCMVDMAZpbZtA3oGZJ/WgQacjfSN3ZCnGLUfUAl9aQQfXqzFbdb0/lzAb+7H5OHk9O+PZQQ3
/BMA6+uvNc59fW4QhMzakRjc8OZE2gqIulIdX9b7iawWqU4JSpMZv8qzO/58f2k7ivf42rMOxxdO
c7Nh3XW4/tqflWc8YxI56MFV8LVNtZaDWW4GwzqdAJViATx+HJ5XbyVIdEQfQJ4O9fSSRo+gTVNc
WRjtqXCHsNeIIsppn2zb0xVBR6ToP7YPq8Rfo9ibUZb7zRadY/EKwLkWQ9istK30Ffs1p1q1uEGQ
H0BSPH/a5xjTxZly0mpQkAtGT1olwZc7C6yv9oMzfBrqAuldDZrzx/sHz/B2hC0w6zK+cBg37T/u
G9VyBOLUZDLF+D2OgnN+uLtlAAoTQICx2gn/MJa0b9H+R0w93tIEZPjiLC1w7YTxNS5VIsax8x7s
Dz8SI1BmcCuuWGEDbOTt4XxXlXlE4H/oagsTbeoD3k6Z3N8+XTEF2lV0CkbUU2kPSwE+Vs4FDtY2
QRKdHrG54KKAM5Q8WHgIXON4MyxRlk5HmBQAFUu57iV/YCi0DtegOA0HbRTYn1aJRUy4TcArV220
jo5L1DTXxB5mzkU83ttWmjPV+pBwDz5hu/tLc4oDbEX50Nr2b/fwAEZDlFCsvoLDOlIyUinY8DfM
KOw/U1K2ueyMzlF721dJ7mp6owp9x/FlbNfPaS94QeZK6iVL75+ntQ5bqya2wDWmzuuvuin0Whnl
5d3EM1Lr82bXQTzSXFMwyAAnNCZb1sQTabJGF/mrbSMFkL7BFLXPMFpqL51K668zzU5MaxiAjFbP
1QSf9cl2Ma4xsL/Rzxisylv5UbWGr08qRZ8N7tQ4ZBqoDBtNZ6i5kJvjG1e+R6low83SVqOcLAbA
Z1KPy4VGVls3J5JnfdLqswyiPlkrdJqEhE4AavYSpoTvNHEoELxWEfJYHT9wDScPSsAxR+5/Ly9e
F933ARyuGncXLbCmyHl3h3vBlBY+gSa4MJLduDq2sF23SUZe+OXB+zI+zZJL9BHLsCFIUDj9Awjv
Z/QPaR3358eKq+/Re7of7qDJKV8/movuSeWFZ4f8kk1DzVr3Sud8NQe4PcZVkIiW1Ocfnw9H3O4Y
6Sgm1WU/Ga7SDa5bHXGm+G3yyK+mIEh0D9T+aRkAiDKamvbmha7g93HJipKPn6J2CEBKKy7B+eCj
bS+Nq34nD3lEuRKlXfCnxV60PS7rmDm/MYwuhDKNggz5Z15SI9du4nDpPUWN+nhuEXLUL+6kudgF
VU6NbAfF3gsYp+dGFR2eglwh9Hhj0SkdSeh70ECGwHW98qg1efTiyQLn2bmBrlIMPYoWp8jH6vXf
wQVfWe1znIh6IT/uF/bchYrxs3JwijqGTJCy/nytl/ZJxCXkP9LTEDAW8zlFnZylgWNMqUlJlDZS
Qr7wdPrORxvKfS/gChLEC4dS+Yh6XM/lpu06+Y36/QDOtOA1Ax5F9T2a8vdo5lcNRqBfQdmQeiiq
2jZVS70UrrwRO6Yj8xz4vey+/5N+3oTFkrgw8PvBJfUyvi6nKRzBRGnoaiSBXDmxG8Sc5W6Utih1
47QJQPWJw7ik/2rmBnrv3Ga4PniVWNNVcgCHlH3cR61LORQVUTmkAsBs26lMv4p7Hu4dUR5VyWnN
CicxHwZ285kEdwcrYUsMfQcxp59Mvz0Mx7yp35v7UpXruHKRTo5PUIg0P7h4Qz2gOAaakbEfLulK
zMrD9BN+x34+eaaNIq1/vf8QYJvlEhuZhfQRsz9tKB4EQPt494xtC1Iyqv67uGQfub2wgp3A6FIz
za6IAPvgD72tGmK8U/grwtDB9boFnQ/qniYlpF0eQ6o9weeV7Y67Bxbzow1LbK3VC2StZ83yRWk5
JHKarumbKCb2JARoaCe34qG8G9xJrMVXHLU4gWMSUKbzJ2r9HM1yCIkqxJhHljiPoG2qPP5nWF//
4FGZS0123AQ1h3npvucysGqIYmNccaKA9mfxsh9HJduUEZbwFgfFCDfxUQ97rciVKgWm6n3YYJvG
Py2UT7pACHNBdpZrQmpqv0zkXWQuJiLDmCcj8qXNXOQA3/28M6ho4Wf8GEkWgkAN0BEzzKz6vp9J
djmMidwzE5GmDaCHiDOoL7/yhaDVbOc1RPMBKTQLoQdwnhPzGVFJqU7NK69IW7IYwlSjbVlPDnsj
h4y7PFV7pY1CTmbC/ZAbMK8XqAhh2jy8SYPAPmJ7rvBGaEJh1ha9qkKz2eK6y7QtheaKA6ZHDxG7
YyhNbE2FRuFScoc51d15NPdx3F3ufrNV0vLpdcZmg/4JrXPciY94QY2dmTzoZmjmCL4g6rCoeRxo
pzgr9qRFZUWZJkdHa75EglZ1F9puuEF4/U22QfE0tmB96mPxcfg2Upmugwy/MZvpcIQC77d5mbdn
LbB12EXGFpKf6hrTKEwhbZsRX/ERcBylEDVBLWrGc8lYAm7OeT0O8qDZXzaeO3XpGu3n87a9xJWO
17ww2e9mjkGCRLdTM7phVVUseXh5diz8+PN6yi85WgwU+Pew986BBZoj6TF5FSPe9KME6bOG2TTP
Ac30bWF7JBeVQFW43rMKlOL21PQgRwXG2STlDGanAVloErT2EjhepTouvP1YzriJeFdHubRvkW5t
XbBbD17Y313isgfu4ILoyEn94NSKtJTl5pfgi4eExlLywJvMBwqM9RUxH3vp8jqLqA5e4F35SgNg
RawOoK/CKWxx8YCLRIDhQZ6aJd6FmsjfV0Ud3XgaLX1q/zYvKmJAp0XLikY5PdTiAb21pT3BAwEN
ujGSzcCNLDgxcnNj/7mZDTnPI4P+BLr0A//kU4eYn5gyd7iuZRW62y3nmaW8HA+SIpmOB/iQudZb
Ui0stM/6UXTXRPAp5yEWcB4fZ6Uh8wUUZk3UnIcAEtNTCJZBcCJvY4ZKK2QeNtJWV9L+F33/Ge6E
p9Nh8TcQPvTZSdweLZg5nJ8KR20j39FEliqvzdUirqrr73RNoznkzDJlaedXOY1DAay8VnP+vuO9
uxkWAW6tq+/oXencoJFW5y79BCsvHK4O6I2ZHvHQll2bwIkQefnLLinX+idZWP8MWO6kIiQlXmVA
Oai85z6pXL5FgKE2I2DErrUESLCN2RisdIj43CXbXcb3Xqy4bKHcPexVFk0QZBzveushYvinD3gL
n92zWLAbH1askpbB+H7U7jl+AZqDa7hm71jszo5VMSxN8xz1Ccr+ZllSMrWePx5f0SOGDL/Qxov3
7bAK4MEYuAhFYKpFGtCfAGdRTazPX7QUD0hdpKJOTVAFH4DI6TzNgUTpRvAyr7cGe3il4p1KIAfp
VKnEgraIpqfIuCfEMNhainqxmxu2EDDZ6HdKsTzNQxCWG40jM1gNhMaV7hx4XNvG2IHSoyApsiIn
Ps/0TEuDxWMUoXVTTFB4RhGmppTbnahDwdvL48o3YjUy8m53yfM30B0OWvIVAkcBsNTt467sW14W
wy0kEULcnjNmyuw4JUJRft1H+bZeurpkhofKPnZA6iGpBqiq4+WDd3jk2xtMvNiKgIMddzNsrTYw
WMdHIMoOS994MqjNVfVn2DrpiE7/Bnb8e0g9SHnbYSZ/NmfY5efbAHwWPCDFNP8qT7ZFmzzzIXSe
V6/TZN4FkIdzl7g3ze+GoY77xgmGocZuvTePQp5Am9XbhIW16a+K3Kck8j7i7ua5/cTAey9i8eLU
FNApVNN3FKgZyuT2nb0BlC+pgY95kp47hC9LtAZ8KiVaynQsZkCttA+p0GvajoXX1lIkJXm5t8zh
6JfgTlJuSzuDNYclfHn8xThD9HsjZ0iDl/bhcUZ8lhj2Eu+1FcOPHHsdwE63d153cvYhFg8i3lZA
xk1UIlMBW8LJEzMkRIZV0GrXCspPuWzfSc46wm7Pv90fGf2AgTmmbV6hccxuuyPm6eUkOvP51/w+
cgLpyyzLr3ghWTQuydWgjR9kGe9VrXMnnebH74DxWdHW6SFmarbspW4osmlzqD1uNvWtc6UjEHix
1WOsnMjfGkjVsCpk1yF+2P6MuE41wYTVzQxsxt5z2ITtCUu3KxQwNvtIi/pIXi0l9Uu0dLWr9s0r
p/vBXpkmHYC8MLfZ55ZwXX/VUirr92zTrbVxsDvA0m5uerkPMLBnD0cXgYa5oYg2/50qqRn2uQAg
08iri8M1KXfGsAZvRsCiOwR8F8iVAaznjz4rDfTq/HMKurQrwhZiXhKxKKNybblOkicmq43EZPOH
QBpQxXnNqR9kpnGT6/EFm8HxjfGEHxyyniWfg2BGeNYvn6xrvUuWxnN1pzXZYzY6vQ0FBYigzwk6
4HDgXI04E/rUOHibWydBmPnvU3vx8v6hpUZtUOdtwLZLrmNIwwhzEkN8OubvPG1KJOV0GnDAta3B
6kSgZKMQULGQ2ynKHF496SMGyR4vKpCp3AuD3V/ZN5KIGttFxiOnkIylwIWjObdE+LFLNE60T6su
02kwFjpSZ+ANAKl6RNU4nLNlf4x4IbJ7mFP0LGOdNwebFx1Xio7x3JErC4TJ2q3hPXeeVRhaE0UX
uYif8B325ruz/pks8ZuYAvSeYAho6u4xN41SUBvxbzE3teGmECAXZqztpiD/Bkp20/kdNpab8Vba
ZrvnhXvh4f+RAdBYuUAaMt7s3t0X5Y6gcE8rzSHygDpSvzkRhkA2pitJ0GTUrC9zYs0P/rZwcTGf
XzA4qCdH5Jvny8aDTBKOJ1TcRPtaMZiWZXvhDHI+k6qvmtUemOh9ZPx7ZclUrsRHDLut7MTa5dxI
kWwS7PnHqUuuDRI+vKW/7whxsFZGFaywMRmp6Z3gy2wGeDXXspA7pwb/0+7sEENdyPvFngrX2LnE
hPmCeUAZGYDWtsDyMip0BOnO8wiasq3KFb+ebKzY3rzlHzqqGQqQ0LsAY0SfYc9IfkjJtuE9x2/R
LxLF0ybYL6+GpQeB1fvkBmdcJHZRxlyeES6viVJgXtpJqDTRPtUA6hw+0Ns7eA6IJfobi9Bfx4Jh
ZSY3DoL0HNyHBH7Dgn0x66ueVCl3e/RjOyRSBWozSQatfd1cVKe5rVcjJIPonyoRN0gEJ59A3LlB
t3+Dp099x2Xg+KXzmVhMLwS6N6VsvohYDZwkX5XZPhLMrv4XHflMPSfsX7sJAyH2osmsZv7yVv4j
7U9MtF5s0Q5HZQqlWr9fYXaBEygotPQrXfHTf9tYClAQzMw0mlzWAP4dKb6MxjCzRB9XBex1zzTG
0hTbdgDR5osCz3Qsfgf3hm35O3tg4xAOYsensaKWvzZr4+Lo3bKfrOnhpj430bQ5vhCdrZLt4uMO
C7R9TpXPvpTWZLONflNyW4DcaE+OUrv6MvgwciR9rqTHTEqp2tSn6cvICDciuV58aZsX8EDiffVJ
SzGlRcT1sODEo6CuOwtWebJ9J1bCCcwb/cUG88op9NRCNm+ycjipqCALGNYserHrgC32y2JgYl2T
Nt7I0SCuI8auOahsoiblpDOLBVjc+XLbrk2Z92r9hBP71y97iSjQAVcUDkWnpxPeU05JqKuWdLq6
f3lIcYw8qnDo2alHmcdQRCTs9CuR75sbhmCmU9G2uNWXliFibDctDAvJ3wD5bW4LTiuOK46tEa7M
8GTowtomF4v6CFHekWEhNboP2VnJYD3g/bJNvM+K/vCrTxb4FC4mStBE/uFkeSpyxkRNXh1uXZ9y
7Jo92Uz/FU+Vqt2upraFzNUuYpmeNWqu/j9urBn4HDwLVvwAqDz53Ur9E5kKgdZRUT5vy+v0zBE4
RNf8udgGWhzmN5v3l+jXJpI97/R8Gd5tLe8H3ICsgaJ1N9aVxP5hMhov1Du5Sq5uNhJXaVeOE1QK
gngio7qUDV7l52FK6GIIp/E77HBl8bSPvecGzLFHtBIuPA6D99llP/G5aLqjLNbubCBbWrGVTbBM
m/IMrzdR85CgaOPzf4Nvi/Dnu4QEZo8+fV/Z7/fnhGHi46Wbg4BAXkRFwhkyPvNar+Te3DwvfQGR
hUkRH8koXyUqN2f3aXaZbz2Y5Uacm6EkYwr7gBQl+OJJBEWkNCljvwfzFO7NlDZhnppN6NEO32xA
6ONfyAk0YnWWgyYU6EySsTgsZypuj2qEf2CLYnodVRyRSzs8IFzwtIIZQClrZD5Ui70yKse6vsM/
7ykfLFEl2IPs5CgCYExPYbMWj7/L9H04vMCx8bbXjALVAgkZETWUAzuX2Z9oEu9Eb+jLFcAPjihl
I5otA61gm+AFGaHsFQ9HE5JYkbtkhcqoCy9I6r6A9lIDrKdpDROmcmwdVLVBHt/XGh61m4I6ru0T
/jWvCrAcJXTrHSxNocWC9HK/WUFgyY5xu+N1pnMTcxXN/gAlII/JpVADBYu1Lwg8izjIikn25QT3
c7QhPkYlb+9UxYEKkJt6lQcJfn7AhR3zO+xbDtZSn3qzBF9deOj/ls5io4NrieCkAnkMB9oyamkW
4nCNaWW3aJwyQinJ3aaawoxlm1tlUoiFfnCy0pN2iSsvSdDGNHHT3ru+FuVThlG5I3V5SH8Tw/gA
Ea0tQyg5qiy4Zwg/S4/Ulwjvm+53vxyDJXLQY8ZOTGtv8Fv3gI6XHuEXn8G4gH6EQ+HEx7+5i7wD
rcpIZqk4MfquUnrGiv02yKGmFW+y+aGtYkziE8vO+PuuGSReNIXPl2Tb1mJgXWoG+jb4dhmjBH8W
A11tzVOslzdoFnNiWWrmeMjdsgf1cSaHGhgnpO9RXwV8m80P9xcV4gRnGAtAaMKUhAOs6lYldaki
34t4JPaM/QWYuxAb9Wog+TJhSV0t+3cEw8EU9TjD+7ZojPBFtHvCc77eApikzJUI7gocu7sUSETE
2YCWvDhmwHvKu6+8u2VX/1QhidjpjfyxBClONi6/wsWIZ8a9Fy+kidrOD3QHWmuMfE53WQ/kZbbA
AOOCY37y0S8VDdMlCusV1MQThN4SCsUERo7HyeRSwdKsqr3RwcqPZI3lGQqBwe8Knv2n492Px0f7
4Y8APAj2GmgPM5EaYegZAzMk2W8OpEzA+6JCojroX2W7WfEba3KGSRpcZ4t1HdLs0hO9ltrW6gXI
ooJrEUHzeGuROkAstTibxHiIMwaBD5XlJpZ1kjJDjKKfF4G58ecnehmm6I5l7qegstOXlUZve/Ns
5k+sS0PHIVuVMftz/u26JezqSCCOpgjs8/uAY/Kd0BL0mQLRQYmAED3Auxn6/g2Y4q8W7ZyQQMdJ
ysMtTttNBgqPSzMxezpkpg8QSAO4pRntusZg8ylpXjnCzCAxpX7uz0r8wiUnmSiUlm4LrQSQDdzH
7BlQxlCOiQm5GhFilQYayq2UwSDAoDG1LNiqU0NISbyP1pHS/3/XHUGeWkI1paKXWspNjaJCATCM
TwBQrYDx00EZTk6GY91vqyVXqHGUQSgUDpASBZUvQHC7Ivl/jiclAxFhcaTHoJc/MC/aDXGzhRwN
jrBWlrIDKcm1Ifzzo/fDhM+JAudBBAODYKT1CUtr++q1nAxYiWFSsRPP/bJ3cfXKa//VPTctyb45
M15JE6DIXRd098TdruUyLDPkGXzTJuCQUmHRVupZr2vt4/L73FbX32IlDVeLOwR7cTCPCJP77zCG
ZmeL6NrNyq3rca2doAtHbCrCF+6qP7NGfA6LDMF7DAQtgkJqORhUNnBDRbped+4fGXuMaIjURtAg
3tDjZmxpEIrAIqAZLaYXuerrAjvPL5mm31ZPHHddrYJvaBii2tAbqWXhOVltOhgsH2px/LedNtB6
bcqye9pWWMUP3nlbU6UZdwIT1xY58mv38RAvKMwVzANzOXwdKRhRmxQcFMu3Y5orTvjShMySjKID
ibIVuZjb5XrmS6yw0u1mO1vIzMSUvbjq14nbQ/Q/77Ny8/oKnaBKU1H8SZ/lkzZo3K+7apKXfwIQ
GY55SettP21ap/D8pkJeFRtf8HQiJ+tSXagOcc2IFfPMv4yAqv5KiXxUJQ3c4bGMWtOXsfMhK57u
dsaSxjT4gV7/fglg5DHSa1MXB6I1rcteFlyosem5hNpJr20+ZsI1ZGOzlg3tJtdgzLNUgIl6rWXk
9tw4Moz7A1cqOQP26caYC0oLv7RczkJJqgJqcAeN3/PcOz1ZqlDhN87wo/kuqKm4iOjFBhJFERmA
q7xdVPfHZBBWn+Hqhpxt25v+dgtKQrWJcXZjsVNtKOop6MpNqzYkfWF47rMHJOo2+AK2sxmYWT5k
mkPvLgpmoU9ZrSXvXuHoTR+voJZraN5np5X9LXv79fOpOn4izILOF1U3DWaxR5an6va2uw65SGqb
zn3xIPv0CoRDEqMXBiAP1qWzBeMaCz2bhgYpZsp1o7K1qjjJnGzlDsb60Ol3I5juud0EWy9jDPD+
f7ytpq6+QUBfKiyv0w5UrsTnNe7wdaH/4bAI7Db2AVfhv6w/XLatcRiVK5kNg3T7Z3SdUEfKlEzx
+9bI+4+FmcMWnIZO+198dWlK7Dxweds9A6ARcqbuYJgfakS3tqHRCStNY3S71UKzq0XYGA8Z2F5d
av1gik1QOz6MLH8KjDtrYiaDimN0abD7X9Iz9PNr1WzS/YsZxvnC690btRBsyqg1AaR6hPv2Lpv0
JjVOqA89yf4njZcGzQF8qy8O40U6LWQbT8IMHQQMwxlkb71QlLUB437owzMpPa6BId7qyKkh5qrh
6gwhnhvQIqV/pvb09odcCpkkwAQAdLVB3SmfhIGmLyvg2oG7YmNQJRVnF5apbM2gvEpFccpZJweF
VR8Ck2AYWssXMCIE0fMwS/v3ODjBROssnIfUZ1JJ7Ydz2Bowtqr27ZzQEayPg4x8pFbgk/5IHMsZ
ItLa6zlxhiIWkyaibxCuQojjb/uxqP8rbm4hnBsoeCoVxRZ+x68dYSXsrNHvzN5gvy2MUobUXOTM
UjvyAqYtJ7VsbACQjQOM9lmGSDVKjaez2OhLZaAVnVgYkl8NV7lW+4ichAunBzbfbYIaHSzjfzRY
xySX3r/agKLw+Fz2v9il4S7JX9steiGXqcLSWwy3Kne1Mg9Ez7uWTpC15uN0DtonS3Zv+2dECcsV
3iuTIRGs2YUVejMgRlBruhKU/4QaMAMpw4HQLkDbUF3hSCXRj7KttxOGWLXxN4jzwQ+rbRU6Mg3M
HB9KlxiHUh15huZVu88DRTKO6tEU8CDh6lMQLFDqTC8IX0vVLwmrpJxdKnFCdCiVrDBVTROpzxU8
uiEhatKhJ9dfJpBJhSkHjlLNBPt1EawbKN/cZHj5SYFTsUQXoKOFcnvt8+5q7vxQy+LDg5UxWfS7
ovxIK1BFTis6kfK8yX7ErQlmC3fKNiWVFYFJKdTsS/IFLY9u2iuCfFcY2WOKV2PX5+nMkTTRU2Y/
xD8UKHKsMG/bLd0R57Dkw8a/KdQ4W98G71/jYXQxAmO80gXaW9kPIqaH7MAAtlZRIoUDYXfGKWyg
9PokxOqD7RxC/JnGZdGCM8f2GUxoMkeOcXVgP9Xh+3zHaiSFVf31xA8bc6ipKFMZxjVeXV+Sx/0F
95M2DA0cnbryY+yeBcAOniu7zzkm6twB4dojj++a5BGU9f2aDkfJIPNMZ1dduLJftZlZPBKeWfcg
NuzAoPvDF5bFtAm4wIfR99MoC/KHfRNuKN9/Vj4ReTe0VodiJNNJt7+MGu51gRdVoBQ8/l9/1y0m
FjZnxDKBwqUCotoLJyIXaRtIrz4SWK74EhzSIchJXUlHvH/fwAH20VTHcjZvXmkXvE8pxor7GU+E
ovHYQ+cwdhXGDIVI2Ld9stDXeCf+rkZIvAHKxNuRFotQlSmQGrUETJ5Z1tY3kmEcVAMn9S3hK67N
A5PfcNsTT2QPj8LcgloZSV50Ja1nhFE7UuLRY+IDz40gWa1QkxqhuY5568eVodcRBp/sLQ/cyJmy
FA6lhA/9+6txV2D8/VNdEfcMr5wKHeSq6pcyn6PXBdRG5lZObIxXOF5fhkKACcxfY+O2EDM0L36B
mGVY0W+x42rScFyquH3y7Nkyr5YG5NaCaNMDmIf2gPIzPQeXUdTVcKpJVQzX9xKLosZj4S3xlX+H
Ra+/drLz7kHul5gKedUx53jWAiRMY6Y0Dx03XhlkxW/MkGIm010bmywCm2aNhc5b7Als9B/sFRMO
XHXwLC9Sx5kpZcEu6SWZzskQA0OGFZIDxTunS3xm8YjGPlrDOwFOd5Ayi//uA6JhUi6US7pMxdPI
4PMbqFJAEKWI+exj/Eetop5ULt3nK6MdVkBdT8BqOZIO0/AMqoLgTTRK2IcBq8TcKzYAJvazsAr5
FUa3iXzs6iuPlHGduMqpfDb/SdKHVD0WrexLROqdln6TdZifbUnKCOTQZEMhn/tzLj1eCguKe6qH
5MyTgbuNsUh3oylFkaFA1SBrxUe13k+oSE32ltoAZlHEwv3fzlm87mBGscTexFuxna7/JWI3JOZA
DxC+TZOWWpu+HPgQrUXtc+uBg/HoMmLArWjghNinf0f15jD4iJShcq1jJJsfGqHUq5c6B5igmW1t
x/FDCDS3e9+6hAl9c+wc3RagLaVsEBdiYCokVb3HeZFTtOa2G3g5IAcZsYj10EkFFpfMios6H6/o
miM31NEuGIu690CaqwI5MuFQ6qtMhqilBEeL6FbNdzbgZcx8xobHrq9zF/33VtEgr2QGv5nOfSJo
29BAftPmCEuxXANwc9y6XSkCDiBGrkgETUwR+DreBVZnE1CuO43kcrw5xlOQPgwKe5OagM6Oa8v9
YmmFXgW5I/lkMDR8ODzjffJ1sYoCe/+nwou39W/AkbZDr2UZaXrcWU81MZ5Aldr6Q1HlOEQJysDZ
GHhCrGW24taZxgXjYkxstd70/VGE2rTl5G6IRjLV3C3CDgUIPMaR6DZn+8dkGz1pxd6i5IFM6p0P
0qgXaklfCYY09T1UNDF9RkJ634wm4V0fkwtOA3oMjWTMwsZA//x2UZRuryXZEoca5Hvn5TFekScz
LihTCNm+gvtPaJLZmnvjL1gebfr7/F8mmGhrmLOP/2tkJtj5wQfdudW2BR54qVMrE4ataEBVwwdl
zHvuS1f8vKJiy079fCm+Wxcr8XqrZf3C5OdFU8I6ZZmUPOBRG8pf0+zoX8ssLKahB1jl4kqyIhRf
uo5daGqI6kTmrrvmtnN6IHpKTcnEs+c9+GanycTNak0qdae71YU4PVFc+CG3poIpI+311O5AcowH
8k2AMu47QdyR9N5XeiHX6EFBVV2jzJk8/9skpRdoyYEa2BM7bmKf1PZ4lhJ+NrZlVPrrpfyB8FyR
G3NQjG08hOl9l71Z3rCAvFK45Fbg8f8cQf7fmCezfGOGmy34JPiBdtvrKnCA9j+9rYisRF9XeD94
w4mphnmNz5TYRZ0XmzF95WMYyOKEcHdSD/NuMPGv7c2PGQuRMRsPwdDVlmU9pnL396PHGZOS1a2B
KytxH0USyHekw/bRlIIc+l2JLM94WbsifkArQk4YOwARNcJWuDAucVdhXQMXo7lstEk3253xOKWp
Vo72V2Og70xGQ1wvKAh/ZnV7LY9u8F8viGuc1AQJuslqn852PN2pFW83kdIQZ8K5dqN4uGl83quY
Tt7CoBj41bDj+Ip0nicy0KVkmpEnqeTMkBhvPXjzfsOZU5obmHOgAvY1arUuW50WdpPeGglpKLpn
ZDrh3KuIx0ju1h17UGtYh/tvos0yyB44/Pmu7PqbWcYXY6vv123INaDTZ0yWGucu26/FkRwaJE9E
rIAdQz5KviEtmt2hvhOxVah7DMnI0/DoTwjXPsDr9tRLHbxUdwUV59JIp5YflEdL++cDEzXsM5Si
s52cCm+zb6QtOvMuhpzAyFxzjvdk22SAvt56eNBHi7QZXiRyJoveyjs/VzicqvKXp05AY3B9HIRh
U0T3WehGjaPHXEFsYtX8uculzX8ImtM3Fmz4jrOEofwvbO86PMCfFVprrmuxttR94fyIxuV9HfIP
D1fGRcbMZ919k+OT9uJoI8R2WRubmo2i2ZsRtYG5DnlD24CZDYfQNWrMw96egEDYPhEGbfmRBjfg
DLTcxkSrJq9JQffOypxbXreGr5yNVwp096abRYRWLPExhC4h/+6WY0pS5qab5v367byh0vroIoU2
eIVMbw6z/V3H2KP3Cro0K+ww4aC3RUQEkd3s1duMq/htdS0oHHnKjTynlqFQwoNjyMhmSL7oQgIB
VE8LVrGJie8TSXHL4dWapj/0R39N7oIbRTKXS8dvU+5G3FbXKCD/I2ix9iUPiQNylwTj+vpEJKLh
S9fzIatanq40H3xCy2L5CziKvfgXHPyosYgQnGfXYBjFJJy1JAgpdMx3i6RInwvw52SWap7jwqrS
88uEaHRnQHlLFrLGjTCmlL2aalRRW6FYI4ty2BTXudHUnlTfHZO4uLIbw52vCEKdCzutS0CxkmEI
QEH4ZQYhgj1Z9bzZA0/5MtZ8NIepfaY13Rec1KCCrEFr91NNAe/96PVSSfWDosuQw3hj8f9j9xZu
BEK5BVbOZmI5vw94lmyQ2dDkIEHyGtBxJ8WUnwjdUAL19IzwQHHKbvGFpsIdh3bXv5+cQrYaSZDF
Ad51Qs5NIBkCTSxSlpkJdiBLMV0/zO/0ciCe8JvfVzMiMGLZ/+d30Ugi02tQ183crWN1k/VD3qpx
pqoD71gkyjazTTSN0f0qj58hgntjKGqICVMlwkIdQE+oP4Kb0xibFq0pAlSn75Fa2W/SVA0/nTZh
8dphp/yrUzm2Hil14xlopd2/5KpkynRtSBk62Ne3tJalcm2cVflbnfhfjIDODDkGfWqyqxJ+C67o
VtKSLvNYYicnLd5vtQJaB3yGa75reJNzgGDOAreE+CEXuXlXKa4T0/a0lExKcs20Rt7sSy6NijpV
BZgZdOQjb+8UY5Cj2t7jHweZw3ol9cMjcJwNzq3gB8l7h0i7atm7TTnNSQBzZd+5LR2yXlsmGH0G
FDV0ISi7D9s/RQzaoVJNIS4ZNwpzsCwxXwz/nWER1nAOtmI22qiKwO1BtSdPJlX6M08aDZd4CE72
viHvo60lazBhD+yuqNfCVkTftublvdVZzPaJlPPIdv45IH0wvi75iKQp1F6LuLZGem69oYWJuooN
P7H/IT0fXIRBzIwadIK/6KlQdD0bXP+qzjEfRtJT3ooaiPEextudA0K5WistfNLyMMlTj7Ogwnpe
4aol2uoj7A9MDES1SPwA/SfUaqDKuOGBGJjrq2ZIMoUNXuh1Q928ptOAXI16GqfuQpyjOV6/PCWy
rZK0mGKjQpNKtsysJj4Rof5duzpb0Q7aW0KlB6RywAAAJe2qJ3VycITpfaf5/ct9Ugk8/YE/jsuY
mNGVpPo0NP6qI5zrddZEyauITm5DBS4q5Sue6drNzNubbJ4BkojxOC23S4cu1Z9L/al9pwLRFSUI
v0bxPHmPxd2nrL/ww/NM3LYZklExXDjxHnwWuYeWfkQ3OCPebDPFjYOGXrWUbj4G2HEcqe5I/oGa
u8ukdLPb8GLb8dD+Yphrfy/06ttLimu+P4VUWVnu5rdTY3YjRPcN0LtNXq8ahIvk1DlQiUFX7cGH
BFrUUs8M33su+Oe99CtKfyOCBU3lO+b6FTJ9CjPMBXGKF8EaBszy/lK9XAE4NA1va9VYShtbzWyy
rXBgeithiN54ZEOUy61gVMRIKba/k2t//Ul7tUES3vkxzz9BoADABgaCgIr9onxmT0msx0rQociZ
YycJnkhShktzYcKOID6NjJNfa/d9XO251Yg4OLaq7631RDulrNFjINN03uuLrtz69JfJ9PhklEct
uPtWEvods3187zxipc6CB/ffSA2XYYpr8CaXbJTv9a3d6uPcDRujDOFXnqghEiqVyF8asNUITfSS
uacpQxJqkyOYpIfk22ZM4/lQkoJ2igKve/6wflJuUkyX2L1QcnF4KpuFHUmcICzUBDSvLkm+ChSK
de7W/pgpTOEF51j6AoG9oAeEDha4Vd8iU4mB3oYm7s/SxQ/eLLXjhqfD5id9XCWrbh28H2Ed3eey
JgAXUK0nPZGrdMRjjNUfgXz4WbYJRrFxiK0C/YVnsOAjqShtcqtg8slXXkbEqNiJh7tvo8T7vgxC
gRXjPJNrDkUiaD+EXMXq4upAouXK72zQpNag9HAKDUTxMIffQNzIDBD0X30LaWvCA21WSFfvHxjK
oBJZfEp1lpMQLvvtP6EuCjB8TkninpTsgzd2EYUn18EGrpeHMyNkbNj5tRLceVFjj2W4epaFhcU1
NJchmh5f5OclX4AgCL1FSQPs/JE5fMwRsqd55jJsokhqHPWnY1qc+gVKngGk0QunAKYnScgeCdbZ
sGAE6gf922+BN+0QKC+yqd35Qp35MAbO/CvlVS8TPrhy4eihexouRwyLAGZAcoWRGKuJj3+bhUln
HJEshKtdbRszZHdzmqfUlPfn0UXnysiUwuG68n4hbL89IWDoAJ2OnsIAF4HyeN/z6Xu5EoXE0KHs
JUbvusanjWjVrSxWOSsab/KHy29J1JsiljvHlltht6kM1hQSjaKQulf+2Y/P4I9ydXypze9rtQoD
g9a6o2fOU7eZE8rJHUCbDkD00agbLsF/ryf44wcNpd6oZaM3BKjwMnZM3e5tCorIHz1DEgY4oTI0
8oKYmacOwmud+nqOIu45h6V1XeLaqeJ4CxHiLE+zm31R4V1P5Jo2IRta/XkyZdVfFLZLM4NK3wvz
y502F48yfSaybsFcn46WOK9ulpXcSkyqCE9jzi/F858gTxS3pisbdbgpOFJEgzniys2cn0Xpot59
Ym03AYHXt58xD427ySS11B1BWamzIB185boEfR1Uue2L/ruwGIXs/HYqGbptnMb/l+IcnyQ6LofZ
V83iD4OImVimvzJq2piP3AHXAHJof2z/p/7ASLy90bxKLN3uksSkC7AvoLbz7aKxobfJc6KqCmxn
0fS6tuI/kAKbUPuFBuQdBCL1CTvDHV2DrBUj88UfowY5CIR+p1jwNkTIHOTfXC5kEcCh/v2RbD0w
gQu0yvmufp4nRfl7Mz74635IFdsw8bKYa4ujXSghYyOXkeHZfRwmsybkKaOjJPybYNkHizCmlmAs
//IMTkLsikVs1ndAtAo/H4ZnSNG3f0YuhEloCh0sjKmPUJOWooz+92m0rKtUl1UAoo3zV3+flf5O
sBaZJflQb8dpHCoIoBcMxW0A1rDfYlFVWBbm9Tgzhg2dlh6O6JJgrVwMXwzoAwcR+h1R1XNM/zz2
W4sB+5AJWq+dlHBopH3d9W72O8GPWZke4ZZt/wgiPPLWuUOx/UKydG2gjEh3LMucOG00ClO8YMT+
Sr52ys1Kp2wEiwtXepAd9mK8QkXZEz4aME/bE6oO/PFrws1BznS+6XAAEqph6jFJFhtpYtLN/ERU
na9kJ8/7K/SI/7A/RfG1d7/n82AvMKBV7QivMVeu2yjPzYZvCeoJJeVyr3Hj3+I3C3CgBtq+8orR
iigNNcS72+4PZdJ3TVG8HfGuWTKeqMJZG87EBqb+170wFbQDVkAWq+fAkNmDZkaCx8+KZzw9kwvx
skwOb6uZHksAnLZkQX2+EkNJlP22OY6pSNfqCrtgRBIKOjcYbPmEZkNTBUVsaD1tOuX5C1yAdmd6
f+J1HG+ELglAoKpmWlppFJrnsltu4MampWbEVbE/9ZsAsXMqdyeGIRfaWig063M01CVpG9WjhICy
6vvYuCfeXO/xwsODEMFLBA02f75t8yOtCJF6x9nlwAyzsrnygyjRDhG+hOYxokJ0rDrkKN7eJdK1
6fts58t67CRSvopCiVSl/cerS1CWH4+Eu+L7H13KPeD1G8OQLwp8SOsrTofFptYeCRQLTK/K1Zh6
DwEY+9RruYcUcVNuZFt+Rux9iNWGa7+v/3kVG4ypUMW0YcmQeqfkrLe8kn1lFOVH9AGx8MVog6qI
L+5kJ9zLqlmAXgBiku71FBkJu1KvdlKRGMvpf2Qks01ROilAjZTfeNFquG4jIS0JTIeaG3F4JXHJ
RjmD49HFU1L4ZWXj1S3acimOa8cUX5i1zKNuC3WPKOJqvVXXT9q4clx5i6aKoijE5ABESfFzTkYd
FPjQYSBTpP4D7xPQCuvF6Iy5e8v8OX+WhysvXIqTVDj5bY++D4TdL4aYAwj2lvBYZrClUGH9pSoL
97RklTWeL1ZJXW6EuU+SZ/GXRNBC3bsjyPpVTHRu14+/haCPFB9K6nciYqeninqOghMdkv7uGenE
j4FdulupXkyme0kllnDWlbyWiAxopYX+HiU5ZRW5qweFVWG7FUps2nnE01HQnr7LJdAhaGke978W
ckx+HxqTwX8yfUN3ctKyxCRoM6eqSCRZ073Rtzwz/teN5NHGKUezbOvkckBHTB+HQQEjLwcBVm6X
Z3HYzIJSCT2JBbDOcG6vfXosYcej0Pm4oqmvXBQ2gj5u+eEFbHxvC/8SYOinyENtrsLcu8/9pAoW
kL6X2zsKeqBI7HMfNcn9nWTFQowjN2vRrhDWXF8KRPEGO/DLX0Qesh/EZyzZfoJfbmJe1IS0YRE4
DPv66Tk7FtUMigz3ixSOdENbbJBY8QtWyxCVuMKlH/kqqbS6tmZDFTP3LVwyuC7ZkFvuEiIktqa/
avTmM86RyK+yQSRqkadPOvQ+Lwh4SxeegLWtqqkWd3IWNVp15iq7zYx/Hv7nPq9gbLFvxSs1EvF2
w2q7FuwHwNGKpCrMQmcDRgcqzoMe8Jyyzz/x4WKKi0/mp84oXvRWuq1sfVFpkRUjuZUL0N5k0ROr
NigI7cmlOzmorL4vRI7JqwzF72mfK8wYWRYkjY7UZ7B+RFgo37ZF9/532ZU3YP3MHttFEsiOZdOb
dJLiIkGBYimFkHatvwA57+WzzHIhAqPOnmUmLXqasFpeZ7xnmNm1fai/ot+OWToVbUnpbjAImtHJ
5unwDjXUQyLfafaD4jOKsZ3j5anSZnarWlrkshIbDhMU9l/31WIdaUYNQlIJ+rSLX8mhHK0gcIHy
J1Mn4W4gxrInm7Jynx/lBVJhoScC0FPyylcAQK5HEs6KyMQBWNmHuvl17M6rMwYJ7mZswqfKa0pI
fPgE9JawTI5MCWW0ZUWenbNnByW3u1LP+x4Q5L4xsYfduKMV+AI6DJT4EbwDIeZIxJGXcCzj7nJ+
DqiUdPOFiHDOMPeYhh9HHddrxcQE4oGDbAm+7nJBFeRFJByhvl7yQghf8y5UQj4W+6yDB/G5dA+S
QeOgYpVOvkAsQtv5YveIS1lABk5VpaT3bmWeMUrg/GY8w4xIv0nj5t7ZoLayrw8Z4wX+1cFaiKug
OiXZOIiVBoVdtSXWnuUA+tz/04Y1p8KH6y6NkreXe7QaajlpVHB8zQ/BVVtAgmrfhWF0RMFraK+Y
cqLsVVbV8dD7Fk9XTSt9KoixEG+E8WO2WAnscPjxal6SdeBDOjdLl/ue8ueHoMK7b8HyZSxGHxJ6
h047NQfYF25eXZ0wZZZGG9IyuIzJTm95zJMyOnHwL9tz3Smhx7ytFVVw1D+9mrVCLuVVOWBgm/AT
n2wCapReTCBy4g1+/BNd31Ej6VHOlO909DIER2om+eLqARpw96mAlFGTHd+dEddJLpPHi40sNBn7
RCteUA+5pHqJYZnetqoLLNjThGNQKzyA2S4Z7HBWPYI1/WYDI/2SztddgU3oLc6yydtbfq1mcWle
cGVwTwdtjRnlrcMiX3HY7kgtDqTbhP0mOJq7fDfHL0CLRmHnBKbZCEKTDJ4vkCHjCWo1KN3M9HeX
O6FJ8yjNUPm6pJJfSKmgZsNK8Ym78ME419d9eMMQXmSF3Ykb3KSFMphyi7XOQpkevgAu0orlofwE
h96/MuMEiN5zYHjfdORWLM3DO2WIXOHLCxcUB6f90JaUDYQ/GJoBDdFKB5HQKi7c/oJ1vDzob0JJ
TuF4CjdxSQPVBfL8wZie/PwqkfGNDUk2yBbNg9mVQHGKnCu5p1WqoiwcpG/OjHzEgVg3kQFqXAIW
vPk2n+PfzUTMvMw3XiV2E7TfBzJPJcXZXNEJ21E2sHyEUYOMJBMEaZEpqv3+hsCRk6yi4LMElFTC
QbMqbWGv43algggIKmuaN/Lr33we1NiO+pGY8I5fhxfWu46iB2fhopW9roPlPybdMSd9wz1dHwk2
8FFqOJVLskhOEptHOkwzwfiJd1cFgJCN/E/ml/c7HkuENk0Upx4VQhxPIM0eqDd/44U5QajPXeej
0jwROLpBUhUwcOcIR9fjTfvKsxKkJ2NE85G7vkKmhdVu7bcp9I7sIUYINPV1TZ8NV5rTunrE+7hZ
uw51YY2Gp2ese7MELkZjQExJNNHjMNzz/DHIU7z/x5cEsmJgOwPeQPn1wdV4DjwciyFhn4DKthJq
vppK2hLluw7Y7F6o3xMgqgInnqXu6yTttYE6kf/7woQy1x7054vObYYcdlibGkSM8JsXbjkWnEcv
BdHhQfAyDRTEXgnrKF/BYSZRoMzxifXaYzTIxlueSKPkxYcmWK8GspwOiqE6iA/9tt6XDYSfZXrb
zbKwsfJTMe59wlH9FeX+C20hgBUNLLJy3LIl/zwuzfJHiugsBkhUnmimgaNukiV41jbOKx9jTTkQ
PCYW4u2HczI+ZCXAFP2Rmt+Y0cWI3xJzLJWHEkkaZgxIeeYQT/bx9psjuiGjP4YREl8b9UZ0BZ4+
z+mpZoAN6u88jdR1SZTkwIkO30y6DWXiULP25FReTMg3ojKYfhRPSCpUhkPJ4FGr0IL69HYQcl1C
JfebM7FlfI68xwETizo3IPFJzY8SH1qmpdwpSDqBKmWxd91GbuRA2um8ouPSGpn6gZmqooYCqymy
Oh1zzDFjMOLNoY1VPEMPgIdNeulq+/fAmAF3GTpV6VNg8Qqa6z9GBGBjpmSpJz9FYLFSr5KG13zo
9A7vta8H53WcTnHeYu5FCiGuBuhIVGWlVaNvM694AEiXiJAnTY/92qBuS8ejvU/+e07+0Wup5rmp
8yZFOVcFMq3u1Bpvs4zHAItHSBvyLmm72ZzfPrJDo+BET1rd20bjOVaDLOG0tQ/JQxoCQ4GnnJ2E
RlALE3frwFNSLnU+Kz6cjZjkIgbg3cmaI84pOPruR4jY3JXQCWVscJ4vnA2Uc6tdDrK5HXUWOZr8
3HWYEq8EP3W4JXOXtpUL2tEkvjDeYCAbwi5rGB6UJW80GrwvFhecXnGVqoT23wUwp9SJEMsejS7K
YqnJb1RlYMiYghJhAqTDiknswp+vYFiOyaXq3cDwIR/WDs94WdXjW76/7jBqhdtyeRahu3dS0SZS
pOy6MCNMTkCiTQLIuA53iq0sO5464KIcbudog5+ohUMnU4IvYROCuntn24GCctNGy6iXU4ZrX1/0
+5J3yQY2zWb0l2wYnblzQQYxvPMfwC3B2y23cIwEQQt6hM04uzFAVtgjZofuU6QSuCAdy7NVUOki
gGmBPTtoI/ro2mkqvBaVX9EKi5cJU8YVsEZnQ5MqcdmL8JK2wTbXc8nPb6Mmp2P/FuhEG50WGH2y
lt1xl4UwSXH2GlHIgmKAYRXQrYS4BrYywzbsGgUSF+mxtdz9fTkAHCOl0o36am1PiRUoIGC6M6oL
UMhbv5h9BCXeuVlpjBWxEoAoOZc3fHp+DwlnoGEsnzUoVQfMVDC4C7c7vlznZ6zInoTS3dbBgJgn
rkPPRRA+IE2ER7Q+mLY5bsbltWjRvyHnS3zxhvbGuz6ZN59tAaeyNG6u+oArhw2+se1dP923/78K
TURA+3vDA5HwU4ovnZlfkhn/SKF+M2YV3szDiOKW3D3PqAb8N/TusM57w7bj7D0QbIQZwAjSv6G4
Jd/H4byM98Mhqsmr0krXs6UfZD0eGsQZZErA+dVo2lhGnggFjI1GaWb++UMXohcLD8U/JiNBaeDD
c7zogUA84iOaxezTRykipbzx64IJqTiK1hDt3VoN/IuOtyNiA7BhPEV9/OonS+Yse97k3He1m2KB
j1+nYsxERv0G4r+lvk+JyYpc7vQV+mSYw5/6gbY4mWxyCJKBCCyyJHymj95BfbGJzt5VLkxA+Yqk
W0YUikutfG567eisi/++unCfHd6dUHMvKOdqwhGiOkrgnNQozI1RqA5hXZW2rVVsOg/CtDZzps2s
C+/b5FDMGLScY7dl1fisQsN+lv9bpLwDmuUc6NProa0m/jh3DJf1dtluOjt9yu8UP2uVQobqDuyJ
GkUzh7/vlruB4xgOKZOlqXKi+dtqjZNyVcK6zBwtRQ7y+Zx2h/MyyAJGSEHrdeX5zysWLBYF3F0j
hU5br1vdc+EXdnGJ52/0ZBvJDL9Rgc8FOkyrSeRhVJMgTIuKegW+qaJH8xs+DEgRudQYupB3X6LM
alI7WpYrvPov5jwb1axY7q7G4K/hFCKRoObU8tepGNu066WDyo2UnUM9iP0JfNMT/BfSu9r3XgWI
S+acXp8OV0G2kF3PZ69ONq28eNb74yZ5r4+rDqHhs9W42LSTDKKsbin8l/4UPXbBShfR9YsO+DoG
jbPijl7LI9s5/TQuMnlCGkuY3V/kSAk5emUR1vN2h6MMcHqvvIdreveWYTsvJdFyUKnr+Bj3BSFR
yfsDodBW6uyk1Ngedk/IUGFiaqAFc47SuQSM5CPVIQi/kc2XxNrvoEXiPnfp/goZdsiyY7Eo7A0C
d6P+9sfXwqxl1sLkJCimxTb/Fc1qFiXQNFN2vFtH8EIfvvWrXTI6wWMgbQN5OVZmgaZTN9iIDbtf
yvUnYI4ANd1cu2fnit9CAPmyDrBH9sLa0oC9tVidksOnlkWb0VJwJFCLiktuJdj2oh6eguXH2saN
TSv0kTPcfWc7WKZ4En4F6ckH7uZbbbAtscTTi21KSa6uAokPFdbnGqXUsD8gtaY7aojyWl7eJ+Ac
yQhVuujLMpB8KbI2xFvuOdBzIbboguv45qeXI+X82OeBE+8Y+JSlF5/ylps8x3QAzFVNcX5elUBq
E/BZTXLTBlB8Ci3OUNAdzsqfaXoPsCUTDfq2JCdpRl1pc56ymtAAT71R1NznHjtGZRcAKuJdzYKT
ymkf/VI8wTnV57BwChcFEKre66jQ8+GWKZGGx5nz6GLfTGm9inau+BoYLTklGiVbOY2WSHOzhfpb
gLOKqvB/TpYMJJAsPFIihnrpEULlnZJh8DpV1ZPNhGmFRNv8nivuOy7PzpBhBPdvnyyNcQ0rlqzH
qUfQCSgy9lW1cq5Db7P11FbY1s/uk7vE0Eum9GOnbf6yBaklDd5emJLjG++G3kNCi4/W9p6QqkNi
IJNw4tNzB0WaFXBsFOUKRnN8nUzpP+JhyHQVCjTs/BEtnkRYPvPXS0KhCCrQKlCYiWBXBpssYPPs
dBlrG/yMMH+CGJkFdREIOAoMRs+xilC8ZOW204CP9MmswjArv63ScymC0Z09wuDbqD5ZnwsdbXPD
b6S52dj8LKpHJLleGgSI3kRRlUubolvE0EE6+SxNxKSxtDoMdr2n1jYVdyBHeJ6mMGecPsX1hczA
CnDaeyxI2ZGkaJdBLYeY4ct4tLKY6NXVDw4APli55xtLet+b7yeC90ozBvu6Fa+f/xt5w0XkwN2k
NZNNHg5mwFpav1En1sdGq+VOv4Xxze2rvawEmDw731cG0EZAbh5aeFkUb651iKiVvKHLolUwVnQh
vlMYfHSOmF/GQ0I3vYB0gwLa59zb1IqhPDI6fNwQsxj71L6zuq6ESxmnD/QB2oyQBb1Q/Dr2nzfq
W6c7XCAAxzEASImmHLUnYMGr0ooY74wOazMiyq27VRQdWheG5407/Rhn1hCrIDxue6+olPzVJA79
Awhn51WMCkLzsjRZjOygK10ztn94cSySE+ymrZHUkus7NLplpirbTDvbmloOL7Xl/Eq9DIipV+Ee
OPIaP1EdfdLjSz8Brv0hDM61K/5OLKLwN8RS6JmK9kKH6LL+hOWTHIJIVMcZhgtJatmi5L6qHxgd
wpi3VLRQuYPfA4Eqz8ntcO+yvjPCCdVAUW1Mht7s+cx5dpGAeFoPZ99vAIGKdAvP/PsrEQazkhBt
zaE3gm9naOQyS0VKJdaHAv9ZiAtx1b/k3l4zDsmJiE8a52M6/UYE3oRinX1wYydNn7FXY4cEzuQC
bRzar53Wgr8sNLNHoNsu0IbqG7IoB9Qe0gkj2qBeJAvONCAiyhyH/XXn0KdRnHhqjMmy6HGJhY3t
EpnekvVYM7C4quEU+JYUKwqQ9/mxYYIa4eqCVFNVnj7WNm5ktptXRROjxbUODxBIFe0Y/3Yz5qna
HbNfOI/IlE5EpId2xejqApFGpZtX/iULpQJqNMdoVvhzKBlGTcBfOWnc9SL5xRD0Js0mEzKYKR+1
uMX7DisZRQ0OVK9+MSQ2wAjgRrMIwrQDXwL62/iMm6VdiUukKBwm4dz7lSGtJ3WmFTOb6+6JjKWJ
2N/gHOn4zdaLlZfujmWiNykeLuC9lzHMuKMw/YwUIEcXnS2MzogokX4a5N8QC0vxu1sIZ0PwG2LK
2H0i5nrM93C8enJd1rTOaiMNKdZUjxiQdcJLyauwGz0yWDz17vjWrwsRevxiBa778BmLzcwuYOwu
JgEc2r1To9+n3wdrI/ENWqMgS7lQlHIE4QR76Umi1GXeKVrXGbh+o42urLTX+VAz8Umy4DqtQi0y
wSeP9vPOjLIfL1cLSs63t46W/97/O4wEd5R6ka+U5iPET7LGs77jMo5k+6BROR18FBwnCK3TGNbr
TQdikx9R1YCHDaIQ7iyt83WRWdcb/B52UOTmFlI7B6nv2YBchvB/VTt6A7i2Ew7p9n91CL8rbjh9
YCdO1xKeaP8eKvBe2kYWR/JAx95YqhptJAzj3Ozx9xF9PYiDLwTrUs8eXe6eFhScsroTBPpvtTFQ
BKevGi4DR91jbtINB80rwHbJ4ITOKfo3JPEN4WtiTZtlK6r2r0JdWujaS0opi/AbQaRlpCqnIu1R
fVaWacb4WLdcBihWEfcmAkVHcgwvIxwSstS8/cAeuPNNCdavzQ/61EY2f6vw7+9vneiyoyJs5cha
n0/iStekYnQlGF05BKVLh3VKAprtUGlq4Gl/GJ0pA81cKCjkmNpZRIcSW0TNzP/XVEx+Vd4H3Wae
qRexEVgqLV8fcGlxmue7otFuyGBoByl3z6/v3vfIUSknhwIBTPM/6v39kmEQnxLU/6ShIFtpzvn8
tyAvTcnu6MYf+rAN09l4FuROmva4HeZ9/qEV28e6Ha3TO2cJ6ivUT2kaAgfKbThOAAgteU+v3LmP
N+8heKnt5RhKV+6GRxs0AXnhLulAjR3Fxg1knsKTmi/Zb/LEsI3Oyd1VFLRLgSBPPBqgaHjvVxYy
qGnmiFBji0n+iSM2zbRuctOuGmTgL0BKjvrEwNaxf+Ro0+PaCQgTPpiZPQoUAF771h0/tgSqeNhC
FIodjFXse5VFV9Yj33ujoAVSfPd9i+q2r+bf2U9DsTcib93dPYs5fzKg16ga8SnyduiG+QWKC/72
zYDV0o06ECXraKkEgAnngjm9Zmaq2itANxsIKFi1uWdlxH39Le5O4rUfYaw4QQEmuLHBJF+JFUhe
f4hbUs/EoiDIMqF5HYaH4vTjwkA2eJXSv9SufAoajmyStoj97T5HXgf/o12jDg44o1+rKKtPDBPT
A0BB6BFbAJ/ViTAxwgNSvnb6OIXE91ahjVgiab74/Ml5qE4JqoT240AerkkTCLfN5huQWFhYU415
92nmNG3Zh7CV3m+irN/4QxNZypbHodtWAZRy3pxLg2Sd+4j3bNMZCAp1yARemEv+VPOettngZOx1
CjHeQiBJu8FTsJOurLSW3SN6sUNcvyVXGGZkzOmvvfWxY93QrFlDkTNvdwz7wxE8mxaspsVpjX7c
12V4CkHqivXnKmpq93hr+7o8tTZ+cO6cdV7ljTG6Yx7TMoCu/JFgd/HIeR61b5QwB3PNY6hoIYSm
3aF6NO2d9ybUBM+eI6Nbx34YnlVx1gtowaaI8PJX27qSiwF9g0lEh+1yvhgIoc281O5nMD/F4P+Q
3NfIVw4Tfb3df+Qreqe92XGqQviJgugEiJmI8QraWA+AsAFhOTESU4HvJ1KXZSxVevaLB7AV0kzq
ban8X6xZ018wGP15xvPCfRsXUmgzWxuQiFhtvj1ZWXbWdYOkbDqtoF9EQ82YL0zPel3GzqfOFLUA
2ueIEMx7f7KRgBEOaysJUwaDw4qQAJJXR04bHCd3Tz8pHThGCub0vppfEE+QTtlMmoVl/LOR97qa
/v+x56rd3JXKJhj/m+YCqp/LpPT6iRIgNkVD37OGNZVr93fhri0kBcSGRxZNNEGBVg/YfDBuZDq5
y552U4hwjY2EjHBV69GCrTWbC/SI4d0iAlYp41qaZK259sKZCQwPRl1MBdyyDoPjBYXFCngtPyeM
79Mqjqdw/xVyuIxSqpxzX8G1IE5mJgwZmPilYN9eHc4Q/YD0fV9IrmINsTwbIYB6aSAWYiFjeuAK
ZHIlglbExz0XVCrjEAvWS6hDTy/wZx7VIKjo1Hi2QSN4yjFoCSe84QgQTyibDRV8+lhnOwEzvwW8
Srf0mchqfL98fWyR5zk0H6N1oeDZHhHJmWRlDd/Cg6cHgDujmrzuMSQ9jD0lUjrxjCDXaIfhsHPV
G7VakuYftCn81ci9VBSaax7WIgyyiJhhEdEAb0qqDplz8Rntc+WSLOyJVZHVLMWIm+RBUodEo5Ih
3ZHGtnYVdQvHewmo1X0v5qJ5lIhzWLpf289s8BacnTVz8VkrWB3lJD2zp/u4EPCP8W6keckTIRgA
5k6ITBJpeaHZ4empgHu4KigRksVkjNrqhEeQR/qW+nAb/mtGbKTbEYSvZmgf/YFwbtKt1hlxANxv
8jt2AuOaYaSbJXGiQiK6//iJqyRldcPLr9MAJDCqIhxvH89m9Q/RuXE80QHW0w2v/I0vodAoBiqm
TNggw/jMDk5H8nRL2i39u0vxwvi5s6L9mwBRoZ1F8kLqphwF+bfZ3YKasSCkAny3v33sH4Pcufyb
d7di12+qM8ifqOBxllen7iCknIDyAHGNVEzaFzx4Y7M553YWf1Jzp9NoN/dGFdhdoDlL2DAMCHvw
gTYbyQGT1P/XZe53cOYrsbUQTtw2R3tanePWY11rOp7KJAUBGY+jCeu4k8i991tiTn6ZJSRo3mAr
VHFI2A77vvU2bSb6+gchRIFfAFWYmWjvgwJ0ciXDNOXmpdqm/YfWrHNSkedi2Gd7dLNq1/V7xISI
sOQTWQrG8uA6Zy4gqIETwgbMVBzBlvkNQmsXKlIUfNMrdROTGI+OFPcA+CSKRv0OtSIp6zCKtYbV
br+i2la7LtCiRKo2kjlToQTWwUl7J61wcDiFz96MGHA8PKwXSx8tBiWtBu8WQlUvr8WRnfVC662W
bh2SwH6ZjYvefUB/iCgYwu4hMR2Yi+IL0CVjRTU7LH48DSaSvM1n5mljvs8fX5YepCvW0+b2FqMX
OewIQmJVbuE2hZ2KMs26R62qYOSlSqdUYJccNDeQU7SUxn9XW5mReAz8GCaO9POi7hCZm4CCaCjw
KcKT6I69N07lLPUrtB0yJbk7r986FBcp/CNFjUM5vndBhDLe9jcCT3UADNn9FF7ST+D3Yf9Vp+w4
BGEhX6qe5YWwBXcpw1vvr41J3VRTJxFid+d4Gaz3sYNL9LxdHe8URPvKYky43wP0DXAfxpJG0/F2
xBsyUqxMrXAW0zbZu0XIckMAb1nbOZ3tVA9qDglZNw+neluYVaG3oT5zvSMcRtoVjRR8cS9hPAGs
1BRBV940JR2OmFdh6Ffz/9xncPDUC5lAHJnl+wi2YxA1oqeMZzNz92ctTP6PA3YPtCkX1atd6CCJ
OB2WT18GDgIIKbcT7nT3lXRB7XdC0eTCosnjLeEp9yjcbxtN75EpLwsaTLUze8APAKezfuIaiHWW
6/G3zKyzZQsW9wjQUK7FLTIqmGQW1L278xjceCLNYUH5SyfKFY8lqHClTikwx7UqmiQJCodpB/K+
/KlhWFPMOnC56Xpsn4MAaG2BGu7atLNPGZqd0yxhch9XivtKvmFDx/di3cjw0aNa8XG4s6k29eQr
a0VbXF3GjGwLIAbW58202Mz0rMzss36PcpdRr7/pKxJHk1PE7V1rCCIffkUA/Fscln673ddvqF55
rowZ8xYA0rWAFkbPhttGUHN3vIfNGAZWiSAEbefwVwUsOySjEfMmbqu6QxqJGPFnTM70RdelfDT1
ROHVusMfXERwdTAkqE8GuWcBWr/DgsdGN9GmQXNyFhIfrPGNQdX4tkwUSwqlJD+NGmldlKwXdlvE
p+bXuCS2a15LLc3D856KyGJtT5hIgSbuZTvfxts2Xe+8fzPyzEvMQEylnfJkn3l/Ovz58Dxt9gnG
30UbMTQ53wY2TFmK+aBTlVxJMRKhcwen3AEBSBD/48ccQjcxbYszQjb2xCaBbtSB+rMRkDXBKm/b
AN5aXFSlxdZz3kKXLTG+Rfojm6GOKeZE3sF6cfBPWdEAQ4Jp92HlEsQElCQ7S7ItakRqdM81KrTP
EJUg2c1ard6IIPEpKUBU2ojWFgWs5Z6K4QscAH5wVlV55BMcevsMDTInY9rO4C5OhB8ejm3c/3/7
ccWt8VEG5fOVxNfJw4JpuxfT1Z8ofiiro8MqbVTJ0xMdQVaKyS+NRXV1ySd7YZA7i8fRSoYkt0Op
XRMWIfa3YEocVxhisLcezzTXAZbqUCRbsWm0vyP7fKmae4yUqr/fNW9QMqLZd8Wcl5yWURKyYQ24
6gN0hz9wHroy87Jt/KwrN1FvBj884mBzV58yw/uDlcvaUM2XhCGyN9EpumjF0nGTdP1lR811D46O
WuxYMMyY34U+6HL4EKyisTLF6Fd3onRIKgGOcMRvCHexkbXyninj65RtmhNO+pP4nvgFUKqLuw2U
gIEnGmeIAzGxb0+4jeUikSorvkJh4j8aAmfKWozTHwI8kVeAiB6ysJfRfkiK/TGgUES0P89vmoyU
CqHVJziWfg4CyI4HCkfEiRhvR+1YPOJn6v3u0RfxZENfTxSA002BC7EanzJAJp7p6BxRbEIvVHwA
sHmoMgP6C5xSX8J4DvNAn0PPO0YXWxZSQgj+FULFWMWKfkOWKzSo1gjYCUHJ7bq5htvftqJxzYQy
O00PtT4CmB1waVzAV0VQSerz3u3/7b3+7mIkKY5WgYdLhF0kVIdsZQnxKctZjMdG0E/y+v4evoDt
bGI6S72rhBfyFyyfB3779u9jC7M0B5EZFPqpTaMVJ5T42312kVN/0f8zDZavRBMnTtNIbLZ41JYE
arQbPHWkxIZ4be0G6Wxr0vBXsFxHg81QvYfC8I4w3+Hbu1bssl/6DMWltNEaq57S7KY1SD+2LXGn
YfGbnumBRdUP54MIpanax/bP0OOyaljpdfnb6OQ+sedU3cWMDLs2vU3HaDavFzaR9djN7ZIVmTzK
8jmO94zB0HAXiSN1q5leths7/oMJKywZOzeH5OsZeTOuRLBVzUT6zhs62GdqxMsTJOEss9MqHNG1
P4nY6obpzQrS6OD3rm+2DkWgkKhDkonSyjAtPUSpur5pddq53uvQTridavb89vpWBZchlpqU6vI3
HyU4xOviKqI97lGej0qiuJUbWho/6a7t2pAWW1IOAqfzkLQl9QZavwa3P9ncVmU5mY3n71WzJOZC
GlohHFO7irA5n3pZaI3ovncec/uQ/jUgyn079IX9aff4nG4ImMt9RG7J51MpKFJSH8jEX5J2jC1j
/sCm4Pj1u1RAwjApqkpatYR2QANRa1n4kx9QpbbmMuW39uSfJBI9AwV4hJVjfRcL9b3mIMm7IwsK
Ccy/cbmH3W1SnmDD31F4qksA5INc5s59rnk4GsgeQ8c5p0orTYwhIkyZce2BpDQxjZfKRaLwvhbb
vTPO/WQF0ZlzD3qArXv2+VMDdu+QYb5yak1as4yQfsGp723DoOs7EilSbM1X8/MbWhlsD1Bm8WQ0
V8gAVC8MCUj7bk2Pd2HG0Hed3I/wj1anRREKllY/6aEoBDdaBpmc7QpeYXr20aHABQQlQiJbwbiW
lP8OsnXSRxj/BTK8AFbiB9e3h0rlGHBjGH/vt22nLnqDMQmhnT345FldaQume1b19ODI3rR5TGlU
GFqLQymk6q8to7PU3YrVRywJE8KJ1NG+VnGsBwGqyIKotBNmG9YBnhlEyaUAySfa8DtUPEFHjlLe
JU6UOxx1HZrjKyYO2PX30BmDYabdSalThofZEpXcYLtMzgPVw+WTYfomLJ/TFP+5GaLCbdw9rFgZ
2ibaxnUuSrtmoqOeCXEPwtV+pm9YbppdxHLpFUOT/dPRiKEmCqM68IXwR/DyS40rX3DAF8I7bp+l
brYuxma0/OBN7sQOJ0VdjnlS0thLBaBS2Y830vyURQPaoAY9Ie1g9bM41ntL2SBVRVewJSx6JE4U
2RAAXlKFhJyMx0w1AKR2SG6JsTsSW/cLYxLZ14W8NhAdJhjVr/bcmx2HJvJQoPA+6HPX/Zyt7Xaj
p7PDXVl9rwm3Zl81Kbg2tNcVuuECFfosxY5pabRPfx+K/P2blvjKdXprVCKuUemxSaHjI1LwI/cN
NAwis0UZ8xievx8+DfAtlH6vGrE4gMzadkkWDnj7tCPjYtGp8AowpkA2L4h3AvX24VXHwiGAq5VM
xt3Nqa/gGPcankKKD7hJkkMsOHM6O85+mVxCiEiwoTCxQ9KsIy836OAFHyevjdGO7AK52RUVJI24
VNj6lpbv4WQ0dc4caSMZLga9nX42u0ZcYp82IvyU59sclK26335VQSnBgWNDmzZgzhxqQDx0n5ii
3es790MWUWpQHSGRVwWRBRL54hpSY0RlZ/7PWYjEYp4OBGV/48fVrhvDXm4H+SPTAth3We8YRDSW
Itj/BjIJwUoT/TR2HQVjINxZUR7C3mI5OIKi2JOsGiUO6CUs784aYu8/YRnipbQlzpCXYj6mUxDy
Kev+yqIG15NFl7tYkRnoe9H7GBXTeasEH2PiaztVDdwcXmxqGBixD0YqtwlVi2yiYzPjWLJ8xfHj
cy9qulcwr4HsTyJGnGF+BRe2CRNhPkPMqiqm1dgDg22Lh5ZmCZo5jIU7YJTC+STeQ2xqanRbi3IL
/pM6iG+yIs6Lyks/8wsbBfoseHxk3PezchnC1o+rTYROXoZ4Ub4hwxlKVGfgctWHFU35REWRD27g
0ZDc+dbATPnGlf98R2ElXQdCduRk+Jd+4eTz6LFUuUMjJh4azjLZz+KXbHF3KDOXsj5e0cBgYzNS
fVzZmkrfyHe3KU6EoEJa4Gqv4YffX3BT9AqLt8tU0Nun1GLI+Oi9PjoAXd4mib9w/J9uLjNne+vq
U6uCEFegl14pIiZP68k/k5Jpmvk4nEbBYy2KVOpp7M9YZafWboHeKqiUdm00up7NhIYmOaXeqVNZ
7XozPspwlDd+hIO/9ukHZ6maar+dIfiPG2qtVppYcOo2W7hYD5emra4cCffjKYu+pN3Z09O2bBTg
P+MSM+2uINf+LP9n8666ORAevuRJy7IfGDNl5SVx1/htdkgct1rR73UsdsGjuuRfy4bbPxcrypsl
rM6HuW5lM/vT2KyArMvUggBDYIQkEvSCIUzP025NIbr/3fpvV1fwm5N/D04eWpEVV1M5qrORyBTD
8om+DDP3DCoV8rAyS2QF9oSvO6m0XPLTjGLfRYaOz7g9MpL8Z+MUZWTZbRgSyVIzSCsgY9FnfpCw
YhJkwiQrcHh28vF0Ugf+EUXkoFzpgzku0KUMBVQgtTriaa7iB0CZ4FTbB8hYSrnilyjmEn4YoX9v
LQsoJNvVFDopR+m5EV9VnuYG8Rhw2Hq4cfTrjV97R1ps75FG1CMhww1B3vxRGQC2uc8SuSxdQ/e7
lyReQJDP4t6aUGOvn0CHkxl8XyFMTTxE/LSyJmTp8Ih/xFEVw67prl7DuQPZh43Hpd+e2/cecO62
Gd11oDFlmHpnF4oZK6y2mkwyvMf2mrbwThxR5rXBaPvh/QvTE/jbE++FfmLI6eZTzr0hRUZRoxoW
ex0Lr3mE+058sNKPvJBYURKbNFB/R3EeYP1Y8RiQU36cWmO8CX4N+IQjnNBuW2OG5K2qGRWrBjzW
EBHzakAURMdNYmMfNYp+TXdS6PUm9NBzT9wwg+DlsiozbLc3bnzLCgvMzmsxz5h10K+kRMuw/w4a
2Sv5Wkzl+zpWBnD0OLkcikvybjgMBHpdDtpDkbodWC60khmVJ9n0W9E93UPYJfMHgeFBOJ69qRpT
Hsj0G0Jio0eVlyDvDrPC5cXcohXBWZttNa06agFkPH5VNReOYfulZJeOApDCT5dpPtmdIRXyaeiS
FmJoY5pAMo+t0+Euu5vXVvaHkrNGjIwclAdyiI0XZ+dhw2aBPbuVR1Nw+zu/sn7S6fCRbWAU/uf2
mdxtnNgsifKDZ65GJqJeHet1sjO2AKL2/i5zSr5ROsEzdCgODsexwj3dPdgefP7zmh5JnMX6fjN9
lRsxgQVaSN3Q0SEZrnA6kdGgkTN1zXErF5fUdFfisIJi411PEa7YbkETZMqXg8uYYKbRRqcFey5z
00OazIXvtToTaZOlGyU6Xv/wTvwBncQR+T7YrsaipQBX/E/SRl2CL/RxPSbCxbnty/myd2lC6y9/
25UyaBkpr5ju6q9MwfPtyjHMyc/4v9hZM3ocWew4/3F6VQjHGphhY+FhsE9E5t24bstn5/HXcfQv
tPMsP+ckDMzA63Ka3r7OBlrNta41dygz06v4BEv2g43XMvg5R3o3i8aJgcUXmykOJxNV34l5Yf4p
62OuYmhT81FSXFs/tqp0PHFWCxBdYMcQ97upvBMjP0mqRn+q0/uP0DHqVcV1UBtv6dXoXmIRKsPC
y+xfjgUZOb8W8pqn7PHh1PWUehKjpr+cG0Ag9QZ6TueAZ23Hh1Tf5jS6WtAml6J9/KmrmOyHfFJb
o4fw/iyIOai36PV1lrYdnzUcO+DOr8oIjGCA5JU9sP2XTLvUGLxKjtdiP4r7DmuQRVLcF8/NGUvf
tJ4ovcoOOb90hThEoZjJtWUS/FOkCgeE15z+2crRadu3rVIMZRRuX5M/zRG5cVjYO5zJzy/DjEHV
ZgErbDlHXz8SQH3Cv7yd312ghCcwfBTYxklu6j0FoW5H/QYs1qKdze4bHQx9o3AgM6PdNQoHGpY0
PamAa0aVtGWuvGT/buEwG7Aa+IVSYjX5ojLNwLMRP1JIgeDXjP/+kRkHP4FO7CvKM48q1nKVe7b6
EkYR8jWQKERty093BEVGj/5LWrOC6gQ3ym06mRmPsItcJItqtJqGJlNmqruwI3SJkB71F6qLf40w
vYd1OpEr/j69ECd87HMe6oCppRpwT5j3aZJp/YzReCLo6bL5VQYmYbrLmX1r5K5sGM2JMcBH10wU
yFb5VtD2kILQbsyub7A7Ukt7xcV9K0t3hDJoUn2GtBMc3hM1p0qLA+mqOB/3UWPKsFe7N42iSdcX
X90pN5XshVpK+yLBulnXVP3bq0JNOZXiwmvk82JihHndT08zQqgeydhir/PXRQq/VuBHI//U2iRU
ujVc2VS5yAeGQ8OBQZbH1JLOQ0VIpjLLvYrRjtyu9ZDeCa9ulUi7Y8SVGx+ccaaIOPpHd5fnjnhS
uP1poGDS+OeAKOUFq9opbORXkzCxFwdcuZBmGmdeaii6HlxCMjSwftwpKN7SKy8+xLagT5RvLoyZ
1Gv8fsTTxmtme5hPs1mUFuHbXCRFxeYgh1X3cBrOnVyI6NFoffq/Ev6bMMofb26Dcpe3EzhDP2mM
ILIFu/ozzr8eAGXiGSgVIYjkaiSRVQl8CIcz/rlMerZNrNloy3RjfFE3vaYzf/canF98hitpAX2X
coOssIiFYEdDowz+MmhoG7VRlMK4wxoXmi4oqQH7z4oP7k1Xvw33CP+nlRR/QmVtsW01UcUUJf+Y
WO3SwHHciZ8Fki/JYIWc9B3XuN79ZIp7RdACdkoRNuUchDPN8JUUdCJzOOyxqfKrBDnNJBjNBPXU
m/CT3yTQw9KFwDM8JJowcUjY7vgnQCcNyRPxgEnTxjz0dR/t/xquHzHyUSUVhCcbfkHZMk4h6u8E
bgwM7ahPzvcXegUYbGw74iRRsQ3fCeybFBU7e9EiR5hZ+49WXZIBLaLnorFcZxB7lIoC0vNL9X4e
iwjKMRSSPTeO4nWguwDne1W8+AiySBv9b6TjkzKJT8ZzXuRxUd2pE9aaQt0EUwCk/DOED80VsE5y
UFp0A8WLViVO3qu1Wd2E+QyCmh6T5qBPYAu7Xu0o+rMKRaLxgWHcxXH75ym6pcpbV3oXGXkXcWBg
i1NDXdyFnLi6VQJXBWD+OjYqIjfXiUjVbFmTYp0uIvkVfjPSvwCYNGBsYVjGiCg705AhLj0vf6LR
bDGeLDmj6E4vCWCVk7Vvxd5UIMQH0B6BarwxjqkY4Yczv3IbJgX9nTCFdpkxn3pWssxVub0ci1Rp
QgApgGi3LCVcuyEBVB+BmIQntKPVs386HYGHVlqfgRmKgsfa78Nq1afid4HUTOJfFd1P09+Tolzi
0J+dwDnP13FG/oBCQb0gx0jNgO9YUxsQO55PCYtW5qbc2diZAsaqIhOS8iNbLC1RsDhh0H4ELpYu
XpAxxwu7Xow3IJH3EbitlECPK9Lsj8kPmTVsM+5TZmfirl4UrKCX+/zR6iNa1kzJg/ToV+VbBWCh
OTOg3VRMtZMCWldwsnJu4ImkOyqRTLDRJbH/6iPTRluWI4lipaRIaIxBoU1WF2wF0doIAEMvmhuw
rrDeWB7PeKlnbtmZFHWB0gyKtLOPMPh4KLUzQEor32XuK133VLedRfZBD62hGAk1hSGtOxz3pI6A
vM129HSLYfJJQWBvI0IJUhMEMhCRzPHXT7QBejRUPTW1TFcPBUgv0vavPbZcIAeW0JU11A8cA7Ek
f5abTZyiZ3TlrbaiYWBxbLdWang3bDPP2KTYckPkHvBGZbb04jZr88lz3edaOHFO3X02RGoSkfWL
sGZ8InKzU6TYirZK/oggNcEbJoYbUpJ9iCZtiztJxz/pttahBGm9dyFq7bCB02evEnedl4GSBW8+
6FFL4v5Y0kFr9h8IFINfTafInRMA5xrgiWMzJkpDLqKrwgoBo/RZk+CO4Nf33EsUO0bjDfkODvc7
23FlKNY73zITfp0tHrw+q0VbSxLyLTe46RHSL2hyvbqOUUp13Ny3mr5foF/byLJMPEpBgmKQk65e
oDI4iiiQ3fa1w6M01dIGOUeSVhnGmOUhYFE8k1qDFXDRUe8own6yFO4o4guIYnpmMJ1JB+s9o42e
BRAo7rIAJ2pFvBIHQdVxryjHlfnv14+Y7RtFRpIz+DsYEIRCvQLgvZHBKvcrA08ZAB41HrJ0jEgP
m5enSY8J3v/njH77zIM37jxGhE5J9exXYOTi9qeaX99dWHVsn4RBFzVvD73/eUZrrRQYhoLVK280
CyUrwc/JHUsE+yTObb7KTCr0SHkTIHrRGafvdskFaiPuzQathTKiSR4Yur5sHBXSaFSM7LWeSiqY
RJYn7V9iQFuE2rf+axxYLoHo2xl4ku/n/uyBVKy4I0D+z0iC3Dcu/YOcRQkkdlmV9Ox/KgFFRyTr
jHNC9wek9akfYn8dKT9aUaxfUmxWWQvif6z2phf/8U/xBGcYz9q5CwgEyoBnYzAtiDM8BmFL1EyR
2agZDWpmYd/SKfpdZVnFc4W763oYKLLIn52vEVyt/lt31c6/ZeDOoQL6ZxJ4iquItCv7d3K79/V+
ok4hpjItfMJhQrY137nE3cabsI/VEbJoUoQozzVIc5GanWoXKk3l1U6bolctdeHuPVFFmf0cJrxi
FGuwGKJz1xQlP7pAjmmqvUUu2Gc03TattYp29DbchPxmskb0ID6RUZvjeDqca5StM0YHmHPlb/qc
JZGyfyLo+alUndDBNuM8qjJNowiAW5PXwZO49A8PKuD6UH1gyASmdsLgYjYDlWgn7J+333n2oAMd
9EA/m+fWG/jZ4NeIgtliBzsptERnNXrztIC4gck2/klhgJ1x/0TbqRV2YSwiKG42SKy/iq3MqSub
nT0CSubUQsuuh2NOlqc8f3jVPTknCJ6UN5KsletZuqQ2yfCMN6u9GK96wnjqOvWMPphLj2WeWnRg
GIBkgTrYf6547VpxPM+XKYuO5Bb+O/CJ8x6pv7jRJE6lcwOxzYxPRNMWYG/kMd0r/hm3j8UzSQ7b
lkUQhOMLjoQ3tGE+pcUIWmx6mIqhdHmMOWNHO9iGk+6TqUR78b590ZnJ0IZ9z+vqwpD3PkoK7SeZ
zXOYoVJJioKlv904Fy+BNh85OgxRkAjnBOuEcxRT80598da5jIHVqT22xkeT57wuN3JLR1djYmFG
ESsPaTdqeuNNJBCdqyPdgvgifzk29GK1r/3p5TGFoz+paq1x4qnPvztFQvFXEbBm6u375Kgq/Eks
q+SUcDmZ3YhQ94r+y12fQcqYJAheYq4XmH4PBT3rznUr7TZeXrUQ730h/PaSxmU8lrDLjTLFmjoc
HPvhkADxIdJOBMNMLb2dxp1LhTnGCJt392qcXrdPtAQXsln1bhhb0opC5YmP0xjczIy+hOrxB9Ay
OLWY9FYurkAiui6Fx5ZD0okhSWoDZNq6Ucf803qlU8gBLENYiKBxZBLiBBsPLChDQfD1xJjlszLV
d8oZRFtnl9TjCAFH0tQfP5aJzrNBdQPS52v7h4w1wFWdJt4mk7dE8+0JYrfO5jvmQJYwh5TTyYLy
nmzCDx9PX5JUfZBne6w/ssaaWf0C7QRi9WFpDo5XV5cqJW04fcPEbkZle3+WSP7iDaZzi5Zm7E1G
UCxQ3ifir4QxOkA2dhCH0TrJDFANud5SInsD8uIUs+fzDT9RpsLgyyhrjxStntZZL/ddp9qyXe6v
hJsbTXi3YrdNnM6kr9o8tQGT7O7hEes6xkBIgOiZFSzsRfXH+FM3Uc5lWCKI79hOFao98JCacZ+l
t82CoGkpnxxZCP8YFR8GiJL6ah1wHceKCh4/qyvwaEQPFLNneNfic/c339MNphtNQeAneLiMaSHX
m5nagW/V/dv8kT6rRYclPCzbpLr6x0iTNKIXRmoAqxNUJOm3xfap31Jkfy1GVVHh0A3yGUAgETX4
zb35eqRViqpAXWE7vnas2o3Bt7onNn5OjkhDxp874pIyY0MLXS9cEVYJzOIFoYODtzSjE79SKuYH
4llgitHlQnyRcEVJ8DedHvUxIOZHg5hRJSYy3IaeWJWRlMOBzKXzQpPQxKpn6MFasdztWujTYuJo
9vBjcUFLIF8LFRO+XoG8f40/hF7mqAuyHx9CIqwucJkeuU2VLm7RjBf4Qd4/edvBbidF87ENZQyg
iGY99qSYCbwcJP+4Y3/NHIi8l2INUuTFFfmOW8gAQW04yQERzLHpFIVmXQpPZWkET4mZFjx91uN/
KidfIi3A3y5MkNbTObChip/DZ0kgq686jbWoyDtF5n9y0jo4W9NcwMq08CsTYEHW+WeC/Fg/bk9E
tTukqutmmLv01+6TUlTMAYRF1a03Y3hsAI9Ege8d2j/Zr4x5/eXiqYppPTeY5wGYnVgH8hPL7T+3
Pmjt3e1FqpqbHuh4DWBawlIbAjz4dNJ0x+iaj0SFNdwRybOwQz80aU1GR5Kiz6p42UMxPDuwdCq1
Ys+/HKP/wQCnsiE2IIj1B4SdGADvIde8IzVc+Lqc1KmJNkNrP8uBpK00Gt9WA/cgVlAJNGdHOeiv
4fK9XDoX0SPz+vVvKibnri8qfUdRn2Kx6gHIzfHzh2yF5YgKxAhwATFhUgpoLUi8xiYakas8PO02
E9vBDEADpWm2zBwNlqvC1iB3qdQkZ596Q01slW0PUqm4QlrRFzMMDYvyIubNAHq4cxLF6kW6akiQ
gZ/jxyqQiqBQgUDc0HUPa88HlbN64bij43sb1wxS9Z+hXm/gJhuUqdSMgeqSZLy8ZALwE3cJinfM
aGgNrK8TYeUGbApkQqEx6NVlsuTR26LIYsCvYQPVJsMZfQWR7rb5YYFWMY4s8aQ3OJuhVtMqPFwC
2L3txsvGywhJ29xZ9ImWQI7SR2bH7yx4yzUBntj/1TcACOmT8UGTXYvqsij7K5bwIoE7F/SMHOwJ
4E4yT2BEcigFENKHBXTdqnsRXpM3jEqkORHKIXHiW7g3T/IlmAUlzgUXpFtoKZY4/RizkC3/Mdgw
Hxn2QP6stxfXtf4LUJIAD/DSgFWK1MB2R6pXFRFdz0AgALo4ixjonx9WCOqjaFkp3WOcJbIgT0fb
0/jBu3LvcrUym+bTvUjW5ItuT+VgvqX0T45a70npcZ6f2UnnXeuLs8QoaMko+5FSQeRaYdxXaLdp
580Th/8t7u65z690NXKyt08l5J0gw49yY/D6FB6tmaaPvd445cKyKy+apoT5RTxxfCXxJvkTJPHy
aKPwOUPF07Hwslgpb2LFaQ0+W56w/fU8utltn4aU+DWqQf8lip4kOpbAoVXqgLzWwIRpbFyJMJws
KuotdPsIz6Vb+trglz39KGUw4l6YgkHfh8qOGSyfd7dX07v5Lm/qe8SRklP1N+WeL/Ci2yP0aGmY
RxMJPZmjGRcz7ZXkGm1ndNy/MMk4mz7H5CFj2CNWgT4g8x4YTP7yr05w6hMGbYpYIMGagnXNrFrx
RsJAkpqGItnYqmeiSqOh/OoDFPcTgMkjBtFSgSifVHtHtRJvi0u0wLt4p9KpdiOOnu9sApo3ATl+
ONN+nzTtGtsKZdEKr7uC8RfhQZLs3LEpQNSUNvPFUAuemI4fqlL6TFoflV8SNv7tUV+4i9nSOv7X
nvRBlRMmeN+oOVgWpZIWdrDF5rFUp9YJ0CXWNm1dEbUdhhIrLdvavk+fgCgXJA9LoYBq8SJ+QIEV
23Y917tDBbt/toED87tKMbctYCTCZwQE6nqVlLA+sX5WZmiPO/7VUsduMoo6mzOz2TXp/LGWfr9i
iCKJI64xsDpvBin2z7KZ4+j9/LROD82ILMSMQAsqlhO9mtUJeCS0JW8UoSJ/ena/TZNFsJFvhLu9
cVIzrT0GBil/AnremJEgOKpwjKbEgxQqLkFR5rjK17PGfun571Jlmt7RaCNLU7EKA8eBfeAR+ONY
u43iCWUXaWJIiVnpOCYoiBEiEBqXdME7I65IdZfvFYKIJCCzbGjOzEI9wHo2Fv/th6u2KzPAL4Nf
8bYMqmFVxNBep0Of0torSzcXlQpteAg3EYpAgqxaOKaPHryzd/kJ83RLb7/2K6pmOFDMWyDaPFyR
Z3H9Swgo55CxS+54Rxc8jGuWzPS46lICVpON6UWIjxX1LMkbaTIhdPoF0bgxfNQp6s3sbN2TpeHp
FoWn1ZhbS5SQlW0IfGpBKKIPuWMbKV2/S5gVNTNh+0BhEVirKYIeX4MK1FG1yghMiJ03zvCsNAZX
4S1Lq6HAoxZOoKpJ/6c8NI2RZ1faNKtj8tuKiI7KUTMdksgYsxxV/ul2x2Yme/ji4tE0KNzl1oFW
bIBXUGfpiVUtDQEBq3pogjFIr8hCUxLQhmd0xXIXMr0aSCa/8tewcedOBpYwECSWJPaboNABqDiV
wR9TlKH2Tv9TksDuNCDBJqT/sBj/IoRuKElGe72z6mllX7H+2u+oVVmTZbj+6d5M8rHV2wilockF
UgtCruUbEX3plX3wzSras/z/hDzETQqqJwn2dD/P2VA6sbCEHvkaWmYQti1OBpBhGmFN8EvM8mNL
hXWds9ibAeY0X3ysTi1r/Q3FsZI3BcAtDDBuqK5f4nY9aviiFyFlultKMSBHuSrUstT8oabrrZ0t
qvjaeF87I/AJTZ0l1r3GAdwgXFDi2HOk6erHULU2RPuk346rIylqJ+XIcdkzEnLpVX7/ZCirzzss
PMAQn696uPpY4YjzNE0gBXnDppSHRagL0oGKx+UnPDbWBEpIJch3SmFX1ugoV5z26wEXyDnnygo9
fan6ZqdhpEsb9Lq6XQkZiTnasWxDctMdIhB96IZYvfPJL82olC0/oV+Ft+QaEqo/az6JI7Rvl60g
r0kX6IRWt4TNC1m7Cxe4cFDhLT3nqOkZESxkwj8J/TEUAD7oPnsGrRG9WCovDweL6CbuYkJg1Hfi
Nz574vZw/VwIxAGGH2wDAyTr/z3s010FrNwnaTCUlQh7VfOi8zs9l9/qQl2zWXYs3RyirpZr845h
z/wHUGO6rGLwTiU+8JDKKIa4eZD76++mSMaXW0ehyp7baWJUCJO52Y0yO87+tSEw6zsqeLbVBIoG
XdSOodzeYTM7AhwBhGe/cPgc4T4qS5tE/isxIJTZhLR39sDrkY2bjm9TY38Y6IaCzpnS67RiW+eg
/9Y1evoJ6MP6pO5xSr7ZZBeDqfWI5KmzPechmvMekArVW/h+JIDNqjnrTF00hLEq2QRw3AYFFe5K
5oa4tFE+t163Ilayx2viq91mDu639e38XDPY9Msm1NDH/arzUuUr+IPG9JyvSwt2wpywR8o5Sgur
s/m59MdkncT0tgEMRSaLig9x3xnsYH1ftGtrgaIs6g2Jpgmk5hD5RhpUFLzwL7get5ozZu6vbftG
aT7MkGOkrn+6OHTm6b9di4EnN6N5qSGUso8loF7o/YkLDgMnulHSnJyLegg+1MBaxS7bG1rsYJl6
dEQKBC+NcDhHQO7PiOjxRdTKrgj5cVLoga8O15hUayPI0NQEeJBfp7Its+By4G9TPHNCWBMdnNzJ
TpCVKxoeKqLSNtVMHW8HL2iBZumfWT2OrYBsfeI75yueAwIar81EQn8q5ZZAzodPxhnKWxeciipp
x6X7MFubk0j8G0ImGQbSyUAIOAcK2KgIzBdwSzMOushVuLRS8kb3hA4DtygMlyMYmky569eB8EN2
V7qm+PIQ09QSqio91XvoLVIZIySh+H/TLDTpUqMl5x1lBO729VTdoKz3ZfDx+RX9YMw0pvUJcELo
21RQfAtqf/FHofihdAjllCkY/gkpl/7vYmSZAIxSDKKTjkurVUtRv84BW+hVHqTBorZJwcDQiVKW
quezRmFhKwPWrqtQ8GoJ6HidV2F08zJbk2CC6nW6WgzlUbkxU6ANDkDVteJ9H0+cZES1PM3K1evq
Nx4jphBD3eNOtrQ9tfTEYPGjS1EIPPap+ZW1i5K82LyYxPCv1ESFOzfWuRzzTFFnyIwVExo83HLf
SHeSQuC9ajWmGHX2osFqGGk5dYXuf0xYgopFFJGAdiweEmcvyWLBRB0wfWXtG2Ry+4X/b+0HNXNG
bnhUf9FYJ+Pk/IyfFCBlKSPMe6sxxgo1Y7xiSBuiA2vMV9cLY0DoyRd7lDBh+dBEwsBh/hlgj8+H
SPJKOv7emS6KSkseomv3saeEuX+ts2BwCHC5LLK969rWbxua7xWAH1HbMQBRTgrheK5UnFYvbBNc
RACE0uSO9P0Bi+r4HhWX7S+pOY+3vq7MYPzTsFkTplnTElAArQxGMvD9MogCDC/YaSLyCLlZ8VHt
o5RbXhCBNbrZSdFmmifs/WrKQrIeKoxHDXaWSfcCCkQvhzl0WTtum5aalbDu212rFpsuAsGMdIMK
U8V71DmPrE8YnQZg+p993o/LxOQep10Bf4V0e5eR5ICNlmiBoJfLlF8olmytzQkCDSPUbnjpfbN8
YbblJL8IiT4eJxuUjQEvHDNq14qzCdtG47aGvmsdk1+iKyXpDY/M9dyRBN5+KZrR79wpiX8gsq7K
WagGnROf0o7MAidSNxZYY3XyOC5K+wlyTsx+26NcCHqWjjl88AE+qXWD8IAo/T7lT7XfIMQcNAex
kBseyqWcyQHtfVBcjuBDeq+usRqopLamV9x7h6T8iDTkdxw209Fp+ZyTj4aUiDKQxKzTpQ8JV7aD
10d3uZlVY4HRzW/bTPy8pZMHcTzli5YhMiPq4ARGDsiyrrdrrcReWBoa8s92Ydl5dJfNsi9mGYkA
hZR2vQNvzGxkv2LsC8cLF20qYoWFxRUafNGgIYDfYwgt3CuBsqSZ02RUb2YkTC+M0VZBgxM86K1a
6BBfGBomjchoz2BCJm6uZTItjPvVcYOD3dcKWnuxlxZDGj3UBNY6XWnF7Km6CgScmp+c5OGcHKzS
BXeRszLG6iQPPKplVrlzXwuZ26D4oBrb1OLyk5POpQhjgOmVoGk/hddCFc4K1Fd/kelZ7pbReZww
xvHdU7L8amiuY+wOqhfjqKFMggPAG6QAv+op9Xa1LNrBOkbjousrxmtam3Ez/onnY3MIW/N0Hxpy
TlPQUAkiDQQwMeasmjMvprnfU1lIUxhPSH82uFL2CaTIDmv+5dJZdPRz0W+aZiMcV4cExNvWjC9E
v+jcIEApsfRrUxCgUTyaoIzSNPaBlk26DTWdLYLa2VsoGHt438cq/I1zzbWS8FQhkU3DJ7dYwz3r
CTzl+bgwcQoAH97z1IDiugtIxR/4e1o1egtiCkBKX+8Wtp22RpkJT3XSYFWwVQtH1lm8E4YuepF1
ZY81elX9DZJv+aCwBj0JTbpab7c8FD0bk4sff9hFiPeE7MbXHU6xYl6rteAdvdYtrrqtbQs80N1y
xfhXx+asyMxeXSNz0dLYeVRdEKO7eqwIsdd5Owc5cfqyuDd0wSZvGXDAhXyw/JckuBmz3C8A6SKI
xSncUA6DFpREwEuxE6C9PekFpaBiR5B2+vUNMFMIcuUzNN6UsT9EmIoyAkVnkBJ1rmqJHQ5VKLma
inyyJ1Dj03cLJp/MQgIms9LUV4Ke612HLkFk/u8oySJsUIZ6p+AW4wsTTi6cTp9HDK4MsWS3XTnM
Srpyr+ButIA+2x5saIDzgzSOG4k0AKFnbbgsOdXv0/BcgKdjYWIjyZCBQCXi5+LIhioB2cGX9z0x
2clzahtEMQ+wf4mVRKICj/bjekIlR1vYnN/Xu535QiX1fWsFnqBOU2+csfmqyU9xcQZxD7rR94hb
YcV7YRdCnBYzY7Zjx+wEqnihoAXRxgi/kNVg5iyuWmoinnueoeCxAqUAkoC5KuE3YRSnKD2PT43X
haJq044R8i4tTsRGsZZaY2xcfomib75BSXSmsycvjCiTxMv+vMgGm20yKY/HtpZQC0tVEMi8cbpk
1D2f6T3FA2k3QYSlbhKZkOXeIFZNr+UU7CkbxkSM3z11nVaHe8+vtpFUKQuk8XqLvZOHAbywN6ne
wmEVIo3p11flbpRoDTRg8TSKWd2bH8O4r5+RiCnYZSCDLYmAZpw17lkmfcL2ORI0g+iTN5FxS2Y1
pALoZD2WtHGa9YtmuDgYjDfp54Rqa4D+ThUSjOpZ0NgcE8WMFNM+0x1Vwvra+AmSWq+vrmH7s0zF
GgSUq0FBA4T6Z5gjvBVL7JRxIfGU9bu5/KIWHNeKeFHUSFZUVNtLuZGVclnwtLLh+H8WgqTUFQjD
hW9sf2DzawY3/zLsGT+yHBT380O1Wmwpn/awwzb+WRKe2CRIgzwMYpCXOMJV0EPcU1RlHk5dRQi5
sMlVuMSJPIngvamHeMAJGiQoKDUXZwj/yPLC4BfQiwXnysZhEJiXXjY3nca/zc0cYTqS8gFWbbSh
VOYpf6C7kvfXBoAAM3n5XhrL+EFUjDUIr09x3oIFECdzvqN7wQrXbFnVW8tVlqcu14KYJgq0H0Du
9icW+im44siI6xLLgQbsnUvU29XESMVzp6i/TlbKv9F0L/L1aD3agudPMCam6hYb0mhYipz+owek
Fv4mpPu3eC+S1HBcYjsjStT/YrQUa49BL9Uju/6wbHXFCaM94ON21HADlOC2L87ejGQLX+0Y9qT8
UKUoTrFjHllsh3/hod/ykjtyADm1kmpvtpkgWhNsA4dGdCPYPzDKD+Zsn2rPNOr70eaqLECHqGUH
rVRYwIOtJicZW3HDRDFTaAlm86j62orWpJgQZ5xO4qFHt+HyddEcBkecHCj5pjqFdzHq645S/Daz
rdpxggvauT0LNQdFLlf+0jgOwoIl91piU0rm8QboN2BQS/P/qbS1Hl6+8m4oNtQwFSALGc5bXCn9
OzoPDKn3NoFBL9sAO46+PQnZFyN04UlsDpxHpZxUAp/sc5ktUm68pGC4SoRQ9Sua8PvEVLgAvzEk
qCuF8VWEZInXdmVkJJYKc41TlBIgfTvJB7ki00XcwkurRb00miDo77kKe3qUM14VomXkgt0DwZqg
78/v/G16+JCicAj/C7lrmQUZHFlFOa0GsUMVZNwQ5DaFGwUQffHLjqYTEWpb8HIgvI7Y4/IGqNNo
1AfECMB9CPEct9s4prZZ2Nh9cBHi7ZVQTudRSroTySgGXeWamY5/nSCxckglEDnNWu+PD9iCPp1y
1GBd0QAd3M4+fAntxQXO3mB5iRv9SZk+PCS6siJwWDzLkjlZ5AooQBH4hrqkgTBiSPnvQuHE8LXd
zyfKP29U/ZbF+HY1iO5gc3DPSp24HEfnni+ryjEeNe5jBbKNs1ooCf5FUbwZyoe74O9BZ02A/KRD
I75/QLg2g8OudmlDzSPjLhggmMV7WoVfRruhlfY20EOkeBCWrWTpc8OSVWhl54cSAe96MZE6OSWC
0teOjyuJi3YH3M6osY1neoXbx9kS9Lt7+x0kGSinvjPR/HbnTHeCD8qIniEloT7BnsIXu538qkPq
M8hEpkLNZb0DAhC1aL0SWRjixP0+VocW/8NDCiYtdtWKhyf/ces+/JgW3zIPxa3zUROqWoWM9JZL
HJ68JeqhhORpvup+kc8qdSP+AB7Pq0ApPpXxgUjOzmef9Fb07bHqhiUhRHKKCuQaKgzamlPqY8LP
/m25RM///PY1zbMyBna+dYD6elWCluUKdOI0joQjYSS2y91zmrD9hpo5qR4ztGO1MzmHn1jhP5MR
FIkYtr4//bj8UFJzKC7KrLah2L2ZbpzzS6xlwnhRiHXYXqu768jbt8ihnosYWJ/qtdE9bLPpBJUg
aBDLfmdehC1/gDhpl49S6sW3vn5e3/QAADGtYNu7zps+QTGfyUy1qfyu9j+SshNByzvdfv5g0wYy
fGBCioxhEkJLnshVoC6Be1i74yli69cuHI/HWm+zmAirR3hnIMV9ogfkoKvKE6BfZhJEIK+WtHmu
tufEQEP87/vSwYwc8+TXHyVadVube66acQBUY0rXjhkTUEK1dA9lEaX5iysqBk6tdLJ445/zcVOU
+uSXp996ITJ1+MJflTb+IIl1VJFAYnOgHXKCXqq3X9yhxKUkdt2B5OEw8PKg0RTWmRS6RrDwXqYl
ssH3lqrKMwG9VxWBgPL3mF28X5h7/iQMKDSKGxkeKb+U8OxUX9J0BEAZ2ku1rZNdjsI7O3w5/2WE
eiHTniqdDmSlJTnqsZO7nuPJtnBw7xYTYj+h+XWkfRss3kBF2dVG70rmm4eQy+g1TJpwXTLmMYm3
KFYW657ec2wFx2fGxPPtannKrztCs/ZGMqpzZgWtQOkHpJg58MIOSux87YqL0EQsVJRipXx+ujp8
at13FFwV9sGIsMvXINZxpW/3QScwy1pvZlWL/GYF3sJGxt9ty/aej0Tvjl1TMjndF3dkWXVjUM+Y
J4L//ADN1Ut5xmrkeKYVDscKs3tG36ECZNCRrWk5WrByTQxqqPdJdlqZkF8kR6ngyAsKCWZZDqL0
D8zkxEOwRAbulZfRsJrxGvM3qXCmIFf/pkidAdb6DCjZ0z07r7oiBlbvoatSNVoZhGTz4bB4nHQz
JTojGYHm2QGgYUnJILfKqshpUcaMgP2KvNvpTrXMX65FgVMwHM29ORo2x5TKyYuvRvVL1nR7iSWq
Phu9smXr3VqARsZNeQHJHVqal3OHhYBs5WFADK21NMwNt3c/C8G0XKx04A/XcTn95gCKuScGmWfU
HQ3vXb4jlauvQOVcR+qiTAjw3kfv+lz+Td12RRQkx7mztTFbXO3/VIjdRaaRNDoOfQuC1ZahXByx
RHQTKbIyHWCQdo1ZGKpCp8+cppdm2KFxTUZxZV1x1IKrmCt7SebfsgNlnye18HApxKgvSl2U95PG
Y58ocSzTzu88SsRLsRodLQVSAr/b203FzIsYTZSlM0wwIjmQv3t5ljP4tFog2oYOh7s4XUsEN4sn
ao2BWw4wZ9Qosm5u8c+pPGo5/l0qKR7O+4RxZtXdryqhWSfJbCazALdn6QPWekP1gaEjL9EQo2Sr
+6CTpwl3KOjq5sg3iik1CVylQADsuzucOsvsI4yo4UjajNL4xTqLxTx7YUtXtHCcOYAaBcOm5O9u
lNr0YOqiMd3SsB5CTS7QRpk6iCXQyLvtmdjq5SrrOHK6kTs+fpDQLNiF1omSj7Q8egqbPy1ZXJqX
TZXBRqWiKQeTrPgdZgB9Rn3GXdVolVLeS4swrmAuTEobjAINHyaWQx3qjIOm05kItGdJie7wtYVG
4q9fUb6KUMxCRIsjZWa7hKBjAcmJ0UrJV5K105DeIXOTCjzJcc4rAUJJ+hfQ0T/8Qd2gmlCWiluh
Ddk2H3wfQmWUTfLQ3RkfcSmtRB40E8xhYJBTpqxGDl85YmHZ879PMWwbRWy0VwUIl1aQjgkTJMdA
1ep5aX6xCJWPWsQwZdwLAD04HCCmSqTSbJitKk+EqrV7B9aHnnAi4viHzmqrfrAPMiNYUP4uNPDA
jHeC6KIyZHdWgCW4rE25O8Lc95z3u+EQVwIDRdIulrrgHgbbJjMlP8yE+36hnxOIbJud2Wcgmyu7
XDtSfTor7plhGU0lx2dXCTN6+llHct9UYSmjo0lWlSnJkabKWfl+Jx4tmCPVuSUrndEpZZComjBW
BTDOrNFpMkDxbeEYSXtJoUhPiQyWZhvf3vx1kWTbDy617s6s2cMhNp/29YjhosmxxOsKaR7I/coR
vsrzmSjKRKsG4N/A0NWRW76xQ5bX5p5dH2EpWNg/hZYkoUCSqYtaf8WlF6M6oTbMimNhUAdmszoX
iSQnjaqFxR9yX1Z5bR1qnJ4aefm6eG8RkzWnltDJ9zoZyE0D8HJDHXbYWlK1HBZSb40ufbPzqMOw
NyAvwpa9iapllnQ4wPMFm7Df4vDv0AYufzu1ejVVPaqWv4SNVgD40OfeMu3kat9TF+9wuyUbPDTL
gsv/mKcGXzJqN50KGd9XsO1KAh4vaugeRQMl3k3VktahQwg/EhnYAFx9eMSI7Ul5HMl/KMf2Hta2
PE7tYL8xScmQSLG1uqbCe+nKWINwJjPnCIh9MgQgT/fiSsq8KKIdojEpMNy8AgHrWR3gjpUXk9LV
mi1kb0CUPOQfDN8vH7Hs2CbQsIGeNJpqzyz3gvblsBFBSEkXktByHVVn/lAj6NMlKocbJEtIkFGS
Gn99ca3OwJ7GfIW0su0lGxvp1H8fqJTBJzbKX3K5xo3qHdZfJFJL3Ya+TBAxw0f0T9JLxXxECByS
v07sdqkYYXX9ehTJ2njW2WkGVMJhG8FY5APyaigjGBVHubKvQxsO1q+ZwHvz6t4If0zuZDzNn9Kw
JP1tbAtfnwIBBuNsHB3af3BUnwn8oHSNpQIS0VA+nOPwmIgNWvU5wgphjZGzzzU2EJPOEv1Psbio
AvqjcqOP/LRlUNhlA3ywk+uHQa9SfBcEmpJzgIQwJ/pbTC0EG/keQ6GS6BEFwdphv5NZkjmsnzxQ
rlS9Wctxb0d2Wz0dKEsICdKbBAK8uu/yt+QXh5IPQ+2+/XgbpgO6VlZNdEi7eA1xnCsPelJVb/ff
rmBRIL63GK4ip09ti8I/tdgRcGk/P+al9NWM20hVG3bYWcnzTyl2ki2IOm0DTewB+4f2uEvkPpmQ
Pn3bGyjnrOthOWUHNjWfMmSn04BZNUqrFGzQkA4kQ9YAYNgh2sa/pxrOv/qGM4qh1wKH3R24bhpL
5U/d7eorYfxdy6j0emx0EP2caY7zOFIr2TIqf9KyQXxNh4basz+LKxBzrLSj+2tc3zMYrdOygiYi
udhjDHAtF9iRCJS2xad1T3QiXEocydp85lwzodIXYX+BA+lRXD0eiqXy0sqL3EPgMndQx0r6rtfF
YDRwb3Dl45PiBsW3umMY7632COsz2UpsHb76XQSexzBpSvOydmrswGStowEeIJoufVY/hy6MpHZk
nvhIIKcew0od6xJtB2NPmYUULdXPpci6YIXCbjxpLs4Ty15WYAgAP4Zcdsd+M0Ea7kcWAoER5agB
3Vz1/10+s/X35eTiHCnsHYTmqYksrf0Wo0H1zue4TtzhB8iTfP3QIrCfsdQuIoUygSgb1FQBLxgy
OLxnR+542S1orhxM5hOEm7XRNUMspzNTnV4/hBN9ZUPC/UWiSYhxis/tFZNpJCs6fRXZKQRrbHKa
iCGU2oFosZ20XlELMNc9SnW3YmDhGDn7BseoDsZb/Wl1DssyOiwKXRs45tIsEK9XmnnpDl/AQA0J
GavwZnpfVWe1JZ9QMpLPqHRpEPrY3XL2YkMokzfC3r1oBG6SSdWaNVgcs4KhHH3+rssViOJ5HCCj
l8hIK505eJVapMpykhO7yNwqdxkvrPyEGdC/vx6bPkfrbEFytctrfzlGnvF+Vx0qTcHrA8IozIvX
R9vTiUYZ9CHbumxjNJ5SGfJ7RsR/BCnRPDSswSW0vFFJt90DPZ72Yl9MsVp+T5rC7o8tI42/olHz
dllQ6A6xJNCKdYZX9BqMz09O6Ajzl4zhTYyZDyZ5dBeDTHKl2HeCPA5Od59V4oooOTlYZZyV+ylx
/0PwLxobZoKq4+XY9XULskglEz1f1Ao1S+t/BOjSTg7WfFZVZn6UZ3UJVEeq69eenL3DNOmARvXC
E9cEDS1ce6rqLkqM/UWWZ6/idnevRJFpPBbwPJufchKAi01aElz/Q1IO2U4wmByuNOMFEMBPpuT3
/WkZ4VFXf3S3Z5LGZ5Ag2skrNjuOmoyb+aO1duQ2/L/eeWZLVPyQqzb+87DpLvNmxP5zsAKGNDpY
S3B+4yyGs25Mwrtu8XQigJINqe8OzMokUFs1MQxuWRhHtPxWvUqEh8sY/AcVKjCKvuf/0HjOQA1O
9RKuySRX65NpTZZryCobKuhRiYnyrsbeC1VbpWcT01frNIz591sz7YyI8TeT50FWqW0HnBzQru8V
3jitjpqs223V+S3DK9IVogoNkZi9n+nZppCTwNFYUDnFME4WZsYdXC8VAnvDZEVGEonr+5DGbisr
bYKRT2KU+M9jFgyycQd40pee3aCb8hZZ88E6faNtK9IMGzAyK6VEZI93E/OVC2h8dyGe6J8yF/52
VvzYNo1fO9nLKgJwq4/VYpNoXg7S9qxh0nBs+mjDjxCTQi72y4oa1hEd7S5ofyHc+07W8lnRQdyG
N8WXmmG/rFcFSceWk6Fcjx0ShTZDuVQrhWiCtUD5pOhGCXVAK2pZEwLybKxuvsswWR3ce/vg7MMF
7v4CU4g0SZK6u3d1oclVGTF22qiGOTN4i4ngCMBwkTfA1b9TI0UXL5LZynCPE992yoCODm6D4mP6
O6bM+bOuRkeRmlBqQk/+ydazvqZCPDfZcZ6LqnhXDlCkCn7s4bqcX5A7lvq9FzSaSk0de7T7GX+C
cRy3BYnN7L+hflwQUv0VP/mnIf+cDw8cqAgA9E7S12cbk1SK2pg2+WNyXGIFw6casDWj6ZZH8WZu
LjAFQfLozSIfMNyn5K+WrjAuGNf6JBWPVzoX4EAIJFjqJjlA5TBJdqpvUCCrtGAO3vubqZMucxud
b16TL3/X+X7R6ssL7ioiRcli/S87fsQxbbIFqIgFBz1OB9b2c7LK5/GbMIYnE8VeAd8PhqMco+Q2
1OwBduvdvIDdNf5X49i0NAxCOQwqCSvx8mWrRSF7dzQmThKB7n1SpYIzZ2N8ZoFTK99m3iK2UN4A
Phl21pNLLYaZTnu2ph+7c6BsNo0vhlJ6xMnDO+cBGpqKMTTmd9piA6NQvfO4HyRbQVr73KBDS28f
Ke8QJZhvRiJBtcKeZTK4j9olLQkqHieWIoZnij1LJaEqFDYwy++SYlj87deqMadR4pTWUbQr7LlH
7PzXEfNa4iBA6aZlJqegONyITo72krhDEPUw1VAG6t2H97PGaMNU1CXexEw5IBahtJSaKll1Ae+6
u40Qn4b4RrBm8OnlB6CDPtWf4SqvNlJ0e9KNJUoS1FMvstiSH33REKKEt+nMgN1lpoubLjR5mI05
DlKEu5vq7X86USPsCpa3mpdxjxlY0/BqEuyBAVgRXLUQOep30HrLEQbKVRi6GAIBG9ZLWsbNz6GB
WGFBLc+nWGA/QzZ4bKq/U+Dzxa0+knReA36PS/xV93Yk3brSGumO1nb58psRQdIxbCZuIVRf0poD
y1BPU5ZM3gTFMcmf7hiLOmu0HBom1vCYrJ7G8t6DzMGIzz8K4BEe9cd76ThMS3UrIugk8Jn80Uk8
8WlzLP2QKxSyAVb84sOpKV6Z/KEEcrwI1wND8tlQhDxtQ0dn/FTitClhdlBfyS2+/M7FP80ou0Um
c0chhOkuC/Ud7lYRMcJ2k1sBkNaegceC9vzEA67AVOnfuLF6JAcB61qvAcquGgp8SY1F28xASNs+
vsfXcu1Bq6xevB5wCwbG2XVfD4fKYigaO2n09+pSuehEeNo+nnu7v6i93xVIYIXFZ9rroOWTuCEI
X7smSuU7Q4t3O469D9tFo1FY09tzDwc4VhY0RvUDu5mVsCh7tOB6fPnsQmImKphlFB5AkgOVCn/N
NmSeEnLs+ymLLTkflsnTVTJgo8RSbTvn+ostEqYOfRFlUacIafSs8aWalXU6RJByOMSTw0ykKyK/
WEMZWwo2gMKqmRMfSI711dv+VUurjcG0qRTn92OnW4pXn3j6Gg220VC5f2iVMGkv8Anp8AEI24S4
gFj0GjixvyebkqirzLKWzQ2e/x1X0lMIJtk0Forf0qILNedHWXSxqCf0divqviurjikhXgUBrbmE
ifdvw+6wfqAGx5FR4VmrGR4Xm9G3xfwVviq+t8uQmEhr2lgprnldlfDRuIgYzhLzPqLnccGZuO6w
nC6RApHTguqqzXy9PaDHhZ7yvcuSe+ENkFqZkEu5Vsg+xQ/y20X8XjhBH6/ZnVFYsKyeIddg2Oam
U+kRYsXvqXukaQ0v1kCvV7a8lwD6cEg9NMoFPuw+9Mfaa3UZIJQdHL/zrB1O8k4cxZR1pn+cYK2H
9sFm4Q7a1lDhsxNSJ3+CSU10cJXMC+dVU7zkboLZntq3GqZvtjo96WNP/+NO/Ur2hxSh7YtARd8L
hy3Dg3w8oybkz2JZwsGXMLrFfMdqWG+6g4wmVomuTNWrvaD0WZhydDxa8pJEHc98EnJ0pXVBfuly
ONlk9M/TkWfxjNvKCrklpXgO18IVRTFR8F3nzLJ0aHgdsS3R5XFyl0++Iq5llhiaDKuuQlnGGL3E
fEanKiJ7jD7gGGDDP65ww/qXa2zgqy8FnoLxyLzTCQ3+FdmkiI+s1eoeoGVndEipWliSEUADRS3c
iofaKs/c7afLG/yqccQylyeFwoLtEOiJV9ab/gvZYE578L7yee2AU6mMHSHzyt2V03jNpEK765bc
FkK7o/nr7g3IypXwdAeYrP5pY7M4UHManL5LjiwrfwEVY0C6PdOCGqWwKyYrrOpXvbWNR05C178b
5X5+bD2ww1+zdnil1+rFMT8H8YG+u9MAb9KkP6DB9lAlD6WOIm7FccLW8zNIISzaAZbnaldGvk3R
XiDvlrLxG7qQA+qRNPDqoT8DlOdTRif2G3+p65+w422y6N9VtVvgHTqGYiP/n+g3msSaIGRTsXSE
iSdgijqvvpAhZCpAxF4v3GpxSf/UIqHfIh/elmq74EY0QqP4XvWKde8M4oSGzp60Yf/5le8I9Op7
ITaXUgZLU9kbZmvD1mHLtKw7I4ioPhr5SCyCSnfLqHJuNtPtIRMGPuMb2IV3UBGmiy1fofw9ZTd8
iCGecesjAcZGErkkrxqVr68EBANLHaVmsXHDwv25XZ4Xi63736Zm/EJSE6C/aBy2jIqjFEM9KCsR
KMn5r1G/JVOrkrjCU8SGt+658o2WULxswnuJtpeaC2Pj8qi31iTTqE6Qf1KREfw2q6zhQwHO+ggC
o9l8vvQl53K8Q8Df7gaWt4gmY0G1Ji1tsxPRsNbyI9EleEAOPv3ORo6eex5pDW755ltEXHfa/fc9
LuqoJpJeYNQWaVV47gYWag8GexG8sBmgL5hI5AgO7MN4wMAz5wM28I0koh4PoUMUGjsSIjxAzJHH
A36IHIHLv9Rx1XZGyAkXoWpKJznQWIE9fPXN8Ubmc4VVAwnCkqLysAsyt7Xb3806H1hUtMRId2v0
nlis0EEWAf/QIMYYJT5+/yCdsom0QzXfaRMrBhDJBwEtb1n3ZMCdcyq5dO/MoEGzi4Eh0kc8Z3nL
LS2uQhHea6GUxiXUXuY/UfHhX4DG7VrUvTuUy4itp1ieLbJfbpJYl4eLhWgj9CS+myKCu1DOktrJ
wH28M5rx3J9oU/V9NqL24ayiYjrd25vbhBfDc8DETyfkUKOseGGdXddk+68DKE7mJEkL5v5Vu9fL
/Gkr9HL90qQsdOIQp7hAj3BJc9hFqYqCrhDOy24SDH30clS+KMRP+j6Mx0V8R23at7PX904OPef4
cDWbtiQqc8eVr7gtGN50tWAKB7bqXevWEaNpXAVTDo6yvknN2PEfBdmHfnBY4I5LQqpQg1aTaHQg
SJxus5qGd6Qg+5lxgywu7iccvwDFfyBJRTjTpHZ7VQzCZn84t4UZHmVEJ366y6Q+IP5QCtwfcmwd
J7XHiWBV5MG5ghrzMK/OuOY799gRXUP6MuCx18Tf0HXBObgMkkNUCuaozRo+x3N7ZRovsCAFuYsF
aVUFqRrroDG7AtqHI4hhqEBGTU8vNmSbAqBsvPc+U+DC2roSvupX1/JdBLnb7Lr9AZBwH6ToctOD
twZLr+JGYzRROo5iImXTSr+6M8wSEQqV35WKkyP8Tt30M+p7TiCSXXslK9Fjh88To1E5HA2SxNCk
80KJc95obnKHnVwWhxKZfqg8ibr6H0lkobK0l+W6TRPbjMDfOHllq1n54pSG/iqYBqA7BLngi6OY
RsIOHtQi9u9y+3jeTX0nJs9NyYC7G2gyQiUd5fH6K47IBPi+2ATyswtzXe5CcZAW9MTYHY4jrlH+
MIuMyRzMC5lQ/4c5gbH2d8V4i/x1ULBrXle+rXJVnaZdAyLzRJTiIli/poDVRx4CJ6MI8cWtMunh
5QaCl45wKtsaj++OpXI8DxBImqy1JOvwpyqGAz9p5jt5M/iZTGfP0teg6Jm1GNK2zLtKWGGexjDr
HrXSx8d6SV6es+9h5e2ijguWw063oLVCE75QUvT0bGWpjMbH+M8jUOJPAxsdqszsz3srUPaG4NlI
lg8K6xKZrwhjSpMTn25+kpKVgwyQVo5Aptg6lSfBJsZLDvAwh9sDe57H2dMu8Fue0KWNV9auCSeg
L83HZFf3tnjVbQ==
`protect end_protected

