

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
GWT/RJdN/UcIKTAhVxs3scTnM63xEPkso8NeqXOmx+sudHjUMJ/qSt5GFjdXAqexLlRND8lEfssX
Q8fYY8TuyA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
J+phMqmkYiPgvjvEjlpcdWdxzP+34SmYIPyc3dLXEqt+h9EhMcqfQg7r/svpEBV24DU6CyKyCXke
3gZaY85pXANGRT/lW2K8drptf9l9vYajWMSy/HjvETFYNanQN5XDicKd40/UNr4NV+8K3+zJSD2+
6HJJVC0iWa6RgWieT3M=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZrkwjC6jJHChQhf/EDIYzNRopX0ckXH4NL9s7GZmKhZ5Xuu3xV3LqvLjlAq2T+/3AXtko4HEVfJk
jD8rEKHAwLnqMbikHpL2pup+LY4/a45y7duxNC07dpJvYX19IW6mqYLKEJTs330XVwBLE1KOyaGV
xhWwwqThGo1V39JpBwMcpzmL4YnxHaTlERiq7vaoQpYAMkwdoBVpG9MMAn3CbeZJI8pLk/zNkztm
rMeS9pshqNVtzdUse3pl3EDxWMB2hg/4/G9fk9okekAXBV0rv5NMqf0xPrBsTvRJGO21aW42nO++
dC8am+sI7nAhoG4w6z/WxE1BGkRuZGX4CGhIDg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iexpjlh7M7dlTcv5seskQPlqyHreGwsr94b5YKwilWQsfXW7U1V2aK3O1/+pXS09S+pTH0rKoHNi
ofASVdK1RB4/i9AYD0Ihai7zYaqt6eRX7azypmOnO0M/ZZIrM+63BHWcDodlNlh86PWfwaKQSqJW
hLVuOmY14GXZev020lRZWg+2UhI/Cl3c8nww44erkAvCrpxmrhaZg0s2YPKI/KBqZbZHwn0ufJSY
5EPF28uCCS1urKeejeaSBUmimEDyf29zU/xFd0fvevSdWXaFhwjT2mOL7DranIxEzj0yQrN0jiKy
Towa0uazE4xB+gMrElDuwpcw6ZUMyEBsaW08mA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DVPBxTgKjw13z3lZMl+QMKXV/uHfXNCgMoWbgQb15TKXtTCmkLiaCYkk+UNjnupib1FZuwkbZs4q
pFuDW3Z3x3poQoD+4+Z7IIYAmkcV2VNFgSXWGO5qpHWhRfkulPfZcRStTLiN9EUcwXJUsLi1Rwk0
oFaVSUr3p4Mr6zjC18beDCFomH1w+aZiTDmIDtnqdWVtxtresAhXiT6k51hdPESOpe/yPCGrgQj7
cckAkNk0Y7ums+FtMhs5xsfKLV6GQGr8vql+qoCmnMNbYofWKIq3pY2FrW6f7ZGbFhW+vgaVatOo
wR1vGhSucCD4x9efRbKZpd3HOhDW/vOAo1pd2Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uIb1xi/b1sGS9N5+ge4ctTMaXcuHePw5wBb1FVa9aecf3hzk8F8+/rWvK4DX9IjVKEx0PLXI6xjb
IH/rGtJXdtbDJdBaXxCtQZnZ3bb8a74BAJHYm3BEextG398AX1ZCOiiun/unyz5EkREGrSg9f1qp
tvP1wCaUgYbP8iAi+ak=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qK9lK7oKxV9h/658uwPcMAAwYeLmnKNpsdduH0hJUA8HIiT0JfF3YHf9Z/+4sugCSI1ARr9LlbO/
o+J2NPNqOXlyDgJW0FGjeX+G4wdX5LlxdfSIcRGs2vzyXQiAWVbMq15jqJGV+qheK6QIsLI/qwOR
naZ46kfkwSE8kQXhF7WZE2kD7kLSTF5QPnmYFPP1wrSHpjD9hfcjmg2768Oxg74FqPuAHl6cX4Bj
Enf4+hzQMQ+IcGssYzesFwyeHIqJFbufwMH9hDnmz2bOveVtLUI33QRmIvvIjsEuvmQwCu/AC3gG
UyfxcM7HSiPQe9MbxhcS0KjoubQbTx7z04URRQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504864)
`protect data_block
1quR0ylthX2gq8ZT3cIO5WOB15nRsHoIhESqHYx0YXLQm/5AON2a5KFfOuch+OKdNqc0Yq3guUXf
lNWIMRWVk68e/+6X3xKDKUE43hinOK7glReCAkZmiGEacl1ALUCxwZsE4PK9alVSAUP0zeh9qj3p
/+nH/40EoBF1K3PRyY/uvbhYbyiciJeT2KdHK8RewRki6mfPJvsVaG0kSP1I9Mk2ZNJvrfjIEoZv
Mtkv/xEk4HAkLQl95jUENKBMqlMSQpGK3nqJLpIRkQeaRvrCrKvOvBAh/fMd3Fnz6y+s5uSQVO86
ICYAfOrANY/nonb8pBAS1ZzPYjR3BKHK2XKyW0HdPzBwhIPZ0QPHpRDAiPck0rykHT+QT1Ie0Vd4
h8HxRCXWYJC8EhQB9SHbJL11gEYnqiimLPHXpMYnPyfGfwQpBBKmEVSX4vrA5QmGnlfQ4M+B0/oY
1YKuzU80URsSdF1vZA+cnDv1ZeJ5ZZPpjMFbrkg2GoHM1HgB3WJ4ynL+lhCk5gqouSYSo9+CgQvX
PBtKpxYjivOXC29CYxr58cBBDUb/5wzWb1EpujI2Y35t+lNfBKWCCNpF8Pd0D3L8Flz749JYpoLl
Cpoxdt+luK5KxdWW/NZdS1y4yHWp17e7kCNi+EZ3entaNhpw1KwDzzSYoN8Ut1KOPRelP2E03aOG
oaLaGL8OkAYmfc7rTdGB9gOjOeWLu3RTgPwbO0ZQ2onl54xGipCU+qHWLOpoaxzV5+xl6dcHy8V0
n7neo/iyKKiOur7R5Gz63/mbjmGwaAGHz39qq+jfv64G8SZ+B3J6UGgYYTimEJ/FcMIarpLknamu
p7O00F2n8ozXJs7Cb9fO9AyuzkFXzKVUVwqm9loVCJqaq07NNBlkSzBwqyBHl801YZEA+qMDWAkL
o5PCzho5rpjRXyxkC+dfFZqm6P9aK4Y8oRlB1rDJ3L0NWVCCWbQKa/I2adeLOR9MSkdgA2eCAhJL
5V7PsBuGYGr0KxdXweKKH2EKymd8FZmlw4eDdCz9TjKZM17dQY0CqRm0532kBgFo5AEfhyUglWAw
Mogi8YW9lHXb7bzqLIyf4ubba87muXKwywH/Dopdkcr/7jyB1+vv9SxyE3C5dBO5368oqrVo40WD
7eCuZQ95u98SYm1RveBE8bjCla+OcyuDTTzIYteTF4JJhrB0lEGXq5TRWSo7Ji7kkbWRFSnITxRO
WUSb7AU2knncE6Ybzj0H23FOLOh5dLNqgX+Kap5t/JuX1voFjW6TVJuRSYpZ6wQqMQf8hqAbU03V
iRdTFy8rqd3sbaeO+NZS76taTPq8HNKQoDtvRCvoVa4+Q7uESpUHvS7h7N1noRzCl7z4K2h/VEeC
3ySQHYyiqq7x70PLa5dgbv2ZKqhsfIrckarpnnJvIISupjnXc66c68fTlBC+j1s2+7uv49yK6ZDS
EYRJAaP50uYBcNjJEcbKLkbAvfYCk1+95tA537ziuBXY0lF2qaPNLHwErvDM8ehNywQm8qBSW14C
Sh72FD829d7TEsJ9h0EQLos/YvD14RFOQctavDccTaArfdrrqhB3v02+kuqZx463D9B0eqSEvlnY
P7dkNCUDO078pS355hF3j/ZpjDA8iQhVjN1zoNHXAkSUD9ZF1ZBOU6y96Fn0OPdheWkLmpJmz8ZJ
6YjM/xKZVVQO+DCvJOd9xEwTON+r3g1dGGxqIOY2uz0s5tYZBYqn7URfkxGyFY5qW5fZ9iSRevBW
NykQG4SS0yRSPdl7Ogc6VF8v1QoAHuwSKNUMhf7z4LIoBWOedGI+SpTi2sfFLP3YBe1Sj8QmWpyF
QzHiQv4/YcrCwVlrgE1t0w6li9HAbrQLRl/rKTz79UQ7wcwrgQW6UCBfzlUd2wVkpvJoUR8zQPOr
s+vyu5UXS6f3clUjrYeAawD5JgHpb87R1e2vFGRDuLmVmBHuJMCG9K9+MKFpHcWvjHU48WHkZzZc
oKe36awI7iifaj8ZS2HCBUb2LDQlletSy7nbtEnmZGxlCCEotBWO8VDWHSqo1p+A6FAa/o5mb8Qm
0yCyUsPxRDaA7FvWEs1FXGvTXLgbZBZNYZe4oWkFm8eAbc5MS5noprn9iXIBF6dCu1vQerzDdI5r
msEtY1HV9txwoPuxHx6MHk7ZeyZoliXDx9okpV2VLBpzJoflTTNffejgGHTKcbwn/tUmMgwEKqYC
A6DRK6SR1BfzdcdwLpu2COm2DmVtTdtVSSUxXvIAHbT/fmjGb9Cm3aV2GJYldp4nzZJOc2fNu3aC
wmap2FfKKxFclZNFjcg4VKnJG/APT7OYKEJ08FI3+KPJ5CKat0CtGcAkVzQ8CvZcDz9xvpAHpZu1
GLsaOwPZdy671uzlEZrea9T9ESZVFlPOIyVbCL5k7h9ewVxBviJqQ0AP041/pRdDBwiFrQDolj4C
vfPKgojQZyBqeIIuBzpDoYMyBsGXXHkSJe6H/ZHbUMDRXe2leyu0eCGINCbApk2mfRubf8Iq4fX0
mm6XecYA/JIk2YyWOl57cqKZpAdXJgf5hDA7lpvmArXaB/+N+YNq+Jkptip8AMr9OkSI6E6eb8qL
G6Yvv3q7BNKV1E2YrEWJdIlP8oBoSgb7TAUhccvi69UL+9wXnGuCLEs1QVchZNJqwpVY2GmCP7pp
YUi6tPbchTSnhNR5MN/SpA0q6cV5y5aCh9y9xMPdNIyOxfFMKMQ8i4ZnC1aRZd4lJ8pJjEuZiazl
0f4LdZ8Tp0EnTdGM5sHDYCX1PW/P8Uk6gZkAoSp4xZ76F0wAhNodrNGUVxIx4qEOJpO0sjU6lHQM
h++NEDFQ5HSjk1v2+I+CiSZ/e5v0MTzhGQhGgoJAZYQpc4mkMsbdI7z68GLkAvp+7nB999ny0LQr
64E8OIzcorUNnEJp5n4JnSKq9Dlr0nHk7rp8msNXoOJ6AWTGjb3hDetIgrLrC4+m+i6rAiXl0iDU
JwIOBLjTijNi9HWX8BD1n23RkTzLdSgDNqOQuAESWpE4Pho4cfMy76EWYjmDFzZfXAO/VuU9yE4g
pXGjf5kAUX8B+8ZlTftaRz9iby4dOfrnLjW+5IRTR/f/5CgfGE382V7TtKp1ocE8+aeDoxJDfA8B
hLWR+RMpeQSGTYshdVZbXxpO7XE9wdXqZN+f7EK+IWSpmTGUcG4NFhJQ21wmPh2PpFSO9w2hZFia
s9yafbZVDG0vngfRa7VCko7MRxxb/z5jSszcqNtu5cakVM57KH34yNu2DtTYE76NUX4wwLwCQ3OZ
IQy5IO4wo/9xiF3soXTRrU19iaihv/jDxM9KVjXgFZFcPz9osL8KeZm6f8eP7BGbaX97qi7BVQ9/
f/6BCL3V6/jwMQKIA/bCpd+bX0BrvqnPWmTNc6UewQTBqIFZD5ejlt1MlRmbaSzY93wSUBH3fGOm
hO0k+9btKzV0cf913rBIIDUjzgztXdBoJ4dFhpYyqD56DJsxeF4BL3UlBgEr/rQEmAuPT+m5GYdN
1N5aCtEYOiZphCiLc+ICosUHx/Q5mz+5Z8yASSvlGvtMcPmEgbUrc4Nb2CYeyGxDfsdAwmm867di
vTZGxNlCdphSn0ddjseyejzoyz+eep288JrwWh8Mf7980v38s6ExxWY6H6MhwiDgN2ispavROINE
s7YXpJ6NOn6UutaCO9Iv8Z4Foi5vKN9fo0t1UM660N5lLaNyXovovMzzb65gdmznvSSpoVIpMycA
RuLW8KD+IBc7ZbQzAnFyDE4wtOrvwlsIokknsrkaKpPBKmP+4TU9rHt/X6eGR+Lo72ZsNHKFBBgo
sT03IPdIR5EX6b+ojwrNwXEWMu8xaiY5cQc9zNVVPurLb2fOHztpCBAMeaBSLMTzskm36unkuy2h
tbqPBhg9xE1p78AZ5kolxu3v9pUAGi4uWsxsJ6kbLYccNtG0Ovmo2kon0azyrUhgn2bOGHvzuGfq
M0xKo4Qbv2Cop1iFCmIMfb4x9DpWacvUpELoYEds6/DNPAyrhAxv6BWGdGWzINkL+RlGkbDkF/Cm
/SAvcT7nlN/njnMiMfdV+aAysE0/STrP/92Ap7/BieL4dYlnDLkdPvbEk76fceYYClgOS79gYIzB
CCO6Y4oTNYtOu20NIW1Ri0Sbqs77P/irJd8u9j6YGsaihkC9j8W9Bpbst+DwBrz7N4cxCXgztqc3
7tm/uSCUUNsbySk0eNbon4u8bDY0pDdGFWiOI1MR22fyIL6swuMoZFzW6Nf5Q9PgWn2tzob6l6ka
huOzpvKMX+WEmOYlaOifKCoXTeztnUPh7iObW9eTlH4NIIT7NWJBNHputAqrAtHNZplPsjMfrK4O
zyAleS4Cq9YCXGFAf8DeneJjtM4LYy47ioYCCdJI4C2gQ04/gJmdTrj4yjNLHZ8KgR0pD6PvqtLy
8nHuYx+Ce2+b4P+l4Nhw3/93+y8I0buH+K0YJnJB6GbKM6v407nJvTx1BeFx1hNmReW7eFmtnlS3
9ZBC2pmnVrVVVRueOJf6WxpQCbaw/APncyz1qp+DxeJtZWN2SrV1kRgQ1uYUP/deWT/BcRiP+zdN
erKZQJGQrW9O4foIgdo3wOIjvIdw21HK83La/oQvlCuPFFPx79BhQGGnN/xMVqAUtUd8MILOPtN8
m0f6R7U3WemZMt2pTHuAG7MkY6jTElnM4G/8wG7GzFcquIOi5Es15Oko5DUEKCdBQ96G40meRkex
JSl6OSPz/hbS5P/JUl8Kv6i+RK0y1Y8DxX0fIuBLRylNaUj/ASU0UH2E/Pl06EZJgecO/0Vaem2f
qTcPSTnRl3pyHCXfD+Bsr/VofXct00jCSyf7IY2jyyvnf4ixNrJXaAdgk7Psngk9LZcKzSL7u2P4
gdOFF/VR0KOaFtRcxVlIilC/0J0oj6/JrsAbKfSTJQHL0I1yDeNon3nyNv5zWCp8ier8JjXCtFa7
KqE3iCYx7DbOQPGIJyKaYcYfDXtUMpIE8I6dlApxgxNahOGHJbNzc/re5QZoXCsfoBx+BOT/5NW4
zVrTaDOSbphMt34eNr46J/q5eCZ713LYJGLodsmKln4Y/1f4FA5VE9GJ9aE0DA33eE0EMGPA12Wh
LnYZuFng/kpN8CIC7g7lpkvBPkY4YcUJJoMm28M/egrWeNK9QIrWkzKhWKcu5ZS+1EIT+8JBZ8nl
L+Fp3OPnN3eVmlS9ABpzWhpGbAjlOzhZUYIDJA9jqI1i72OwJHIWYVUpVVNSsMWFW5KNzZgtC3qf
7Z0LQJHHwA/esmmnNzIND2I9mB6unlwMbSBSXbPF8m2YDA3BwKBf/twbdrwWij6PdGHxz9TfcLSO
r4V25ZC+Xr3+x1+IIEX0qNNSqX1TdeYIHQjephzgIblv/iKHo+xY+CWJH/o6n7mk4dpMCu/9L0ZY
Y1NkdpqnJlJcl5syzdHUkfMdVPBfdej2aqtY9QYck8mt+G2rI5clwsEt2DLcCor5MVY5bLBm1Qxa
JqQem0Hz+hI/+DqsVQMqxuFjQgj1HQNQwttSIX3Lbuv/FOFkr2PgfHLT1U7lAJk+/s9fUNxo7uvR
enLzipLtX4QazKhWNqbTAc1EsSWcnxUtDkWTUquF8m7yL5ts8LwM0r9XP7VC8szdZHaN1WykZOSx
RYxd8PJiFi5jf9aNXmrs3XdU6jrZNUmEo5Byx4a2jflBY8kBAsLyPVphVJiMsnc3Tjv+S8wa+zD/
ZBrpRkGOn6PZNmnixCmOeTeVlBFl3i+GnQWN/gLe/OPW3M80fdu+AN2BmCLbae7SyuO6MtaH9FEJ
vnf9hx7NTynBZgTtEEQv5MMVxpu+KhwdIyhL/ZvZlauRqpf/1N3wT4fK3eaEiARNYSErIR+49M7x
+HDnfH3JIM7NWxfgBpRlhkN6zi+J0CYLwmGJ7+GvHJvjuBGYspnufi69+cme5QKjTQkw1IEbj0hr
hd9G9b+E+h7HZzxDPOIzoCuH+hA2G6VYuSMoHn2XsPaiPmI3YDkiYWGKPevNR8Sgc6opAVmK9qzH
YX+VqZHfQ7KR9fN3HHXPxv+nLOnfj+j2H591e2pK+aBl0vUy2iB+P3EiKCS9y+zoMV9mRDTbxXS1
DypYaLXN3GT2NAfZy8XvRgN+GJ+0ZQAvZeFCKxkq7ary4aPeOxLAvga4CT0avkNed9hVIhaKr68m
1Tot+0UBph3QVI2xbvM/CHTc6wJsSez0nJ01IXnVyHdz+OZzMFZpTi4O0xWKBWkrDX3+dKeR6yCd
kaPftAfOHgZPkoJmlZo4zihl3wpwlozKVy7c2X9z1ss5fVAONAXDOB+wrsBtjmod8H4cqNOH4QSZ
ShJg+/kgQMIhVIzq8rA9L/zOwE9BXI1YHzyUYgUtnKj3lRMCddM5uQKnt/e/ptzjW3YiIye4/36T
MyGU+6xw3lT8GX2rW9fR9wA80BFFiFdzk2QuDg7UyDkk1cUhpFsZpCNmQ8FBTrPmvOq2B1D1X7O0
Fpe23pddM9NcI0jwhDruDPVDLVtUPCQal6AaJxZ7fRJcK8uxL0fUh4mKrD2rdgwiHnv4tvYxSYyH
I/D1+pMWaM1N0y66vJevWbzX2QP4o/x7dcvpNMf5x9b53BYI3iFfhKaKOdtjP8KVeA/tZNhPB9JX
62eThkpXwuQZ1z6tAU+zg1cCoDVcpMOR/2vA8qEaY3ztLLba/MzN2Lf/3tR0MXigBOGmquoD0JMR
A/XoPjQI5BNMWkdyyL3LwRaOESkAhadZS3OhS+AQWe1LmvCWscin96AG20UglU4c68LDD78cARWO
2cyfe3xJW59a8FXiW1SZMSi2cWYc37LuGcY5vz2LSV0BIN2w+HZPc40/whEIVF7fHWKcYKYG6BPM
W3QOsrEQ2N5jBoQA/o6fdfmIWMZwO6qJcetxOjHtNEDixZa3DvpBjfGj6I7cyV9w9X7K+xzNzoqk
j4NQJIBiFGrbT3Ui9xUhN73DtO4y0zs4OfCsuChmcHmNQ4wW/rvLfRLp+T7+c61IPpjYgZbkKxOE
PTARV9NJTWKGtBL5NSv7KGhP1atz8T50nEmq7jj15yg2O/ysiYWwrHin3C4vfCtkAWFs6XfIZPjX
9MAGsVqKSiQTEWrjc+ZbCBlEnGxb+HP4dluhSQ26wfhVu5ZVy5iNagIzEzgCxbdK69JqENWu7Ka8
d2N4fXk19SSaKSvizXju0Q+cwd9crdfHtNvBTxRXBEG+ZRNKlfvTjvtDnTYvkHvYHL0Ry+GwDpHo
dSdjYxAfN34uEaCLVGrap9jViQUX85GsBOvLuj59T3FTAjl7f/ppysRB+IpMFtp0zXPDUzuh2UUK
Nx/kMGvyV3oww8C7c7cwAzjHBnb6cBWr+FIDEMQb2C9VCxrWWoLE0eBARud/DTrkU97j3bm9D2eX
zRCk8bbPBuzHEaUjOUQ0v8YWRkbLN7xHhhGptmAnOuj7GP63k2PBKPdPJ188bzp/ewl1ynCuI3Il
TuMvA/UCr1XK1acNs0gq1nd8FifQSx3VQGd09nmNGdhN8uFHQtV8Ko5uIECWVkJBxjh7B6QzpWmt
aYMevnGHPNUAPkko42Ma0uSg5Lgg5GDdbRPr7OqNifFkE0QQNP08qAxWoTkhQQDYI2tdgfpJlOZq
+OJ1xzR+zTvHNUg3d1y2mVFe1VhHbgjuO5dgS8bZralIvDcgDoJ11jDwoKKo8vdmgfnUCkgFbR/K
4XjdHGYv8fACkp1AQf0R/k6wobgjyYj7FdVCSM5Fk8f2qd3uUuVcrQtAV0AGmVagzYkPfThK3pjt
7TSpHVZsxOws/0eok0aagfYZ2gidedU9fefiqplByMz6NH3RalImyuxiqpxVI79lFvS42Qka97Wf
5ya7ONw+dWFMzbPQSheBGZN0P4ZUFR1HQ22pUEvk1eFQy5P4cZmk6XdSvWHg0liIySAks7mqF5kP
neIJefgdxeldoEKNE1UiB/I7uP6HSuMztrE0g4YjYPjqGGjIpT22wNbBf/Uqx1WLN/JGUu5QeeYM
TSXRwzJ+NDj26nfkZazBzSyCWtKB/qkWwLlRiLnYyvEf4bVJvBCNn7RhaM5oEo6brvLIQCABvhwB
/LgQjUmHBYZzRx6nQE1braWW7UCWo314PbfInnK4oei3FmVYxOInBgoErUhpjFDurFsY1ZafS/9T
fauVhejKnRdsAMCGYp6plCC/hKgK6SO+lCosOfxv/7xirwgB4O1FKN0YUdkeLr17nGzVnh2D74zl
lIIP0msqZO1uPJwyqx4Y76Gzaw4KJKyhnjjp1bXBkGCuekhUioG1hzLiekvdOpmUWwJvINetGwH5
BxxYx4yvQuUVwKm+xwDiAKUY+6zkA2s7hJj+YyWGs1gXw0eoRSrRn9DTYLUngxDnCWZtIb0ynbq0
75OwaxmiP4P3to5Zn9D0ME9lM2IXvbbW4wx3xxFd/E6u0AAGBs1cI6Y2k/X7fLmTCm0vhvPIRoup
2nguVce/YTJXm4xNupazhO0uMP7UsCEbRMjUnAxBAOzK23ol3f640qBwlxOe4kR+JnJ5BSSZVvvl
ZboarWrTJf8UnK7MFG+PHf3ZzOwfNitvRAVydpxmf86uE94zfoxr6kaHeyJDAK6iIK5qb5va8rX+
1pCDO10GKV/HeqpGtwclayskwAweckOECtqzb/KVFnLBDb9u3VjtPpKXpHaVpDSCvyv0ZgYswcLy
i+fr1fTuAu7EYYZKO0f4x2wC+Gp+QhKevjG3fXkiQEJe6hSMTLeT1mFlR0ZVJO5zxLnPR/xcDN4i
scmWqKMnWn5qY7umwb6k3njI9KzEXuFfTF+ACndUFwveRabsIf8x+h0pm9nUEulW2mcP3bfj6m9y
32h/65Cmf9BMbR3KewGnAPawHDGsi+tDj+yEcmKS/UrunYZ0th7w0e7ujbD0hkEFDq+qfSk9WAym
is5tkG8PJBayNfGU4RT2qqUHMpoEZjScOzyQ6AZ3Zsz+UV1ORhtGM/k3y5N27gOGhTrEDllWZ7cV
wanRrWS9rWgvA1QUMvAnFd9XsEzJKLG3YIy/uz6dCXWtIkVwy7C0cy1CzASOJWJI9XUezwYNkWHr
DdS6oSIfMOoiGMrMAsreVho+68BQNIg+tAjSta5YEamdOtmbrf/NWJubN1CRedpePJKjJhhUhbn6
WGg0ZcQTTgSYv99xSTeBRBhVcwTM678yrfOFP8Lc6CW+xdMBURlpL7DaBdu+G5Dj94tOXkVGyM1W
oTmuO2VWiO6tkK9Jx0PxnMnsdNSkqbNG8WuMM8y3u1/A5QO998atfyvBDTKsvCyakTvRd67L1Ubc
kBeIT4PGJnZjvB26BSInn43DMF3RMRwLJHyCH7FuMtgvxafS3sFR5aOfFykUAw/mtr9dxdDrtL5w
NmPMoXJ1z/BqONqIlG4vocZQu/a8/iOX0XIQJhUDt98CyUlHrSs54MmQu1dDrkBW5Aym4AbVwo2W
C0RbrhTt3JvMRveIaTv2STVHbIMMv1iSeBJSXlQIYTeEjLUVVH1UvNjLbkluNPddhWJtfdVxTd3n
G/px5E22kjFGAH5TUhiLvDRbDZVZk+NgQAbAkhCW3iYRpnlDj4aT6DB2eCKqdYPJxP9DtZ6cvxK/
rIIyEy47uw+F2P7mYHZRbe1KKaPZDTlFg2i4kwtXYqr6m4PA3TK8my2jEUJBXiNGeUbgTBu91l1C
bT2u8RSFdh1beSk7mxtNy+NL3K3l5etPKmOuDlwDvsKfydGOJr2Uocz9OPWmBlI5QLnKQrE/KT6N
E4c3pg2+b5nhahkV8JiCEaydCvKgcJjGKLyE1PCCZkqId0uRJziG3H6Ab75R5Jd90a8alMlBaenh
kBNNY7Fokmjiy+DAte3oakth+SHXH/OwKyWcFDPnLAdmgeGmUobwq27Jbi4cabbiHm2jyvT1u7Tp
tV7GpnBSal7GLsRrhRA4rlVR7dQ6//InFWPlMfFMZhcll6BbHD0kBsDuYo7eus7OC1k9E9nITSyx
SNhshB7k2Oss0SQ33M7C6QeWmaboZx0Sy9h/clGe0BrTPUZEldUw3z0fAp26rGRpIb9ewR9dGdkY
zCz12wg4gGP1TWjL2wI9ugxrgzfRkVd3zCOOTSLg7rvPDG6/qLdkRQXrSp5RhAiVybF6oXCQiz6K
1d0jyWA+nsU7SKthCbf70NkHUCi5lUaP4J+Yo8VekETX+O2n5z2lZEKZ2n+7QTD9QPXueW3PM/Nd
1N+UhKGgH/pZbRp0nOEfTbyyUvdQctBrpLTXXWEFhja/jI9Y0X5hOaNSQmaSJM9WJPnxOsHD+O4y
U6MzHwa1YpIOs7uvSqQ0KdSIjFM1+kT5JCy10qBWfN00YTV973qiuBt9xdBNNL8z/rZxcuaACZ5s
kozrzyp+mB772S5R5HM6OX7Bls2mgq5hbg80TcLUrP1zX0wPvM4j+HNDOEmAJvcJTMgbJLe5LX6j
yEQ2wmk94o82K7Y8QRN8G5kSbS6VBfr6QbETLqe9aqS18tPjuxtDtsbRrtg/tq1ntVpssE5zxl2/
5/dJHJmYf5grXQYo+26Enre7cWTFN199cbqrSQduDtM8R3+pMEf86DFndGCuwFIlocnZRoOAmpBF
VrDr/T8eZokT6vGiIn30pIZb4+9coxZH5kZAVp/NjoVp1X3PwIYVEArLzgfhpjmBxVFCDDis3cGp
jq8196fRiEz9LLfOOM0MK1UgaEGXHdCOs8aWOaoviQ1EperRoHscJ2vzXGKEe7N4YdL90lswmBNV
ykd7R/LZo1Ps1qqejj+vYC1izh/5+Lxh1sasdVGvVcBUGXVQ28ogXbXPJ1HGy04rh116aEDIRDlN
ExpnCAD8Ar3QscYdKf9uie8OtKQALZuZvmPE5bp3uC78Q8uCrPjbkG4uhtU5IiQZsUyBV4S7uFEC
YSyu9ZjEXcnuwlcXYRXnoT/C6ZHtvWku3SlN25coL5RzCmRyczAhC761o883lbUqm7cFJ1zyuS8c
28lMgBi44McmfFdupKt+662n70346f522jCVrzW4m3Bi/3e8t1cBCh8nOHuTnp45dyUPhDJ8newS
PsltosBgTitK2yChN/LVAtKS7ho1/V0/XM+TkGF9dUnQzX6dBfCFD1Qy2X683Za9mguRWulOLJqZ
g+KoY9t9VV+vTuH7kq2PXZNHbzcrv/C3mj2L23pE3e7Yp99Fz8JLez/Tux7JvhFrx3DLJ7LV/YHU
3b8fo7NeNOUMHmnBdPnrSx4Sg6eikpQSWSLKea9dizg4dxJBmHT7Aj4Q9Uq4jJYNxaCLnNLbqB7d
CELf+M1p9XZTS2WiSOacKlcUq2mY5EeqePSRCsF/VsATg4n5T6KPzYv07F2FeHLJ7Ob+HGPxdbix
Nm9ib48NDaXEyUsa5WUfu39tncZY1au8eBOaugtUTT6FTCQf4TQLmrB6qRksE6fX9C3MT68xqAp1
u+3y+mohY6i3Gz0WkOoXAq3z8zrFGXrUHzzFJb2dNrrwbCUUKkZaYPIIgELa2pWfDxjDL7FO7b+G
Tm54WOp9AqV92VfkEIBQ/1YYku/KgN1qz6Boakb/6BgRxtSTCWldIBg/ogkq9nOhJ+yWc5767Kss
Gj4pGfIG09fLccyYrsxWYUuGGp0aVwQPv6G/ZYtN6PzwC+74tcxUSMC296hNGcuXOLrbqQttGdZd
B5rE8aOkdmVCWkW2tWF/L2c4bn+pX4dDKNmcdZBrA8ZhSCL+Th7MZ9WLeNFpjENtev5WJtj6NGVt
Zfy2jnEeWXeXPrtre6ClquLI5ewqCSCyuQ+kxU40rli6TvQHeNCDnf1uTKJZ8CDmvznV+4N4ipKC
KVrUdNyG6VlBfPfzvZV4mXJUswWAENX/HZ4edH/u+19NaXoo0P/gvQyosmqSRz6nWkI7oT6DrVjf
EfAhFdq5inFlPFKZE8t8PRwAomRK9WtGVbb4rzeXBrqtehsSQ20eIA4eRJYIxxk+mkQ4YoFmKoG4
DCNH/vwXPf3DklgaMR5Lb11t0FvWN1yE5/t50UlI5p8LCvcP4W+yKcqyUjU8gW/0n4yHswO5PtUJ
OyrcQU35NMojf11Bp1nN9OVGrEV08UAeP/ps0ehp8QQ4pSmdKw0ZXh+wTxJCnCJiX/XyEqBouwIu
l0FWL/WtXx/o2cIOTvW8Jy5gcsTKLChSdM3cWMbRhyR8ZbZ5cwUApIgdHNPb4hqQSDOLmYMfw8lJ
869T0XVIWLI33qXb/uVMrdUxEyANpXiaCjCUOr8H8SKYU7oz3vCsCsKmpp+CahzO45s8pg7Ymnnj
JNRpDExDwGbcRB0+wTVB5dwYxxfSlXQiBnoOZaYH1z36GnS7/phPEPXnGzhUmDlVJPAvbrRSo25X
CJr8P4D5kJITq+fgXgINmAbJvEDSFYHkLHrBvF4QVI9c41ViDpiHl5BzxuabsHz0yIXHimB+05cb
AADUjWNpu/EMX/mdQrFGEFMij2ZsAzPS6al1TPAJns3ZsBpMI4rdWbq73aeFNoZtcwB9UR1SNf4q
tkCipzIOnZP9QLi4J9Gv2AR0WHuAwTT2tVJ/IyvaaowrIFKTxF1m16ap7KMI7UOv69iKo71/LMoj
v3FD+/XewBiA9DIdAXnDClKpe7W/i0/WOcrguaiuIX1MqnqtUBgY/RfYPRONrLHICf3DGjBtgdjY
RlN3DpiqAhc6FSC/+ncawVfMvmGEdcK1IW4+l3V2CxHDQPaat4Vh70iWRTt4mUBUAhzWuEu2x2ER
TAukFEUscI2b672Et9rM/iOk1nXOer8XEs+ObB2KUfFPXnYpBj8yHeJBPRNi4sE/F3QqgTmNOF1J
VuoWNwzVn4umFn0tVGoPAMmO/MSjLIt9i7u/qDZtSKvQuenzKxrNb7W0uJjOsJzVszslB6Q6+N4b
dWUMyb2ZipsudvCi9rSLSOWyQB+2LSCGEr/7EBF/HfzOFyPZsyGzKlb3eOm/qxdH/Cxi93HtX1pp
hdVUXB3CszNZ/4oFIYSlRKlRhWDLjTcrkzyORqpV/CtId4+l08cjC6bk9yq3m1bFD/exRRUZjcrs
yCuoGSNBA9HHsVgMmChyvBhCxsB45/4VaF4DgGs6vVglwQOluS+947h6y6LFyCl3QYEknnHBlowG
8qithdQ9R3SEFPeVMUJKm2tHVP2bpN81w56KOKWkxfNO+Tm77ez1Q3sPemXMZz7xh/tg8/+Z4+5M
alcTo6WM3/4KHNpklIFSa2yAPEC3D1wnN3lV8h9QIyCEsbJHu5u7Bejn5judW/SDOEanRBS2cEAe
oT5L++/5CraHkda7ujwzJyZN48buDa4I1l+DVdIviNjbHeNOM8l2y14n17E7BZz0Kc57q4kjKvRd
4eX/5lqZbceo10x2T3+THcxy06e0PVGqJhH/xURtZD+ta9MNWyV7mPkl0hfrFs3zF+5LBAx8TANZ
z4sXQxyqjBzL/BJra0Nw520w0xhsU2L1aDLUHR5Cm78J6D3DTJ7FpOhu4cl0G99bCZG7DG1AGt18
O06d0DU0XqO4ZOgWcub/ES/feByhrYU1lCYrhnofOXENAOx9JdlPiyGIszFJ20yMW6tHnKnr/nBg
jpw1uh8MtzxCdpWjszD9WGsdObvkRitv13hOVkzi827JfFUzgXC4Farf13P5Zb/jdW2SUQRb51iW
GuYcHmyY/itgCzdy5xnh69Nm2GC2in1rxzQHt3XtSBgyI/2jA09cJzm7cTHcyKOZI9yFzy33d4VG
FPtcLPAgLE4gT5xwkYfThP5DYprXXVsbpxvzrbwow4LaT+HOEj0AW66bMqKqMNzcwnBYAfsPA1/A
BTkC1EabSh5hONr9V15gXEADOA+S2t8Dha2Kj2ZcWTqzAhQhDW92cybgkG3Ui8TzsmMN88ArsJGa
p/sWl4tK9F77eiTiVk5gGIjIz9ucShz6i6EInkVXqH3oy5e5+xxFE+DTwB05HMmmfWQQiQ+e5xI4
n9cQtPGlnz6c/bzCVB9vutsBU8PRJpaLICARSyG8gq7IGwE+ZY5AhORyGBm98jwQV8ESTInI7Er8
VburBhXCMYAhsfeElzeHFHt0RO2KYsQpT7H+qnEemz2hDAiwnQAsJW6YxE1vD+3gJczUkB8wUMkU
qFWcuSrRlPGcSH+wJbE5JpTb+Flfoc8W8glKEZoUyppHWTGhS/soe4fMswGZsFmoJSeKgY6z8zmz
ga+/JL1pS9PNCMa5TTmvSCZsYe+pINzvg2aLszF5+cwHB1gLZH9dvUs2Gtyd6K4wcESOsBDmDFkY
Txg8xFtIk0SiM8Vx/ddvgtBY6Q1Lr6yEqleoZWDdy3qCwOIionvMM+usZPYoFZPNI77gzX/wVKal
VonlQrp9sOI9+GEhVqLTwnsX/kBH3PEGwTUPAQjjqr+gVNOEJ/cYXDhClJQ0P9c67QgdnOI+XTdQ
fnSpkZC+FlFK7pDMRdQ4GmfmAhhBl6S2bdX0qpdFPlyzdnsSpg3b+nVBRZYNjs8EgqyYmvmzI5a3
euwviRHMv3Bz9nvfz2rMxVj16QxYPGWgKLXC8o7VONys/cTM4YXgr66vGLsfxhkJkjPKy6elaH7+
O/6gShZ+jUIeP1t+xMhJGFA5fqMCrOvpSTVYK2hrAsA2bH8AXvK4WD6lisQHoLpj8LaK1T0pJtiR
JGs6tA9bzKrDvB7nbsxvpXAob+sIJkYISKUA9z7Lwon5pkjrmYJQNZKZWSSu2T1aw+oGdrttMSvF
aGvMuMvQUsN0/clmV/0mwCIGvPYvFlTzlmUg1JNzlrJJw4gkfedLZj2oQxCvWnS0+lwZV5yfJfWx
KanNTAe2Y0aRKElWgvESci13ZzH1WRyYoKgVzgVfFzkt1Qk3oBKISEBIJTHWUvBg9+m9zcIR8zIH
MCy0wN/mrwrOCgW4KljrRQfx6VGZgIxTJqHmyREGT5ejiXzpOwk0J7sJU4jjn1H6Zxwlw6J20OG1
tq/h5ZaKNHTgECoEYgFt2WMESTZQ0vsqGXj60g0CnIPI6nJEE6dOMgvU+sj0JnMgSV3wPOqX0uLk
EDIqrlpbkjjCtjAu1D+9i00Vbw3rfGma7LZYuCIUsPxDCuzxiBzU4i3pvJ6c3/GHV3dB/5q02qrL
QhFFnQ0M1g+UUEWNvS8i9uFUx3QMkRbaDOIye3P+WXUcGWhVT8oR16rSgV1E1RVB80YHOxPYUBcF
GwT8gmzxglZf4WQ7bB6QhWhjCAdxVETbP7ZKz1wyLnIY5brosciM1oxp3GcRMRpueNcdFodhZgKl
PatXyOE3DR1PZzIm84qGEOreVV+2KRkShKJnaowR9/wXbZ+9rGlMmh2gf4/cwmpsaLnVTh8/ZgHS
U2tTNfz03Fr2N6dZcj7DFlasq6B4tbQZl0t0x8eyyaK1JdtuzWh1XWz8IfN3XktKyBfNEiwfrEmp
J9nuoHwSqbF6BpaVopweFiefZYf0kYqySghoLze0gpkIrtY4tmfNpQMqaUwu6wV1QTBZbG8d/GFk
SOc7N+arIUzmPJzub22M2CD5dk+uCfAIaI8Pv8wrLW3QQxVL16KbNmzP+6SvDIwtASmOf2aG0TMZ
rkN8og61SlPZt+7bJ7jb56WTULB84C8PQxsBg7V5cdwL2nyxIqBOo94MPp1eicCMVfgMRAp2nBTh
JdI0X6NCBjtpTGLvCKVwe37QES+/U6f6iv7MDwWRRCHDeCQwdMQ9u6xBWe1qqJuo+xtiMvF3aaLk
FTGWZ0VYwBNLVhKP+H0Prc/dUKK84N8L/9zZEB+Y8CpedouQ/OQW7ohk9IIAvUVmUebOG3VxwT5c
UE4XrKBAP3HRt+Apk067xZsdEVwawEK2nI/AbvI24RE0xtf7L9EbQoOLap1gWnrgHQEfaS7k9R77
gy1OxTt4spfhblGfW6xuGWd2mleyRM+kp2p3mDUqxe2EgQe5gjrtd6/iQn8Zn6anuGYrEtULjsGH
9uVrXKeV/HcbgMQCooPo+Jkvv0ctcD8/PfQlt0j3OLeeyGQ8o0akDyQUzVo85YKSq3XWu/lj415J
RTZUzkwStohrjIoTP/B6b6WXZJ+/aJKVC500QhgJ+znMtPcE358DN1qbnY7gMa/MordDpBez6RET
rSD8PD06/vMtgqvVwqRpiw4/mpIYL3OjxbQ59lwMlKyOs1wId/1I96OhfgPP9Y35HRNeihmS7Sna
30zwHj59L4VIVrpNWXeAV829N9bdd8h0DgZIvQ1IHX1AUxUfQciLA78+i0rZeHPylJxfyxcx8T75
CdAX7UPvpwFiVBtlbDC2qliPyRocxB/1wN7lkvEEQLWz/q7EN3aWw26YfUTU07M9v2DiFVNLH7zX
xALat4N/m71qyFmrsmD72Z0vlPtp5/wznLgRFvWhfsY4x20ZlpkDoh/GKBpY1aQ4nSY35lkfoQ5V
BTK2ioZ7UTVT0zjyDS1ghsCzpdV9BuNFZQZ0jFzEWrQ59OAAoAcITApKVVnrSg/FFnr8KVF8Fr0a
NF7+4zISzgVu6ynRCPdM6EZ9uaG/SjTWTPbolw//IbDl5bAbFFtr0DpIZSzv7u6D0lrDi0daU/Am
FuBHBb2jlrmzDxervHzjFg6NwP9YD9Zk/iXHHExZrZW83pD58hEXEimGk1J2wlIaJ4h/Lw0C0+ZT
AXp2ijr41Ng9HuZY7x3CJOm3ex0pl9yXNB5ahs8ZwMknCcLRmxDwgLMZaUs3tQBs0bPaxqilrlvb
MeEegNdImNnMUdphV0at/tqoADL0CsIcsaIjQMPtX9rsyszOKVQ70xNpU58vqDGVG7Qh/yDxx5xH
NqAudE+3SkcxVdY14IAg5lwlACmC/jLnE0HbN4usoTGXGJA92d1CT7Z5wwouHjUtA8D75SkXZqXR
9KJ19snKWJRiuxrVFCuAbY8u/x23HB7CPMA58xLPte6a2JbDEHwukfizUI+ZEd0YtE4Jn0M/XSF7
JHJIR+xdPWoWFS0zuK+b4eyES0mxpECHANmMflPIA5fHM75C7+J/lU8nfeS/QQDf9rCdKsrFfiZf
koNG8PzcEN1vKfzVt2QOosM9D5pbvOmHd6enSkYlIOxNAgu4J7Ksnsmq7mws3oXN43K9t0/JsXYF
oIJtgVCfloVFDCHiv/21asE9H/biCphJlSFKpTLedcRXSTNPDClRSQyN745IZBwzhmwtVbVX6RaM
4t538YWImBvPNZ6k2DC69z3OeCKEfWUjtnAzMGgJSoSqvMYgWEmP8odQWxI9dAOYQKxwlGTvqdvA
WFbt51Sz0HRXjOJcWloCwE+1yTDwFIdffC4i8SCN1NfTGh1KGmyzSwMf0UKS2fz7MrVJTkq3/qVy
fzEdvqVsdTj7u03vBt+LaqjsO8D/rea7ojRvFYMfZIsFwa9PEkzNbrejPgRl02QMq+0zoBgOaO8J
EJ3AfXeWuvMnIhs0/sVrl05/TZfiMEPoMMtD8/XryEML4hmSKwAXtFv+f8LUuV7x0VsjAHWT2nPq
iMfCuwmy2LYMXzGxZSO1ZYQTmRIct9n+tYgm6Oe+dxFY4lOUkubWkpIPu0he/uEtsNymDw7i6nRt
8wa7/Wj159xn5oJyvrpK3IClvO6HYqugYtWLGWxJHqzGNDo5o5b/+mktpzvDuYh8lw01tFQXR8Gg
YtVKLB/QfL2SnPddvl1/zlWMe3Cb6fxQ/hUQBa4jHOAYoGBngU4Nb3LsJ3KpZAQz8wGEIWMHeLsS
IKh5hCTceMWzA4q5OCawcQ3x6dCZrnLdto7H4cdlH4+n/fCneJ6dcVreX1KtR6Dw5kpDq1pqBhSE
K4Wv8PAn11uAGfFmYPjXnv2BcRlYcTAjrcdmO/qQU3RNfGFmva8e0n+iJ3XdGq0wztW5xOrRcV/d
bQqa4hqWqX4sDTbkDAAyjB3eO+ubq4W2aAs3Ejhn2rsAaxJZJ9XAB8+8RKZPK6gDR2r3xkMesS7s
FN0Bl9pfT4VM/wPxyEFyJH+fRloGL0EI9xgNbpUU3jj9CoU0Wbk84GcZrivYlM6c5IhC3A99x99l
ThZ5WRsRi9rWO/lHJnVBInSYc49WyoM9BIKB0XOwrigpwsBdkpYCu6stk6/D7LORlujrQtuAyA56
Xp/bA/dMM0RFs2euszxv8u7ib9tmC88tt+FWV0Jl1PX4U5JlATDpn6n1ccydp1RjjlwHjhQEE6oP
CK2pI1mQKj/Jc7qAH1UN/4OpdcUKUalOnJY9YDeculcLAiwgCLy+jKSn/JzJihjsidKuK+hUCj0J
Fe2ypoiKlMf3ZBoP3bGRFfZk3iZ56UhjveTu0vx028Ok3G/eCphjKxeKSRdgj8dTkEdiHOkQGxJb
88Tc3WNq7D+BnTOovZTLB1DnpHyfDQDvdifCDf/bGNyR14P8IXoLMMiWqwVY3A1dnni1Nj91iwew
rVbv2ih/lTU1NvbvAmh8ap3wM8nNWF2Uako3BApQ8oOi1YpcTbpguTK5IO5xYm+RtlclEYeqlVfC
ZLI4o+cXzJJqIPeicQyzytEDbLE3RKxi2HF9jYmd2Cv0ilZt+qzSl2UBPJ/uSs6KMf+ZRbihOOJx
9qU1F3n/RJqvDNQ4nxwejRwjY2gbsdBYaRH7Oj4hAn16cM9A8jKYRBhsFD3AJciVgac5DfWhc+c3
3x8ubMiiIcWt8V+nVnV0z7wQXuAS0yUltroTz6dkzr3Zhf10g6VCdV4aLi9BV7QUlSBNe3VBHAYv
s6C7VH6hO52YkxS0n/sE9qtiEwYXcTDMWbzRQ7REU8ccKnFLbJVkThbuA96OoQ9/3/DcW8GLmQDx
RLtcJ2yKDyEWSDVx5DFTNhKm0/YykRnD/SnZyjFmp0CFWVFAcA4XMXeQ7FSnNgk1cw0hXTstoYYf
pYh16Ndy0R4t+KZJ9tJLIShY/gEcGsWcpI1cucboJzvmeTVoGAW3ERPHzK9vGQ5HevKpsO2dRpMi
RWX74HV5DI1b6lJBiCLjoT66rj4dWPtuIjC9UKhjYWUCrlRB2341eTXE0NuY2qNPCF0vbSeYA8Yq
ovJ5r7Zc+ncUkzPRPH4mNud0I+Dy9a9SIsr8Y/xAASBjfKJI4RlD+tZMiuVy0y0oCw8nAtX3W+6g
UmJm665zakyDPGNsYg1FgAJjA0pR0JJuBH1frLU5gaqUWj5gpkJOHqVuAKjp/QOtv4r4ajXRV4Ek
uB4A56IveBjDspot8f87XTvguiH0v8njuoKRcSTse9ZkQj7veRs6qatsmegnlt8bxP+NAXBeOkrr
HrWPn7Kgy48ZuAv4KU5x4dRvQoMTXiPmwe6qnG37t1RHuILUqZevBA18PGPlK2t21g6Suyplpn3j
DvqhMLLzyMISQVuwkvPoNbukswwwsnUD/ocIadIhcXcen9XYAu/eol3+PBT3ZtuDdco+Dc0U7cz+
gJvp/Ez+lPqIY5MCEVG8ogsReCnR7+1VWCXFpacajDIm8YrfTwle7D0+/dVxL4TN7gMOMzmQ5FZd
MHiX5iMjnmbNOb/pn14yB90ZFye22ay80L+0kmLumODMNltYCjuBwXDlsnKlwFgyK8LukGlY9R+X
RugtU7ctmD1+EXiT1wK5Eu27F0xw81bl0gUjjTF84AisZVWXFV3wxPknkknv497SmaeJvpePwauh
mBUF00RNQuB7d+Bz1fHDGED/ofF67EICJwZUGzD/rDPHoIC38tnR+xr0UAKlpWHF5+OaVR79jDbW
O37f6lThMdNAwm3tqeNI05Lzop71PavNEh5gTPRyr2OrxT3k0+G+rL9LVgfuGQw0QtHbiv3GC0Q9
3L49mD+5MLjzs++lLeyzDYbj7LYraxQ6V+Cti0rBd6JI60lT+H9rxfgl7xyhxthZnzX3g7CMfIpd
vedd6fmq4KFtVlPg+CKIKpZ9Cb3Rc+n1pIbEYx0e1jZu8wi4vWyQIGRUUf+zipdqGT2p9dQoWepM
UKPKTgxQJmHGscoi9dxC1M+h+3zZKXZkYs4jYXGLCCSYbhgdeyaL7dXUdhakmR+mgNdZ/aDD8M8Q
xYvkZ4Dhrc/QAejNRVJVSkSaSkJAeYmLzjr8QsvP9Y93vn3+E4KpupaetFnAqidXD6W0JbKyEv1l
qbzZLa7NOySLnGSn37eI914APOpGTw1DkaFLidXSFkht7kS99aOH8vL3ckNlvjyhn5zFBCSXLHBN
OqwY8XLmrPabvmX52C8Pg8vzHD4hG20IvZv8mQsfsS4TNkOBXBd5YTaJdXU9fcSwvDimd3cNPdLb
Blc4lcyO/oYViszk7An7IWpT5/R1L8a7NOSpUK8D4uiSg1BPNzLlS1CFR8OOJ08E/xmWW1TF0r8F
gBxzNfasMBL+8FTW9wsob+aQqt1duLPV3eVXuR2nEagln0XT7ogQ8gsoLpGLul2harjCHZE7an3i
LEcWH+QD86Qw1U295JNDoWWAkoCCFzQGKzRWaGMR2CrrOTjW41zqUmOif+KOwDb4ylM3CJep2xQX
J45fMdJ7jBauWCrK4k/7dHBjl2HAgR3VL4xNh37bZ8X4xDtoA1Jg1g56vj9pgUl2LSDGVkR8ow9A
H2Pi7omwtrXlePSMug0L6O9+6t89SQzZBQET2wwmzP6wvhT9enSZeloQTvOGvA4LJvLCQQdJsVr4
/10vdWWJUkQV1BM7WTINZ3YFTCdszNmu6QoD3AGn7BBxKVbt6Xs+7xHsfA73XcuYschJb5O/9g/Y
hm0a7MAKDXStdW2loalstB1zbvWFOGM0XEKtHmLwuha1TXZUJMXrx9UoSzcVhvehbqDlwkpzyjwU
XYmWyMcfkNzZVoPntuamUp7AbsQRZKYdJ0tsLTiPvMiWW4VIBsS9Ub2CpldiQMaJ2QgNhj7HzsaJ
mtNGRlPA9nweALFslSCVv5Xeql9f7H7wg8y4QTmO7EZrkB0onW+VG9WaFfO5gRZLxfEP0Z8s7nuZ
4IC+xfTrb/a1mkpRK6SNHAfps/pC74NTyWoaHaUMr5HCKV2MVLqprz5/v/PYEAJrzP+IkKN5ejQn
UGcpbcHyBOYCV/rIS7VpUmibZAN25GDj+96l/X3eKMSrMIm3cE0oVmgEVJV2VcKezPyPyN+Hl9D9
QMKORyEk6Rzucwtx2gj3DgrDnFpHTdKZ221e9xm+cWFkZV5dPrFAp+NhPBJrsymaW1Z8b9AjMcnW
wXH4mx+nXIwQK9FXSGyAFEbAHkiq3Q2+l/IEa/eY72/yYcWKarv/V99FAHdwCzCqipdUF+avxzUI
MT58ARMOpe4m2gE5rC2MJsXUrV8QAsN3B0qg0qIpWMT49SmvW00SHt9aT4EAnXeaz+kuRlbUavqi
pQj+Uq7nP7X8f3SN91A513ih2ZRnx6JfDN2QKKQ974m2hQvfO01HcpDppRhqINuGbaTwxpE7Khgk
IV9rsyY68/cSRq3qV0fDzRsatVgq4Xa/2GtjshE+mm1hfkmzfVhaO8nkwdeoUGP/aVghjtavc359
LtU0+g1YEEryZpvP3pf7W8vlnpyzyJ5/qlYoi0a3OnerU/MfqABdEJPrQW8cvoLVgeFk+jNWMlE7
Ls93eFH3R8NKfPxD3Yvs1Qu2Dtriqv+/vO78oqu3kXFhBvq+2pIoaRdJlgxLwRS+AJve8vd7pDTV
uDdLywiMbq7UjYQhRD9VrW2QxNVzvUOtfclySxGgyRV+FZyCZFtoAYbWvT6srrukBNCKd46LsLQS
WMzxr1eUAiAadVT6bOb8KDOBT1kwtuAjjDTLOKsIdQ/vpyZRTSeqWEXNZVdRXdHLOWJtYC5CDPrc
lsQWPQhSMGkIZM7CBGLn1XTlNT7fFlicBfuEY/MyNMNbPWJAq9ys1xpy7EVsWp3o3fJSBfJ+CRom
cOgoo6M0WGa0cqqjZJrKdHUh1LJzpqh3PqfFVZswtmnfkc+DWEUvSNGe71Dtk37p+hL4VKbzIx6m
eMlU6kSTxTkc7EevXmmQLSxkoVBENSe8IqY618N8flCAYcbnrd99+q2uFoMaP669zv8QLCl6J3gd
c+uTGTaTRrozQ9JalayYdFM86ubq24lIkmc1Gbev05yIHYr42DjBQgPWMcuEF7UNmAWLjC1Vf0t0
Eim3N7UqmHtVlyruB/OG10VlwwwC7cO4n4tUVfqwMHjErxqMrVfEyXuHDD4OIogo3swiMhqSYPnU
CTSZy+Lcy3g/NE/+5mzqKUs4S4zbvw2HL65j0IP8ZOugmEogDAAVSqq0ukkw7Q20ksiPwCqs2El8
A4dx2Cx1TbiRX4hQD8XPSjECw0cOEVENyUYvEBRVCtCBY2oOXKxDfBv1ZOTVDJYY9yj9TxU+7Tom
1FRk+4P1dvfzjBIjYxK33MtzPDDNmzCFNxQUAFuTjH6BSRqwU6tJZRdWj4bO9BcQfvcCjPpZbmvU
WNY5G7Xyr313Uwz/crk/qiOpGQgRJMwPxOJhp2mf2IHpfE/3CK0d0mEWwegZiyZjXepBEG0En6Ie
yn7VBKX5sMrBXSJ3YyPbkyYg/0/YPt0A6os8/v+IJU46cn3rdgkMphn0dZzC9jELyqFCpkRdJCsh
js9PQEm4zTzsk5tB4ryS5QF8Ro1PzhnJiKg07iqqLTjNb5ZWEcOW0VrhpNpc60cd57jqyyM85tfm
Gzi+q7KHZgbIKm3rNxK6vtkpKEVce/HBvPMUogztckfM9Tb3UZ+D+hlQv3eI0foF4uqnLw6WGDl+
PiMcEOUwpn6TZOB2MWE1LqizuSfiXFpDeSXwZyuGoyQNIrGVmyVBtOjGfktfi/LhnNhhS1E1I3z/
Q4tzRzOHuR4M2oN+erP2pbNny1Jcj69u9CWhjC9RUTVIvPAsw0QC/Ba6//lrdnVaJzHmVIA3jUfv
7MsKqoR8HhsyFF2dxcit6stLeoegxNp971MBzq+yxaIrBDx2E9bXilU4fOZN8/WtQ0ogIYvU2EVK
4BdzHuUGwjd+uoem+ekEZ+gUKwSGAOH5B3/jUr0A+uHIVF7R1T+0k7dZ+wfMbZWBwUot7Ss+cE/G
2ITD24uH0XJiGhn7tQ154BsUhiU1UCzLuMUWaYxxkUH/0AkFUg4V4uUikiEy8iz2kPrwFf8RYFFs
ZGe+6k9Ek1QAYnMkCLx8UYJi+9UUeNIoFYovqQA6ugim3BbMyLvFzRNFUIruW5mLguvLQUAvNTpt
eokoT7RdcnKMcd80j4SfJ7b+9bkGV/KMkn4ZVKj8bnFwUQ/Tv+Mqib4VK39zr562fbltBIEtkbo2
2ApN+rF8hR63KHynzBYTuy/Yf8qM/RDn0P1xdQO6qguGEYoXynWd9p7qGofhnqWWqxmnbguqacPs
Mx3PPcHt5eaoJDyIjAfoCk3LULR3pEEjvVakJZPb3fCjCHjfVTvPwG0rChWa5dY5m2rqOir/AjHd
cCb4e5n+KPy0DWJgQJXHcIk2YMGMThlnEEsmyrPt+q/zyPsb9OJZ5RGuCyt0oYxBmgQLrOViGrBw
yOr9do6C4s8UNDmE2NTufFb9p1n6P8VnjQshB6+yOdjGapVTKNQx2lDyoYrrGD/QBQGjkWKpHvUr
OPt1WOmdGzaPEvFcg2seq70eM4FyH2XHpdPPX9zegdoQDqqJ9r+nMUrwDYmM9LC5OOsg73SRe5ET
Lcj1phpl8LVd89myQdil8IZTO8W6u+BBDytyUnt/J2cumZ9Dv7bVBlrD3fAm1jghE1sZmongOrup
2V1b2PB4KpRhj78/y5NlmGq20zMQ+xSeWkVCi6fGHkc25aWIfftH9Yz6AYy+FcLT3ietAfvWdHKy
eyzQWSrecA/J8YupOpnRTMx/I1jOzdPMOdqOuDv+QLsFxM/kZRvf5bqJat/K6Nn6SjJDptMdwu7u
SIonhRYGzt6lRwKio5yAb6zO9/ffV5PmVEoxUIROCyhtq0wUDC8hsNuaq4Q4R8bKIJ8CeB02DXOv
EIhjk1qWXNQpsTDFrfaWqETR/wZEhosczMNteYVKBwoEL2aG4JGd9fWJW0bx5oe4ic+N87cy+Lpk
zkFLjIfVX+YM1ncbystuWdkmWlWVM5qWWxDh+iLGm+f88+5Y/iYeW9xx0HroCp+1M0/TInoHNM2p
ngaVR1kacpv53eploaNkRsz1gkUF9tTjg/ToMhpgQPaZTzKCdCGfoLlMdP/4M83rNePYcYRsyFXy
EGjkzTmzanzId3sloVDOLq0aqY7F8UT78KzH1oV4/xwjjba7XRHClUYKoKSi+j5KgXAdW8wpnsm5
rjzRrxDgzwMAT1kNRq47bUoWsLm/O8QRmBtUbJqe0FMea5YcjPBWb79x4i99KfQbYrJbUDnXkhC4
/nla4QPA1BGytBsWdjHsWCZq9yGdtfIrmbOpbz43F+wFb54/h6tnOreQ1KugRLMxxcca+9XjQvDo
+libAjxy0ASZWmdc9U9UywYd9zO5ICDL2eu/QA7H0bA1hHB77N+3ps1AjVmnCkzYx8/Szeoxn94i
0rkHc0Qi2dmc+C/eoYKFeOzuDG6qPxhMT9jHfokXuA5k9VKsnflvy2ow5bZUxW1ezFl1W2NSaX9V
eIJRmlcFrbMfEX+0xIP05nN63rGPDHQZUkaMN/kMbbjdyYmXfMjmInQCtejJVrfAshE6oAjNgs9i
Zx1O87WDIWpeVYt8/GVFgrMWX1og/N+eWuRiSw9Rma7iw+jGMTcpWRoiK2XSJpwpOz8aJ5ExsQjN
CWdSTZ5/CQV4Isgq1t5IOAxak8u71zJdL0L27PI1FeZ1F5OV2yJN084SLlzaXMIMK7avBqXoWT3Q
nYZPOgTSVWKzmE7NZQfnhNeVySh3cggEQ6yGYHVZObDVycCju3nYwXLSLSZTKnKZygpyJp91MaDu
ZiFyZegDvhIp9uZhpGHwEqOy4OMMXPJu2uXwz/DmiwaZaycmwhj1WjY5L/+8PsMbMyOlaEVSOqoq
KGfN/ItyiSFcD7acyDRH6yBC3PyZLfOl6Rjl82zhkDUbSyokev20vznCOqUw4RUSbl88iGgiWKGw
mHXiPE1uwNBrPZIjn+ilHJx6dLJLjbiMRvMX2MZAGZxOGZkG+WROHFdVQveeCGeH/sZat+0Ksfw0
dUNsI4pzpcUkpE2FFjiIsrgEcqmW/Se5h/kR0j47BD7AcDoDsa1OWQJs8+en83fW2yCCnISiPfqS
eCTER8H4/RdhW/u/ZnlD/vqVLyKxNDxD6SbYPhYgy2a4DtLqctQ61V+iJe7nD7rp1LDIZjeEckic
1fodnFdTCYC7exCB9PyIsN7hcHhxEftVXtZHAGF4lW75L5O6e0NBwCs4pDTA4/T4WrD50cK7l7Sy
Hg6UzIGvzid5HopWpydC9a12NEy28CE2jb4NzC2m+J3nmDGWI1hXkxyHve3kqo9NVYBrug11uV9H
cMiM2srFlo51bpY+CtpBxC7R1Z3qbm0Iyg1NPYVUJyfdgtyyvKS888w3ADoUYJedIoXLzAybNqi+
PdsgR0IlfYTxIIJKFj1E51kxrKMIHPQHRgFG3q+MR0z567vWNWpaSliy4OjJhwjSWxRfwd5qF0E5
D/c2akpwGo+8uLfLUk5Cb2xn4+1SpxcezjYG7Oblx13Tlfom7trRHM3wUJFvAX4/QW40U57NGfon
DHNpef3ZafIz5STuv4JAC/9r7V9kwGv6Wa2CRpHEms25kBZjJILpEU6uMKV370jqoadeWYtLau+M
2mY0NeUOtKTjuuAfmw86zYpp8CBFp+9isl+g65eCveYXyEHzgBP9ao1xDlVs5OkF4OCnZ1Pdw7r3
El1UdfQZVipkMPW3kwE2PXiIWfLqOBa9grfXuu31niyINwro+poBCGItvxfAqjComosn8bEBEFLI
uiS5ew8mwkbXj6ouZEeFHmXxDUI2YcwiG3UTjtKflbnaHYbf+SgdOrDvJfRdFG/r/zbfJ/vfiw/Z
znRPiTXE2Tn+1sj8VBbIAhFuR8pjndA4H8T0wXgcfPgT9WoZhCipFQRjze+XVyy4k7FZDKCtlwHD
DYF0FaUpULT8Nw1Jg8lrLHNGROzb1WR0/Qoh/zha4ild1696ie6ELHw53Q2mCMo2L3sBJjRM8a2K
tp4Es3vXlSGzYfpQmoVUFYGF9iNSY8NB93e+woVTpdIH7g/IdxEhGO7XlCOwuU196xUhmW3ngWe7
V9NcgAhSbKvI3OyA7Dynrpk21QK/yibJ08ZZtoo1SQ8eC7W7Gz7NQ2xERcCEDk/7JqeKE9z3YLHq
uU/QqiER4hdVEpNWaZLMvlgA+cZbwlQDnyUzNecyspLX1U5TI77tLq/ezK8Q6hEfcNZnFxHbOpUt
83CK+L1vZPMSe/VJkg0UNJfdcApdy8mW81JLpH9h3If65wuNhaQ2GdpMpE2pFgMfGj0Hy5cF13DK
M9bXW4hrqv96W1Y7vBVCd1uPUjRAfy7ofziMue0a7BJy/sm7+C/i14VDJd7IhKreUMrfaB9tD4e/
QMHKqkj/FGrURuQayFkgTOYpbH3wedaTwG96Q62+RwYPirL8/VPAY8c0gzID/Hv4XhXkSwBDCFpX
6V11Bhvn/gBBHZGunuwIjB7qjfD6WQ2iutEkCYQugmyNIyuFFXP/R+0/CuHu7NuwdpHgDesLUlvu
DszvpGSCdXhjf9hKVgaeoJuy1s8WrTKCwY1kymvQ86mHd1L1a7AU+rdL285kpdpvUrabY5ltrJCX
43D0jpV2C/Mxhei+602nORx6jC1Hba92IXtGSX9CZE9GEFY3yjQt2IjpooX8hR1JKkL7OasoCjjJ
9GFoOjw9wniSaMHRekgWBaaeQcqc6FC2ChsU315gYccjAG8Qh+KvEtwwU1+YpltIYCxom5EU8xiU
g5Ufx8r6PQC9oo0qNqUYjIBvR0XgGCueKEV0V8KDDGcFRyZyGUxOdrSidiYSJd6KQAh3rbkDPDzM
v3KH9h9qMUbQcvqm2srcJV5WjIo62cuSur/rZBuMRcK+Q6K8hQj1fx+fFLD7ZkY2FGfAsqrGVwve
nRqTJbPqLhdG+XdfOKjMtWitsDMDjvZg5y7cyalY2D+YpxJvJwYh1fj+rcWXXLYkefZOxGJbNoZB
kZ3kb3BIDDZTDPJCRWdwLrSt/hPMn8RodrBb2+c2JMJ+jmojm/9X9O0RuN0HIvgA8asF1ocb3y2k
zFIGfzMhOZnvMINvNxGUyQicawD+WbRuIjx8lbNr+lvOp4zJdFt5SIK35GrCM6B3JRucNMrcq2Ha
kiLFBdgsDwsVqzbxM71YidIBctEYXHu3Lo2tS+h/YZIaJhq5psGPaVkJQZ+b9LOSMiYSOrhAEjN2
U4+FmlcaLvl4ol5fEL0PXXBRWZxJuMAbS75UJgcGOHQac8Vm1Fv6FPPetWUSAjea7guUcsLYfo+P
CT9yIKoItKGyLijv7i5ZthC3yLCp/s58Q45veOpK2oPWuKeR9BooMkp/ntnC18V37D3PZqpox7Fg
bJtkYA1J+2oLVKyHcVq6ijlyHVlA6OUaR7Hq7q1FNYLDUFh7Bf5YrDl184MTvXvRB62mR2zPzaGJ
O0OOKT/IIcIK/c+HgI1ZzlfQCcd1MW8YgwRyW2o5803ePOF/L+lzekU8LElSROYdmTu3N0WDWYYc
j00Ny4KVZEXL6VeiAHxiKPqh2nB+H+mMb97er62R6ABRHUNC1ADgWM/Y3aV3TgRqIfgzWPeacdX5
Gn6CmyCkFZypDZ4HVzgcGFG5cMVKtKDW5DqCF63S/94pessHY75KjchzuGMkyy8fi3FRFVcoJvNw
kglH44T8fPmYwgaL6oN+QhWhkpAdbzuLz2kGGufJwJ26O12md0W73saDoxQH5t2zdcwgQ5XR2rG7
TwmpqkkMakb3rT7oTHp+ESc2w33KJUAO8bpoSsITmunEgoU4iUSoY0cS6uLCqcJgqfqq4yLz0sAT
w9H7wd75Mph+cQOx49OwQqBYUsnLsuc8FN8k7useC6p+TwjSdkY5oqoNh2pczT5NGVYKbyFrvJZx
YN57ZdseQOPYQPQ4vmZItfOv33h0deOt6xoxYkwB/NCzRa4GdyJRL4ZrvEQHkPvqsvebp+yF6gCi
1dTnWlaZqWEqGjbo4KB20CvoXfXoRp4UeTMllAKY9UEJZVf47LAfqyf82QFQ4+SwcZvQ54+/TVdu
aWapMK+nhS155IRG75x6wUGL+y0dru3hb1728VWD+PWtdePEsMbjKaznEGqqpyIjzIbUVKOLbqau
XDH8SXlfTEDIXBOChvaYsEdk2aHok4eH1LlGIzHfk1bhQcoAMBX42y2ek1wrBBhV1/x/3Z2Bx6LG
X/M8okFS4ndkiUHgLpT8dEKzmCDX9tgaIJQHoEMP1dTMOC6Du0f+xbRfYLJ+qxaATV7HQVBdnGAY
i0d8MKZulHO9j5EVC/8eXpiDqBGp4H7+rTAW3faRxpq3QlqTbAGTmnjjqgZD9oYzWcQkgXLovGpe
8lnsYvZsMEXlYWwPuQO5oBvu/pFK6viL9uVX+C5krjHQKjzkNstjcZLPdtTl3Mqg0VJS75Q9MBCT
DnvSx+LWLHS25XNiRRsgWj4qny86VmawOBITKfy3SFHh25e3AeDeUcwqVfjH8iRCMczAQn602ZMU
OPP5htW7BFyoGsrhWl5lALxLutKzYBu6Ygt/xdPGFAUFwFH6jZENfxIl2XiEOGuQevPk8H91fttS
7aWBoefQhgJ+x8XJRrOjg4+/WOcPzdnlk96OiSgv1X33kivj5r1ecLE45MQo1+lh34Q22GyN8PYD
bhULZS/6USu27vLIDeTQobiIFLKpvCg/+syU+fXquNoAYI/HpMsojwPlKTUm7tXlXVUxOsf+Fw5j
HiJnO9ggvlHipUaqWMEAttipUvqvfQKyNs/Qk5uwNBw889B5fVVhNS/vOAvjbvbYhE4AHj5NvG1V
AVCZ2v/LFwdz0+ZM8qBDftwnYRUbbmhK6SKnZlo7hjZaW1Jh63Bej98pVM4LB+cPq52+MO+U88nH
+MvPLkoOV+zDztImMU8HcA4aINR2gyuAO6gQCFJqxn4SZn8zXbN2t/2CX0mO1ZlphHrIM0Cc/ezS
zDiEmSJ9jVWzHEueJcFODD8LoM78YxZA2BCsw+R/Id84cLTIY+uzH1PtL1So53/Fi03toOi8FZ9K
vQGDxjwwwKY5/lW8AVWETB/z/0AIrqoE/4NZsiL0XOX3/FrJJV65kfmvHwRicsiBrRzYbL1iJMtD
LzgzRKFDmLI/oQp1AFn8mA7yuR66feYlMPKpUtVPN0YY4K22ZML6NgfNLrehLj7+ubdOSS8RE4eX
aJQY++gmvm9brziZ/9LWzwceuQ0XJrGwCeVZPzSZo5MHB7WvU8/RF9zaVTuwb7ZR1X9Wt8Zb4KYU
aQALGn9LdXQWM60hBuDAqe8nH4FMhtm0uCoTQz+cPevT4odcnxflpp5eCTHaFNl5wsUdKjV6T4LD
3N6DnzwaBSo0c/dNZKxzaWB75i8T3x9nIH0dNdVtf/IHTcfBRBe0dQxMQUBGDuyH3wmpHQteQ1J7
kyuxgTNdz8/VO10nj2HoWdBiq5znkW6hT7ndqWdMpjJ2hroYw6HWlywzbFFpTOpMB1zyXon6zH82
x9K4GZtDDaKWu00liHiva/qdj+6+ibQCHVG5a0GOu6QYYR8zhWjoqhsPw4AnoeXBDjgqIlFGOYbn
Tk/6RueeMbTl+QmWexehlaiCcEmK5D/PpBgwIGlzAroHIfWExyl4aLERgKiFcU7tfsqy0YPfcjbv
LUlRsLjKLk+pSQ1iVJ2RRrsY08/3ipoqhPOMBjMnPYNHeJW6oeRw4SM4aP5/ntQAyMF3MX3rC+1e
/8WPYMPxn05VSndjd47C2tR3nK2C+YPUYQmodr5n6p0Me5yPFfsGPQQKgn5JjwQDilVjZa6KxN5Q
XUr1YBu3BAccabmK0ViJY0VvuWin7lTa0l1C+HlwBg/rQO0DOfJVwXuta3ozw9pHcWiiiiwKmTKm
9WLEd/wzg5n4POymIZL0HHFdGDbw+WboxxTHSZRi30nvyQBT4COymDQyD2LrQA+SyKCIapXAvoZ8
ENhpOuqRsusEgcIm5z7h0eMkLwYuOo3IKzNsQv16ydAqfuX4upnXmBi1OFY0Q4LPCBNwG4aZJMQM
zui47DtvKWOxTmArbtPDEHSV27YLI7lKMyz+XaSk8MlWZiaTkynO0Aa5cwb5JVkt0+iiy24ByOEK
ws1dQoDXxejlYapRM0qo3hKio2x2G9WTUqXZO0LbkZXRKKDgnhj+Qwg60i75vEEf1Nkw52bx+/xu
bFkkJxlBfR7pVbqauVfoa7TTXWwTZoZTRMNrKzK1WoF9N2lBd7kfXr3e/ad9hUXfPszzlPhQJ6k9
0fk3pvTFQ6UnuW9BEk8rZLmEQFWbD4L9O3Z6zDNzF2Ipihmv44kdW8qC3ND74WCeDllkjFL60l6r
7KjAcVK8Dy1zp3UA5cY/DH0u4yX+K31BO2qHquvNFA7QQNYFhboLtkT4dHVXGiJfr6CESnfwKaTf
L3sID+MpMj8xnTrMb44XVll711qzKaV64INVbAZr+ehHzl4VE+CLt/fb01N5ScyR9h/vWCoirllB
tsWQVHykRNbjuHzZS6Ubmit9NNSck3xU8BlQr/TgD7C8N2rc/GFisr8CdiQ5kp44G07y1l6Fv4TX
tSxoEbAhVKU//Y+XV9orpXNjz4Y6/cwg1Apft+d9nQVQC4S1Gfe4ZI05NOmqI/2L+hOQTSQs7YNa
zU7J/+esn4FyzH0j1lcE7VDOgp2AnwcL5HYrUjnAbTtjE31C7IqS8CcSEmyN/YSRZPQhCbnjLGdN
7htzVvzCTpftzPC0K5+tcH6AwEjYAalfusV1/51DpSbFwzZbXWb93APum+m/twvXUZu1JqGmEEOs
MaGPI7QZ3aKMK1uAqTpzDfKSHBmG9MO3vBlVk2V4tvo9zRXXZnDZxfDP4HpKGqv4oou2U9PgIHdg
kGibHdPzvowiKm7ELoxM22cm7He6jNZZ7Q0AzSvMwmQPFIUqFq1FiwtwbUCDWrp01lxZBEQ+WDzB
1ObNwQ8Vk8OX/UnnQCNfylU4VoW4RwayGESpokvgR/BBGEa91oQ/Af7MzZKsEJkDgXcjbcrxz5RZ
OsPLf7QKOlqhO1oVcqRNJkF4kLZsGpT1BkpGisFaF4sZ3tp8FQXFGlM3EX+WsuPpQfRHPLkTTslW
C6VsJS0Egh6ZVsa5cwocEhFQEtDIvjCn5j7tDpudRcpVpw2XWCw8pGUmHnP6TH2lmKQZJ8OjUlEU
rR4ytuuFkIL85gOOKJ0e19tR16NISd9yFzVcjKg7pOxiWXXGWkuAgLVWMcbcmigwc8/oDkRDoTt7
o5Xt/6dS7tFmg6zahb1cGfd7Au7k00olDo6VX8yboMWIEfn8eMgUl4OtIidIJnDSezulNkyr8uiN
sINJxkgjH7qDgcOyoQ56tCyNnvL2Q6jWkmIyjwA3fVk5g2zQum3ivUxrJtfGTlbdW/yYpaawOuOh
Q289BqNeHl33zV5Xbx23ZX1pUGqFsV2t96/AmGvIM9fcOvSdODtziTWNzZznCPKoP7QXNCCwJGYR
YmaW92nQ5xVKD92uTFCQF3pF6odaVV0zspmbLGcXPt3a4YTEQIaIDP3YvMCey7tEeiA880ZxA9hU
4NTtpMtkKQy6hl5qxc197Q+OqvGDFmNslWJ64cZhPnGI07ZBcS6pWhUCp/pgJPucULfT1Mf8uIE9
2g7p0FZBoJfu53e+LoxRzE3iM4Ew1toR4ks2nh837m109LHrDXsEwD5XNrDHp9VuIEZhVy8/T6/u
PJw/AINyU44xwgVt4kYR6zuvF9wVasCJMuGbZNQhkgwU3o+Ztc8j46pCuzcRhVJ/7sBgearWPChI
200ekr5tajXauCCVpf/jgLlRkIVLgTJDX545vbsH8/c9Zi+7W+mqq4jIKgKMuZXSuY6awJg+AX0y
c9RIhRdHIiCP1J3hrMtWDT5RXOIXYgZwF70zniUOSvv9E6/9vDNq00WsoXxl32cZhfhMJNwdUe7V
NlEkJyRe7vXf9JWZs6RFjlComCWsWGEQYrvBY8iWCksXiGk6Q9GzWo0zdugrgbRJtvRQPNBV4Ct1
p764bFipTiNCNyIYySda48EUziHGIrZCYd243MtZpx1JDJzSRF7gpH28rDZ+26i3uOFV8EK52LLe
K0GpzaGcKlBnSi1exm+LN1CBgu6xNswEHfzfQdzanrQQWDfOLz0WQ0294vdwMS1BC4/06F3ISocx
zTGMCx0nYoRPva8kIrLzCZghO5sHDSlkumvQoqzzZn2FjV7ttcbuizFebrPYymT4pofG0mPOq5cB
WzNY/PFjhGdZ0vPFU07yKNFfowxMk8Dtt094eYxdanuFq4Qe6zYDYYZ7nq9n3v6M9F+o30XxeNda
zlkEuIJ5YLyXeYU6wqoIru0bCMI+QZ0E/RZ0ORIfkfHXBb9KCmq1ng1sMuU2u/wajHSlSEd29qS5
9Gb3ROoR1PmRxB8wk7pNpQZAHmHfU6djON1lHK27Oqxmb0wNAApBw26dXlX4dnMg9Uun2IsxZc/R
nBxFmyoWRJyOCGww+g6+zRTI1sO/hUf8H8IOH/CgcbR87DDr0hF1FhCUU+V0VzvOJDV1tAL2FAU1
qENvhz+1snVOY6bh15Bh/BFsY5KfwX2vSu7WG6djaoRqZkjly1ziggo8FK2YcQz76q9ys/IEjC8F
i4tQ8V1d9jhKjFSA9ga5AMjsvndGAyG36qWaj3SrbFUHb4Ki6YceNNRSoi4qqssyi+03Am7M+4Zg
dzlqKxCttb09AzNjkwmEZD7xUevDJEpriVA4tKFWvZOyDXTT1jN+yffar7SzrRK3hp874t/E5Mag
+Cn37IQMsgb06CmvIMty5N+9VF31SEUEC/olu3sGnHFAKIjTGqntCV2FMUJeNREhsFLCYJREtMaq
IDEMhPp93I8w8ePrAvVUc857oTB/+Gfkg+XS6YP3fhCYEAgINipAppBm+TRnUYeEzZymOogz/CqG
2qc6n/08ztnjTqIohrvh44pVhU6bMU9drGXPdu1g2L5ObDRWZlwUdxabTkmmeIrdyknSq4gCCeaw
HdPn2N5hPLmY6d4SKATDwvaTBcr4wolmhmo9jC7Zp+HSUrcpZeG/JPt4twMw3l27zXjVpMC8bM99
olGNzWkYJfXnmUcsYOHBmVYbAldtgqTvZJZNwt3+bPphJlTwXXMZpQsa1t+wFB93YyWSrxdupNd6
VJU+1Is2S4nq9NcEJH8CqsPNu79YQRaFaYXZmowCUvtQRaUr1MyxEErd0riiMufmRmgo4ankLrFP
glitpJcRm1fJwuJp13qWvV8Qb7EjDEMFX/hpXre1WsaRPcHSivX5gSsnZ12jXgHXGH2sYkEgZVQ1
S9V4t2LlR6HNKXV7YggeEmC1Fmv8hVVAbOqKTN4KLbbt31igF9IteenmJtJrflcYh4lfvtsuYFd3
pGUd1z7wGdCjh1yNNXqwMom7Apiivxbw8t3gq2aEZC5LpMAc7OkgzyvZbn2YqRe1c1WrH9OsyzSp
llAJTapxmCwhHdWWAtgYyFuK3mOGHHBHKGAKU8K+H1ZbZXAluXAnjHY+jw2UDTFvNa21cok/LEKY
JVjr210XYUP/FgUuG4fD5bRg+iAlCQP/eUuWy39oVdAlB4DJvl8cF0n8zLifRSOW3II4B9IAM3tR
ACOaYfvLGnwCK2/8e1lQRYnfkPpwH5qmGqAcMThcEPhz5w/z5jzlvdxqNFIJQaFNtNG/arf6CQHk
0vlsN+cZF0kLPusuXldRdkTzEeRmOET3e9MRJt3IC0fm9piHfzkZAxrIsP64F74sqqLUf+mNsNMV
z/37gH8HCBn5ZlTMtSgn8tvHKMaf4d7erbvuWjqYX0YKzaYGte+qi7su+kF6VfQ30G5P3Fput5gO
cvEM5OG2UtN0E49La9j22GTdWmkZofjCH8oLCILEcNSpZH1zxz25d1QqxzucyvBPkzzb+9B7H6b6
lLQ4HTPlzkFKOrMFn8kO5p+/2qZewpO2Cul1naBnSr/YnkrGRKlPbTGyCnLA5omz7TyM+eYl/QqB
AwA3H2UYaz/5zOrkMagaC2fbTmyw7+x0mOOsddTiNlCBIW9Y6bF0E0t1wXyJd0VsW+0G4Q+Le9CD
WoXpcJwVHThreYHtYHlAN9ztysKAfjVIk8xOioe/Tsv5mYZu/kdhAffuSjNnte1+85B1JQNZHYzY
dCJ7sImLO/e6TwiPaLmKQoKAOWTMlqHq0zLNUmfRhtgYRg/QERqsTqPQrLU44d9d/vrRdUQnv7yT
GX0uIFKyHt1jd0tcclWgebFsqV5IZ4PYtEs9yIl/cjMCPIE/6X2Xpc8dOCBjpssr7AxrnE39HcMQ
tJp7lPx9Ua0ohDMbSm5wowVIz9Xisk6t/p3s+VrpAQvBVnx9Q0+8gGx9p6S0jlmqGIeh4wz+Gqhq
5TG2kvPbx0G9Yrm1tRJV0XYfFVDtc8ecwc9/GDlCA8nb2Zm6ATEPqrIv3EidqoDqSCwPcCK9/lDq
1t2fciz9HUApuxKrq1NndqttiHT4gzVMzyuYOhPqeC9Ifct+drnIh9dknSTy5G+8G3PVDA/FumYM
Z2cfze7uhZvumwkF6rZ0kxSXfgP0ZepKtJ5CzQNYL50prq5utVVtxVRmmviXd/E7dUUT1+uQhBDH
pP7tMghZrOKoZubhCt92tiHCcs0o9//6k22H2RFPr3YW/Czk4wsKp+tq4v5J+2pxyK+gkOoSPOiD
Won101+GKPDGAzNyRTXdANnD1Fv8J8JBt98wW6hDSkRmTqpoxjqDb7c7pLGoAQHhSVS4++V9DNOf
AWLiadnr+HUx2FUtX/zhDotKjnl8AeE/ddetgKmtU+miTxs+g4Wn77VlxlYUT2+y49zZSc/2SW3v
vF7Cpb0xMkTpZod8aJ1+mZRv1TWlAAC8DRAvQqLAVbNocbtZmRG3oxYGOPUq2Rllj9I1mhErjBS1
yD61rPHdDuriJM9GeLioEIx7t3MTsQNO7C8nxgiOEztE/UN9YCC4TWnui5fggx5//t7wKVHKByby
P4luSDYTVsbpwxkaI0ykUINeUzM9S1qdB7RqX5kzWXjyXRBDGsmqmCwRkpGgK7KyE8+KsLQ5AV31
T4DWO2vh0eq4F279IQD0Lu8QFy1G1/nrVOcP7qTn9OdfxrUsI9VTM4OFsmc8/7u1Dp42RkOzU0YY
f8aLKdE2PW0oh2PGOr3R5sy7RkeDCjWXY7fsUoaQocOC/9VNuTjaH2TADvjn0td6ZbWfjpse7qdQ
KJhEqoJ2jMHz/lhrELSuOwkcyPXymUi2XZR1LWUW5Wo7mz/wmmBu2e8Nw1lG3iUtjs3SkA8G6RKD
b9pnKkCfTCWWcENo5r3J+E4d1N3DckzyxjB/Wo2lEN1GvyUBG67PYwE3SJCgKXdhwC2auYbn0y/P
P69i3I5f7LW77l6gaRi1KcGx3qieBUXGkx+XlvAPUL8S94j3uEOWkFykXuXq+V2KRJw7+ozIU0+L
duBVB0CgOLyxaXMrWrlsFwtVfxBtOaEKAVQESCBw56JT/yVk+XNku/cj1iWbt+FPHAKLIQr6fX5O
psLEr81r96tjC8ZTDIhMvbkhKPLR6kmtS3zn7vKYc8f5L+D9I+ppEyc6Qz/xYVhtWnzuXnUsUNFG
1CVBPDkSi+j9sv/HkWoV+YBe+s95c1NxlNGBesn4BC2ZS5B6QRl2ofbyBcVKnD4ZneTzcvGZU6xW
ocH8Dq8poNVf8battNuv9dH8KhZQ9wmce5DTmd8SWRQkHd6yQvttYeKBl/tb8fmf9EmR94iSEjuL
Fa4nQWM/CY+4DxiVI+7ooOPRRGytoFC0hQ43SpRI4cIS5Us91eHhL3V/BD/iVYu5jT2FcbI3qlV1
llO/UOSkESAFWrzTCgUkKuw3pf80xrjHTWgaOYsUZ0zcAMIG2Eu2850238anSz6nE8P2VWlPZcWH
sRGdXGM7N5nlbHdMaP9fZFNYgy7tFjYwASUiolrvg7y+rHBqLOExjO4AV2P409Gqa3ZWmNlZxgDt
W7qER8bqKBSiODKA60na5W/2jo2E4wej6uuiwd1v+W6/NYi+j/eYMfXdku5HbvRZurBHU7uOt4Ki
4vYuz9DoihjN1ONyOA6Ec+I6wbegq5I95sP3kE+3PuM9DJev0o7QAM7NvNHYyEKWknGT/ZW4nbX9
YAMCWoWg90Nv35FnU1TkCHwow0N9yyvSk+3FIWDnNpnGlFVELY4mzwHHAR5tbg+zhrOg81puYaIL
RY9gNaaPIgfwQsx+FFgA0uUwxgXWbZgdnhTpamwHRjFqxEsrBwlu6ihkpYnSsDTLvmAiPBgzGTMO
DZtOPdf6vtgfaE+CAXnq0jWPRXPz4KO4TDxDyKCMrx4eLx4+ZscrQOANbTS8OjDMai6ZpdLyGTTk
InGG/lxheBBW78R9shjTsxJSoGUZlIG0IUCPm6nN1x6PFwl0LfxAO6gwKtNI0SbXkMBZQd5s+vON
G49mYPBihKlyVhylS+ML2Dv8EW6fktfUemQPjbSs8juB2qKS7u5Nvgd3HpghSUESUDztk5kbGjdZ
ulnzXIO+RVuJdfUQrIuLfKmVVw6cXmS0Wiv4LXAtbjdLVkXzBOvw+9t6Oi/tKHYz9vo812gOt4hZ
PgfMjTxKtOUnDFbNQns4pSoFIAVkyiWCcpCyMDSLzVSREbR25WM3AUY7ldZP+H0CsYHcRSoFyjNp
43Z05KNXV0O56oAwVGc2VNNde3B+iRE7nVnP8x/2lhu84VTr8AbSaQXcblHewxRaG88KqL3hbJBX
ky+0rIQ29xQ/c8r1zyRkfdxCaFJV404t3uc3gCE/W/kg6AGqiG4pbDJyoP0AV6sj7GOg6/ZNFftq
MuiC3EDxbvKoxFXnMQRTH9knEULyRpCPmnEhwdkfM+vjSc1iO9DaIBnlTfsmpxjKuCaHG3T75JIy
EN+AoNRyy/JkVApOu5kR8m/yyRXP5/v5m5WwCoIir5XqiuvA7CbBOLERhKPn1ITrIqScbSsmuswu
yz4xmopWU2Qoh+cJ6VRnBdo20GEJIKRfSm1YN6mf0xHa0xyp4lJCYFUG81v2ZQA9VLcJRZVkY3Sv
Ht2kTRU3uW0XsN0LF/IKbZxuTOpCsgtM1o6Gq8cuirsv4lcMWXqnx4MFfEy2zUQBFqtuk/2wEEDh
qoDX6EC6apaF6wCNNFNUsnX1pP0c1T4gZVIXKAlvaDF2YVKTrUmMVKL10JahQ41AZC+WH7QmIFHC
L86v1Cd6VblfjEIhafczmiqjjd898+P8vISpbpOrEp5BX6ptvyeS9DcDRW8aFS1UplbFm845dLN/
AqALUQtlsJ8LAQUWDy1s7w0B1++gYi+zRwJTyYGUnpBfzRFDJd2qRLZ0rXX5Dm27keif/wIpRLS1
h6ihUqMwDAvhmuJcxpke+kFRhCBjJ/a+aM8WI145/XLZfQ5u1TWkfp+1UhO7WULHzfJQmkq5oHIH
KOhzZvXyE7BWRk8N1AFohUEjKraMpCddZLbGrroyiQGD9wayvPsmTj+ElSnTb1rT0CczI8If2UMn
sJYTZUVponpONwHwe68FQ8aC0cOGZxvgnsdNbmzbjNSuNl7Wly+kDF3QC24D4AKlSsx23Edy6wTh
e4FyOv7dvsVh/QFuf0kMbygYKK+BJhrX8oGO4UN9MrDJ92leIIIhgMV8PWxDNthmj2YDe8zvidXr
sNvBsuZJFnybv61JajRr1cpixKKxQpKE9RXZINJs+GI8u7rRuuifxcfRYRnb4DAnhaoI+F+ram1W
NoNd9sil82uPDI9RQAQkDbrlrbd+RjUJ6A0YQMzTdI8ZWGyKxmNVH8pQ7itgruH+HhVwivnBgLvN
GiXiih7I4vJ49vhGEoQBE4D4ZZ5KUHwl8dK0Sy6UtX60dabwO09ar0B/bu9pRBN38ziSiDuDtsDJ
j1u2Of3nSgVyVPOkEwotrtnh58epw/tUg447q2Ub/jBUSOMa1cRpV9/crleTbWT0F/DKdxHmqqgx
WxzjZ3KGtudueUXVJNvHQXDD+0Q5o23vQ+jZUPAbyu2eicagJTlSxExCSHCFG3yBrjSvwvu3xuVc
ltw9ghQAStjQzEnFTqWZUFjlAe1mpMODKCg4wvPjTurtBtqIE6YfSeh6C7kCTCdSPfqaE0r482G9
4wisfyD1Uc08ijlqvTqx2I8vcAVWUw8B+IsfVQQQP8Lw7QvWXw/OtyVT6UhzzIjgY+rfe1znpflc
wCmpMw9DY3ehzSK9VwHdAZ0ShGh87JN5YPWgFTzYLuNnTiqQ89IU9H1snbF3FAHjyQHCFis/Skrh
UpQT2KjvPeaGZ4/BeIcVR9fiU9HP5/hzyDEMEGEegPzhvV0tY4Ueepb0BHD2R1OIeav5s7BSUna/
1EolPg+VeSisQe+4t0o22eyx3mze0o6YoR4V1acEgKiKOglAZzNMuvQwUB7RXA8FDeWtCg1PZDHV
2ZKQiBRdGfuUqYDiS3lxWvL5+Ov1Kz1ZcDi2q/EJ/8yUgSHuSbkBDhZkw8sNZi23mdmE1gWqvu7x
HgGYqYa0xEvQahc/5VCtVGhovYxN3FHwc4zv9VEFLytLMRkGEz0H0HV5z4Q+Z4BTAsZ0cu4l9m80
afYwEG3VWL29FARJvHlkKL9A8yRNmIjactj1Vjt6xYkDvS+nvLnEyjIoYRsxabr1HTeCL/+rs3C/
2oBq7ht0NcXpliGumIZXvZCqRHbs/WYiQ8Uq0EuDYMz3GDKyEFu+jFDZ78vyPXZ34Ym3g81mSOxt
5SdIaBObAWqAHjv218vULy1sXsawNGKvSAQGd1X/I662DC5icWoOd7WDdom1KreAzOdk62LLCVv4
sixs5YfI/J+7aeBp3x7Wsm6Xg+I+B4uVTFcvQztARpjAGPCnhlVqoW5vJTZN57y/8CdHs5ifq4VD
/HhJSGtT4szPdXtVa9A4PEaHibJP3fDEsNL+PPnMK/TDu5M/Bb0YT0U8DABWrRg8O7hElTz1jpim
DyBTjLinWDI0TMHVvIXvffBqklsZ0OLwRNwgIADMMiouERZVgVsI/T6pRnQQsbtfm8KQI0rBv9FG
MA/AhuZaS0g8Z5Y3KyHZIi/zv4Mz95WYcQH5q5qm+f2xDjIG9SUxxME+3Lri+A0BVAdFKjmMUfhj
qTbzsvY7Gm0Pdkyi1hADxnfXCWlmvvlo8wlNgVOheDT9x2Tsqq8llRzwRcUTREs9EjUlJ/OjU1dp
oI0TnB9yBRsj2p5DpYpiGRFEZ/hNsVWOmpJt1Uuo8/QUF5RhgWYnFWNPmeaBOI3YwQichItGKmlK
oH90u/GaLu7EigDSkW6uYfEgPjVUNvMvDRDGupsGTuluKfq1CKeDkj2z/BtfYawHrLqZQZIgzz2X
930q8gM/X+O+DujMzZjBmwCNj9RKo4fcrDRPWnQZ2/N/z5cO7SFRaUCNIVuexHyJV+H4rO4L5+iq
5PAqfFDdnsv1CUGABVPPqc+8eQa0Dzr5oxXPmJNNpwbMClIuKjWfa07PHaBONrSgjhQS4u4oq+db
jDihvjN29SGGCPVBRoHlJEm49gWx0xFr/IAuI8ruHZizgeoxz2KIgjk3E1uKqK7X1dMvJQzg0lzI
vpK8QvXg/uLzT+0Bp0cHu4W9zMSJx5J5peCM+WPGLzGslf9aQpzIvKAx11oCk9NLGuXi6aDDVh0r
+vkUMnhwTBL4UxnSuY2x5OaKtUAy02to/yi6k4OC5b0iggWBKJlnJ5SsRsyPJfehiZ6XVVJRs+eU
bq5bGGxMNqBJz07yJ4FmOiCAK3ZgLOmYSJ4IJF2hOTVX08aK4rA08SmfAAzhzc0gMgXihjBU9+8S
4rbIyx82gij1unKT18Cda9v9JZWNnwL15ILXk38D1/i+tPlfniOfYtPsCLTWqnz7ZpzMCmygnA5y
jZKJDMu1yvj37A1iwGcgQjmnnsR5SafCKLWzBdTCLf0YicgcKHA5+HxfErc2Hv2R/HMW7ausMnWO
tEgxrOk3l6wZ/8TKUTTlllxXNLjQiDJB7Z7WoQwmWNX0mRFwCPybvP1rRHAH4sy1mevDfm7PoCwX
Xxrcgu0abXA2Bh3oziEYjEszWAoir+wV/LPZzhFfFfC/vJTA0SzJfDGhm3s1SDdIx8dXOX4bfanQ
Tc3ovKSajjM+Hj13giDQld5T9s0LQT0ivRXT8MxABxj0QbW3zheGPrz8d+Um0/V6jFV4SLqmYHhS
C3FL9Oolu5mVBpz2MZmfUv0QDh9tQU6jxjHqESBGd9AX9ln8Nd/clzJEo3mTMHvW3jf8FRSkZuwg
NJt/Krr7oxDlgLCXbnXPMXTm6RZ/lHGsy7ZCblBqVTIJhxkt7ZIN3sMOOrpYBm7OdZeoGkazmlcU
nzmNwo2K1NE4VsPjqkIXzh/MhMZcxeFjtqrLb+bzdv03kPYsJWW1dpzvTuUz0RR0e4DlonttTVLL
JWghLGX9MBUONgz8KHin+WehPMXf08rMNt2thfuxwSkMBp0hoSC1B5djYTqFJ11Pgc9sIFo4q0Lo
yIb5Km288fGgX0kD+VTPlFaCG4Py4rQ1wKFfxkr1uuBapDe2i7L5J8TAjld32Nk5L45M5wx07cb5
ixSt//mIkDsANqLP9O9IhIbD7Oi7/feJNMOGr+02VkAyJbOBZtSOiIexgZ+ga9mZ8xLkrLEXFxYJ
yS3gS1qV3FVhmg+711dS5fNOhIdZIabWpczYJIvFm86QeCwY7Opr4jUthCYSIf/yk7KRb1NrSNdA
KrwVEKS7dqh1ubzh7T9cT+zD8rLdf1YD0wIc5IM0re/qBWl+rELnK6hECZQ0A2WPbnqzan5p0xsX
i75OGbjYp9N9iI23n23PMzCAItTquJ1DC9i7Udiuh32qYSZx8F3mpM1RtGyKGjvOTiSNZE6s74U2
M1rnAiTEdaGD3p7d7suCJ/UpWKX1bquNRXaYH+53JjMEQ7Pk58Z934HK0wOo5eQ0gTLVG6dy3EfD
ZbN0i3yRdE6Uld3ZkjvjSth7o85k6w0NiYdiy+X9/UIa3SBxcXqz97MRRAnui15kZx5/770Bta3P
MDiYssHRCl/E3Usgs8qGsGWOYasXFfBW7V8ZukY73ca3u+Hf0OpF1R6GqIREFs9Mhh/5Pzby0WPA
+xx9JJd5pO/iuZkb0EhlGkW+v9Lnb2J0HAogHWMlVwST6eTo3tycRjHY8zEmSPThS8OEKhKYcwXq
bMZbcnLw/ijahsrJUgWbOB/Ar1FgowCfgUh4ODg0BF58EI5Abao1Bth0Kb2ih3bLHNW0dGMC+XEj
gPo0ipN7UxT9vSTorc7JopEdXcm7A+DmbyTNH+L6sKUqCggMY/6FiSPbAHOvKvS0+Aya94BU5O7E
J96bcvEyoik4mTqt96YXCdAy3M3RJn5JmtCqZyUDd4gKXp61iOjZP7ljg+W4LQ2KVthK7rehnaQl
iZHXU7XGDl/MNiVQ2vNvTlHoY4zT2QqpkmC/Vr5hIbsLm7pS/ubcqbrVqyQChoFGKKtHinmhDZ8b
nT2zuVQX2tV9rPnwbTEP/sdkpJ95Jv46+L+tiY7mXEzBlKpo/4he4D7rDuuX5Lyn9MnQls4I9WXA
UtaVSb6gAO3NXVBTcY0Qa6Z0ijxohLi9ydL8YmV46r0VmFeIjfPsQP7djYlU4sd1+nKHvCjhg5e8
NwlETONNF8dFM53E+qxU+9K77OUKfFEnanB6AXhGVSDj3QqptTmICfOvySh5bFjk3U1DWUEW7o5X
089G4fIbg2N9irX+Z+eqYujMyrLDO/y+LZwR6EercziqvF4TRAG/fB++PeZcH2rzH/YweO4ExSoG
IjrxbGlTkgVqs8ZBG/xiD5cRjXNF3u6ktvI4+OFVfIWtSquz5Q2Imc1cOp9SO+1EmXic4VCf1neS
5HfdtlfxYFoSMnyouDNxq9Ao03nBQBThkaBjZFIeFL1y24Z7RHb8LSz5sSh4FJtD6rTa+sI9Y9jl
/VlzDjtuVsBYy4H19fk0Ou9gPpO4FWxDJkOQUIuoL6SnENWMLxaUvrEoI9TUR4Uv3OwAg43u+qmR
ERHOA/J60icCrd+ZlOqFFSjGCrc5jMRomWPAgeb09vHGISSQxcySQNBDytMQNoZvvW5M/BS94oDd
WVqZM8AhEW4kXeqv8xgZQlX+T3+gjtbpcqwMviW8LY06Kv9+v4T2CK5Z5kNev1qhaS1Mm/wNTGBq
+UK7tYwmrOQZrYYOqjWE/E6HhbPvadwNv7DAxgNPARLnWdGnF1fBUewxb571l8U54SpUIeRh8wMS
YAQbFvgNs85qwdRwLpBTTNhBsvcB6pnANfsEkt+K9ieY5yRwmeOL0QPq/eH/NSOqImfVOn4HM49o
9tbtjLutW3sLGkYRC1QVGQUnZm79qBTANnuqT11M6mn1tnRvVKU+x6wfwbsQHa5XNW6TfAl0SKgX
AsjsewPHPZY34MgEi5zK/pOatc4mxb13W4haGrgowVa/AuEtn2WVsUR9+gPm98y+SaKNMLh4kW8t
hkzpJE2g4zB+BV1u619VNMr3Bd8x/M7u/9pmtSRSri4ZpfJLT51MxWxKJOwXimZNauFMQ8g+swvG
1puMmdthdInfUWJEejSGuUiferUtG7nuq9gxBGISytjVOx0yfbRn45ud/WNpXzk72B5CPpfb1sgS
kt4IrB6dD24cLfit7GssF/DVLp3wmAJGdVFxUpxuQRA2oQqfU84mcZZOVNWNWUNZ1eNOC8KyCY0J
A8OIQL5ppZ/fsNI4UchnQ44lrZZVqF9ueW6sTJXu9Eq2FTUfCoGZH1cE6jO7soNngk4GuyOlL1OR
Z5yevzcolSyQ6ztQ6h42Z/sJWiv+fUOYJIvWbUF0LyyQRPYYLM2sg+yLkosxDo+XPp3GUTqFC6NF
hF2oAEFbwvA/TXD6nokr+K3+v3hbeQkLKVpFpO6NxK4mqdCFxOtkoytMbGt2WJfOf19HUbjRFaBd
D8+bIHPpcwmKV6ycZzBC2MM52IOKL0hpDKcMAd0y65sfOdbIKKipJKZh3qGDGweYGcFBVcNWow9N
MOhg+cBBS6AIVIat46Qi6HRuVpd6cSRZmvu1vvS9Hi/Pn4Cp0zfcoEvJigmV/KS5jfHefzSUWLcQ
b5zjYRfXx6dyUXZAlUJQjz89vRy8Qd9+TD6NSut8e6NAYTwZ/IUo0RrZz/PCFykbtcMGyj+aLdaU
7sStD9+MgiHzv3GzXT8PdNnA3p4Ns5nzHcyU21BvSTCz21swLGXl5ta4iD4ivPmp/uH6nZP2Hs1k
aRCKzF234dwqIRRcwmBBcGFdvCQUyegY6gH6HRx8Q99u87R8EQt30E41M0a4u/F70pidQgnSeKHA
YXzTbUKia8VtKBmBElTbu5prk+ypuxl3XpI5WQvoM6f+6dcAL8fV+/e95MWJ0VakAX5ukSmzCg+X
3rWDReOhd+seSfIJrd7szCX1KIOXPzjhqS/lGRrxvGAs5s//czadC6m/d8S+w0R3uIQOymfQUC3+
zk2krGmDo+6wItXjhabkr87tUFuiKYV5tLS7klDug9AHnk8N0OTf86W/StQNwKqcF2o9cEvagzQd
eevUZDT+qVUKP8X9rMYY3KL1DNF5a9mY7C+f4uUBng/Zw1YienXMUy5dS4epoFt/ynCLhe/6Tf3D
ikLNNmnnhMPOdYmvEEuIMOwGlxJ0DWTWo3mGpYsYhJiF58s98THtmkCkxv75JTxVbG2POBY1CSot
hFtfmPln9o39hB7cnguiPFkI5kRrcuGK2i02b2ELEtAy8nrJDVWdHNpSZPHqq71lZhcRSl68cZYe
vCd8ZZXdgP4GrBe1w9AIaXitMhSRzNcKWJqJxDkgSua2fhSUHI+4zHWBhXgKnxThWDX4RE66VeWV
ooaewAeM+zQuDS16wpqN48b7r0GlSXeg09nt0yYHuWsV3DWS8+lBQxgqrazv+/Z/vkQbB2E/9HLm
yDh3hX9m4brR97M4RnRLKD9RjRMHXPLKURHumk/ireYnbELQ2BPsRM7pyCpBaiMyEum65wiOcrw4
a2VfnnPLPkgoFP8p4ZuWKBIsV5VfpK+S4/8qjkErT+us1M/FV1iowuU5YWem38rXnu/aKAZepDd9
HXg7hw0pKYXzlEPow57Z9p/YxR9KoYQg78yfGFj1YF5vBACY3Z3zAo29/ycX9a/s6pzvPxmxKlo3
q+2prbwVlhTzo7aEEad6vKJQKs+HpIdhWzvNZ3TRuGvONtit0o0yuHXKK2HEx0mZtfSn87kei2sh
0hripq18NJocOtua0pr74oM3ozH6/a36x7yHpRURzU5ZnW9rbYjSx07uOlQuoS5jBjc4EGc58Fji
sGSy6Wn4ss+TXKyTATwKgpQ3Rd8auHXJCkQ34YpPlZqF+micWCKug1Y1LBH+OorleSE0EgqkqgaW
e0oolnAfT3J5PW3oNPamnW8kRjsLuWe3IIhTetItWkgo9b4kTzKpah8wYFv0hZ+diQINXG7nup45
7nRumow09TmPaGibJH4dCul2jqvmsTdS4ePIeYuXss6cdUb2u9DxXhOoBN1XxESX5erAsE81Xdex
vEZcyEaQ1GQJGZsCCzkVcrMRKww9Y9mSMgEJnnFG5ZGDGAqAKF4TUJ6+GHT86DOQpVI28FscE4Aq
O8xTfvJfOs27W05QVZb7N8Ex9vUUzrtAwtNO8u1dmaBrPhEQOZCT1l0f29MKReKemBjLmwQv2+ts
LHcFFdjhKc2N6ssb3OtC3fWJF442p/wkkaH4TtxJa9PAnWZKGPKikajcIO+0kOzoyr4Ov7nwGjmP
ghqTnEwaHL8L0DpIj3WbUuRP/oMy0aVwcyvGAxGEmgE2HuNoTOtz43wOTP/2LLM84+q85bpdzhor
t4Te4g3QY1RQl9LvGQhzdpvxVPRtzoIRYt8clJ/FN8/dhATYSnsriE1z8cqIYt+PdY3nNUSx3Dzr
8gMnzE2Cvx5pybBViQmrFmtliBHDDZAiPOdScLbQmTGaWMaBQ8+sij6tRztugGL+ONuR4BYYLec1
g84LXzP84rRYatNK9HQ/ZhvJABcB4LIbcdeFnckNIx1avR9ULDYPnjIh7W5CiRcra/yanPtXomZH
7VY3a13xqtOErFUJMOh3l0LhsXyOR7bp0s2tJ7lmq5aYLI2KkCXBsFRTiqlKXdy6We9ADKMEszRT
FBiJKSdzLIvq3uTvc5i9Xv9mtxRbzVqyDSAlOqBZdo0F3JlPTc+yk0bvyFYmjNI79JHapARoAubw
YKVdho44QAYQDFValzcebSIESr8XdyfAEaPE9dIthzQyj+ODqd+QkxGoh5eRDR0qSP+BVIQXaI25
11lzt3X2M+KUiuXvhklnxbZSGfbrdlK0jtOz9GSWzK4QHavWrFiBNoac1ly/6TKUIGLRso4UtYzg
QBvyM8tGETzFKXo4CKhSaeCnEROPkuWEL/Xobu/XtL2GXieoIGDym3DbaxxbZFuyPfADiVhW1J+o
70W1b5unj0HXVvHcMuFYrLTgU1cq0gS24B5QAqEL5nCcAm+lewaZ7PCm5hvmpXS3APTJmb+gaiIG
AlP983doccny/rvFJal8KVrUPqynVbwnymqta1DtOjommJQp0QnHuxWGgD0w2UNtzFYVgAWhHC3i
A/FphrrVmkOuq+rpKPUT3wo7A0JcYNoGMEwZ2oZc7FExVQ8UFUu1cox+AR1G5ovkUY8sAbfNfs6N
459oVqZUv6eqxKWmvKemY0s+K0US+CLj5MdFFO7lZQlslySe0S8oAZPiBjit1f9R3QsAmAVIffm6
GN8dwJ5YJgTQtMMm6rpPrw8Nl1cw5WZOspiDH+BOdCURQ0pM3r1wau8MMBk+Wrqwdzf0mwSQLwGq
bkq25fYFR2i0vS/gD4Xnrwjpb3JGSivlR2DI6v9ojxKnEV4lYVEXqWn2grSnSjkfvE4+/X5yaOHZ
6xEoHaFUkPfD/ifadCF16KC4WX99h+EfoyDZvuXny/dKMGyPAbVzu2N/qQC6NqkWCMcqD8O7WuQF
2/zc+8JNt7W3TAE8arZd3sm5RvjwvmcfKr1dvwfTuuvJyo8/hflCh0+oXEKnoiclAcvXfcwgLzX1
9OG+sTm4RmE8f5HhcpNKr18lkSsQiSImPZ16fui4L2ddiY3pCtpaoV0q4EZDiX/lIax9D+MM54vh
Zmks5ULgWNv5NRKb+i/ZWsfNT2V1hvt4TPmcDgmW8hE4Y2/OEaEIeiEtbZjKuQVlG2An3iCNdjeT
EmL+yozztC/hT36D48SYHIjpATUvmRYA7GQJc6P5fkeVYqKUnA8NaLa27C3v/DmtRia9U+ktSro8
CkdltVfYzhaaAN6PV1AKXZ7vnUAy6+6SxqT0K65gVwIAQD7h2kD5CqNRfM+/wcEqBTQm2jHFIeNd
ZE4QFG13quYeTKyIuxWCD85Pokph/8wtohkPTdOjpJwqkSJz97OezzlqGJeFD3t3Lb4P455HsjA+
HFWfWMLPA97siRRmQ1QtUUtFim3E7MKnXN8NLM0LQ8PbdhJGCAdDeFvzkj4x1JEIl/BWGmIakbBR
sJr0VYp34HuUZJshHRTpAolDTiG7ZMvE6efC3gSDUqESci65FayhSYpLaZLI9tdHd5THC2gd0DYJ
l3ZMYNZeuvlZ/W0tAryeBkJGExqPqPkE8RF8nPGv3BRRUo675LiyWNns/XUS6C34owPxumMtROAl
weLDv4dZ9q45AR71XDSG8wOe1h0qgdYJN6dEJwWB/4na36uUlAAY7czQtu0LBHkWWNb1qQQM3Ku5
KBZYZXctD1eNTHhRlzW533XbrE0SAwakJZPViYytveIu443vcohMfO9IB1OTe5723sMLYNo+eiZD
67G5nWra6N741TIoaE+wiLXXg6WWnWcBStJwe2zuQhXqBPTYH/f5iFl/a+zrPg/T0BWDQgzjjvmT
/L5AaEFGILu4C7Fy8rzPILpZQ8qw5KXvU9fgqFo98/MMXyuPSenOEnbRiBE55Mz1vGRwBu9Yj1QP
OD7of5Qv/rImCY6JaYcPspJNlyVbzYnZs9pFtPuYjwZU+xPuE0nQg/qmivb6m++iSm30BAf0Bg40
zcO0/vFpzi0JJ2kurdAKkK21iQXlbB7/+qV1JNv5h51D9AqSje8xHQyXEjjQH0/cLTaVsuEmO3XG
D5+TU/mYi/r8jKqjV8fzmngxewPkQjJOH0BTdh5InFolaVOp7hLDPtlXjDCX1tTr9X2PTxU/xxTU
PDS7V0OXdE7+Q3xVUvcQQfSTPiggeupjJ1vBz0zBl2w66WCtRaIlB04vltvmt3rEtwf9CmEiE1lC
jFntduU3YTU/HOQhIDUi5G/c9h2V/xLI+UjLEQXG7uoWwf2uWXCEcWoCmayqv5qL0nflLBAbAQwW
8N7MAXjoBROPFAPdT8CcqGPNEz+gYAPwj4O/MRcTvQnWmL+Dd4xV+UFFmVMArY8FkOU7yqyFJqVP
AgLwDqfyCbCHzqkB5xwZSR29zXEqjH2k++3cPSfl0Fgw5xBEoMDtVYqtHTh9t97Wtl94dIX50PzD
Rh1bFI5BeU/hECHt9HxZoGbrK/wG1tG3kuGiWoYd5t0eOopGkgSA44nnT7EjRE0Z/fxuB1Wsd8xW
nZ7eRY/aSGvLKma9ZTYU2U0MKEnOjkIb/DhFQEeIr/+CEby1fYhP7GzLDj74HSS5IenUGWNid6U/
067FtpDppxPA86HRUhHZgEa40jVuB896cCG2+XHX8YmBcKthlBFJvQP30PN6Ldl0iaMI+9HXC3D+
4qNNYLDH/WMwZFGSB3ZxdElgs6J9iB0T42QE2iz9JQx8I3BcbJCYZ/1V3i5jnFFcYxNqqilQ7dKn
dNXbeFGZDnMmoG8GjBbQngXfflt9cYT2bQHrLuS2XajTmu9a8CwgpV5dX5ooGEBzwis61gaMCCZX
/U2cjf0dP5tKOfuYWyfkSXX1yareYhILHx8xVupQkpF9jggQZRJBlQZpIE75b7hL2NXhBTnAdiSm
AUuDhV85Gci8O4JJ4nppniLsNOID3jqhzT7jKqgtL0ORk+GJV1uLK34TMtSeMi3yxg4vRmaUiJ0s
Bitk53MO298UftgFI/CP+K6tdMQMsI5OKl/IEFk8ks6XkIEOdiKjdE0LAHBmsebV6ktj+Y8zjWg+
sxckFoniAEI1Sg/+OcXOElhgL/aDmIz1hquvQd8nkQtM1m1ahpzLGrtlrk8yUn3184C9NIvz8uL1
wzB+/Qd8Y+Ki0HgcYPSydYNatei4Lzs47i2iQ8gNPoshRXYjeNbcIV4QiPKSNhHC7oCL9m+FcQ24
TjY0V3HoJsc7zhX1zA5qFs/hYHtiZPVou2DJlO7dOVNV0xEsQxa6hA5eeg9ValxwsKvxh7eYDyMj
dui5xlwOte1bdDR07/wcBysX3R2c1jXMlGuE5qp9xDeL7qxIyqg/7TCJ3d5OrcpCvj45F9faWn+Z
LbQ0ZKMOLmA1mM3Bm6trVjghakKoMAATeYB0Zyy5iQ/TbJ71Qw339v5v4SuyucTL0ffYl6Ha5uiK
U6IDKuQsd2A1/neB1Zs26FbgaKLzn5R50gqX9jazVqOHOC7TUbkr4wbIM6dUFK1qJpb9EqDbwQx+
u4q2486KXgUDa9imPK6GAU/8fKR7wDhjxarD/5eBbJIJEt60ExjjKaYPIT2odSuxKTrHGsQxNGCQ
gzXW/1C2Cpt/CLusp+qkPbLRsYm/+jlaAMHTuD5TlhqadCPOVFVckqJ3PfV7VP9yAJ5FrzCjXQQH
eD0SnNZ4ADBL3Hcj80uHJ8oWow4G3k+q3gLi9EjMCo/OVXWY/R7nNSe5EGKYYH3ejh9jUl1IHMUl
hG9/6dDnp7eYPVhqAuBe59AKaxOx/HqXIzTz7x/HxSiM37pyfza4U+xM3ukyL+rfUqIVGaVJvmgd
+T3Hf74G6ZHrkway0dkFNwA6PmXub1B78gpDcsN4W0QQ+cVavUWc93qQulIDdV8KsuePNqRhBgNu
q78CC9qCvAKSh0WhZ6bhggfVFmk/NM1xuFFVm0LM9kCtcz7agfN4qMJ9RKBy3NLI1S+FAjnD8izv
tfqbr2C/zniMDCqyE1S+sUTLlV6iJjVcMqXe2mtJd8SP+vMu3I1+VUrAcPtbqipwGwvZS5a2M7MK
dA6aK0VpKyMRCVIA5Tte16EcHJR7h155ZvbH6RqKxzoSQjiyegj4FX18ZP4Dt6j7tu/UxyCzOocI
N+lSfSA4K2d9DgCY68OokXGkaSwiNrDJDbPfvl5pdUYrr39A523cxRaPqMf3wK0JFm1WeJ7zLmbs
aYELEgs5yYNbq0qWj7Uq7E7wOY2/yJ4Q6NNQyOVGUSFxli7n2b4+rwZCCv5d+kwduX51AHCmszmN
nhrSIaw8YfwT1/eusXdB5O9BLeyM480RWNrClapJsaprA4NlqxMcRhiBwuLj0BQibkzxKifEriNx
t7zbYxF+VoHlPChKXef01HUPQ9kyhUw4Ix3CWP72CAAhKBk9gRTfWEB53mSY5C2HvmdRQa83vtpM
9XB9elg1N+6E6U/QIlkaR5mPcsc/kHtrMwxev8zcwQMd83uwx+Nq/RqNSgdou/MpHdFBn9laluOc
SdKqpjQ/Lcyzo0HXBSHiZC/xco0VW16ZhLp5pA0OYqKhjEJqjoATvfelyyNUrtRVuJgJ1hKmYguz
VkD7NOHgQynxKQ0XL3/a3flq8AgvOIVUGMk30keNWqGpZJuT3+gdvvnP4xgJvrzMcVw+ZeV4s0jQ
rQElgMgcSWuOaKVvPmBvxFkPsvdGQIVMr8S8+3eYnAlBXx0VAvvRSS4di7VdYBT9ZUfzZnIEM4uV
GG+D3RD/9rzeN9PyQGgzQRwffPYMZtc5oMOGlsqqpqYBR/1WWRUWvjs1LttXrxrgWw1UJxZGTS9g
0R9ZYSsLSnPl6/ZBZ77FISj5rnvOioNXyjaLIfRvyzSRveJeV10uVMY7AI3RIBQ1J+eQiXmQ2NCr
AqRn7S2JYYeVrMvY9V9BXjZSWnZD69jVX9+7RQij7XiReNZzeBa1wVI+mLMkvxFWotg6IQvqqk7M
ryUDI97vdPZ1QCoQ4YwUd1N/zIhZitDa2f6BtQUP/Oaal9NBs85ib3EFyLKGGR78ettYGtSB2rXT
QI/XkrCuazwzxcqZR4JBfif+2V/+fXABZ2oEs+hzYeHkL4nBUd8Yyoq+8jaZ1vDKdUcGGZf7D99Y
Ch5D8Xy5laErso9OWNzXJ1vc3YDyJz13jNrXKBF5Am+94dn+bZPSmCoFALNa0CjX6DeoE/FTnm2j
zpfwwQc/bIOB1i+RKcLCHO83BTyWjCKxbDYfWOISIUkBEHEi3MQU5F5SKP0ghK30Ng9gy8CGrr0f
a3GqKYPhtLz1MJ+CHu55KvSYSdkFh0xKoR0f0u5Wa3RwKFJ0xZprXo2d/vyixP731p2LzIMEZS/9
1rwo9PKHrE/dcxWLMGGvQIhJbDMxO7aev+Y87T4+2e+TjjrIZ+6uvUqWLhiDHyCAfKAvy0vV+7ku
CsFw830JGtIBaflPS5DIJPvYPR0nYaMAl1W6rMjfLTOuGr+UuOVa+DQTWLI5WufyLWMl/DvgEOIh
WDL7MY2RSEv+JiQ6vXPyQory0U7EI7yP1LWgh/AhChqqsY8t9CkTN8aO8UrbeIZkO/9CDGo49yqG
o60de07W+ZvWc48YE7PVEfFEfWypuDLml7NYca9lhbC+cduBh53E/r4ZTwJagZDXDAEFOAbmnLWZ
9pCZ3sTjSYixN2wZNyu0bWdH1qXYrsR+ARUe0xRNlLn8TOzHJZzPhgb4/KI2TsGTlybRjHqSgGCi
y4EEZZ9LDDVaroZroc7YTqCvIpnNfEhv+g8ukBREdHfj4AsThGxwtEk/rtQVcUbvlE95yrygfeJq
dW2PPlvGcjP+aIYv2PVZMd8abpOhv2miOKqt8QFVkBpUl2Jb49SC3XjLOpbe6hn/qRz18CpTV/4y
bIDGy2x0lWiDreAG9OoBLhIxZ7PMCoU33Fz/gav73UBY+Bou30ldQ+AGR69v2QRaAf4oJ0x4xzi+
N6L5fYCZzDuHRHxQFqWOadTyLOrzt+AUgy6rPhqbVXhNGlRPyZZnhXIZDt4+dHK8Li0fp28Ll0Su
X7soNcqtcFUVIUUCGwWn4kPUmhAqZYwh21Zzg9wRBrce3PfSno/I/A7AgC3R6o+b/lphHvXayhmC
2Lls5EA1Fmsire/cW1OUyAeds0uiAMdmtWPh30w41oAE2h+79RNeeAY5eTtZG8UDBfytvLf/1Z0h
RKuFInsBsjgpVBDTMxeaAAXlpGYUXax2BtoOEDz/yxD2NDIFXrf/m+G3rS9anBOqr08HPIEvTSNL
R+A+bNa28ukJdABIXUsGpTvrzgcg+I7tMJXFQxbXmaC7Yd9keZir7KtMXxSlKdW5kLii9KBU1/S+
2Kod554A+5P1QcFWuGx+qfx1nHcUrwfyJVmdFPP6d/uxGcE+ZIgNMe02Elb4ob1NAD75ISK0WmvF
CGwE4uUiGiVzVC6I6gXQp2BdqAiFuPwJzhlPMHX9CCnUS2qU2q7Uzg/Xsg8UtQSb5fC3xDpfwref
Q7IdSieie/LrddaPjZdrDVQfMy0iNkdyYMurD33URHitowZscEzVAc/+NQA6R4iR/yQKh4ot78Ju
BWGtkrUEkwwlminwnEBhck0Ld1eNJQxqoHSSdoPt24x1xGgnaz3zrTt6wHxDT+4pZwsglWXvqSvb
lVKsiPL7eOtwoAbeV6EUm5bLoBZwW9XO9b9bN/R4e/VkCxoDROz7E089axuo6c858frSuw/7IfPn
33ALoGKW4+ePfoGRSXlMTjgtY2g1Lljr8f8vfnrgpvat1JEPz9HvgUZ3XgtMDhVGnCSln68yVkFb
UFuZfFGvt8gDh4HVb1wuwzPnFONpvW8xAFVzqaAFJUws9BaUNL+ABsB9CamX8yKaS66VpyWG2v2z
7RKMY52LeGyiLiVh3VU1wOZitmJL2s2PL/PG+lGvzf2wST8tpT9EgwlaFGfj2twOGPy4cGwLVByh
lf/AHpVhrWFIXPZ5XdBenT6OIzENxa05+KPufNRYFzsjYv0iE6jocd6tSUr3RXOhGNJun5uxb1mR
VMLX4vLf+cPM5JFDYiABnfo8woL1YgdCKEAEFuk9LIRElj0Kp+qmXm85fTZyqs/1Nxq5w0s5uKmv
TA1bNuuUQA4IF2yy/r2VatYaQ7HUUoka5DZQNPZgNqa5yhowVTOg1hezONrBAMQ6VTifMhqWca1s
/he0xdRS18FnS7E4191E6U4PhQSaJaRCUHYB8P/gwkX6iNM3F5ql9zkWS5UTrRPRdaL3OzeCgQRp
IbNvnllczEYF0J5eFSVzbK6aQjvTtCeJMLV2h29dFXHIKdy2+9CjBgyXEo7N3kCBIEZRtnAS3RLD
WluMGDe/pTYy12+9dDUrAOTZoOX295OUYT4nj/TSYNq1+uRRNc2SjS8ZujznzCHJQcBaly7OFCGd
INtO72lyptA6Gy7Jxo36bS1NmKHevUMIjOECGmb8+TI+fOEWiZKYhSyt3hkFIVo7/7ohIfkH3U8B
Dpgtsm75niOJORwBK3i6AozEBgNbvbwaqrc1OUcQTgAI1eZcs+mqzn+sDBMYZy4aaWTJyUiYwTF9
EZIXjwc9b63fM0XzzN6SkZAzMH6A1A+QxGjf4Y6GsgAy8IQwVVh8djpjwW3OLickoGhL8lu7n62z
Bni5b2iwuOuNdzWWDnUczz1jxzeMJ/36bLhG4TtqEA25MPP4W5JrCtOfOErB9erbSfXMR3ce9V05
2kKsUvvynLM5PdR2LwLUCCH/pZb9XSXRNlKGz735r4IZtR+ALuqb4ffgI3B8IAeej3FOCUtxaZCT
VdUs0eaHlWfMZaojQGGVwcuHiNu6CCjh9hKFpepoF8wDSKy4j4ZjB2aaHoAL4Z4b2Hb5OHyNFs3J
5BJPu1wUuTftkESJ5xfVu9gtG5P3iFWlatXze1voxibNDhAnZYCeJ43uS8wZGcuYdlnyr7rsKTA8
UgWvFsdwEAG0jtrFtSrCs3KsLrJI/u5vALME7hupQlnd6xLs7TPoa0mv4LKktAmNqMbamNH2MgE8
rqBKdJGOR8HIZhuMB12brGDH/r/o5PqHK08ZRNDXULuvqu/562t6UOHOX81CbBbpLIHFP0e9P1rZ
GBzMcskC63GQCiKCIcuFfnwkY9Wdyxkt4fi8Z84TYKX1qKZNfaRAL5xtPBPbWtfU5wv4pq+MdiKw
0FTKyiqtkJE1PvyPSqcKReKJn/7TmgbHUeMYc/mmEKL7Gqz2vCqZvaqyfqIWTOqR2tnUiPoYCPjn
OXkIxJIh0ctUBUuImHsMx62ewwNhBjD2DM22SGy/TBqIO0AEjCH+hM7ZQqzrbSD/PJbVtfpu1o7W
psk4tut11l5K4GqLB6XvTka/tJnZwKwGiZ6oTGiikh0RiwZXIPUFNawnieFTOwup9x0nIHTC4JoZ
EMoPm/BNTDzZKCpDiF2uA+wMrfvl5l4OERP33rhcH77yJN6MfF2EYZPbOKRzv1zCzdwCKkIXgtLL
U7jgf8x7pReLnwZ0hP1Ca1dJgH5f8OIggCzvlUxrpFAr79St1+FAtOwT70OarV4/B8v7tF3OtL1T
gBPJBMFBL4AKLe1qW+TwYVzZf5DzEdELw66gKdY1SoiFxWPu0L2a6dVFjMBaZgHEJV91TI0fzaZl
w1GbxA9UBqn/42k9HRk4cXvkf38dUFyRm5QWXL8nV+AKJB886mSrBliydAbKM7W1bW1rzRYv3SLt
PUbUMhO6UwJMeN20c2m5VotqMjTXxYUBft5PklUEvnbqvE0FR9xnIf3oKmyGgD5MjIRf2EVGiwVq
pQl3PpSUXhfYJhwbcwNn3UxKR/8vmzyu6mHeQPxScK/54OBpbeLk5TzLUPR/XtwXsBXD9SmyVRAD
pGeiL00p35Pq2K192bJK7S7i4XVPikQz7NGFWASg0rgwGJKeV90cN6RKLbBntccco9NmHZbTn5h4
KQAt9B7EPbE3ah7d3oqEaqVXszZGML8h89FKCrS+fjFgv0ARFl/3o31IEsMM3H1usQQ6EycC73B0
UVAe4oN8pFYnECjtTHIm2TIP0uMK1p1rTM7Hyda8+ugIKb3hxZwsEL1ITeyHi13Lhy5qVirUJMvD
xE8nJ6qr/FbVFjZKgr5NLTWsAehDNVIJScdHF718Gm61Y3KqpV9Pe0tt/tk9dfHl3vPWNqwrwIDg
S1lv7mUUvhCgLUSVJnn36tEkX/dGoawmHqcbEfGZFazS+rfapx4uvhNNL+oxZhEbL8nCQKdpQHCM
WbuAlkjqYlNS0yqnZYFs/MnXxyuZBgkrlLHVJFRO7lyXBvb1l5QF53bm6retdhtq5C9/Sc+8kFWs
1jYQA+W/4i1MYQxt5ZbCzrkZ9j1uM/o4FaNTqV7Rf8OlIwV2cg2XzSpgiyQmCPSP/deZNbANJeMp
9oiXhZShYqa77tauEX0hoa/0ms4UKE8yUZ1SBsJSD7aATd4Qme7fCYhfUyFcN2Ml3+WhGBwNHccR
Sj/4P2kocZ2iv0Hw/mvRGkrmNiVJDooZzH+IxwIYXSWJs5NOPwncTOUq69LwmLdsF+jfi8GonbiC
zkJQ8y0s9ZeU+SgqCXCF0x/WU/p2qqaDGEOc7NUxmCYkPhSxnrnxSfpkr+b9o2laYRDD3BWnYsIs
isqtTqR6YXH+t3flz+F0Ru0KfefjveBi/evYdySWVLjx0XJQiIMnD4b5EiQ4K6sO5ea6SrY+76sc
P/vZCLpg+S9iy/LvOO67C3HgxRO0onxhAdJp2MTxtOFd0e+fiXE/St3tLAgZtnt64K8Cq0Ho+9LF
hCa91s5nbEKb4mUd/UUDpTtu1ZA96rnG8zKWgg0oTplTN01MmCrp3H2DZHFs7Gd0gPUA+E61zFsn
xBj/YLyfGNn+igJDu1RXTIo0SFZ+i9VAl8fNg7GnwvfA7fy/wcQ7obGnpI9pjXg5C0hCwtMOKe+/
+bZNanGPFWdOEhkjy6V6vDh3Sbkpuc6PjoMBueIPBf+Szq6ZttNcCIXNId4YQrxgiBtQcTZwbCKP
ecsKx8aTZqnmr7giXvSEOYgvGw84fvW0iGSgf4kYjj5H0w7RbCmnrl5WBrpVmxK9ndgtysWuPvrH
vAveMCKcbks5KZNp5jcnRxa8hqw5Pl5sI9WnOmB6FADBM8fTG+PPgEmsoRCAu9oxBjN/PiXh4a9L
HtfhTD3U4UYLxcb9YKi46wYohfRNT5r4fFV1qdX3Ua3NeFPVFcvKFPVwubKzWxRd38y46uWiB+Rj
Uj9J9K7VodwkP4L7CrA911n0sDdkF5Fsr/0B6iY3gAk6xQ5DgMYrWugo2IgtfO4ehJlUZCGb37hC
Zz/ifo1K2VfuAIwvOjYCY48n+73QC3SnFIj3AEPwNFqXgftVTWLzze8/qO38meQey+y6ZnoNYD+P
FGuIkwM/5rPQjvq0RKRYunMKfsdrI/2N7xXePRAyaDwHFOhLRIsIan6ilzu9icA/S9i6rZPoL72v
ALLXYtfR12XsjwSpLShWpkXVjSwAlzp8+wcuWAwNBZtXVjazhhl2/CwRNJNQSVdXmwl6AHOMU2uO
LDEFRdCZGb3L8B4PN1Gito8Fuklmxka4W18uv7oOFEXxJJ1EetxlW9HHro/yPC7savlKtOhOqZoa
8EBR+ZfrJd2mEyfgjNE+pDtqB7vPd9V3Nqqh+vMfbpKLNP102pvKB1wZBTYinEPLgl4VGc6MqzGy
khyO9B34Sm5cL1s/g+0s6UhxndzDXekVXG5K0/sztPSDaGR5HVUVhgOYVaPLZ4igrMnyH7asH5dp
7BaQYCloF3OteKENQwzw3lbccxK4XHXwMqpc7cvzvfytmKAo/2Zduzq67zGZ3idCxpdKNAwyThWZ
2KENY/fUTWaJGx7I3LTDU9/H4uF1Y35r+5ud3f9IVlV/78rCYWDmOGfmUW1NgcTXOl08D8OjWMDp
YnrrWuY2H3WBa2Kskv+Yd86iezDNTvL20znGNU8pijaCtai57Mam2OBhkejQrVbPCThVob0iVFRl
qvoNV7s5Eso1VxUEwfRjNiLpXIJ+tstu47ftRlH9wHIpoapud9DMZYt3Yws32VBzc7g8l/SuhL2g
A396TkeiiJovsjP2ynDGmSYXR1Ye1nQYk8t4P5ZLCdtXOvUfo3PKShQA+H/XiGQ2H+nbzAhmO28O
LeCiVJ6oS18LYMkEIZxFXYzARiOZ246JxZW3zl4z/yczBUvPPiEo2elMO04y4EzCAMUk4S55PPP3
Cm1ZEJiZfzdwOUhy6U+gyxFeILI/oG3hCCvWgqjqVRC84r34JrSaiKZ59Eq09u+fgl7d1Prys01v
wgWPtryGivrmsqyHyZB3ypl4kDusIfvmy48XeBjtNL2ODBChaIcNWiljSzvSgacJxROCuBImjiK8
kvvqo2i1bSBSveVokYV2etXkQ2ZQv6aa8Ij6mp7XKQNe0xyAEfK7D22kqyYTdHR+fqUJkk8w3VcE
9pnOHwG4aPOM5HAburjiABm956IJw1fmppQ5Wo4s8pt95lhUZQ8B9at4ZZcGsvG49LTe7tD4hoXd
Lv4fcwgKKigsTXH07t9luWiVNQ3PZklAXiBbTUnDtCSIqGeCr3QZH9vIKe0iuGbXeOL1uQX67u2U
VxkmrhhVB2iVhXmCG4gBSgdWrUSOyxhW2ymaVfrql/rZFDhygQ4vObMQ/Kpyi7zGkym7tFw0txl5
Pvf8mZ7rXUYrV7bcWu+RAvL2diyxsu7L/7G9Kj7orI/pxTYNAc2Xy42FgLn11ugYzPDT9U99u8Ly
P5dWRoOfZLZUftvM4uP7CSfD5SzX05ichY7I4giuSrS8nMp50qh03tWciIAyIJAc4LOx6leyA7kW
3/uOu6z6+CNytFf0YduQN78pz1QpzavilyKyxUj1zud/c2r1rHXlL8QsKmo7efvOm3ynF8eOgo/W
iby7JYpotC8iz7PIpZsDeLRi+zU9M6MqoyLm1N5UnKW7b/XQqfXvsoJA9+mdeCqWFk6Zcwb5xFzy
vAwcXr/YXXki5qCnsp496TrJrqR0+WRJlzrPDEw7qN2JKPlTBVVDa6o9S7zJVac/qfrT4+sqTQDV
0RBLmuc4LVQYU4HsUN7eEkzXu5wCpfvhIgRcKctTA1NehnXOgzziwEseVKHWMZQ0FogMNfgpO5WE
lnKfpR0gJHHfy9qvYZ+EAax9T+cjawSBYKegyWObeGp9PVDJlWPkZRGcjrIa9Z0NxBS93vHTl+4M
N5pfYhT0fWC2sAYCg2Bt8UD8n0eEAzxj1k1ubzGJ4CsRM3HMhXlpJOtKy4FxG7TByLxhUC66emgM
fqQgHEn7V0FSBsLqqpayWAwgGG9XPSZG4h7HucsaVjfVGMeOyqZ6YbMDVU8F5e51mSstEo+hHy3S
ePsUzX+Hs5uNhM7Zf7fWL/SkGbnPjOT8siPxAXeZ9EeIqHVpDD+BjGpz0uTs8wT5n3JEVSQjOMa6
oLHchHLp5pJ1EaUTEzo5AsG12g4wJox178l5RRDklneyLwf3wnyilohZPMpABJjcyroF9mZJWoTu
1zUhTNZlggPP3SpbvAPxU1PpcnlpFDXHec7IXmg+eX/Bhawp3f+KLiTXkVMWMf+I0OTWfu+zw5V8
HMxY+BAvR4DkEwJPs7BRBYyvjU4DHUx665ttWO12cybMCCs4gMgbGnaTTr7FlZo4qORrL3uEsoo7
Eg7DG/gCGThJ5ZZtNB5HZdLAk+qnb5MufSd3mTbTMMf+axugVjRoLQHZg2IdDlCXOevm71K89Nk2
aGpRj9xbEBsRELPl/X8gMvTWpCWnjiYu+4oCt0N+FAB4dBfY5P+ClVy+Ax+ju2p1wIB6EtnuBqNW
OV5+xMQ/OYT1IySc5NWb7cjFOYnzn1RPZH3m++58p7ILv3P34KG3f7NbQQObFA+/QosKMoW8+qXQ
S8AE9Xt+z4IvtJKzgjFASwBKtMAvRnhjbXl0TX39QUyZVyZxbWlpRmL1w4bg1Z8ox47AWaJOrn95
ag/5jgtxG++fdSmTG3vmgzcOhuZnaBGQwKhxtCK+31/fZeKqjOJNgMBftkZszaDyIcAr0kyVhRHh
5IVfMkM1WEdvH4Qt1/5O32leHSnIOE5kavx7ZO1lu/0R9RC+ObtNYptWeiP84vlphL9N82SUl55o
BMGCS3v6FwO7o6stF0YGgR/lBONGag585sT/LybTAc4GKhJFF8laZKj40wcAUO7uQM0/mnaYD+5u
4okTSDZ4zFJpFcYFmjW4fyg+3/JXiMET4iyPEtig2Lt8VJs79rs8P/hFcyfsICsTaDMRejMeLZEX
/p96mrR/y1GNz2s1yQtPMKh+oWtESDNc45RQzQxG6ukN/4d8w9U0ILTjELdjWg2j2AtkHn5V2yjb
fPBKA0SxkFk8E7DCTJMtbLU9CGx8msQADMCAbl4ePoqZixYUeM5yKYVImx51eCq5VMrT7KESmOO9
Ag24s7gDdSfTvbJ5YaqRc0VBF2b6WfAe841fNRxhM+AdxZ73Pv7al/LS8fivqXomlxLy5pqIy381
jK8c8GhC0w+5c+8FJpgTtPf16IPCu9PzklEimfgYMMxn0YK8fGjB5uBCh6gMuzsLz8A1G/isyebR
t36U88tS50JtqStxamhNNH4Gdp5qTwKHqRl1RazoFrWtsoE0DXYPBmfjhF5YLDpaYqwsWJ0mgLqn
q25HpSNPO9irmiBGoew8NjxkgeNh4uoonHSaTZ8tf3oA9ttviWS1KKbwJ/7L2Jwph/rSXMvrV/wi
oJCUclGVu4a1h/X4W2D6YTwx1K84IP5ZmKqhCm72rkdXnh7MCJ36Vqi8+bWVldm4y2jdOMpTjPT+
clRH+lSndxiR7xyxj3ltiB8uKhCPh2PT3EhnE5vikzIRqAL8cll+Pc0DkNJZkVmWJdjOjmO1Y/g7
HoYCQqwIqGkeXXELXTSzZ4L5ZnUx6889U+pniw6yEimUufT7EQRDahh/kdfSGaqkT5RH9vJgFXbY
tYUu6Z+156e3GELUZ2A1IVnVjYqVXML5rVQ7psgn8x0IwYFp5G5DgoGqEoKjsPj+6G8nrlEDzyCG
xb67GA4sWggPLK2EUAZCLBuwoZ1dk1yk2nK3D6IX4YQmK7Uo5ScL7zNYBBVFvtlJ+sDkQyrY5oZd
Oh0vF9GuKbepI26M4lQBqvU5eFuAWz4Etfzv1BiGiaMYeb0QX214UY03SMQA+UVlrsfD2l3F8IxT
Kz2TjVhQhCFY8K+3bAvTWSPwECiOVJVqAQf1P9IXAbFZuG4F3ISjHyQS3dg/ofZ7uZP/zHD9JR/v
bCVl9Bo3MrYSmAQlh6KlnejeMol77GwQHdUSdQMB55OMr7HziBPXRHm8YCerhOVExwPoW1PbYL6J
05F0BIfLpmjaa648Ej/H5stvflYyejLcqRIsYwqLai9Lh+it1S3TSmxeol3epLpmL5VJlDAmjg27
QCpFsu4HxbdUH73V3ioUvLxerxOMrIH/FJ3mnyBLf0rS9Mb85m969CJ4RUq+VZA6uoD9yKl8SaNm
F2LYCFdLelGax0a2C3D8Zaict9sQllc8A5xjCwcCGo8ZjP385kx4B/aPNC2oT+pnZhkDGIYEZNV9
fCu1m5rJpmLh5sR5gIgX8u6H+iiuw/oJKQJ3bE6tyEZWM7FtPz5zGXrJC70bcG/boNsLyrhEk7D7
GsDtVmOyKIzeVjh7PtfvJmdam008kI1varI6Yr7qAr4GScmASpNoIQkdHibjDDYfwDJJBrrtQ5Ez
nv1apjbGIbF13hqZlrAu/nOhVSnPBTyyK93cZi8f4cjScJWSXEF1pa7vGC9h/axABpNrD5uuqe36
gnXoW3jXZ1i3TJjE+45jJMu06o4/30xmfVUkUPHDx6/fLJ98SrAyxmIGg4f9P8tDlwj5dB4PGk4I
pkTwZGyRVgv0oXhwd5c+kqfRcb85RIl7DSbqDrYWRDN8bdCrW4mA2ScTyshak8eKAxsfy6H+QPJQ
Hk0fUGKu5Nz+RUS0YgCy/PjvXbN3ZzqCu6efDOldoyCxRFx9W+8BxfeAEGvYk3jgZEVl6e3vQ2FH
fWVQspJjgtBrZhTaOphngXMx0flzNFJCufXyvztWSSB2Li98+FbFXpFDdxtiNiTDq98RoWu47B+Z
+azSA/FdiLU6Y90lYev8pqUXWHtlz5FPA93X+XyTQcsfOB3HzfS7VSa9pzKQeFX0s75k2F+IBVf/
6UhG166K4EVbG++IMupUnf6sy+pfCWg0uWLmgilPFoQhrM6P49xxaqR5ZPCg04GuhN1WqOMfezuP
9DlnNTnGnr/AsktBhCjq2RnBQEzWyNGEv9GN4ijok35GWNhyYmCUQYhMXyi8mGHpc+wsfdQQNgmm
c7/0NCfndMKwd94dmGGCwEBtO5FPf7GByxMbTzynUiHzJ4DLteM+HPSwbQCwgjO/gorSLyVjzikl
BVU/UHVLtRmA3S4yVRNuZtZA7WTTpQTANMCPxXAacvTgSMJIne/ClJP1TSGbJWy+DNjOPqM/OA1O
5ohgf/CZfvQinX83QMe41ycabMg+Itt0Jw1jGn1E3itfdu99gWhVtJ0KrSPlRKSi70ywazy8I21Q
ze0CH4DiGppJBUqeOLPb6W347xaBhBTzt3g3i1BFgMWzvnfVqxBG1nnytj2l80WRfwctUmjez4k/
lREblcJWI6s1Y8DZauBlAg2y466CWRxBMXhZvNntNMu7AOT69ZaH2a4vDBcaK/qaT0vhqQyk7TJt
DPaVPE03NxdDhT1MkiRQM31UdYImixpMdasgBoAlWWwWDq631GCkrb2yI2GHBT9aBeC7L530kxMO
ZPmsvAoznH5YKs2xDNRNDmac1yiZJIns99Khq6kLrWdVas7qONnMX8yKgR3PffHsEUejYTGkBSdb
vv0YwMwokrh+sz16FWSRHA5fSzG3WhDcN31UI+evfPpsIsVtjoXclPXAmZ8stuNyOTpf+fPMEulv
ttZMLdprokpGTtbSJWdiR3eMhIHveOFu0nBUvlPyiZQPstPPSLOLPusvpOJvgdT29qI1KW+kRZzi
m9PFPRl8aO9o1UFD4YldJK9OK4Hr9pl2J3yRjNzWIp+SetUAD3yVN+Azu4Alz798QRzLi10Aj2tC
nK3yiHfAm3XIC7QXdMy9DnQ0DrANXJ6UrZW8ERxQoPgJHKb5IbJJM+TuRNkhfZ5HS4P3KxdYyqxI
IOxWGYNZmQOUZV+ARYwibowtv3lP1G2vFQ/hsOuVLhgIWcQH/5gsllqm5od/RItTHL/5RAj5avoi
OskJIpAL1IxyV8WFrMMaJ2XWX+WDoqge3mjJBkwypcDJBxDTYVhdT8ejRcQrt0nZyJKOm9WHmyO0
2G4VTU9XnkjNyN20U6DMcdt/nrcpZPn6Nr226H1Xw86FnnCcbcDuvnrlayZ+WIloLuTTy9oOC2R3
Tozea9ebDhDcY6UDMy/dsFZOLoVdRu1sioW0IxoXRPC5Jze5zRucdD4vyuFr0C2omaKxwKj2Yi/r
WxQAKVBKbBWSPkpL+CNJph7zaLdAnuP3DHqs84NyFuqLbu7Zu/+ePeHgKaxfslkR8SjDj49c1CGR
TN6lWnC7ZZtrcCRxCLRK8qZNeMjEc4sj5E/q4J6uQ6jlYnPj5ZeC3cdDRGTDGh8ehDrq03fC+Hv3
4cDD01Tl1fiQDqnez2RoaP6A/jO6hxjyUMXNCzwA6IvsZ4sBXpTPbFR0HHyWqvueusjuv9R4jMP3
/icMVvK7n9B26btvAygYBaiPi2j5x2aZJxlVL5psqOFfqifEPeNbwgaVwG23iQ5GuvO+L4ewDphT
uJHa6Ql2ikBX6LMGcGiYhDOgidl0PYMJ/wS/rHClcvFR3WHJRbAZS8cwLAihM3rIGala8Wdq1PAH
asjIHyXnt4TewtjSXoicU7m14sCnvZvP/tiLj5M2Q4L/7sPJPihZtP8TW1Qxpyw/upcWjMgpOkxH
jhy/VZNDls+LZSuwuc+7uhb3FiKfO4nYS6OmrJp2IjPy7x/wtTqKnFg1C70NBS2U/jOhUrRPmDSv
IY/6EG0BufEluKd25L0Dvl5ym4qPLbJ1RnAug2Q2xqpyrZVyTqoIY5i9+rOlBJ/VR6dnF662q5zo
fKATEt/uulrWMiP/BBZ97SsPuJyS29+0tr97Qvsptwrtn3VzdAAo9+jI2md9zju7GzINW1dde3ln
wELR3jXjeiR+gxLvd54C6Ga+Hmd424qv8qEfdSCKFt1VGsiXA7yAWs9qhOwFPM1ZWsz09NYm9yLL
ME2VkKfnOfv4IJGS3e1F8WkraMZTTaBP4rn7P/cMp5vj3rWpzQz2g+9DEOkxGnTzlvS8klE3tYN8
VAKXEj1erKdL0TcKC2SFvaDaeR7XMKuF6YOAxFGpYDs+tGZp3anNvMnnucyaPK11aPtM+029tZ1D
Px18MI4tH5Hl9xWVPzM75l8yWTKsKBndEpnD+onyNovanhA27xf5eOn2iM6oInsG0OjHsOpRySdb
0Mm7QdCz/cToIu2VKb8/VAHSypabzmi/VtObNCraUFrQMbPIBq1QzNoLjUyCj9n2rceGAb0D69Je
9SBehL2bVePc3y/c6KUmcgcPvbJpyY1VIN1uljax3KLUIhRGZ0Nwkb+8rZ2bH4Vbt2pJf5nAVleO
K06rvgmqUxM2EPvKBIQJcNyf5lI5UB4La/bwbboF7xS8219YjwK8IR7D9qL/kCn5gtfWwUo/lVag
8EzIQky9MRo7Qo2kXjypTcS2dYz5SOwa0E5p7XS9iolIDs58jlSHdc2MHmjp6KZQsAUvarTKj/yp
Mf66XNYPEyKM+1xChemq+IwAc9pobJV/cf3OWg5yhOESVfpVjCk/XsrHeLJVJ65iKQ6U1Q4HTYEc
YcBTGJe6pO9hbpYP8TJkfp+h3JrCdbG4wbfEV0EpHp0EJDt+q6ib9xwTpa2yUIRsUeO0z9b/FbVN
fiI8d+K5Yb/Y8wPwQ+ODAXutKP98dKiZtjBtFLvmordzjkCI06YrQkmc+WI5h2ebd8vV0ENnAVfw
IUXH5M70Rf8VKS0TEfpHhGUjcrpEkLhVhqKoD0zYvDi5gyVl+C7fOwycrGo5kqZN7unD1fNTAhms
HlU1vmboLlI4H7fMGYZiTDBFWr3NEAB6plqYEoC2lS5yffHGsan41nxs/P3FvO5WItBTElt+HrNA
YC5ju2tPb2svY+ffH9C4C2B+QRvjP7ixVnBRMcMr1tyBFxeeVkyr917C5BphcX9rCAFfLhwWEA3/
N3vR3Y8Vw3NEO6D/kEjE+xeewKofjZvicXWAbp5aVxnmqODRU/kH/hpi2rohFhJH+v89kCssSupx
7Rq5SgVZh8muao3A8A+k5GWyhOpZoVMnYrd77l3VIK3vRldrKXWMb/GaLQXMA+7VpaogkJCMh8TV
VIvVumTSpnnPJVRCDSx5YL+Z4J4yz9wE7qQ5DLl1dAUwYzNkiTy/AZ6dy/k0iZ3hq5f3HsWrjXPl
50g8uS7JVxXC06PSwMh0iE8WUvFZgXv9a1pMxl9VbKGyaCVkXqQpP8wBPx9R7mgEt4MKDOI6IU+y
2E7uJbPttyhpUfmSQIdBjXWgUt9j4u8zzrs6VXmXoQNJ5LUuo/sssFUqMjBFGjMPGq95FpageTtY
e8JiHiGfZBgazRmkgkhtiALsVFODuGNZ1mbKzbN4oRc2oOVHUAfJjYq0eQDrESSjUMFoOL1zHRSt
FwCj+WJ1MWDsYltc2crR9XcsshR+wOYcn/CzvoNp46ejtot6Ukv+hk9UjOAArZ23h4faJqt8ta/d
IOz7MJXwvZZBfmtN3nO/NP39ScH2U/SLtAL837MURZcxULYbU6UNaEsuFIXPugL+5GasTmlbUCuR
f4e1xiyq9nCQVzBMOmjF3+U8UczM8TfgXxtX65mEsY3T3NmPHghWexoTC7CYjhBiY7pDEQ77Kgft
gwh8tfJeRxMZYySNrODFFpJRrQCR2E+i4DkQOMq3SxAvXXu6+/UwvSi8Iy2XcamkU2S4mk09AS9n
3suj9T3by+GzvlLFvodL1e0JttkyNSKc7e02A9bXVo6rDa9nwWjVYOLY6UakyU9VdP0fr2QXeNNi
g6UJM/WTI/rbxuHONYA2BsR3vT4vnxucEmuvrx0QuBNRBYBZ/HhT/xu9aQ8iQoA36bd6JwoqZLbf
6RFCwfdGvB65IqTiIYD6K+Worzu1DSVdkWFQfSKKw2jyukZkfPfma+W8fMs+yEkjT/w1Ega9QsdJ
PPILa7TLEk34xPthMh8Ry7gxjB2aUi3JGej3cYZHjAfBsqoa0uAvsJNquCO/NHktJPIjq4pU1a1S
u5qqU0ZZYxbTT8n7LPb7GD6P72pkvPBiQhPQmwIoIAHhg/iyd1efw1yR+w3u+qQXh3k5X/BRnOEl
XXIdgGCQp74mE+bNxO6f3HuQMt1V+6Ilcyq08qWpAZ/ysYqhL5Y6lWcMghYkoK+8YAmlA8jSzHj8
uaFDDpemFnIIVq0L8HCzlBYF+4Qv8liJfvhc3Bp/SYMtnqai6HtnmDmGDwdsgXqz7Y/c4zw4lJ0U
vVYAw2GYPk44IhEHKolvTircxYksJmyVJP7RnTiHmgPtt3IJMMBFykllCNWFQDvhe/SsYeIgq0JS
+x5406L21xUKDRkwrAruHNQa039apf3YkMyU7qvb0PvZx/IayeP1pYzixHFy0YC1x3CdWkcvV48i
FJhAM6M2xWZJBoroFc+Ldnm7gIvayt001TyiJlM2hldQ/fNcxYY4+Lfm8rjwHBtkdrYaJrEafEvb
IhfMid9/jpAlJXUlufeFcKhtCxTiz+jsdkVF76F3RTirB0QhAsdf5+khui64xn/gnLjFT3r9tD9Q
6g34FLUpc5dj1GrnqC5Ms9ddiHghL2WhzlgaRiePOMOaTZulEWktN7F04u9ppLUeHZ3iZBM+V3tT
ZHf1maOMCxdGUAJHDKGtu9FBAKfFimbKIhrAvsRvbDBd4Y/d0cT4Q3iGPn4Hb6qeDnR7AuOSulG0
eITD0b8uRKllXu/i+o2PBolYLrUtjwwiemFKVcYKdU3DxycVE8AcWMjdat4s5ipRLBIgr0lblz1c
KUIeEDnZMsio+M3XWqB5HEXLI9mQ0eJf94Fid1bUjkpfdKi6TpuE9MwGJOEagxSXtJ1Lwsua0cqF
Bn7D3N+oCiBwuyBfrPM5PRtQfbAotvVn2ZfJiHCWhFYr+W551zRm96wPoX23qH/ZwVik+mhHcb2Y
XWrI4dPqEQsDcvc25m7QF6qyzJRx4yX3OHqBnNfZx0yITO7x/EtOO8WIXbE3jpif6Tcg1obeQpfU
85OiOHAXraUWxvmCUuAV/TwPuBC5batEPj83bMyKAZ8lQWZogYQyh5Ne42HZM37gMbiG7gmX6DyJ
tPyRXsjSKqPxiTaiCniXpBWZw10uQUfU+B8qYk6S86ybSxVByeTyhsck2ysYK485g7I1d2nKUmdl
ky8niAP2kyMulGmIOytPhIMs4nFpW1CFKoX7VAJOA9B4/DgKJ8WKtzerNPJ9ZQDRIPxNr/rVv9Ek
4USHDRVhMk3EVD3LFm/sbu12qbpXoDc+KuFOBW1GfjdBdyKEL0IxnQDKU/HIzQAgs4OtcJ0t+dh7
IGQVFHsMyYCJ0RLdda+hlkbcUDWtUQqCT7rnyHwmPBikrZDV8ZK3Crf2jIS/ppXYO+NXutErOLdk
IVQyuSoSbJRMYbxZuOJoEn6IdfUk++pqfqo5NZLEzg7BWiMM5qSj9akZkP+05Wd1Kt0wDsVpiC1m
of45nhL9MXihWzLFlBSP3EvjF4/uwJh7CGGeUCMnP18M/nsCdRip3UujFG941AIZDGZPWcdSGBkc
y0d0/lI+edTQTO47DQEFZZgnRO9Xnn4+i9GiOX0cjioFBxdL4xuU/5PtycREQdt6oNQ5uKlZu9lw
HKZYwM+b2VbOIb+qDUcHTeq4XyLj66dgzOy7wSf6RaPOomdcaQOEam+/3XVkvXvbo3LOAqFCkzGu
Pp8f80gbahxwm8rCh+unGLvGAGlxjiVtceHLVvTbl4ucWsvTy+jYQl3LBdWNbG6dXZ9SzdpIvfRF
CNe+EAjUJlByYTyoJuX7EFMbGtNAkNGLffPT/JHs5cDr0XR/pcgR4+5HA08mJ7aI3XrzOuQQLqjX
oazuwsYOIxHtyvyz1KsQaS0sZtRWM5fVHG1RjKBWfDI0SXY7GkFRriWlE0/EQ8gKD4T/FNCc1ixU
5QBdeh4XtjgnDM7bexRJPEtuPC8fWLFO3aqlhdvOb5imrKEtBajb7foyk0OTfmLftk8We/zv32o2
iSSQzqpqdFiw1Q1bumd+wfQpUeeVdvE6TH3UbU4DO6dOmVLrA3MVpDSuov+5BzmwM9g0RaoHljYY
XJOtEVFL7NvJMwSBPWBns/ALFr2gOGjhjdXrvVE3CUpfDYBogeGc2Mo4PT4PtxYhMTi01ndYCp8t
xyLx0OeI5rMs05YyEW4icMVD0qPvyZUqBvmsuuc3HrBscqsxFqn6q3VtKkIdRJ9Q1gvuC2b6JRwD
5csSkrLVXiCuNsTQ0u4Y/jDtrTP7UVoSpm6rl9rdIhvkxdNXggD0/+L1guIepXDeTcUHt0z52WFk
2eDbHBSJe/ZGYv8ESXdKKZhN0vTCa1wFu+n8tSmMiolwP6qrm2fjFOWseuidU+DZYWLWDlr+O/FK
Up78oHeDF/KAVkR5SYAvxyT1lo+7N5Gi8Xj95h0wMHJLmxTLvGVMQkhITPKuRe1OiYq/Dq8HVQmZ
t7oKPIYH42i+0R49UyN9PrLrDn0nLhaVUh/DEAMlHasjL+IU1waRhgiNJdo5HVu+whz6QBW8d+F1
Wbx5zfXNADnwUdmM9uCNkV9XDHmotS7vRKaS1KhIeW7qRy8IW4cpaR1CVHp4TtcHAKFhzQ04RAFL
e+/QFojaySubM9OCqbcKx/F+hz1Um16V/Pw9UPIk49D8ZspGVUT3KmDkasWqCh3EfWPKqwxvJHa9
mz11W8hutm06GK/9VNzvnPobTuQ29wElKb1ysbpngfRRbHJ1Mj8ziMzpmf2crUDBV12U29jQAQ5p
TGK8eHDzo4tDC/6xxzdEpUWnpSFA7Eu9nyPSO3Zea9tPhPJfdWo+GwCDmqG9gL/n23pMEAZJQ0nf
kUzLWkKRWW5TFD0LAXT09nzRZwirdHkJj/8WFHbrJTdcT8yuL1BxRtMVipMcBRV/hBIgbvJH/K02
XGzXRhVB4IkKcWoWXnAY7W3GmyswfZ0mzqfSUUrkC1XJFuWpxiM1GE1b/m4EiVdOJbweUoj/b0kN
YTlWyY8SzrV9xf8YDPr17PjVPrYaZQ40EO/yJo1OpFYA4uEgthI77OyySu7V0nHX3lEnX60t9Q0h
SgOvNy/c1eknVxna7WaQKYCPBz6uGhwDGP0Xvo9EuC+bWiEbdnHI5/khwKn+pqNdYY85KpbL1eVF
lW3tf5wCyoph/Q0670gNWSrAp2HrX+YLHGIdoRlddoTomQuimOD3yCvPk1ciynVAMkHKdmhCEvY2
snI0y/1Yrr1FRIZzqkz8fvJpRLHzNcgkgTqPq2FWQM/Y1RR9jzkHmpqayJmi85qErUJmoyjW77zI
ieVNnVCzFMSjm0XeRdRsLGd1A0aezOMujuw+72bfLFVJo32GQwkrgEm7aUInOajbW+3dkw0cPUOB
m83Mwl+tPUqpxz1pmoB+xwfIAUfdrLQd7Oob20ead83dAvedItsMpiAlyVVJFSa8uhwBjC7B7N87
H5YsfoUjQzu8GGW/YRtMvGvy9DekkcS1lOhE8AKfQFQ3Q3PEKWzad8+GgvluGx3+WtF4hetwTEko
sM0b2dEWZyPpkyaBrA3neUOJVcc64IngyBwGIHKdmFZ4DvVbcg9ZRoEj9LHpOyhUd1EUw1ZNgwYb
MvRRrAN4Jsp+uT0GQPkJ3XYRN9u26d+aeF+8niEVXrkEWu4zQgODtZ2uPFc1buTPZC+s4m4Nq3Cv
4SRqGYqXLgYPINH6nnFW2B9MieJt0Z4RWIeyOdKEHORgTYNijwSnX3zok+HmTjoTUq4PdmRP1Sel
2JQ3akdyZyQNFXTRgiot39b0FXISdfQLXLHzTz5SCknlJMeOhh7yUM8bTU7tHm1qhNrRl+QPVPyi
yJJvvcFjsQeCFCQky5jcZcZMyWytbb62PnNTvMFGps5DPKwtVJhqh8kv4X3GUFf2IM6j8GmA172r
NF1gZkFvqdf3zdLECC074CoiEkivE3yZXaMgkAqopBGB2727MeL8n/iNSwRE2D/Y7zG0mr1Khvt+
2EFfcW7G3SP4nzX6UDgBxoFlkH2icm/AX2Xjns2Mzbd4UAnNG6useeqc77Bh9BVY7DNcCSUONjsX
svvehw/83EDo6Kyk76M1aS12iXuYxHmX4pp5ZE+Dv3Wd0KNzXwJ5VpPZ5R82V1bO52KNGNoct2Oc
4qE+erZLjm6ckZNY1j4NSOT8wbjaE9bNVR27A3QR+z7J6HgQEtAhaMyIaEVHN11czW6LVvARmfVH
zP/IzZnfXBPHx3SN85NK8pEffSUxOUhilxgJcwzbpr2BTE5WZFBJqTZzto/WQSwmHVxX3OhNtCIX
vuJ+dYhr5QU52XM+CxNY6GEPKZu1HsKc90r5pp16upmkekPI6nG6bAQr3aDekMQWROfevPPUEJqb
1K/T861MaDuY9qnL76Ubktgvt62bldl8vs7J8gD5xXGYj5R4c0NcqPxAvImyMz7scMSBYGv0Glib
O2sg5dyTMV2kmGo81yva5Myn/FOFutnpLh/ECY3ceuXbMCXOJ2+OQpxP2YiWSvaxaDr4eh/r6FR+
P/TfclDj9XEDSWZS0Nmu00yeimH+zs/Q5VsMHwiPhWqGkD7/GjlnW6W4nmnp0xp/WB6x5pJkF7Dq
xS+qF9HCHT1AoYMX3Iy5fZjJu2nxNnCKUW3cngzAaOvkdzbTIONrWkucm/ORz2pm1Aep0tliA7OL
p2H0Z92FonCWTJO+nbBK/WuXFZ/+L3Ah0qzjD8Q5f4+oY8M+w7SLN7A6ArkyomSz38YKzabo7icc
LnI3sEz0U7SF6zRgd1ZNtfGbwgyEkUFGGwhkqDddwm1DPezEwEL4h9rUk8UPfPnJY9XeU8GS9YC9
PYmrdZTTjIM0bW3i/XpBZTdmiecFDixsWVzwS3HGu5zPXJYDypFcerHGdHGjIF2NmZeAfsTM2FGj
R+4QrbACkVtKqF8PHYn1uvzGiU0fDWugULhsvNQFVYN7UetfQFQtte5akaJrMh8B4V/Lp/29CmOP
g+uOp9+wvOvrVHyl44vgXXH7Ww5vMV1VKfjQglNEi0MiFBm9PU7/q5+QKMUxdpW+n1EsL7LldEz9
4D7l4eD3S6eR70JoomrsHVq6TSTcM8u8NG7IXNilxLf0eY4msZUMmCNf3wjfB8Xc9ElkkInFTsYG
A8Q1WR91Rq4eFCsr3A+Q2w7/uw1y58iYo4cQs/3wl/EhU+tj4PUQqbmxu0ijUHF6p0LBbp2pdNtB
7l9MT3WPtVD6uN4fuMpB1R6+MFW6qoIwXIzt+QsHbtipTuhoAvX+dTFqkeNy3tq8xCAKZhrgHgkq
rEHayYpqc1crn4HGdHYH+V5A/xLpA4CDzk9zyO0W30sI77elMfYCL5V8ed+dqgvxc4uPDQF1uAgk
ShnYEh3nDBBMCimkc7vGiqaVyDc4euWbIUCDWVLpacbH0gVb1eAXuxh41vHz+ylfg0R0cbXrb8Aq
VcBA3h+1sU+qTfb7IX71YhTJcvMcoduLj5cHigcXsCT8hv5PPXuUa1QH8hPAIQoYsAmvXsG/UZsZ
FIltOmFG9v5tD7mX+/zd/U79xRfr4V98t3eyDO01HU83VIiMLJ8Oxcskz6aaJzRUuSQ/FN6YAKXJ
CAm+f4twgMOIc/U2Qe/GhV6SGDbkbDIesTruvfyAHiOqlw69vZ83BJzvAh2MqJqx60kRphEEN3Lk
3+0cUMEUFVoJHo4OzDBZzr84whBWg2SLp0URpmRj3/f+q/V6Mn27Z62ObD3tmnUbn46LFwqnUyZM
cGcNiu1XZ75DhP7jKQKzXwYEc4vWVR4s3Jy+UWxtKHosZmT60jd+hubsZu/kDIERn7ZUT2nAF9Yf
cabJJmxwHNpeMfw7Gl7ovLnOxohqQb18hdh6SKn5Ycq5v4VmYiiUoIUVZbn176gk4l6chq38NwdG
TXyO7wY/5D+kDI7jpbVIXKLGWsD5LRfBi3P56bieRG0pANLQSVwwxozyIX2JPx6iMs1MdY3IvE6o
TOBp8DgvIMdhgdg5EnsWyYs/B7NKMtqf9vcIpcE4HHIi8ZtI6THNbFJlCEeVQxqGo1elH4o+5qyX
PoA/YwSdC9ue+2GHHwC+KfvA56l+l5t4DpKLbQM31T8XgZAe2LoVP/BSrsQY23iVW7QxnXF9ZmAR
6Rp+s1Xst1qmYj6U0m+43q0rppNA5xyImfet8c6scgMTPhte8wg5dpxyUNnrXoiOel8UY1tJT8/u
hRRz7kUd94afM7ZiTyQbVWUlhwrQ6yxxVf9t+xqQNDZucBcw3+5WUWCfR+u0AIE3TsE12D6I0dqL
I2NPhWZumdQWEHJpawENGUpM2/9/aVBw+VtqB2lgI+iFipZKNKSyYglIcUzGWt7+/mYl2WX7KHeY
KmE7rT6oJ0iXhN9Rd8JOpuluuYj8XYSCZeVTn1pNmDK/VXQQub5i+3R4SU2Lekn5MoJ0BHR03TaR
qCWV+KTxlXGWxFNIRk+i6PeUUsfY5aSa1mDwykhKYD9F3gruyCjAhRXR7Zfs4E6U7z/sIMWkkSdR
yf5bJlfCIFvIQUlaVmekWGNMySIY0KZrQuYijHH1GEXfzawO06lAzp/z4GoxfbNlWrRExs7KjuDF
I0OtjVH1gdmce33/+grw/xOTqT3h9bW2zXFcoznhuy60sMZPJMSLOaEf3IBT3xpbHJ3EjlTRiIs8
rY4rz5AgnQ0eSRy5gK5XsjSnj+EtAQOB51ovouNzG8qKz7jC/LhfVrroFoZ3zQM3Cn2Y3U5QFDd/
KgFydEzIDwKb9gmFviO+/xKkD20A4h2C1WAlSMZytejsQE9uvEVpme62CkUzbKK+oAcowwQ5MVTC
J+rgGE2NmHZc2mJyzD9jfwbUMdl8EwcbAtNf0r8ytSxWqbyZ21RXfeZtPc6GYtKqJ507QjLTq3xD
oso5/K5uH6P2Vpde+wsC0wtiC/LWXB55BQmCdJ63B6uTqwIrMx3zaPsT6+ht+GhMY2zitt1dg8NW
0QBSQ1Wz/zSi9/dEZgFc6H31hxjHekfWf4VENGxHeFMgKb2h0/yFDTg+vAbk9GyTTtetX8jMh1Jx
FNRo7R04FPrkZ0rLgAeJtpvfGRLguFr9DweKy40CRqGQkVMYRzKIu1RHCJ+qLqKvRy/0dUJifuE8
6Z8dM/LVZySZ+92qqimZjIqOxj4L+AG9zniJMb1L0V/tr7opSb4zQrz/mc8BUIAYmGh6eOKCqOHt
C7H/Uo648KVmATjnJqDwtOxAxiFGKwgCpFMtvM9mXQ/zwtVTn+GYp14UARL/P5nzeJm7+gKQup2h
3vh95lC1YuS5igGbKlSeq+QU7RzhSS3hvNfaUOWd4rr7M4niKmwwb1eoEb00d6I/2+Xnk4mQKPjb
7M/UzGaIOUEsWNDXuhMgR1ZlmK1Yo2D76BPWQHFvAn0hAJWCQvVbsTs++Js+ZYB/6nVJbpOIazdV
nc/+lbnW4/uCZK/P+kv0edvVBPK8HyJ6K8D88gzK+7piCysijHmlC7y5Tl0fONs1QAMHkkYuTtRx
2Jqoi1UHyNhvepiefBZwrNWHet6Fn1YVnGWU2LV15Z8kEVp/n7YoLLhT0V0Xyxpix4UCBHoggX0h
JYsSZegUE6Zr+xvtQ28/ESRiW26gpabJNakTYcFtKW9S2wgPsQ5oJSoE33xN3QV30mSgmRsx1pcY
ZQzI5D220S8N1Shn/5dxgPW2MrHh5fVVhRdqIYQ/sdPfhzQiKZb2eo3OOECMyKYf4Wi8DkLCpG+c
HOQbgImSxx2GMjADKEl9X510TFNZhy/AMQVO8fkgO401GK6vpOf1NZkXv0ip+L1XpBfNr0a4T8JE
lTiv5voYdn7ismebnguXyzlAijJyidUqA5PvqxteCtweDWL4SPa7jI6FGI5X9SmOoCMn+JIBRTPA
EN8Mtmq76KqaXidpywxqEg9dwUvS/xASP8EsfLthtNej8FFelM8zEvfLx5rhY+hQUMji4OMYibZ0
tRo+/i7XOVFKQBAKdr2uWsy127gr/pd93c8fnczZp62S6XPPIToXyyZcEbKXhJxQFScpQJEE2W96
qxwU5XIYh3qDqUZQ5e9xBbWfAPT3YFDb66M4NUWg00NTCEFHv0u6EmxHt1IxOJXpr+HYkuOe2CBL
Mp3EL7D9uOWCkbEnjsLzSCjBytvP2iohUyRqC9HKHAwrkiffQyJXB4Nx3VKvRI6FJxtUU1+gQlUi
UCd6QPlfi2Rs9iUilvL4kUoM1LPwhvudkdLM2knD9c2KgExv8UfTx4/fRhaWEVsar+OiYZNDJ7r+
RQPtFvKMiwUUGStqXgeKT+Ehe/aNIsNA696zmZG5ZUaeQfBAToQI+56ozQZabue9yAsz21yp3VQG
StwckaabR43QnKGp/ZywiXhjZJ/RXx0qM41bEDgLhdSoqAykifTRwvM1ltbAbEq7ABUCLclepXAK
bt2sdjUszH9VsdfsQ7qgq18jIML3FOEfAiLLhIaf7SyCUV29Ig/de0c329kEl6px/jy/eh5Qvkn9
z/dXKDQCU9siSjaIEYM3hUGrqRCt7Et1Ii+Oo7/Ktj2u3hoLHnzFoDmVcImKKO+jDmMktgvM35i6
3sb1FjpG+zkcB3Ry0RrSaMlMpY0qzDTO/2wOSDRjYFAXsFuiXpMfcou9Cdi/+j4KZI0GiZ733lic
QJdvyXSt4u/7c5DB/XuwWnpJBo2TNrEyChkD9/dTiDW5VBtEy398f1e32+ipwPMrgUT8guwwWcGV
Pb0LrTog+jQuRReHZbf+a8/mCCnkDkqR1Xk3GIkRaQDucRGpSsfl7m3y9bE+1voKuOgfZF7A23+k
ZeI+2d7kzFCqqCN2eWeTnjf3EzCHnXUgbWI3CfRBSs0ryOtitWCYXI+mQ80sf6a1ftBEclbs2Msq
tR4ggrL7BYhamshS2ff7F2eO5u0K15sTdLeuvRUVk1XN1PbsR5XJzBJ6wav9pJ6kp0UhMcjfufaO
1PY9s40TIjkPR7oo4noYu4gUcVCcASCfj3u2WGBMbCR1sJydvHoG5Xg6teKBgDI68eD9pEJk8HLX
HfHYBWAZgF0j5JuxXNzTQz2IJIUmKSqLdeV0irOWgSpRNYh/2NYdEJbRTPTr7lunXTkkiBKGXWYc
/C6qj5jUQgpVSD566NSCt3kWLdNBqL7Bpw+wOUFRDkM17Mdk6nnokbgLYhouXFzXkQug9i76VsJX
rgV6ehswDAq06/LUIekTVHFXRpMsy/c16whFJJFdknWNC2LAnb3a0s8lgCb2aOyLN/fe7S29BJ9N
m/xaRVp0JE8rc3XLyxdWENY2gby7sG7HI60k3tzzE6/eMRJyg+AMil9wYGXIbQdfK0iOeg1/0S9t
Kbwxf/FY4u4k3itCUIBJdMvzMRP9O169kRcKswbMNVtDm2H6Q2iok+h0oY/Sw3ZhMQDDNBwR+b5B
Q9Hb0ndaTwIreXsD5TN2eRAPrZGwDEVg9O/uDDpFibrevjNdX5nLPKAf4TEb/OQG/p/9lXvBiklI
W6N+F2arfmMXP4D0qNTpxK6+CzEtqowrwwLTNqbNPBuYY3W8StYU9EF2yYUxUnj8x6VHKt27cWRq
3Ulg2OluNVT3jeVBHE6U/4phQpS1iglZrgNq6Y5Mp/q0pFI5nqzE9fcK01wTJRIluv9s8e5lnYiu
P5u1yiYMlqCDTQfJzDQjqxruWUcr5kNFVRw2u9bjcollYkwV687aFC08On71/PVu6vcxVrwKZrfn
Fdv/FfXRhN6/jLMTaKFPRpG3ydqTBG8ZgEeaBuf7I38tX0JwqYBFtDA21H0G7/G2+ADdaa/XWb0+
vM/ebCPWlhzi0KIDQ8zrQfMTwiuJOJH0Ul1F3kxp+9K/sX7FtgANbHPbMGTMAftQIFPURzDWQxlS
SMT57PXXUeyr79LIbKCw9LovuzexjHLIMM12FuO7C0pqdUSgg7vOmeKYW3ZQ7IpmUww3jyD7oe4a
uBvjy66vXUNP3xkJFEcxtc83Ui+BCJaCrcPo2I4GSADKGAcOokvnfxmYFRvd4knOFRpHCc5hgdJz
emqiJvBSTveXQ+iNqKNPSJH0+fOMnxBW9OYf9sDh2ANGI0InLCQLVP6uwQf7eWT1jDbUns0jBFiy
tDGOXLcQUhZoJ8TM+TEZE4C4++B1aFwCp1fH6hr9F97LLQPG9c4HD8YbQbtSnIuaI1YMi14uz5mt
r43plpNF4gJQeGKGCfNaoXac14EaxtsOoPMi1XSHODVi13y/pxzo5BZNzdzs4zDFLfOY7YgvlZIQ
dYYKw/NY5zYp7CKrFLmBAR2M0kCpdCvKASktzmXzBVkB+XlmSgOfcMvmN8liOGMSELNBzAYbAMgq
OESSUTwQhqjJwf5tJw48NvGTHncIOxzfcJe9Gc4XsL758mZVHetnxbyZD8eC9nYpA+6mXUudNtgN
inZTPw+BB/dnRg4veNZfe4WHtqcIoqgzLsUWcQ1OwJV+DYFQGMxzzL/e/x6uwFvuMguFYK+9QmnC
2s2ip5imnV3JU9kJp/9pWZRHiYsfbIzzrClWth69/vfW8UkblLDfAdsaNyh8QOfcpDyvgkuvbR+N
vXZ+Zif926SlwritUNzsx1/Qj72u+y8JPQa8Snpto98FyaGtoZTRiENYKD8YeNxM/QCl34462vod
FYVwOVRQDYti0cyLXswVG4GSI4ebu+gTBd08wxwQ9HzFyKqPY/I0d5vNG+9gEVpVQHEmQEgd3l3X
QEkyrkAcY3klZeZt0+HktEKAN/Gk8PsAM/7K2ndQtQEm5h6WukFMvN9w/d7DgCkW9411cjK7haJZ
gtHTSgTQojVhVKx7hjoIGet48T3ZsxLKgoy0QRZI9iDv5z2jKbm30wxV8z9o1YscauX4DnaOJBYM
Pyxl1tQShpH/w9sEyFv1C8B0M/yucmjR/OvAyN6DcuTriIwRJ8FuUCIbqj187o0ZQsDK8AnJUekJ
JbJd8BfAOgtyvSxHe7TJYuwOcVXiz8uXCEGgrJRsbjUN/Az6Jq9WG5PCHPfjt65rztHRXSCDEo49
hK01lbHfOGb4/rvoSfyXLvUt621EvY7XTJM/CzBqkpKuzEisj8pV5joXforWFoiFG/MuL3u9wCzL
vMkqvcQm0BZt0MvFHgBrdDoEr/v26dWyQktC84IHCVq2mUtdCSXPH1FwQyDd4YPa8syJSok/WF66
Rrk5KBLGm1wlfCCDLv2ZmraC9TWLhPWKwU7gIlYxdyC1LCihp10kr/rf0sh8VVBhEdCwW0a4XQJ9
YS5NzE7FZ9NZyIc2WAEjNUOtVzMDI5U9zoC02hOS7J+xWoFiEUphBL4naHX3ly6HIn0vkisKrco4
0ln3wmGJHc3k1CfIrdEb4KMquZmNqAJlZ0ErRjky6rxCE/j0R/vAAiy9dzWQijvXavgOyD97+1cY
czPoI3Vy9J22CBdi+xQxmbgVy8rM6yzpYeBpZKhnhpLccOic5UqOZGySW7NZgYl8YKKhfF3AvFuj
VxB1bHRTFh7V+r6Hb5FW75pBxDB0jPrnEPUvU1nJ/qwgxdf7rhe/79798DKy0RXBXwvYd1YXB5aO
7WwA9/Pv8fev8uSz79VQpFxmoC1bY/C1GbS9GCn2EbckQVrBSYMlRsl9CERvmj9cnk8lZi+y0ZCq
/oNEghYCf0H0XDE+90YPp3eaFE0ubni+h0F/GB7GXpvUBP/O9VRecO1TqGJtC4AUhB65W8QrWyP8
UY+IaRgx4yxz/He+qCfrPe4jXUg4aomcN+o1kkniT1kH6F9x1J7kKNMu9xYLjB1evngCdXxR4HvG
86oO8ItGCTG3rsG1bhZAcPSzzCi3jBBBRh9tfZzKw3nUVuBTuciGP7GENLjYjE1NBJsWrCf/evYc
reTWcgcNrzpzwXBXuIusSjwymsfnOm0WV6QTh+LQfckn1NqDs72KHSX8eXpzH2isUIhP6aB7kzdj
+ll92sxlgmmzR84meIwn0dobgDE9RVESIGfWWxrtxWF1+TYd3wNl8hrrsEUxN/qRxsx9DHu3z4Pz
bJyKszfRgvnQXPN1OJUKeOYn44iHwB40uxj+V05mdOXzMqeLjjoHwkwkxCPyPELlvPgaNWpN8GiN
83f96sP1QBxP7I1dsGpSD4HhSklFkMaUcOzRciORILNAzSsiM4jBh3hcb+61OL8zOM58mbSqwrgi
U5xFdT2+k5FAK44d2+tlme6q5LeEVCVIwa0D0ho5LqzdCLE+pvJ6/3NL3Zg0F5ue4bHBL0nQD8vQ
DScsYKALWE9bcH4ZDMukfdwXPyE8qYo4MEFtWVi1xjUY8WrhmKTuF5JlxBC5iCh20NN9dyujWF0x
Py9IAnpxPGDYC0CTmQGA/SycqbqJoULgPlbcJj2jwhbhL/ulBGpYil1BYt6C3DslM2P1mM0mw73j
1qXUFZyh6EcRCoG5jbeDQEzaV+w9np0applXkzKd1RAomkstme6W15O2yo7wsByZXXI/bGQO1tqY
ioshy8Wz9v5khhHguU0MGKGPJ3RplMQE76XXkFfU5S2Do80RO62bZIRVMyqyO5CqKqFDWw/aOf9C
yn1tN2UJRooVM7PBFgn3/RLykbRKotMtXcbdiM/KRuu/qKk6vhDSjcLwZH+HYCbAmjvxV8i+Dbmb
BjwDlZzJNjj2aHjQIzFxFtTx01wY4AeIDAg78K5pYZD5JkcHqHSJEh3bKSAxLe5BUp3HpeZvgyjb
pOWkkSZVBioFlpF5KNUGNfdDFnts8zZcHa5TN2hUv0ziN+AfEkRT0GSbcB80i03N3qUdUvtgDt/R
ChInyJhyre8WWy+HunSFXhmtirm7oK+c4UfvJq2f5OQLc8CWV03vEQfHn8OLAKOiDM+C6LUXWOz9
0wXzvnHKTp2GouRpv96ZrAAFsyLBfSpd6RtLxW4QL1u62UxQRs0rGAt7ABA43miKar2w7iml7vO4
KuzUCd3HNNOkIfq6kz+7dKiBZ2Pk0lp8rQ8yVr/2EHpTUuoFI4JRoTclbyYZ8dODBnqMpTNsAxoW
Rh4baf60KIwuZZDlyDjIt1XhyfkSFu7R3z8kkMgo5k/RDnr1EU7+YsT/16s2USiNzPEOfpjNcx7h
uXln7F0UrSwI+cxlLjFEXjw1cu0QQgVCqyPQ2/zZHlK7vtbjf5dLLmaxdU5kgEzajFRvC22BmL8z
ULknNTAw8bw5jOoPL+nnLsGihlx/Z4LtA3mhm/r/SI8Kv/zOaBgL3VxrsrPsh3AytUFp6xu11RQ4
TvTnX4R+fiDN7gWyQTsZUo53lToERWviSnD+AWcrcM4lDAeUdN67tucFIv3i6lc7KqfTqGRU6P9y
OtSaAr6rrMeIcpDSVXj20aER/A00eObK33fIt8tw9vtvs2SYavl9Sa8U9nTUnt8kdIIfp5K9E3Ts
S4lg+ySaZ69DdyUAtFzxrMd8260jMAwkjOP0WYIJMDBlItkzWMt4rdaklQny9dyLhm71oijKk+2F
U+kzZF+yXZA6rjRRj6CBXyqDAnzBNM82vAG4VRQh4RdaWWhH7wCD7sx7ZmmZGzdYZB2eutYx4omh
TbNmvXnV5tbbkzogvLt0ZiZ5EEGcwhckIK2drV4qRSXflgbXocj/1EtE7Zbf5PlGMVrniLALgmoL
5oonzzxArCqTkXAkVM46+LGjsXxgBZHSUquY0DRZ2yUrWIeXhE/V2IFmh2SmxMWZQUSbAyBQoM7F
vXr4EBe+mqPhy+HfFcyWzd6fJoCiBQbIMX5Xveg34SGdYuH+J7R71KcKXNG8v56t/RKGGYfehcmL
uB3kYC0zzQgsfuV46ujoXd+IPIvFygPTViD1cM6rkRCQ/s+TGNFBrMMrwCdyPRnPmZDxFY91ilfJ
A2oOvH7QJjDXoBdB3bs2BgD/aAddZ1Y7pdXzHIzuF3SI1uTyymzvmOubO6CfL0QCWFgB026wY76S
xuHirbemqjpSDz4NVU11r041r1bntezjy4+p7e0tWEWL856aaIIUe/vTpOHhSO8Rh7qNCVpsmEVX
l0lhwIAIDjmi9pZ9bx8ilYam3rubckPgsP1EI4un7HeUcGojsJ6PJdu+VA6yJLr+nw0i0GBscWP+
oE43Mgula43jTuTs0krFZ/JbLSLplRG7VDWUIhD6zb/0pPPWt8xJlfRs+Un/v971Z5bAgJdEXADL
gxVrhkowRmXt2/RHo8+doOvAJ/bLPvGr8BMw2fnHMWJWNTKPecoTpOXveTyuvHOoLL4sfU/cm8Jx
9Rqgc+auCr4YzxzMLYIyb51E5g63t3KeUiGr9+ZrTIPBv5oQ+m2QV+OjoN0s0q9nac5HcuyV1CJu
7D5Vy0pft85+CwAP7m53W3g1Hebe69uUdBBlYsNStcbTxbQoFUbdndUFOOOfQN3fjk7F9HMiSIIi
dzmVBPJsO+e4Xl3JVbT5P8GvhvJHXR1W/x7I26pap+0fEg0cm41UrIVeTuReX2LC2ViEzYx5AOHX
9NhTnO4AsvHvxQhvG8XvklXaDdk5Po/OG5gRaCReMm0QQxYv+JdkUQ4M36gqIY3GWYrUEiDUOUS0
1LbpqGbw27pnNAWzeSD/GMgV3zDnlkck8QnzXj5BHhjFX9OyLbXvuBoTSTuf2rKmpAK6ldnLr6b9
HLZ4VOf9B1WF5p9xU+jICV1HAnQlX4lt3FqRLns2EZro0pN4CWwJZB1MN7l0k0RLn7WpES6KUezJ
jeDjvTXBecfcqMEBjmIvHqGzWBvAbjmPqL4kqcfBScoKIT1Zf4OGcfwHT+/MQfr2x2/Qc3XvH/qI
MDrkZgT6Y574EeLnbmzJSzjNjlG0uxnx6Kb8bN3xbVP67AdhUbH8Q72nv9rvHb5h8VPIMKg162UB
QVAgKH2xon5k6eBoG87jIE2YdK4d7AsVSjJtX0rz4wiWfVY/ZgcQYQpt54dJU6eS4ZCLBSQaAduF
hs9ixA0/tzyf3XGMi2+trFrTdLdib7Ynpv4+YAR/mCMGa5YWT0unjrbnTNFnbx5UY3zQB20ttbWu
imdGZmkdaXeqMznGE4ewoNwIOSGHVo/uZ8VqpB3rhHkk+TMaF1FO+GOQW3s3u0M7Zba75ENN6j8A
agK1TUD7cuDCNdJqmHoDHARBpdQINn0ighxWIqdhJVMJpeIwg4aeRK6/dyCPJUwCitTmUb0iXkXB
gBA+aR6Qpnhk6hcOCOtt6uG7qG+X3bLNigvV9Z9oSOW9QrqGs+50nh9xzl6MOnIUCG5jZGH7NJUd
aDFvf44du3QlTdusgcIiMnyCPPz6V0ssfHyxudy5Rfiny3nYEPu3pEU8XEa3Ub3TUvIX0mT7Jh/9
xJhVnEEYD21FQHHzvvSYjk9O4b4OtGsfA96uewjh0H6Avvb3IGVCUuWEej6vvpEmJ2ZUcC43Xqki
ZYDhyviGHAkuUSbUbvtZMdj/OloHpI9qANYDTihEpMF7EnzZN/FE8E3OQcxGFNbfEyq6wmTA1LFv
r2tPEOtn2wQ/Y+3WaBoHPIPG5BiOzQ1sVAgOlhy5oo+o8GS0cXrtbFXBLNIiJRWuUbMYLVKWCnek
UxA2wiCHgZ7G0yVYlzGqIp8GA9MfY5j8WfwjhOpwS87lAvp1atCvFjwANQvczcwmjkyvTHDKtsG/
3Q2ehkyLNYv2FrudzX/NNm5hM58w9L4h25r728LRnpNP5haqowbfCijOmdhoLBSXkm7aFUGEpzxO
SdAtiQdu1ZM7lYRSL/WkVEhDjyG8jvzQDX0SpcuopVsFqtEsQg0aUQw4dft6SzUKAC8Hnk8m2CJG
KCrWV7vOMaNn1KY8q0OBJfqUVsmj8GIU7XY7TQGfohksdqtQ2+AEw4dSD5EnlmvaG5YJcSs1jg27
q7moN8Us/+fgAGpadxJ+1SEWHmlFngVpKRct1at0s8W5LRk6lePUgnW05oe+8dQJMDhgzqOdVQ+b
8YpZf194JqmYXTXsh9ujbPPz2w2xlq/VkRAOnz4ImqYpcZ/vDpLwguMpi0qbyNekQepWBAikrOWk
A22IZ3UYt3wbhKV2QS7If4K20SD0gpLP37EHvnF/ovrdJuft+8AWOCnoomebTjD3AsaULOxxvHeW
8wx70Oc19efeYKyj5GVqw1bjAKxTvfa7NM7cWZSbie0NCuFjUSUCmFHQB21fqXxApuYQnNMNKs1r
I1E5tF+E75dH6Mp43CiyaEkhs0bvxVbErXIpcgOBa9aG7IjdDspKjQuZVxEQvAOK+i1Fo/8umGgt
n/EBgMv+hVyBR10ngf7I2O1DIbRZuIjQMC6b3Lqms9p2vrvVyzUiZsG0qmsABGfYzpGVQfUmCseG
bW6IYOPCD+XLDokaLsziQBNZ//RNeRympkt7eJoBjxgjN8pGAdU+xM8pk9bpdLK4vwawHTf9U5KL
TZaeUQ30uhROx7WaWdfLxFw8WGmlfABzkC9e/WtFg4w1x9PNxKTD1+lyf5KhTh27ZkOWI1ZfK8hm
I40NjFqkwZUh4mepsaTC8UdfhCtb5x1KLSb/g0eEB6CJ4krvq6LtfKkakTyW72Os8CRnkkjjEObW
tGfUvMp8I0bSDr6z97RWMF44iHP7a4KSTYUG8+EQkXQnFmYLIMHd/+l2pzbPoWcoba0DGhzsu8HQ
aGoifuEpHD46vqGt5o4osnHzxELiI6NVKD1azJJsMPpqA9IqAqBHEFePexS6/GNy6u7wG26JSpo9
ZORqG/hc/dzeyJV6qsAApZi+udOeH193+3qVqpYaXtqaFgJ3rGZyyTCN+BarsZiTK1R3d3443m7t
XUVQpSMlcaZucyPVpGV4kO8wYtmXSLfTZNnGYByN//aoJMniLAMELz9uoibR+VLtDA6M7SxcCUCu
TWXnxL7xtbmBqIkwlAkLet/dy++MNO2xL9DPfVk5RY+yuryNCVTnFJfAkxUldUMOwbxPvrnQKjiZ
6w3S4Jq+EHMYyWvAVAhXwyDBpmNCDzaA4QoUM8L3CKVWZG6PyaDPcv0Bbatkgw1KSVb4gR+FUhdw
bRxBmOgKJuL0uSon8NTqNZDoEOIVC0e9wAI2Gb1WI0iIKCvSCa0CPcxQV2mvJlr7cITQ9KDmhmnx
LChaRhDG2CgY8Y6yUOtvSFhiZs+euy0fJjqHnhyiV8w6+7kL64MyhpWg7+mUtgW24HTfl9X/F4W/
8HELvnfrakl7NsKzrLX4fG6H8mDRZ39mf4bsv1jdMaGR8F69pAgRVIGbSRbmplCSYS28PiErs4ih
InspSDNHZ5Ae9tdluoFQBjqc0zMtZpwBmDBLko8ZqnYLIL7dE6eLm5MUss0kojr/ph/mcVp7e1Ki
+wBXFmtaa8CAqoWBg57eMxjndNjIhd/MIAwX9xBcuAuhY3dFM1rEoMzQACdHYrvE7vwoK7Jywzrh
A9+Jl560ix/zQW7CM0LDrUs8pZPT52UR/FOXO8PLzYA3zMxaxWRou3ROzWITGE0X7t2OFmPozZyB
d8t9q962fn0VX+z0CBTxX/W0vX29UlSZOnbhTC4VkUM8C4wjF9L9N6Fid+MsNRJLOAiNc5OS5+JJ
Cqj94gUwxTwkvPTzmryYyU2+Q6XrnF0v2vmwHr3tFyR9WIQmiikfNMIRHcKKPLPvHPI3Zh5dXhLd
0KFOMSmHSk8Wre8z66FSxfKMpfUH4NwxOz+T3BgyZnbB9pMbUk9GTt5evSKJOZP8qaOqqcLp3OPz
dfnotkOBILj+tSE1s0vyN2Um0ynxuAjKauz3+nvNGGsOFFN1paGFdIdrPD+Iepj7wFJ9DATmTjwB
41oj56hMU9W77doWRiQ3JVFVzb9di3zla0lHubtt50K2i+uAd4vj3gLyBMUhTsbuMZjjxtHtFaZg
6dJDKE6L9SCKSATCRlCM8KQ3RIemFLBrSAe2tkMVUJMlixDM0B0ZIvnS8mOXQGV2qRtsnEyVTaIa
vU0tDW90WABLItMXdVJhXQEEWKcfTc09WjJiJc81T7fI2aerW7m8zGodAJfSH0nDACHQD0hFoRA2
M6u4TC2ZWKAcHWut5nUbipOFtXv4tP9QuRikF5XAkAVX0+xu4H9kg6OrWUi+y6JlNt/NxD19YVz3
+2w+/116AgDIk1P8WngJ2etSBDCTLI1hRnyHmSbn9Pc/Ju4/cBsWXrbqkLJ+ZW224A61QrH06J6T
X7KWvpJaA7r2czgArnD1/pZk7h3eGXqBj5HxGHIXYfB3YFQCVnhOwdj1BMCYKITcp2rngv5plmq9
Bhz9PSVlwMzjirRqEPNCXG8JlLnUIx1XKquLVyTwZuIEQFWZEsqzHkjEgRN4tV0SWbpCCeAsjNBk
TAih1qUuEVCI3d+rxUZOZPF2YhUxzXwlEHjmZltQCK434/pbPY9c/BRb3QHilJn2SUlQEaifISwF
t1AYD9iVZU5Tzr2bFQc0LF2VrOIaZms2rVGrykqBQ/atsEvIW/y3KhVcZtqo5OJsGxBraxLIeazk
wDjj5SzGh5eGFxsKZ7TxORGQtlciWZtbbCEmhko7iuBaYxqHICxRXrdfRC7L/3ckMPnhPRZcAy6N
6oBzx7PrGJUNk2/i68vDY3SHwB8r37XY19F0V0neI4XlaFw/QHnN6c2X6g4kxYB8KzhkuTtZsGMF
j0uGYQQTuQHQ/T+7GsKHFlAJBMEBiJpDE50uHB3AsxCZxJiFf2qLM2TKtFRXn9U4Sj91gpFq/QDo
Pzm/g60RafqzzWKmW2Zo84o7wbZnzk/KRBCsDKcm6w3oyRSY4wI6ekc+TLIMW2e0QE+lN+gPzmKP
W2gEIy7RRVLfboFpcY66zzjvx/gE9TBb6pTMKd1ZmhqINeP8QdjogPqLIWNQvlXukJzv1Z+YstN3
7C1i+q5GYA1VHT0prn5vcLdcoKPQmNb+wN245EnqqIcKtS39+CJvrcBLbXiBXMqPbSGye/fqYrcZ
J0YM1nkot0gP5avKHxZsHFOPDEqUCZFvOb0nrsZ1zOdwzYRnC8OTN1j+CNZkor+S2iw+gPZIZa2y
lf6PdoG+fgwbEKtBAof8BCH2aRIpD5MHBeX1V0H2pFM6tDj8DcZcRr3x8tUEx+LYL+AvLIGp75Xe
8BF/yREGYLqH0M8gonlX10aZpUWKs0An9Tz3YB/xCF3p/W4BCARQxQ9uhlc/jotR1ZtYu/hZnPmc
ts2r+wnVTeS2AThApHJUXgb9vvQ9IhV72QVel29BXcp3d/TH4zVQeVGItsTA6ojIXeB6OuFl6xgh
jpsrFDRsdY2c6/wlnodpkXNf/wy5UQt0ALbRNSOmt02hw7WgphsHNWUEgJQu5VO23fbYdhJFbBLw
pkzMzUmES15tZzoqMHOXtxjrWXNBs//curi2/Oj9qubHx2KRB2aB40O0lYrYBhNwxrT0fIl+Kvam
pXvSpTaO+FLzxVB1yBaLtZ9iVahT48j3wke1HdvMNLks1XQGj0VT56y6U0eLzorMsHi8SVwT+U2I
MXuc1XPv0dxulSZ61YWEy2aAwfGByXgRTcvYn1EiT5muOPd1MhLN/GV8uO76+9AcJP+8lew2Vi7o
oDut1Mwzc/0lHCPmSt1OKVLL93vkGzVlPJP/KoMUwGOK9D4NodbmQBas/mz0XhnNxEU0qarXh3wM
vU93oFoBZit7zq6iGEavYBT9rzvHDXAjFp+/x/wgbQAtaxZpPXk9dDxnjE4aGqSglJ4XOM3YZr5n
uasi0eC1CrZwqp3az21D5hHaztNVfyjlgYe9vQDn96vkR7EDv76kNYkFXFmnyoJ6TvEaQHPLccLd
sBAnNmBW8p6UFw4ie9FeMrF1wgmuJPFVUhK/Qgg6mm9Eg3hEUyN2K53NsUwUUEEshaMcVVLxvab9
lzsLpX1NeJXXHFNaMMmj6mrNuCfcs4JJmgR4fPDAXRDr1YylpDyHKDXSTtYncNQoBCMEuK1ixtCz
pv+F8G5DZIk9ymeGGWQy93lqhkO4YfZvZfVW4bLO6w/JBGswBrT4V4pidc5Klb8TubpPTpH1HSKU
i0lBLQxjNSxZb9mcVplvV1IBILEqjldJJDAOgFYQEvoi65g4b7zRLL47UzK5mDTMBHxZK9NR89fp
vvrkx9mOcX5E6rzaw2rgd1RDl+53plXxmmCJj7DQvifg4tEzyY+Nkx6VKXyHdY+LmCBmZb3ow8ML
WkG9V2B8ifJuLv/+Fe16b3FqcMIZQ27yeB6b1nHFPN7kJ8lV/AXpHR4C2nda8l20fgeKsL1zYvcZ
dZB+7O+vkte8prh9c3dvwn3Brm9DlG2TRjCTBdVnGXwrUQZPntEb6QiCNpPTAQhhCu1C1xb+IY9H
UJWZEQpxdq00Z6+BBVPjUNfvd0QM83DyNqDbZ4RqrUg20TUmKfFcmy3gkgOelaffqcScSyKt8KCH
BTKwsxdbYwyKLZlQ2iQNLqBhyd3Dtn73n1SferTuiCU3Xm6YAA+zIEGA/jMKiuMEaEfcaqu0OQYM
kBxP7kfUBBLKUlhla5bon8OBwoFJILlDigd0bS68jzHd87z9erfmyu6G/EHZxMJ+IQGAe5gI0/lR
be2EPQF70pmUPWTKrfC1hAe741jD4z2cXTLO5rGFNHsEJh4L2Y2rFuHZqBxxpnFKbM+kFNK2Jkf3
l5skBz18or+gMsxZU+Vf95Fx5RL7JraOWhXpXLrtXCqlnWUv52ObAAk9GFtbZDJVJHiQ4pHzJSVY
4i1GCE0izTWlErXH9JVdYIin8ZK0ju3KIpKgF++NIJV5mZ/g0z85Ud6dFy2+1zOpsSWwXS+oMMm7
nhVu/4kCjGvDzrB/kes1+rkLgWWYtduWOv05ZF4xPkCFjZI7XnTdmFvnozu+V2780ygXQXFGz3zJ
CAjl1IJLG4nJW2+SYQJnZ7tIVVbWRi8bUvvIVMCsY8d+7BLrvrTagkwubWgb1lGd2J8fDfkOVdr/
8IxWnZ5I2RsUcJ7hNX7eREh22orK4lcEzJ2JpEc5xxJQui7h1PVNH118TF4bBlcDuB3o/uLetidj
ekXbogxVDORiD2ptW9yQz/8kpD7D0BIak2G9ojnJ/Qp5PRYB+jobLnh2PWUr1PNq0cSBkKS4LQdk
iXImVa79Bbc43Jf1Bec16AA6OC9RVNML0dry3hcSKB4l56rYyU0c1SCl3Lwp9MLJFkEk+DLmqWpp
NQ6hgYDlk5RfAu+ywcTfeFW+HPrkpAuNEIiFpm6PNJ6JfPAGjTnTb5n3O8S69xXg4SEqjdDnwnZD
72C8aSmbxqjF5YdjfH4S8ArcFdempoj2apna9hi47Xaa87yyJGTZkNFYQArvRF5QjQoE3fbQ07eB
72o6msoNCYQVac4Tvnt4LtMp+r0HKqxH78VbgsI3bZjzMVli68JD5yUXJ+JvCEQ0tXB0meej7ENy
MFpyq/CBndJVmEx0WixJstyaJbx7njxSjdtSXeyTtkYrC/0qxDSIJTHUAFEDniusMo55/uv0gk7b
czmj+U3T1cBM+d94QEvIjXITUm2m9bZcCDk6O6zIQ+DgBhfSxCdY5VRgrIayQA5YVytiF3Bmt5KI
eFNeo/f45MPBPfyKd+omxy2EOWOslOrtHtUC7l0Pefi1bOBqmHqN4igeLp+7QH3uQypZ76V3ZSwt
8SBcbFvwrdEUyuKXO/ww1b7x92/JC7djGnOUUZqVKnXIMaDHs8rq01KrLdX3o/SFgxQUKl2GiJah
U0Evv3jH3Ui9JF42hCbynzsjM3SLFZTHn3cIa/j3R62vvi/GEkmbWtFU2FLScSERsgH+uE5RMTZu
CRgh6T1oXfrEYbYC1Ftjc7nn+kZNT0T2rd/oWw1aJLIXbbSWVLwXAziwAA1hycjwCGa9/wTKVphy
uKr1F6bmUnKqx+LKDJVHR2DHmzeMdVCzLfWztnEaBs/OYIb3nNnXxm6HqVxgNMo1Z0qx5bBnZ0qp
9/NhKONtrgDp4Uj0O52V1YUXPM+fF+KFB6e5om13vLWrqdFA3PauaY8I3c/q80I7DhP+DaBAWnpP
UHwvOw4uycqyTwT+OQCU4Aaq2rXQRHbX0kJ7BOMW676nsDy+qn2MEsW0h0daavyyvU2Oy4FYFF+2
czRA9gPNUdsTBPl6yvCgaqkNAXpR+XrsRby1KefyWRTgHWq89SKF7xxbLJSmGUSgqYDenyt+97SC
klysk8vSB6VC2MsDFLMU6jZZWJ4JiPHUMLGXisgZ/7yaJdirzXU+6MbjUakWCATfabrTRipjPjX7
t/jHrOptN+y6Xb6gt8F9rf/43pRPEng358mnPz7e1vyrfVYFbItn84nxMK8olx4nIco70HrpR1ZH
n604oxIQyDgz/VlU+yRmXSZhh5+UK23qltXZtjQK+XhKKzR+oOr+hp7NAdKTvTYPWzh5K882XwJW
a5Ut/N7yQLy6gOTv3XePo9lUgTvMo3CO83T7iNtNpnZSiT54vlMhGJ801nKT8HnWvu7HuOv/nF8B
OVJWRGyNDMvDiJ0CJ0xM31pPBpkEReNO/ONlw1iSgtEHPtW/wILGEV2pD40JU1MJYKv157u2CYTf
tEh2gYpf9MBELARmUJT1q4ovI5XTZHlRVK1DQIeEyTcYb8vziPRTXqIS6e7asV6y1otWOB6P7hGu
a9mPf2JLa3Fas4rOCsaAQRQ4e79GEnzVIEKdaqpEQx74rOBxFI1obu7CGeLxHIr2a8G8yAgYo4Mu
5DAIbad6XM8f0CFaxqQCqS5/7HsLHfoFjEX9vZTLWjaj6VYebO/2B1c9pMmQwfRoTfu+RZXOXZQH
/4EVeD1pVp/TZb5Pe0szvVRXBfIJn6U0W/mEhYYyBKolMpXA+UJplEMFAb4mjCzi4Rhm5Yp6bjtY
GK3hofkrBSkp9nNplyFWzaekxHBzg6TNIzd2Ont9U7jx0LcwJGGgc618imy2UL4SIgdNSX7jeMc+
4Ge2uCYJ3taI0pslQgkTg2h8kdukXZutFnDdnbitB+BFJVmxkzOb7AXXG86y+YfojHZe+J35Vm35
32Sfk3R48vzP7p0dykWaWSCNTdRD2669GqRAdUG4jlK8XfDp7P3h6omerFigyu7o/+d/OhUd4rt1
djIxO3qnR6ix9QvdlP1MII3kIOdEMylswt1WuvTegtSJ1c3JQoLN/aWKLLVkCrlgdRGSejdGVmdF
SGHk6GaK3GWBymu4y8Z4QDcMigDN0azXY97cevDI+6WVhpVlMnEraQ70s3MxT3g0kQ+w4ohxEFI/
RYjZQfRyrk3Fe6CwyjgjXYhZ4+bgS4Wwe7kUPerB/kKsLBihAF7UdrujJmAt5d6nOHKxjp5BrMH/
gK12td4lXRkjMPg6d1bTINmlg7z7XKRItKnguMUuBhEFDXZax/4KWJJ6GqDjNOyNVXMJmABA6rB0
0PN7YvbmJobZTf2tAwa0f8R71hG+FuywHxnorF5L3DEUJ13wA0pm06LF378y6wd8n4SKW+XqdIsf
lsD2xLaq4D289nPMljds1qSxB04J+DaLZ5la6NL4/m5nMpc0SYOsP8qkdrol/uXvF6a/6Zw+qvhP
7itdlaXdJp1RThYhqr1TWVRirjHIm9ABFtG//cYHbWcyS2d4NlmQGAEiBowpjfmfvzeIF6gFUdm1
XwoEFevfFmoQlQZ8XyNADmvnNCm0VwD918P2hOzAuCR8Y2d6C/ZBY0NMy5QfVmBIPzosDmdYIu7j
xpgydbd7wrOfhhc2fjdLf9NKq3AK/T/djq87cZRHOMdsTqT/DZxDjGD2nUE/2kdeYi8g1sJ4NGl/
4lUES7WFVIBbVPsvtGYkuSQQA4b7za40Vp3yvvqr3M81RdvmL48vr1Sh00Z5odaqJH7osIr79QMA
4joRb3S/1JnOXMoEQe6gpUfpAfs9zUfuSZZbrf3JID27AFcqxA2wBL2no5wx6YdSmzKem3TNEVKb
/NnCfHloyXSOlxBrROrtfAztIHkIzY8DJQ+HyDebB39TX24n/RgS4i2JWyybzN+ZC74Z8NpBJ7Ry
pmO8rmifjBd3cZanqgJpOYVBkU7svIIYEKXWVjslPx8VFE1EB5/UMXiXTmcMnJo94YuasHzswM1S
lTYP1QWOPXyzrON1z4XJiN2HUQKN1Hpv8CVsORCXXKOVnt/zdn8i2nBWKDR2sgzsMOHrIjmuY1AJ
mB4v7mBaLryHpxbMZBHedl8sRtgoDQ0cW/PLpRMMd8BrWPdkTmpe4CXjhssGo6oLnTLyMi+TSXVR
uB8q64JHpaiTzBBop+IGJjvcEVDwShtie7Mwg+VYLlCeX14+lKXDvQ0EA1dATdzskwmI+ibBt9/L
rcwvVBRzZEt/mE/R0keUa3GwkkFnm7zRyZPuphaTUCTwKW2aRYjRNB2oyT563d0waig5O0ud89nl
+i1KN9MYZUeUP9eaptWoDsW2pUpgbFCg2UE2CmNgaH0HRrC1i3OT9dIlj61hqqkK+Yia+jmcQbto
S3j5uI99UWPGYUAEHLNFuo1yLkL53dgGQOdS9k8+2IdJsIry2N5ObFg9Z/p1Q8Zp8pwjsUePN0dy
eiDIaizJLEi3Cw2wFmFm32/mk6NO5a7zUlijJ0XJ/ArbkxEurwpTYQIy9GhbKqdJUlf0hvkIxjKF
UIH8vYqpYmjnatcMi27H//sEvXxOI/ZTtM+VSLko2xHc1IQjigGiDUt2uZ6haeU3sSGcYVxxH1p8
3/zyeUFjSj0P5mXuuw6YB50Ei2JCctfXs/2eMrhCRixIaQlfTtsYxpwpFRzHQ4fvgam9JrMpLfEk
Mw6bVejjYplVbSyNRJfO8pA4shgM5jKvTCKp+DPx4114xvz2FPEQMhwUmKD5g4/iUG+QpazUZe7p
pZtuhPhMIOqHYr4VMUgQ6TvwYj1jfQ+hFsLPVbo6/htGMebVIpfBwtFNirToqr3c4g0ur+jh2n5p
Lsc78LwSSTx7VScqmXldCTIYecQI3SvjH69f7r/3YekCpr+ysssLiWVZ2psqySYDp+qHU4KG8TXB
zSFopdzY1BN/j3EQItJgqHDgiqd5D5VU+nNAIgGAIBEbwHTyiY2cjpwawA45TQYvaroz/kdvgxG3
qu+3PwEqpzX1JPCf9qCL1XbvdaNYm3BAqdmLrX5hRD/hScFTGvZKzEvBO/zPRBiGPOVzumZ1bNB6
2mr9tOhGM9ncO4H7hL6jWN3l52huWTDVraxDPh/F20z05LxeLksH7bBasPpSqxIiHdF0HUEBcwxI
5jQELsF02p9Gyl8Yu2xPT33MMRLQlXcsB5ShxHcXOHN7EDcZg/w0oXXJs0+zcuB0N01Ow98P+1gT
vFqp2+PpFb/PTJsw8Pzudo1H1bDR5pZbi7o/8fAhTQKMNQJKFtjxHkyLqVXApWG9H0E32b76m7VW
pB7Z273/DS6aPPyMgZ57TVdzejZq9pTcHdG5fvg9gSASc/2FW8SkUi7l9WMslLKVEF7dy7W/M5rD
zTAKkHcQnFLWoUzJaD9+tKc/+TfoTjpPBjKR1E4UVm6JEFoqpMwVldyC199OMKbBytl43QlF8IrQ
2FaNcGHcq1C6+hNm6dl2E+mkMLQU2x3wdt53tB/J6utGvvm8GEaccETLY2HONVtrt+DHYdRs66mg
eui17cxE7QkLhzbnS03d3D+mWvvD0ESFG2alMVIqfF9+CfFcYUW/Xcsw1yq+XnL9pcFmHnmDHs4D
i1h5vER4xGZ03SpCH8eV2GOqjILHZzHzjF//tTbcEgKZ4MenJ/998wI7amiIQlUVfh9Q2yUQu31M
HfN7Qox5YL7loVBt3jyDO1wkjrU17ZCrF9NZR2HeZazB+rZfLLOaiOQu7ZrzicKj8y6O6lACczbc
V8QTwVyqCTMptmlF3RXfouOBFGbTJr6oIRA6dtdXcbEZaYz/L4cutciDDR7kxR6syqGYDh5s/Bai
IB5zIwoh237iZy6j1720wl/E7Df6bcr69GQS5zhoyThZ5Sl6cId4aPHmEjk6el7v2OWNwGgdynVH
2L6nMb5/MLTSwORHN2/O4icaCoko7qxIbUpeBKX0MPG6aDO3IZQwPU31JhM/Mj/Ifw61RuKZoQLI
iZCuU6zpOG5zHnKB4bM/Pq+9pcMG1rSM9uORXDQ5gvdRyh23RiT87xwtQKyeOL5YJ+XPWYf9EONG
cRijnNozRdEVZXvC1oBzCcIari7/TOln9xLgDFHs/DS/jMw9DHzAxh26tOpzptzseIXqtt54i50u
VrMiMaBGOObTRxLpZV1sRQk2x9BLIHvyE8vvZap6xwy96/8LGW9tJXv4aOSqDJwLkSlJL7PaAxue
NUZfuFShzMem51xZ0mRhc8quOKiMm6os+pH0y37IeZOnyxsUFD/ij7QCZwIHvavvVVMa8BFTZoDi
bu81zDlUmLHnatBBazlor2lTASOUydBz/olstyxh1WluZ9scYPC2wA/r5EYr5IEoBgg9OE0EVv34
OZyDF6YF+aKJg1cW7tAsaZSRN71Vv4wv+kgTaQxjxO6g3jnO+3LyT8GPvE9lZ8whVLagL2sHaQ/4
akqJV0qNmHHUJ3idKMcWsgXHSJ4SfZQBT34bMV7w0ymS9Jv6Ojf0qqhl0/j/bUJ1yD+43AghXKcU
kDucsRu2zUiFjRpbsQQoFW8UIUWn09zGrj/oyaMbBw4n+z8p02R7lLbnvjoMgBPnakIXDXiSM5h6
EKd3sGUug95hq3/2jqZTekDMdpEH7n1SlcR1SpYwjUW7Uxq1UbgQYJNzbD4FggOG1oATR6OFhZgK
RDqwP4S5ctmsTM7MUkYn/bt9xlFldWbh1z79/m56J6zGNmWxygxl+VdtZsie9NIftShI9VLMv7jW
jKwamiuGmWXqC2dkPKeQxpv02/bY5DJsHDGeynqhQ4a3peaA3EsW4quUdl12U5WlNs8kR+CjVEeD
MNN0rd//73HLU6fF1Xcb26r2iiQbtnfmU/BRuX85iDBhV+jOT0PQ6r2FUBbTkKa1C0ENCHPOMw+o
Z4X+meoFHPJJOX63KyswVWstN2LHJUpvSHAJC83m026DpgQ4ri4cCHOZ7Sb4URMZTnOeGu3mqWRZ
fk1ZE5AXEOXKsxMaN/IDgUPvfQXf31aVgRUAOCwNfJnLmWPf7DPd5ZZIRGVRqTpzDesR3N0oBQHc
EFtCKrY6xqg60lZ9PqCWts3yK6CBzKouYfreXg1zvmFBjM1jE6usiL/QSukPC+aOhx8GEFGjFeF/
rS/EidIlLVP6B5hhtaSavmVLtJzDXPGguewbufKCx22VQSYzdLb3YozQMLMtz/lgHif5PPste7Eh
EWZnlvGdaJ5ZIorar+c7GnpE7NmobcW0qxaZAE7JDTWCufkDTMsKHYqF47zKg+8zfj8BDHFBGkC2
CdQc5U7jLfdeiPa7cScdKLKmU58SXZ3AfuY3yLl5xxVkQPZxSrK9P3UkWwAHjPaZU5JeYAQztZc3
PIpQd4eCzu7CPbzH4+9I5EZr+1r5vyFB0H1+0/RvEeP/oMD6GUGYiUzgNxu817/2r8wEwPpLaVzO
N2rLN12LbTFCPpf0VF/Soc3QQV0JCJUJeHyrDMIbSIObqFr+8Ejgi+Pw1jehQAnmmcPdCcHLoblB
Cd6Wh29flKCv02KvZ1ds35HPobEJBugexgKNBxnEh8aXJCG2v3ofFGqF1MCkDekYFlAOTTLtDbBw
5JaKXwHiZWwdxqfMsbOPrUaKqYRv++leIkSNsto7p9pakgs6rTyF7BgJFzUfB2J9e5aP7TgOY/QQ
fpqb8QzKgYI7+CFx7HQdS3zVj+G06gQVW/jRKpyn9/lB5+5S1kTaeSj5EJ1+whE51DGUmzbb3UGX
UYBaBNx/RYyDOEDXCTL51CgVcqt5y8ryE388kOHgxCEk/8UhXvIfPqyECwh+dSOzJjfrGyyVuSAf
84NwszomxQb1BWTKVu8i77pLz4bghBpHCRSqCPIiYY1Z54gL+Q59dRSgDilLaoMOC2t9vNb4jrPH
S8cl2GNSHL/E6ZE5MHQfaj/0U2k3pbEJ5P0ysnEkBltEdjhvx6zaSmHqNqShGzoICUNWHh79tnL6
wNC/aDEh5sfSI6ZHZB6yA+bInfWMV9nT4CqBNbhHNEZoe9JyAp+ZDdB1c3vgfMAf0mhx5OFI2II1
7xnBljBs65EiuxR1j8uSLsCeNkGqO6EnFwx/3acsatHwXjPj+QnFG9C/lzqvS2xGVMpKh/gJYsyq
uYSAXv9ACFbAcrUmCJIIueqZ4WzdmIbEG1jzoOnsjefwoQ5Uj4UW5xgiLBT/XTneIw2hwyDIB2d7
zv6Ekj4VMiStUvg2tTvA7+WSna/ov4QLT1bRPXXCC7TmJAzH07d9+GzQVKCDc9s+UnwdtYOcHNMp
AYjUFFMTHEoZRd+zDa6jwPHWXWz3hFiVprCKIBmNuxp31ggrhZ8ULp4vrojEaCizWAr/9hxGZUlQ
qno1hquYaagn12e7e7zSDTBAHdnY9x3ED97tMsIC3hLbUO/41oQhPxCT0gRlh8STMrxgdx1AlTZU
3tYRaZqpOqifkVHmu58bC3zkTy0pYqllv+31ben7w01vd0wB/xbpy5eOaHZ5bLAbilud5QZQX6uw
sy9TsaO1ywjflI+YlbXLZ+13Z2OuXknXMzq1CPSPWCqSH5BIciOsPW74dALasgBfZK1sr1bbhJkO
doCEf5gGSZt0/ieolPQhcf1/vvxRKtWFXBTxv44FIdOQMkHVIpgGlX7VSsJa3QuYDpT1aeNxTbW6
MMK8amFeAhFEIypLmWNHak7TsUwpSiHfvpDLbU27k55bflYLiDZeiYAvb2fcUeWy9jvl4/M47ZWB
CH1zQZgJhMpk2+I/p4o6Zm6a7wV6RNpTHZffOV1fhZdY4N22EETAC2qZc45N/FSw8SXaPAf3EUW6
mUsFQwCeRZR+HVDSR0VtsaVbF+J9ZbjAcifESsqrkw2Nl6JXA7bCLzrVKkkRQPgTYgYoWPFl4DGD
m9idgFFd5/lOsY/QevaGlQflzSlKRfIj2WdHWDcsyEGTVwG8PCQWGUbiIPMSagHbx6rWFHRQbqKX
kxkbpkr9VRfPgSY0Zrg5ArM+SyGH8HgAcTBq7WOMC9DQ8Ac9RD8gO18JZMuTWwfH9+9edVAOb5w4
/AVvr0ex7s6i3sEtHVh0bvhRygk0WMEhhWm2TVYGaJlqjdALVeVPGmvSShimu6/47PxXogZm41DX
5ZO792F2+A8OaGDSHDmByAROUmLADjVwzLUtnbMqrOLYZaLtStAhPRIYUPo0rxpYDist/jUHDqFG
4IjqJl7LqjG4TGKqEjwzef74BsY2TjkbmP1k8fjVl0wKTHxiGSWsXFUiEolBiATPOoUdFRArnejz
xmWu1cPFslhBZqYSGMliyIR/i6UIR3PoBY243xD9Gzfw+4KK+oapvLuOC0DirYZZRbDAkGSBTNVJ
rqhhcDZlcMqMbEB7b7iSMiVa64TfgrkcP0G908qO2dytaayFrXeXDsHcncRJujlqXir1y1P9P1n1
y1s43r6QFrkemCm3+AVvoaF+BWJve8fR6lFrpHui5d8ABnC6+AZVpjUbxaiOpU7U7MbYjjEqiGJ/
JMxTFz0V1ZV1DvW7hejXqkCm6PsqreQdEydEEskG0XNKTBEN67Zq8TXMTGcOZDMidpfZKNaXVoN8
1/hOIY7qRczOuxGesiVKfM/iLVPItuqYj6EaLySagTVH+CjNhDI6pr8MPPhFtMNxOnpa/ddMs7wB
LqEBj+FFj4RWadxVbpyIKqG+vhZrdcPjiXeALKj/l8/Eyb6YP7wCoLojDjv3T2U8IUPlBVCholdz
tUuS/71smGLQxrksoKvUuhGeewF1bh06aVp3tZsYu0QckibqsADsBil3NoJwcsMGVVXPh/v4eYRZ
4ABpk99+I7VFGOTgtj94K5lIsyI1O3WoskA3sPCN2MyHUPLUTY0/1FT6sr+yenJvG5dFhLV1+nI9
m5Oxm/ogFLulfejIeOj8p951jJJARnoNyy0Z2hNSO7JOaknbTy2a5Af7seE9lL++Zxd0qyX0O34U
EAg+s/adAKtc43SPnuRE/OuP9xw+6cbfxZX5nYaLca8z7cItizo/9iWUfxHqVtLhoS08Hxjup8DL
xtC+hQlZ19ug2WNOKl964uaYZdimaa18PFFFsFMdgvMlbC31D2PE2S4SCbvGiZ0ewmKrAk8BmbpP
7iz/l5ZWNc5+2iZeDeCDxC4B6OXE6VpkfzG0ugve8gOtXs5s5Qe/ZBSArkMchuu/j3t98vk2AOuI
PHdPtZgwpSD4cbYioYBF++U/KY2NWtT3hFRffTXuRF8MFEw0hm50+fpktsB6kR8DuiisSUTnVBmj
GbVmAffMbc69rL6oQ04xSLwZciv6uLfA2MjSZXqr8NIbYTFpuuZBLBsEkiVjQrXlrIny3P4TAWE4
0CJXjX8TT4aDR6iZeiV5kQ0WH5D6a7JbE7aBkqfHd9ushQiw85XOBkWqoin6l3h/V5pJzl0FA/Wl
znky/Xf2g9uZSTNtB6XiMwnPnbugSXfB8dNy2EYD0ZzDmwuu66zwkNcTnzQfGos5gw1I7otmDhQk
EJQh1EQS8h/6BcQLjZjcibhUe1L7dSKN+B6Kt8uli847H5euFSoMwVEAuCA8lATskqu8iWSKnjoH
VyQCcCIGUKOi25uF0BjWzAvEwrg0bk2IkqGAvjq4qt52K/E7SovcGUNSCUcap4JNueL/nKt5g2nb
SvZpYafE5wQX2aRwvQ/QHB45ib/euHnKyQErrylC3Gm37TpS6dyIwPSZbETKj0L8vmIGTJjHp9iJ
C+4mPs3zsFlcJRfRZxuzNRwi6M9owm+OW31JU3gh6+sdxdaqwkk4+Q7K/UFdBVYCKOJAMXaho/NJ
eF9UPhgr/yyowel+TgMXVqGQt5msdw5coX4cMod2jKauPgFpOhHK/zeiqJ3NJVcW/c0biJaItwRB
FOzCL1ARpQtDAEQ+tBtjHN0AGQL8qrpses2Z8aolFB4izoBqkQI5fyFaWUWHY1ihvYgLLpax8CQb
nsylxV84TTyGFXs7br0clwX2HVniNheeWo+aVaa6APikdbytLO+Vp7arIJ+Z5xqwovyeMtgq+99W
hzqXk6b9TG6SP5cVPWOb/D1sYpECW+5ErpKpL5Grxd9o896DFZF6dF3SR7FEz+1pgrLMyX0+FijI
u8vJavn7MECLHoCe6KmX+zvKMFXGQozB3bc66+Y/vBQ85n+iSRtw6kvKPEODN81hP++t/2YVku6K
otL3AhUrgDAxCMkNpzeVmxHIGDB4oAgMGnCgLDoxcZRR6ZDaXeF8eT39uhetyECYEaIstD2meUQK
1kaXAlFvRgRZSnqoa4MJautrR+judyGtrsv7bwkzZvtaimvCD7RbTEkbCtFpP3+yCdlM2128/NiH
O/c35BtYtnlBLpH8HUqGj4/As3Z9EoXNgtW1rvVJM4AZm4Csxl6GaF8hGYXOaUHWNB6jYVHJpf0u
tW3eE95qA/Y8CsTKlRnE+xBx0t85mNo8VLjIoqBG3ZkoqDmJxfGRAKtc4tE5CDzrd/peGGSyMeDb
5Q37y/WWNr5N6SRDYqIYZmayo66Hzqt9FGjdNqJuTfP5jzfKNOfIOhKyOPBdOuIJBn52X7PVbMvw
N9vlgiqoQXvFQY//dnJOHFxVkLaamr+HIeB98OneUl+3WQU+Itw4R10YFnkAA/EXMqbSnyleMEsn
NkYJ6C1BBMEN8j7C+40EqV6k4BKAX+n5aNfIYpa4PTSydQ2+e+PchcxuS31X632+Cao7iveM3QCq
pNEmMSjC5cLDp5vFpxfO0EQD9UDXxXLjxuHBBRRquCYKlXgl9DX5lw7FjNP+6B13jYL9Hzw+D2Fx
/HuX03cHy+6qUjpf7eOo+PPxgBprjKs3OB0VCzID2WIvr1qtFDiGV+VWFSlKQqBNG84SgIIzQfh6
bR/I6GSgDrnlqdBebHIa+xwYPFCjDwoUoMPB0HBZi2y9tEDrf30th+P/5qLw9NQTMLGMw5Nc7G3F
18H67lHFYfGGRJz4MluBhCFZsWl8K2x2iehvKaMtNwfdkteMnUuLHXtSlZNn4HVNAVcvK4vLOo/E
tEraHnWag5LbT4rNGp+WQgrAeOX8rLm52PE7oAW/RqbjqGI+OVjKeX/14gGWekTXy+Eylgdci/jp
MdvCIeKhdMliFk/h5u1+ATlNLNaef+BXA1xMsn1e+ifCfb/10suMdyQqX1csuLkoNdG7RWeVM72D
2L5YOP7oV5R22qU+0rVMh9p/rY6prFLbU/hacEF5p4JjAhhQAKCsiAzTOUc/SWncKW/bz6Eh+G5P
ECZHp5W1EeoiiEHBiO2BW2GjOjYCLfl+U6NphTBD8wuIyNqSyexyJswTOJpTjqXojOelXLxB8U2E
zHtLMWQhCVp6irP9zdcXkHvDQLsynxwkj62LXKsO4h0fD4IoCZRaqXkVuc9DZqDrTIA7Q0BtpB55
l24CYQyScUgp9yWgpbrFK1rtC5DdLXknqjOjDmkDpWHa+ZjkqY2ARRaDJk1P+kduNSsWmVIpp13W
YcEusdOLDv+Boum0GsLqnqOu5ccMYYWrf1pf1rdCGlTWht6He2wASSsWXXd0MDcQKMP8rVIx6GTz
6oUlYm5RU7HOjUfmt8ttiVbHeA94YUhdH0RuIC37R8KoTQCHB7L+bygUCj1oC0hMAxNbzbhp2Smt
fo4ovGKm3D85+fOej/yCgJ6GHqWJdT2dsI1GvZ2P7I3vVzFS00LJa/UPq9YJGfK4UC/Qirlyytv9
BUyAXmkOFjI6mz1L5WoKwNtS5eF3E5MPWoxZUyyaMkYylsuqqGGsqRvTlj6hbaghzTX351wRjr5i
xZaYSoCs+h5zT5Ya9IYUGRkUEZh4djDoTfzZbKAytRhrfK5OpVN/Sp71sEt3QKH+NB+RX7CLX9jZ
1JFWMEJXdJ9bTaqpYGuSiPU6XpI6vKefdtDQmmqitBUULvxFFC71iuH54PZ4V3OeSdAPzsVB9Oe3
hCbX53eCy6rR6DbjE2tx7rO2OVGeZbxlTUDCwg+ebyRQJ8xalPDe06KTt0Xd83b4SD7eMG4rdB8u
HflFkrXFgaWa1eeAKqojhSeASVGSts/eQ6JU0zCeWYwjUQTRpQEvH7fOSdIJgbg1ZGmfNpsoLe/0
zeRSQt+RrXcJSTsvoHVYZwfL/OoGtbLB8M1TxMHOw2e410H0CE4y4ujxEBRLyu0BV8auBEjYLolD
1QBEsw8nFItD2Pg0sKcVMYk7vGGxxa0SHqDLTkNBG6/ho4v2Vz6oJ9vYG03OqeBOeiz/3m1VdvL8
2hdZTF66Yu89DafYxmSL7EkA93MhNWjAoXdGruRd0Q65FRlkauXzL1yBzQCZfRU085W+IL42PNrO
dVN6b1UCnyvQkkuyOU7ifR0EdjUU2d59OjZ3xpdam2aTyydXjbMxWHt/aOhrgz/X8ODrg7nCkI+b
f65tcMoTpYXeqlaAMzNXQWll6hdfs2mgo7RwIHN6vDJVFzCwsuUO2bNsclGlHuCLSRqYVSFeWU3O
JBqKjoxp0llOgmkGxMNuUC1bKHN9/G36XepTUPnY0ZuS5IqRRmA61qXyc80QMjJQxa2SAtzPq3Ag
KuVNPylYwLeAEYLw5qVFAiuDdRHYsil+1M81c+NEXrQFzLYJZod41co5v/2zEGjkQ9izndQJmYFH
8VZgupSLOP72qQ+VjwHujeLuvuY+PVrrwO+7emPnZHhvM+joD3tG6aaziJzqFADBDaH53FDpgmdE
jYP0FDZLZoiNlEUqtm+GRhJzXfn0ueAxoaRN6eOulEkMteCVDq1O3AODVxwgD3UVs7+liOSrEJpZ
2LUsRYDXU/1ky+pfu9mxc0kBjr/xnEnMqX7bwW553XKr1S5ibTx8R1X1mgHSG93XcCgpXtcSxtzG
8QrK2giPqbFb5zi7dkJF0KZyqlWylWfnW1d1DNWbG0oCVq+27NXbyQTqYwPal4aDYYdHwNkAzNPy
UYG5aNA2SEJMRZra5LOfd1lJWjtDPFv9ieF/uYAaDl4ELJaL8G7zXV6lxG+VPtp5wa2xukos54kM
45zZFts50SMpMk6E3zHeraKwkGEOOlE+f0LRQjHLbDlV20cYecbIrbtUQ8Pe1DcZUR1ZGK851DQb
2VYxJExF/5gZOtrz9FYgmKiicmeJ1E+u1FoTF6ZCbzKa396fXL30fygXVt2upmiUiZurW209MJ2L
MpKIlCm13J912N3xTXKQcyA9SAqgeDqc9BGkp7lyJD4qL1+iAdcaxXujQzR//wY4V55TqYvbVi3w
j5zM9nk20L9UzbPKPLAvV/ry1gyoXoklksJgdeztyiKiwhXE0eALUAtfgHQ9R9wmNSQ2DI0hfyGs
O5bv2cNQouYLCP8HhwkGAp/57JFw2/z5NmgxC+JhAKfxfRCPzTR5Lw13P+5vPhUpmeGpMiJro+gB
738fIdN7y7kpRdO4tH4YVN/6qFjXcf4in/8ULaeWK9L/jo50tYERbafhIv4Z97UqbMgGfrirGe68
z48DeyXext8vLuKn3A8q1JYvtfUR5PH3bPWegwHoACwEjzJ5U7lPoQnwsKwb8MQgp2FdxdtZNpLw
aaR86+tVsSOuRrvByWdcwoWIAPz/a76n8iXBb04PZJ8vRuy+xxPtqBNss3QueqzDRJIzrGfCSnXC
1qc/lNe+rWkGJ1DG13Ef90/bSk3R8+7IbRKXSekGd1YMVe6ZcpYBCa96bq1AffrcQdh3MSUb02LX
lsHwnzFzj3SODZ1PTUx4gc1HTbX2hETJGEmx+VWMxk+wZO3y14RSOCxQBrDKxIYhbClCjIVfPT6T
lyNc856wM5yhUycbcDKWGksBc+kxYKE714wwMZR1H3cHhKDsMosGl/X0EfNSyKgwD4CuNW4dCjuQ
LjqJAxEnnCA0qbC6+gVzQ5FENQugBqfHoBxq9oLxW4lao5jnAnQtehwHi8zf8rI53u0T9UKV3nzB
ewougqfV2TpkROdYB4oe7xFdYGxLgDWJMgzyMhVUUy6pw+WWeu/szBJTUtuIbkp8XYVHXg86yFV9
fBFkcBwtf0RZhtPuKduqAPbbEhg/H+2hEtaef4KFDvpulUTLD2yBlZ6stQUyZNU4SLnpR+TsF9qk
vvIrKFKfa+2uGXTFG8ZytVEow0QgHONvZDDxRYrpkuGtKraRcKKZZUG41Gz+Oa36MU2D3K51km8o
n1qWW8BJ582WMTodz7LKXiZBOR43bgXtMnh7qS0QKdVgBs3VxC3gMYohyOqqQW6rdEcYViZIl+P8
BTUn96sqq6p7PJJa5WalWdLwdG9ev7LyRcxcWbaJa5GU85iyMpIq5048L4UwDrpwVT04M/NdFw4n
cCMJmNAAONVh2/z+5/U0h1r3nwb55lKTvfba5opdFElSlW7LB1/fOawifEFSUkeW6NFVPckwFg/J
YUVtb6caGbOE/oAICnCfRjnvCwTFgz7PcPAcObBOzCIjEjy6NRbjMQDd3YPlIWqJNDqFBnY8ZqbE
RDDJH6j8MU8AHh6qOR/ywPbkpfcbuz2OVG8nR94MxC4OGyZdDvRwdQlE5xoK33rHFflfdydEOleG
gQVLKHem4OqEVcYbceG1Y/DKTxsFQu2LSRVMM1ZWeNHtgnDvqh3PppmoTTOXKk4NcZfDt3fEE0QY
XzGhdF8slmocjBVh4zk+WOydz8JuYDNHxBXeTDG9UteERSf2e4Sqx7LxFKJ6rwNySq5wH+AA+KUW
dqygJmintEaI8vFiKjVM2jGOAIFoFO6JhqUbGxVoo0zRVvNQfsztWf0wXjTMQalmqxlQWNpEKjpj
6v8c2CMnkeFY57R+qBh8XwAj81H5mtPd0LOhMCN9iDGtniygvtB4vcIKC1dO7JVXZwgzO4j98koO
uW5PbmyCiZQcLnUb4RArV3Uo4HSKsnmAkfOe8tYLbTLuem9zT/8jLHCtniJVAJX1NWjDrLN40uJ+
kY3bIimtZ7kC10nG5p968FM461q1txwGLMHyfaw5ZK0zxAxLpAaNEXhGnqwZXyLV3YX66dpohHZW
Rh+2BllR6mvmArlWcbJTvcLa95suivqs65vQckUNwNmhh7jnTD//Id8NW4ceMtBZ3LV6K8a9+yV/
AeF64uczmNqGQlSKdfb3kswsWTnLXY0ElPSnBupuChGFk4XlE3JWb4ranWzyvaSuwaj4lYDggVP5
Kliivby5O9hcpfNZHgTzzn3FknR0OViW0ulXzSKyqHP3u0YBN+P9GlAQ4Lj+WTP+JFWz1A2NqdX+
l5I9BT3hoTQvUQunp4QZC1QQrTt/umAJT1K1te/lLzTXhsqUiWrqJWmQalDDrouhy9km8qAjckTh
Dp1e2NaxO5mIGGnRWdUUbUdr5gcRBS+xtt4VXdMaj4BZu/nqi1zAZUbmI8UxsoSzjXcL3myufHue
XRp1nYGIJYwpCPJz68E7dWuoclBRGnP9VUJ/coUHqkt/LLqeC7eQ3sZxvOKcHQP3px09MNIh2sJn
nhDy86waTX6plF2Ypn3AUm7jE4q8SPieEorwrzTFZ+6ON1ETZQoItWtpp6qhJ4Lcq6suZ3SJCxcP
mf31ZneSNjvcaga8n9RmiQdafNq1DfOvWq4XJuHr0wfNeS9WDhnXoVVid8GJXNnEXxR150myhGFN
er63ZzLnjcRdvtMJNQCNC4ENULon40nfO+4P2FOkipT6MCJFZaPuDxFz3yWsD311DJJzBUYJ3zjX
OPACotnVOE7eUPcg/SJABrTN/goRCxtjxcj69vZqpsjtHHFbTVD3ygT9xcd3TikRfOsVKJzsiBT3
uDEFmXK6qIQhzmrM7Pg2iFvlDzCgzRs07JAOhYULHD4cZR4sH+lv+2ttsZ/j8hoRxhpE2puab7RH
ZVAN6ybCoI+WJnQviCnAcNNifgJmervohfuMB3Nodo8vycnSST0K0miF2zgQhrhyYGtI1mQ5z18c
3UQXov2hrXppjbRUxQXuE+PJ7rA/1ozCvgeDrhU6Fw0v1+SECegKMLXEDpQBJwwxTHx+kttH8Dg0
x4HX6I7WpLgiR58rID6Bl6sFkqJWMr44gC8ACbVYFh8QyT29GPJomLSYAByBR0urGqbkXk+E+iSI
kjbnXCmtBJBK9C0ZScCgHLz7UgeuXypo5EIKp9li655BNUKx87XGDZhe6rn0nvlR0vuRihDtp8va
SJJyUr8u0iIUM7kb3XMgI5GDR7ZXDJBZX2njnQHE9AB+Hj9xs3uhCHRK/kdZAqNJ56hhJWH0ySnM
AWBLq5Y0tVRGcA6foZWTmXmH8/hCoEen3wR+KcuFjlLH2MRsRZ1QeHNxTYkoypQHtUB/X0r88L+N
SA6fXbtOPNOU5+woRH1PbI4qSUmrBznlqAzYECmhCpaxPLgnv5DeQxOQ96oy1OcF9tzyGsDxcDtH
ahZooYNBYHxVU6PQR9FoaEYE5Z7gj7tq81UuRqG3WrXDOYhzi1leGrQfPMU6jKzTcykeegritde2
Ul94vwKrrdnUNLMFQkchlDi6+BcThr41yCQUpWbU5oqtdVwFQLbNiDbpphCMT0AvZM2i/1dEQtRD
1DrXmEHTVBRn6kiflMh4yOtG70YHB/18RY/mCsKda5gn42KdB736xjeuRV8p/udsUeBDyfRWu1y1
K3pCU69yFZvGIUeAFcM0uVEk1ha5mGG/vjOura/g9AoA0MSF6jX+L8sP9DWw7DQhUsPLei5bFUek
u+JuQpnIJgh+A6v/rEyEM5yPg082d5Mca1+2SJDK36vbgLlmoPbK2vAGoZx8uFggsq8JrySNcDN3
Vbz9Aq7K4RwO2A55L6K/w06X1IIO2ic4kTLAAZVGCIDfxFJlgcT9NmM92idCQcxeid0Lcu65OYlU
JCM2ObhteQDMDEWH8IsOb4e3Hm9cgOFpetLFWUQtex/icewf09Ax8zolAnx7vdst/JLlXGUCKXac
eDXocxkOvsc06idLcEUYqxM01orDI4LQAQRto4hjJGSG2Y6UvtMdVfRZj3/RvZEebN4Xlj5rD8PP
+Zcvvk2WURwv9AMJw7emT05Y7N59aOhtAzFIw7/jo561MljqtnOdq28Pj9OjKm8ymQkY5ge263f7
mLeFXc/i0atq5mNshmokdKtaie9UHMhJxWari5677qTOTd43gePEEwuxaAbkYxXzwncPuwQZwe+I
IP4L2y63O3z03u0AItyvE9TWjKscFvICmM52UsWLfDyvP6AAfJbsCQ34eJyO/YPnRJYO5zc8RdpX
7Cc7/6u9dAIYuvodtI5JktWmDzC7t+l0qGQjuXTidT0CfkGP+/dqI6oir1WsHayP/cqVIWduJNic
lZJSXoGTMDbboXwvSuSquc5jnZcZAzZlaWnuAUgjj4kDKxUFeg64S5U+LCH0c87aDZlTaCK5M172
OhwZrpdvFS80pEsKkMbWHW3QHfWgYk9aDdjoFd1UKZU4ADI6QvMGYnlP3hYzOY5LaGmHcc0fDkVN
wOBK1vD/W+Mf/EJZ8DYc0xSZzPEo0/+pGySRP43mGPnswxdncz7GPwEGrDW51F8jVJ61Sk1WltDJ
Ku3BM1vMU14wfM+bpLMIbVywCdiDJhPR7sDhXvJuh4OtUF9dPMn6mTp+MpYovPxJheOkG4r5ALrq
fo7GaC55cc4VMUpcHkTOLdXbc950AUKeGqecO7avu0Yyl9/iXg4ZDev/cVI5SUHCieJdaur0xiy9
mXB1+9BqQ++8qvCg2HkWLnIsFuZ6xz7XtGj3nowOt9DMeWh8VWfw5oVSvvGXyB5VuRs0uFsn8wtL
4WUu0XFZvJYMVtQihvcXUOACZRX+urJKbvFDIiqWWM6qd78IU6poYYrd7MFSpxLM5+V7WozBIc2o
Hs3ZtYgMxYtQcxbD9Sv7n+Wgei0nTJIpp5JNCq2ITj+v49FgrGpLNMufRmwGTOQZLqNfLAF/Q3Yy
L1N2bFUUmmBueQ8qAnEoR2pCqmVxakQJpRIwSElie97T8JK9mrlIuTR83KxrF0eBFat3iisxExCJ
BKM+45DsaeQRfl63JCB3odPQPI5AWwnJug8Q0DKCU2dqLA2FVhcun9kD3yM5KaQBV2KUKLA/DkHA
G+6PivrHYXn8NkOOp1bVR/e3the3IaigBzncbrJDAHC27OivNbRCmEZbYzagLdNc6cgYxONoucFz
zyymQl6ydYcqP6Il6XQZMc6Ptq0bSSH5YooMstNCQKqySgprQjQiWipiIaixdlM6A+aWcpVGoSlC
zhKr8Cbyx+j7LbQ9fPmhVk59ZSpLVUqKeYBnOtwFZqmNCRR1FdRHbVUIPRAbstyjkNX5cefnX0Ew
hoN2DptpTXtDAJFPAqah3ly+79UjXdVknMgrIyrQj2eNjmqqgmwxJJKdkPgH8Aq1HWHoEt2dHG4i
DpIgbJ/6mz9wdGVGrB0745uZZbRTJVESqLjyha4tAAWDk8Bm93DPcNK/FCn0p3JivxqmBxOEAwHb
9aSYLX1qcmAn2/kE18CxUN0Av4PHHv9brphjDPDMIbEiZopjgJY9W6hvg3dja1EDLggAsNpzwTem
xNCzFof7cKXD5cpQ7QOVfjMcRdo8e8LVJ+s5nd/gn1r+761zVQfP5LH8HfTu9VAcMN5N7Sp40GpQ
ucMJihDYOtohsFU4nYs9khu6FLTych6ogEkC3+jRWT62QKCy3bplAqS9l2nhNouWpP4LCLzp8KNr
p79j/0eEQQVjAbVFSYBM/hWV4jdEYEK2nLYzBvYQEhL2+h5j7hL2rAWcTnFGWJOr2iMecDqyMNtF
VXXLJ3BBEpfbFoH0kv9nLim+HkUDbSyjfvQExgGEa2UxNeJeCwDOHaugKgakFo4M5ip1kXjiSaYC
XBARuAamSOlDx30zrNfN1y9soG3HAyfm1p131q8jiY/Q0ZCcHFtryXXl6dTlbT5g+vQZvGCa5oDS
/6pyQh8mtZKsJIDIPmyt5Slhr5yMXIER0+4Iysxm3b9h649tyURV0gs/MY7SGdvBJaDm6CYn9CWH
+fc7ITbm+iN6UoE0fEyjZJpU5au0KtmFDGsWy6TiAvqN89emgzv/XxTyjkuerDoPQsS95VCiaxuo
5PP28bHRoiMNInU9j6VKQOo8AyYPx9OR/lRrhIScTCsEzJL5ir6UTW9pLltHrQX9APGSEiv/hHq8
MrAqa9LfJ3yFYJrF00QQEnERU4jtyXHwOuc/+PZGG52VOnXT9qmU3PiWuSShPccLQcPn1XpADlGk
baKBjtpl1g4rIQI3PKh1WPrUEWA0xKseeeLBjrmjhdBhpZJPVl+Z9Wo9J7ts0ny5xWUR2Bfv2U6q
9Bw//pKP3E1YFfv2KWDU6985nKKa5J0M0Z0jOWPVR8EfxAvLs1JTMXfK1cRtywbkwD4sg8lGvI68
gDHO1tWpIrr5ruebvpDlgssGoMaiKOzmsI71YGgPPQcv9E2nbX7OzeG9ITVvzV2WzU+q5ES9yuu5
asnizDBpc1Q7XtiwDZE5quWZlH7c/Ne4W2RxjHEgrjiq36zSS9J/OpCeVP9VyE2ptow5igcxOkBv
IFc1sfhrkf5b6Uik16rxRgza533/j9SaDOuMAbrrcgtwIPWniZb/LHxis3mtXBP6WIH/wVSUS3y/
TM5IhusXNyhfL+B2RInAygo1lsLYm9XAaFuWwmGk1Jt7/h5pWPVU0cpa3eA0ef9FreBgso2duLUE
NueqDsr3loGNv+oawrL/KngrSgbxq689rXfV0u0A3KUQH6jHFRfELkIRM1rBvlVxywun5vgOWvKc
MsiCyXGFqmjRldEzc6DDl2FeqPeql7XXWITIbENc40eN6pDJnUOkGNhDBJbHVX0Os4Y6ogtI34yr
WsoPALtlzX3s1mhdtK3avqjhcIUn+011pmjnE5afHVXUG66ewXWKSW23Jmbai7rl5ybSJPMpkkMS
QRolkaLwz3syW8yWpS+w/eChHnSt7CnFBmBc8N0YsNUg0GcqgL259T+sxb+KbU9n1h2LAo+dIhKj
8c9zvr7MiKj7b46g/b39kAdzS1RKR6vqKuOwe3vy81YwrlkwhOvcLxX8ZZgfR26aJ+ErSsrF55rM
xWUmIP5Gkt1s7DZQqVCZEK2djYjD/cMKLiUFUp+yWu0Ia4RsH5qEDZ2ZBW6v5IduK8acm3W5vPAw
y+7eu/h+F5UuHUJY6vhChIXR3NX0S0bdnzHm4tACYyImT2VVOo4SlvBXV4Q6Y2S+ZwSqFfBqF5CA
KV3Y7POxOXmoP0o8oLmvQu494Esk4MVNECtUrvTNWYSnbVl95IADa90Q1b6L/iaWjjgaMjWfxVQg
ItdXJXNchBxQBl/Tn4UmrOX6VJfkiSG77H8C/15T18e0hG5CQlRzzNGWxutEgXcEf8y3hmAGLtl6
FtMszvIY+RSVuNZ8Y54xbZV579T646L/riPYBcP8iSJBG5PL0vGFq22pnu/v75Atdp5nHjl2SOW7
8vtcC0gTww2bLVWrfkj6q7UJqo9nkjMPEnYZSXKaf2krpUOHBki3DZzulmH4x58mXu+X3+TxfYqr
b2VkFbTLZGDLnwTKosDM7nHMywrxVXXOL5itV7aLGwc7r9VVt0pOfrtdw2+y8+KAlur1cboXRVOj
1vlf+Wv+WtSzp4ReoQ2qkuwwuFNwHbgTdGQ3t4Qw4cI9z7U0NPepPwNTts5g88vvyloRMV8ihHOv
u/W9oD0N28FKvxCKZOU/KMP1MNdtvUHKX8AhfEc/YMZsG8lCR3RjPbG5Rkd9Bs67kNcVpI3nm4xm
08mhSboxAXnQBtPnOgBMp6cE6q63YxlHy3TxS/QIcgcIK+6PvL70pkNbBoIZKKH5c4qz8mUA2kbL
rbQxnREBm2iF6tRkmx/Zau6jZ5x82RyKFo9OWypjPV97/8x9rVuXDJ2jDArFea3ZgQVPsBBTcBuX
Bu46vbw2cATAWAW3qFZ7axEFI8wGujNelgqSIAWD8rLjQwjInzNaNM3oey8kY65IBybQW3rl/1W7
/j9NFmmzGcBHR7s+9tdCRYKHLlDjfQpe/YiP4wGS0b8StlN55hwkhGXCapSqbmzl16AP3WScKm5C
FWwjOZc0DmKEPTWjdIPvXx5hHHNMWEzeRTp0zqE/bUFlkosRdenLFXk9jvKbvNvSh8yLGWd0EqJu
gA6NHNk1s2+jhDDsZX4New84zRtwZ/1jX53Bz6Encq4RpyVG3JBBa6HxSp4Jqp9M2/eR/V1iBgwb
NzeOp1O53khmfWNg+JtqTIGvmwNoXTwPN0z2DfI3ETsqJUBgSXr5mJdoslq4wWuMa1eIuk1WabfA
yk3nx8+afKOgBvPgJ/AapOXAmVPg8wmvl8zy0uoZ99UydXwMsEua+A5qfi00WfoGGgeL8J38kPYb
NsnO+ms8J39dHttfq3+ZaHPuZrttCcrhDfvrYBTA6CKnxs6caPfOjgkwMi07Cr9YtxukIcqZqyc+
/lWuh6Ednr/7Zlzi0Kk25I1pZVU7vbZANP552TSw7pZYCbFB3VZQxyyxvZ2IHgt+Ih6DkevZD5lj
TrknFCeHa3IWWN+k2T1v4+jWsJo2cYTo3/r34AXdRU3Pum+Yv4iW7zBZ2gmZKoxCgW4+YoE2sRVS
q4bvUeeI7ViY75zmg0G/N2JzbeRxJbfuihA1p4R7Wku/HUiS4hNPqkmAuLwnzWdY87M3THeOx6iA
WFOff+pTcKSB9CW6yvCSJHmc7tMXbfIiQwzdsW1/1wYrVYxX3T5F1DUhl+OJehawuXw8QG7czG9a
KWaHuPkztfw+hxtIV7p2DM5BR4JV8OeuTL9P3mlmdna33eWZbWpA0JMo7SBwsvr4ugntzKPj/chc
+++5ZpyXwZfqn6xPJ8VzZUPTJqPCW3EXzlHoMwBOq9kzM0MQ3PLqCFPOzRyHq4lUF5DMp7rmltix
TGNT6hB+897tw31VIjxEsqLdGtPvYfZSkT/NZM9XODAzKB2QuRQ40/YAHLD1BlyBtH+1Jqr3V3Ww
chNfIgihuqZx+ORQifno9TSupUed060CUNENO80YcMwkzxpAICiRoDe3OyTEmSZFAjsFn6wntw8g
wTL3QJ09PzSnwQ301WKn4Ea9Uq6W0zlvIjbUrj/OwQul2pGaiJuFl1u+jEzOS/UuIsIXe7+iHGpY
8c1JiEeEDpsWla7Rf74FX2QtHPoY3Ma2oJwEOlhBXueVC0K6Pw0biT0ZEdPpxej5GEMNfTPp/Wu5
QjuDGjcmGDV/PZ0f2aX0EoxJ98zgTRtZqjk2DIzUxacP7kB85wKobMWHOJc/iBMBoiAvUtymXlHt
Xy1CuFznWZogSTkqkmw2feB841q8VPiKxkZnMFzPa3NODMDhv/b+lXOfbF/WeAzAoyXilMu9vntw
u/vBEnpdNYmPJ9Td21cRHuXaMtKTalpKhxni/X0Gee17qpTxBcca9hsHtls6uVFwUs2g0vCvDNnV
i8QOjxD7gLOKz6AgfNEvBvQB7dyGa0tH35esQ4f6gbfIrfgyHHA5sMc8FU6rC35CdoSKV5fLAzKV
Am9bFqBkOz0nZnMjWnUlC2XOc1L4/4iIq6GVcyoSk68gr794TlME7LByFhacsu76gY9i3yW/fzbc
YIi3UdyXC3Z04Qa1Zvflplw1aT+sDPYxwnl1x/z/9Z69pUk/uz5D/UsTEJS6QNYYVZuXCaLy58pE
+8mTTH2VM66eh/tkB9CN00MhFWH/mI4az26FJao4wDuW2EJtxLfMtBErtHMsny6hoaK+BJ/sVS4f
ADrtJPLHZiiGdrWFqtYa4O/AKZ6DZE3L8uErey+3zQGP41w/q4obCP6jgxpIA2WarWWGb2gO2tem
KKXYfDrrM9BY496DnR24khM12rXV/eXI8Gk6FKqE0Cg7c8WlWOTp7KfQRMDRIwY/a3XpK7BMpfws
yC40zVTqK1i5ilgGXECzkIOkRwhiYlXIRGZ0O6UYiPgjWoJgDHsmxV7UArOSD7LbZMb9xdPkQL4u
7d9/Oi6u3WJcwQ0bNymLo7ecEP5fqNccGYNukDPgB6SDwBpFJn1ft7vEF37VvPgTPncTgjrWVRa9
pDaDS6qPlEtfk2doymWvrRwvoHpJC8pckMQzgPKRbrCsBMVkMDlEGRT7F3QvbQ2EjUiWKpo9EjES
m5shDq+e2PTuQbhLnVB5jw5ADCav0KiKMOcvNdDu9hql0WZKdjUNznRmuhY55UOy5iXiyjrG04+H
8j9NtENyEAy4OIWXfyicRBNc24lfuyiR3Pp90woXr1Hp8zXD6CxmYQh3tUp4HSRE9B62Y6HS/0xZ
FvyrjM2dMmfIBp+YcJj5MZVeCOa+S3LV61R7Q2QmSoTxf3QaajBgKXM0Zt6TFhUlfrPJITz360qD
juuU4ToS0AhdaGqLsyUqX52lOnA1sQpgr3h4FCp4Sxa/5zT+UvjjC99Wba/AOkvdYgnb4PL93NHj
w9zBD6QrMWArd842qu49xROCledczkm7vaBL3jj8pmqw8cHWOAHC8X9QqNgP3jroeJJAZdCuN4ZK
ieab46OPZ2SVHo04fO6nwuu8LWmemAI1omtpKG+23H925Ts6lzKnDzNB0I9GZFJIB3B6IBQN64sC
YfgK966BbY2vZZw7AQd71vAAcISo9GqQB8n5JH/nWM5KDyNaIsyf9804aLshdti0MzPg08fD4jei
XV5zRLKuwu+xjfooAwp35pnLBk3MiQHCGEg84ECUAreAITugpgiUBIoyGmdoYakXWGD/uuJMXFSU
1JsZBkaKuEWqZeyOhpSwS8woI8f/BB9+vWVD53HujiIUheBdObU0Rvc9sTvR9IzWSv2lf06Xkn59
LCPf7JkVsyQCF45mCslVTcMHHJo5V23Zef6Mrghg1OzwSoKoywUpRwZBlZXftjvLGzXUoCa4Wx2F
mr7Hmd3nhGh6+aY59C0VWp3KnpTQlsV3TM+FLHzcrpweVSrOcIJyb37DQkkjc9JjpCa/OA7IYQn7
wfuZsJ0mEvl8wlQkNB8/UiJs5xFh5+LLROvsPfEsND0S2/VvSv197kxdHA7MGF/vbag99C2K7f6C
mECSzTS1qJepnE/nyGyAEjSgIrx4Dw83Dz1VkIhQPQ8xSTmIko7pebCayGjK0nsxfBbesF8SUWZp
5J9XgOblHHYgxXeuvsDYMykvJdB6oJBdY/jJSgAAezIlKh13lLZsTynhmJ9oYrfWHlINT7gaxS2B
L0QG0Z6lti3gVQJPh/XJf8SPak4s7pdW+ou0QBhORf8Fb9OEvCeHQP78PsshTtcJiDML0W+2Npqe
IZb79CR3Cgw9Gcq1E5TU3jQsy284JPYONp8qHpXrZWt+sO820HBgOGHxwkFdwRD4OP50j6Kmt+xF
JPiFoUiP+MvvJPuhb37G81u+dUMDUYIxj7WO0L5C3iqUiNV4a/QzlS7BuFDC9Mk1VWY0uBCwUJ8y
l0oV905h4w0IqMPzgz3/YesoO05HFUgoQ0JCooc9Hh/X+L8JY9mcT+e9E0Koyn3AUKv0RS2Lnf7K
prtOsogYeEeidQVaEqX41WsXnczmNzrHXdmoUeqvh3A0Hy+IkK3eDL3qO6E6TddnXU/eHspYWi+/
eElUYOU0WtVpZaB1en4R7mwORlwDA+siQvkRGz5XgkKmaSgdMrXgX6S3nqCbIfjjXwwvSdY6N6Jd
zEEga0Gu3x/ecctap80iOCB5wqXaBFeB1oJxVhf7wc4vbjP7ahFPe3urVnHTy9+nQ4M7u3VjT/qw
1N/tso5Q+boNvbkKbAIdO7WhfuzheWgxqe+zFp1RxvWIUkWGJMqqKRkQZcO3HhXxfRzZ/XdDqltq
3cpbwIibMRXTBwbgVqHKBaAkqIBMU/s94VWqEwGMjqTwf1Y/EA1PLgS0IIYInY1Kz7tE1ai6rcgR
P9K/jCvQie4u3c9DMb1S3V56kKGO6KpeorqNMDKns34PnIK5Y4nV02FRTaSsvCpctvQpGgs56lDY
c1sjsWkulLdb3/Ede7ps8yc/X/TmkZcKRNRYj/JTm7WcLp/WGLe7LwpJqKRufZDJjUW4xja6L3KN
cdHaSDMBsw/gffLyB/QyQXwhe3CjUNLcogDuTZF4oOcEQd6fYcHl9xbxTft8Ba2894yYYXrC1WAX
P0kuNGKVBwmHSlQ+ZccJwr3i9FVEXpD15iAiVXCbMmX0ORH6UchJULzkNtM/3E0pnxozEUbwkwvr
vx2Fc0iDaQKgM2GQ2hHTJExQbzO4amrYjPJM6+Ah+Jbs+LnVHG6sL1OHiGJiS/29WlPeS3SIOs50
oDDziZI5yREY9lJQbFqusD1VkOc5C/0dsDZt60L768gyAWLMgixtuVuugujqkJa3HJI5AzOWRJ3j
0OkoMH/aZbE+1c1eTunGRlOU1z5HBQsN/BfQD5ONj/BIiUYUIUfaJvkzUvJV/3Yj+FYe0u4lVtK3
buIWmY9qWE64G6sQaZjcdpMnCpoRT8EInjUCBgIp+FuGyRVk0kuKPIy6M3YtUFeSg/tZWui5g1kM
Kr22DmqcwvqFCKlV1grvFE2YkzkqODGFy9VR75MfwSbEMMz7MgxoIlc9dsIJinrM9xpRkTjClqLn
dWXGp4OrKO3jkVCLycCfEihxNLrMo/uiwFn7kCALtoMry8IBVsyycZU1tSRvugaLpfxuSdLTsmtW
u7K8EQVC71NZJhBE+eKJSgCsUTAjR54iJpN39DJUMc+HzcI5cs/sAeVpEHkZD1WpMrI5B4Kny2wC
lZaFxdqMwYhBr3LJYNujAYaoJaP3/h6cbnPbR9MVCqa0f6xsWh7ljntf9M9j5Kwzvh/2Ipx92dwA
DbgAzPBUvOGM+zQTXlFWsG0fMWBNcTwEVlrOp8HcgANtkvpSFhUuoU5jCru/BURm9jSrfe+V9hDi
xW7tOh2xHq4wIuXsEuCt9pUBy7jhvJlysKxHd+fYnqW0AeYcMHFbCMCEfwveWj3+MGqrRrZvo7/X
JwSQi50D4Z9NHaFqcsJ4Mzzvqba0k5LaEP768mdHVHKfEgFppe+V68vgUwxE2D9uBEQ+mh1Z6TmY
UzTVpXDRU9HyrlTqVhgbmmyX7/nYa1E1aT+RPJiIU51iLseoB5KMG/vs80s19+nRKzvjUcQSoXJZ
J1JRkJPYRMN2rwLi/2AdhVN4fTyPNJ75ppf+ucgp33yaRx9N4A/zw08fR8MRfGBaOyax2CYNOAB1
Z0WzZk5wwX1JuU7+2vtHNB5uOFYIMlWXPdHOHgiYw6kNnyqOyPtR6L3J8/+tpBKeA0bKn+qBD1Te
7A6suIqCLTJPJDXksCoKkqpzD2gQ3AWk2UHqa8m7Qh57c9yZIYxvhdnwkbJeZUjFNNq4cIW/vs5r
2XkGaF75uf//UzVJI+BPW0AXmJT+NuoEPVzKxecoQfMEPox2nlUHH7Wu8fxEghXwq9z0rvCGRxjU
aa5EkESwlMS2vFkU2GXYy7goEPifgMWwdNRZN7Do+IQiG9Zb/FFrjLVO++2YENJP4XnRi/TG+Wzt
jSwpn6Hmdym5/RHoBsiM6qUqh6BnNRjbIofQ34NQ7ZJhn8ogHplLp6Hui/slKdVxK+OnNB8ZgyBf
+ZhcPLRZ5TqPJawh5obeoSbmGpy8ADsO8firrKJlUlc5ozl3pTFKGLBwvOrW0tPswPXh+tLu7+Uj
GH5DuDV9UbSxFZGDpB/CF0HfFD8fUHc25f3WdQOJVLu5WD7zPDwPsM2h2hDrnZCysKCtVzZBR3z6
hz+jc9jwNC5PzCj9Qk+E9w/c8rpXnTRG6VNg1ILT0UQ+WxaOeLkTASQJsQfIzCbHB0oeEylNrMFG
asTTO8pKDGVmrnBxshQU3cFLcKJ7VD1tSJispYNA/C20Kqa3Aj3XuyLMXx3vNyXZy3F3ZM6PbZ+C
xBZ6zonBZJOhimL8QLitznQ1cv7qYkDggt9DHmRxDEwRmBz7krPaurNQTP1/ewKVvBtCLvqzqKv2
ApOoB7ct23xyC72fTrf46rtZAgLG6B1viKGEUUQvB7dYEk9Y5UbJGEA0Jt3id5OS3BYkPrCr96xF
NH6ux9k6c9vvCMP+OttUWkMvTrmHHg1OWujP6k186uxMA+R4sFZY/uNB+RbLyT7mf0ald9XTrcSW
kITaAOPZA6cXjI4U9UUT+RnFFIXpD8AXpbMZ2yoGjRnuzO9e4eIRDgkr2qHPz/viSzvvpeqJld0r
Tx+xyTjr2vuMA1MbxQYb2uMFB2cX4CEsuerqcC/jd5dWXrx2lOfHRkX7zXAKrE/BAwDIsNzF3zhA
ES49TnvkbXwu6ery22//PyGXk3HYNnUFV6gt2qt1tWi3voAt+rsnzGnzPxQVvhkGGdL3RAyTdCVz
AUa1VcNWYRkT7kWeF0VrWOwED4y5FGNUMB87F6uL0k55B2sdxuX24IOgMrl6Q4vPQtxvur92j1Jr
jd0zqciW2GE8DcDbM9JbFJrl2m6YbYW0tS5uuN3wsubHe7mRbaEThaP1lveeK4tgVOTn5ZZojrgF
ggjQVBu7R6uEyUsnwJiRb+4qIRQZJK6osxv0v90F9xdkIXH9+P/8f94ym0Veg6tcQO11R/jzf1Wm
Wv4I8vaQGdL9fMfkYOchyCvDcNT/Wo8fAvG1EWLhn3JyMNQqwnRnE4Ntnqkdd574bmpaQhhFu1jh
i01W+TNEVvppgBdv/kvuZ0lONtAFNbTUja0Gw7w/AeVXCf/1fbzasTPyqbhZp99P91Yv0an1yoH3
BkdKvp/A/htLVylL9kGvK/HqoX9mc/pQ6pUkYHAjO2hS4MSVYfz86Sri/dGCRIHrDtdwjCzhlzDc
BgjPENpyvMl2l0yr4/hGar13f4scVtJB1TCfSN2ScYf1SzClwXaetjkfZBJ190K34liK8MavYJiI
Nv4dMBvHIAcONi3muE0gpUA68osi/mO22gRrA1IfnytW3/V2EoFKY7Q8BjISPFh3oCJjN+4vMSm4
XNFpZydzTg7cOwW0UkDLU7cZc1y5AExsfDChYjI4mZ7GtmS6ZY4MPzLRKVHCBZJJCptj3LHy/Q52
cRc/0xwig0nbdvyA3X0xeQ96TYT45ADpMzzGUdgwQkEQuzgfRF3egLNxL2h7wyKgYZ3Z6QSDgpKA
FgwqkvBNG2NR3fL6Afv2sUtiagZNiylgZa5gCCNCMu3BDugoyazjmBEbMQmjo+JKq4dVUp3zJ+CX
B98B/gAWCrWa+KR/e74mIFtAX0oZwBlrsmIGt49pzOO1h1VUuNCWfpyXaudWDWjX7OQfIEl/jA8t
VIc0/pAmaL1QHFrZZnw4BrmEizdK+sGz67H9npxN72QhdIlWSgDKbM98wnff+nsOvQh4R2fJkaG9
XOQB8t7aE6binaA5/51H+g5zpZMgVQmu/wTzMr8X0+Q89Usfy6E+6xEjjoTo8lWZ5xcQObG4S1xO
PlGf8oOyY4c8WvUJtThzUGJLqFlZUsZs4WmsJ9x1LtSG5y0CCcKES0HOr4b4q1jvhiOOUhRzoiRc
mVZzs9WI21scv8dbcE38K1ZlrfSc0+Ru07IcYgQyuNTQgUjwEORNpPyn1BwBKws7Nwvbo4ItJKMt
XYMpYtdV9TPrg1mZm3u/pIuk56K1z207IUFPVMJxThsRc/rbUI2s/Nv4fh9MqU+4n3Hswy5PbUJt
0BPQ3nYh/bhmfV7ooQMKFBSC8zDNNQRDuuFVNOf0TjcNnds1cP1XuwO1Od7IYsuKv9l/axwFw/Ob
tCzjUqCNuWwfR7LP+qJrwQc9Ce1uP9jHu4lEeB+hPtZYuPzpIOA0ren9iRCn0y0PyO63cLXgiPcC
QM67xWuRl44aVyG2HooP43RjH1obQK6Sw1STtcjCqLT/u2xkelbfelxR+zwQD1M2rYFE1KF68VFG
P+IhjcKVguf5lpbcqxGBfw9RGNGObvVuDF5mThDJzjK3McsbQ59D3g4s/eNVK+Dipz5thU/mGXsa
PeppNVkmh9Ouo/PtA29xUe/wUXXyQbQ6Y7UIfjFN3i1H5mLE9OYZy/hjoMagnpElwnWbHXzM0JPh
ZEqNrmirJj0OLvdgLsEmMfeRTlmhm7nFL7G2T1sqLoArumkFksmKyUd/rJ5cfHNtXkhLw2RRhmQ5
5aO3GE8qqgLYRMs1ZChgZe0cOxlJaDeC1aKSIFjRvipUMMbVukpLvQzCXvQn/uWG6fryitVyjH0X
vjp8p6prTEgTaRIQxcQeIot5N/6hDCzrbEhs5AcUrWnmTQeIT0BehVEsZXnpu3+TUtcPuCZlMOY9
36r2N/3SH0awPIaGbFRBzACpY5Z3hslXq3DQvwy/04Ct3tUT245nrLW6W1DlQ89woJ1yF8UxNIYy
3ob1NkHQ0vXaCaUZ3b9/3mcv897nP0RhCAKIfCamuvGA0fitNKXr33D36PxjZk+PnYkomIS3/G+l
LSKpjRGhCvTCtVKTItB8IOp0X0aci0Y96pvh8sICGCam0llWoINrFtXyPbkxPqyQ62Uufn1Mxpdr
ldkLn9/EOwC+ymauDAEOJKGbaXspeCZ+10rnr4DJG05+5nLznAknQqxp/eR1/sVAYzhbZ6f6nucm
Ilvh021E/AlU0vfmHgqtrj1r+y2FUN0+6DxsIY65rPKfrz8dTS6lDWSHZmQVT5+Bd0emE8yoTvqz
po97h8nHuuoMpMpVJM8opnuPHhAwnXUf9bCl2Ndq5KyUZ27gD7Q/ylbl89bw2FV4f4WgwZoGUeAw
UgTW1nDEpUEfYas3wckbDAF1lkJZxIaQpnPdRnuzPfaLzK7V4infZkoAEAkagHnISG4Qpn0STzOA
cEkVTMNec7pkcylCQNQxIhr1ZRHu/0OHd0Uqb5nT0RRfAp9mqRSFnV45x4wyOmdQ2lD6PCzJ5tSL
E0YIBTtCuydb5vLp+KnT1l+DJMVo6h0yFGVcE32cyE82VZMmC6nYYxmbgoPTl98fQs8n9jY4L7U2
enY90uVfjTR03ks+PW+il/gPmsys+XioBMy9sJN/0yhucqx45lEGnmFo2MIHs073zM2ATKhwiDAp
lsww9dOOhX0uN5KtSGE/LmW/KfTEPTGgqV+UADYQbJl1pSyP3wcnIw7Utzh1qNLEEdPOZi2o7nfO
3fnLQ/m0e8EY+xEsCOPnaLpnm0sho313401cY8swdOU5f0+qS59vYSozTBiKs7ZlFbUwbbDrzd1N
hhgY8uBUaUTi4Ru0iuqRu4qUazFaGDoqmZZMzpvBDBFxVOJUzwhJV7y+BYrO9TAuDxyRCA7/Nz7/
fXQxsDNEJ/saGackiL/AAH0R4r094bd+jSf8NdKNrIdbyfxxAvQYlda4O7tpJ2fva5gkUXTfrqYG
IpU2lE4ncUdZWSt/hUHWg6yfbTfazFuWr8lPn9xWTZnTTthJkenwUfETQpXqXnSSdstKk1Tpu5oT
mLcLtz9RUa7ILTExqPYJ4K8WIXFmnXfU0UiwZQrWRgvlO4Lyp/TLKyJDmwnwh1pxfUW6bMmjr3yQ
kwWxmxlBHFcxoOKMPY8ZAWWkiU01pt4uYJlbzXo8L1CC5Hw3h9i9T41BK53y8PSFTrQqkDnJlHkn
vjs8BTOoo15rdPUDfm5EeulN+2H8XuDAdZRMsYe4POq54SphjaZzDDIujDMxaxzVr16l8Elfmebw
2IrjOVoV3wVRau/MbhGh5Nc3l0wP6jJBKieHiw+q34k0HTVxEFIzcCQRMkf7WLs+89kmUqHQylOO
mhOfmOGGT7et1rIBb9EOvdWXpCSlxodYTi6W0FwRkbUVIz0GcsSzoQS6x1GDXzlCI/8+91MYovqd
M7wn+cXm8dQ+KJpj5OzBcJmXB8P0zbEXNRYnvOFPFxJp5lPS1T91W0eVBGnWZlJR/8Bnn0UQqZBU
RNeRKIcaAZrp9jSTeHIKtDY9GKHvdM2+zwOm/Zat+EMvuEyvaPddq7CQ8NbPmGtWbVXwYkRsOsEd
noewiFlUWMqD9YBawLq57Q45wFU3Hqi1fdyD/lkyVeA6ObsgZPkzEdE7i0g+mWQQWfPkRtbRxH+F
nCXAaFsAn4w1nSZEeSKEPtJLo3pNzJB3B03rrnOS2JESAfsHK6QWQhSEcIGe2nLQukvBcBP/z/Ks
c87/uymhV30yuZScMK7MnEaCfAiVlwJ5pmgRwRtTcBzLrTPD5wwYuD6U+kxdrYODn5wD0zxe/NPM
JTuZw+NTSDpOVWYyNOKtbFwewhnnRQUR7UfdpF3Xsoz542+JUPTMLlROFVeY6y3jM34jP4QxRywa
nYBZhQUqwBM4wGgVbuNE0ZFWNp/77uAqRlTUxlCuL0H3wmeVfDZSFTuVzebJsqscb14oMb5uIfIn
/pQ2odzeI3KrzbRcMlg7NZmJhnvNrHQw0NLnm+cE8l0Bp7XAhuDnOkz8AdB+pUPmDu6JMIWYwEc6
Fnh5iIdw6Fx93VvzwIPyDHRHOAmPGzgp2u/CUzBsVWUXsZDgzymZZLCkHcqY+GVGF43CM0+syGgM
aHgTpzBx4QidYA7xGMQYXMJeGmg3qZRVdeclgk1HXVebnZWn/uEVDY4TpK7am8ppV8jtTeJhF7GL
Dfsv5XMQi/vRBaZGCcseq421HT4Ij+ZLIifwNHhajC/Ci7jSSJbB0lg1QjemF8a4zwlaXWptv/XT
Kx+12Rmbz1Oht84AoKQT0/BYBJacQJah/XBRX6w1GtsgDn8R2hg4TxH+c2l4YlEs89KhIukB5n8x
e/orB/vG7o262KeDZ38qycwrdloSxmhRVvEp4FfKpRvZOKgHYXXIe4NHbw21/Mfc5opEgtQXUJiS
lZKrmpjaB7F5+zQVbWULMz9XnNEwjaa7hys0l2vDSl58nFL3SkCUX6g1OSaww6N/Fa2jAuHjJ1bJ
9+eTBpoQBAjMIyiLz+ENV6zBhjDRsUKb1r/QlFOlFQbg5lP7dC8EHOcSGygDwwNJY1R4Mje+VOJK
MBAjUgthFgbF3HsVaY9mUI0eJt1Tn2KJDXPwSMeoLbWMkzd0sHwG0KkA6/Y27lPoi4m9XNC8/Vle
RQmyv92tnv0t9CTfLycaXtiw1EAMuMZ5E96fBB+A5d6tXSg07Ga9W2aCE7BV4ntlo8JupBKnI2/4
nZMbqvFzUloO9X1YqQCkYhl48W9yZsM5ZyLsq7z+MCgvfbRHb+4rOvFl64QdzKRxgvPhABTi43OQ
K0EH3MOLUTDjaq6pZaWg8oV/NE1305974v73J0+YE6KolMHY2oNpbhw7Bt4tjdt4rhbGlHKtNwZo
jbOL+Py9NkAyjGmVkt1oHnTe8J81D/srSsbN5/7uG5JfUI8lxsyUaX1qvbjxyItoYXEH8QLTzU08
vzF7MWD0oAR0MVsmmSWJLgZB3msT7fAjipSt7xD2fH2QFns6zhJgLLtCaUra8nmVZBtfpsrekl3h
s+dJ8Xf3ZLHXk7hnnAXNGimyptUek2NI8zBOrLxNZDGwmLFQzVeOtwUiFV/kHkeflwcMc6C+ILTp
LX/MszY/X0NY//+xBpbukGboY3KhW/xcXvZDzR6PTyw+KLvYiiA7YgvP19z+lsg1X/+yqON+fSsp
eF8NeO643cfyHDT8yM/A+C4733TAnYHI1umguOafq8R4TwDwH40LZObbunX0kCLyOemcmnvHHNZH
xXtg5HG+WcWCegP9FvHXnkh7VnG6+qWBM0KC/J3q+Kj6wtWn6SBalMccLtX2ZfbAff0tMLVQ5/uk
KSEDNCKvJYKwvIYRxzabV1LaoSWIiyXXc9XoyoDlmPtUTey3D913fp1U+a89MFdYPuqL7l8TjT+K
m0t8k/mXicbm7QrgPsfQOk01TVSzaqbnJQJXRaxQbRIYBbhkf40+mx2QdWs1AtmhIa7ZCZZQcXvm
NHg8COA6+aPwPYFSQT9DScBgeTWl29rOUjEpX7NOB0LTcR0CUt7Ve/KYvvaq3qtZ7opmYQ5rUTNO
fdelAzTTmj3A0VmOH1xBlWAuozrnVRT0SVDQvQeFibfhslC/HluHwGYN4r2TBkorqTOFnCloNY3I
+4no0G5Y0WTETm9rUvPjSuWJTJzeD0H6rv5eogsl5k76cgZNi1XvphHh4oacsifTKrNaN+IL4/rX
0LT/0+w1pPFTe0DglGkM6USwP27mj7GiQ7p/qomyRXJ3OQ2QQ98luVBT7dTWa50WgXIF/AQrxevK
cnySZsrCg0WA34ScVZCsagZxitcKfAnh0/x7NziG1S8PQEikTXRfU3vDwY5PUO+vyUKtIKas4KnV
Snf1HJjEMwaFAEOYG71ErZMhtxsf3QnsmwP3+oKuLDpnc0g/Kh17I21JjefKA5okUO7ME5ACuDJr
PoaDKy+T7iCXNKfsw9eDy+QHfA9F3KT8GhvMs/XnD79QnHttxD/xeqtQDt2wU8DWyRVj8lm7WzqX
QmVWrX/7NqF8eOS+jtinORmYdEC5oWO5lIHe/O6If881bv/Fmb6XSSU5Efehqrx9P5BZckih1Xs6
LsoTaN7+73Ay+pepPj/cvfZu6i+A4DSe/lSKFe4zZwvw6VVdVvI6U60Q/IhcVhFzArNh244ybz+3
I5WMf3LjzSvI9jLMwBIJhJi+OG9huzO29Rw9iD8rzCt/uz7Ptx5pIVl88ZdzCaQst4pkaFMQoZDd
1GZaAW6P5ZPycXYRRPbkimEu/F7eIdlpkP4fWI9YfSYzOLH9pcd0lnjnM41ijIa6r/isXkWAbTQ+
jQNxYQ76GQVBkwPIDGuz2Dy4+tbaONA3OvdfBaPbAv920P6ZaD94muC1eek95IOiWdcH6K1uhNDz
EwWfe23ncQpExBkkImax635mCVvuVNrJLxw01swlmz2F2sKpvvpArLbLh/RXyrrBGZn1e1BKbDA6
z73Fg6nOGatSoi54EWEVLh0tUG/hvOAphnnMiRoibqPVRGBz37mtq8u9E7/L/769+frY7n4zd8VQ
GGffPKO26OA5yjU8q2twRrLhqwoZmWazE5+/YsnM8Taikygptk93jqFQw7P9dtN/YSMngm2JNSXw
sJpC10/Wp//qzR590Z7EFnkMqURW/AJ0rIf/dTGCpgSVmLVyWDzyPlxnc83Qo8aR/CdqwII6D4uu
Z9bFLY7fjBHjHbfNyvxAqCrOAcUO/kJm7EJrfYwj5UI5YkVTOIv4x3RuUni69lRuZxxAoFLWy3kw
/o+ECHt8VrjzmcJdiuuFg1UtFGABNrF7ooMMCqIimfeslu4XiOBo1+Whs206nTsxL80LgstHd/Sv
QCuLDuQJqH5lDA9xYe6C5qwse9WymFVQCTB8XZnkDzwh9Fl7QoHJc+JW0b6Y4ekRZLVlJDy0YANj
moTlmJLvUl8i3Ki8N7QiOSESBOqotntyxtTWDkJjhEyEuq7IjLi5ar2AsO5zGu21Jv4MoD8yV6hO
1hMMVqRoHccNTKzV3Vb1eyjZ/clW8lcVmXzNGZ8G8TuEFlLnDRk+8knnWb8CP0V1/5sjFjNzUoOo
22GrvI3jZIkNKtRWEKChCm3gyPRK1fjmxtBmdXPOvW4HmMPnBdZHca4XQ0PyT8jE+xJ+a5hk5DoX
+dcEZ9k9Tfd2Ldlpcr9JCDredIMUiFTil64VdXVwLRBItnfOoJ7MekA0GiFwp/wV1gr0HRcLJYzH
3IEOiUiCSO9ieNpoqmuF6wEazlZjAY6F090KYyI/2OQNhPncFZi6pgCOplMLUmE7vvicLEcudxtD
iq+J/JbSmX+tNkb55KusVhykqFzE2dL4lXlTOl//aQpjpT/4bW9OYGWpJvzt7Mj7EYGNhM9Hkud/
9MeEqzeEPXgRwjM+HRUfR9pdBXXVQgDRSpvbPtkXzuNK39/i4RkYNTjtw1TT3B2wEiRQ2xCABTpY
TwUxBW7BGGm3pnGdBeea8jsfV5Yk1d8Lnc+rpIRNZVXHibtPK1AVE2SOYv6++AbETDa4IkYRZWhQ
uMw8M1GRCnTivhifdwNtdJ2izWAHsgQjeR3GKvr61BDng1Unf5MNC43BXgLKab6k+jxpuTyVFfDz
ab0Mvod3FmqXh4htCQZTkfHbIeUJyPS58zvbb71XpW5RhTmpI0ulwGLX/eOWeNwmAnsOF/bhiZLY
94mQhULfwfadZOGAt3RPtFP+E08jDSq7TJ2FmdCU3LutqZJ64hY8J7vMkGovIulqnDaSus0vacGS
9b1iP5h5rVt941KN7uMYWReP8HFAfQTXSSdQiRxyguIeqSk/sbHHa2B9cwWBLLJEASg6ROCx58ny
T04FFIMQK4tiFTBa/29tIaVaXsi6NerdDmXqwaG1QS4v2NLi+NrxOH6r4jZ2JBQjGqa1XakNDeSp
CmQOMM8ARMIWY9Erk0GHiJwSb3la4lBt1wu+Qk1WLtmPZK/0lElvC0zjq9BzeybngHQV/4ptcD2U
LSRtSTdxVyzlsD/TEainmh/9pqWRqdVeuuPzfGCScSdxDv2OfLAnloECdrQE07Pn5xtX0xGt3+qo
NITYmyqKWZMGNyD8zD7tzHOv8cT+zh8GuW/0QMom6SkagHSf80FS+MUi/oPU6kCHi96UvCiTkGBU
jSjKQMj5S2IwThJ1EtI15RsfQu9BEQFzGnuqFkpP9f6M27C87S1yf9JtmhKfHuniucKpViEK6hDO
Bv+3xyoYdP42o5KyfUamj5VY7uz7OL2EGXj0i2APZdX2Wbp8ueVMlTD15kz5mKetutRlyQp5vJqA
4+PgRpTkOBSc4qG7ftvd16/z3DrrSeJWcmdLLqd1IyjaskBrJiWmOb3mYbMRnDOGsIjbXc7A+vpQ
6bGcc8BvvEzHw30pI5pYAMMfVRzpIE29/T6ZhOVwBDmBUxYpQzy8u058pskXY4fi6PWkvO1axjCO
6SoJyvUIgMlnnolnXo051r5xHuX/MitD4LiVmZk+tfBiWlMcOM9s2AtCWhFYOJmu8dxtyxSvzz7d
QFMrennB0AKOefq3BW9yh+2aZ+bIqCC59EN7te2HvV3YHhr0ysyBTJ/Wjxvg+FpCz/5LCpoCL4fh
opc2JDBmUDvNL6yhfQ/60HUss18p8q/VfvFw0z4gdG+9ejknc1ZqC5aEVRXsqneO3lhlbbalX8gy
ZN2/ECcnqD+mZvztQcf01W2K+qasr9bqmBF4IM7uGh4sMSMqxMRLU7fKi56xTgM2Vqln8pgbdHSQ
Fb6M4sMdn0MYJZ6kjZ22CihVtxi/JVL2pYs4wsy68yhqdawNOx4F5yLuCXU3mNWnDSfamoCPmb58
Lfg0JnVZd3VttCDk0avhUEQ4xV+ZKt/kRXR/Dm0Xi8ouQTXi2iPR7RxH/7EZ3JGZgmWcsA5rikBs
j6RU5gOa/WjURKiO/YnA44hXgToro3xQ4ynclpV9wrYJu9VsYO8LvCmj44hutV6+j41Ta54unDVB
4o2SlxLl2EQCuTrGD/Qr6x/jSR+1Vaja/Go7SGwLR+vwJ0H2NDa1g4odYBpxPU7SoLuVqFK8Ekdd
mRqnL3K14BLawfsQo0MZPerNTcOLztifjuAahXDr4Rqq6W0xMTUuhLQhzQioJ8NlSylrOJz3HAqf
boD+R5e4YBzRT0Sc6XPz57Ceem2VC9diewzZEZGR1w+VBbGrY+HXof0iGF3BsISLaVd3VpoMXIm+
rI3XxvBb3yM8D3ilvNXH9CQkRPMSRM3eT4yu9loAdNIVS+W2o+0ejeDhEmWDw0zwkbuYLdXxm2cb
SjugA2rvaRzxFcl6xgYkPUyNY6ctvm+YL4DGyb7C+OWRI+ISgUMu4wnWQRhZ4LyRreMsWyVdxRLQ
ZedzSlDb8gqes9/7lFJ6Hp5PgTICIX52GPy2rAS7LUXWJCq4m1j3bH+vMEih2SnZtmp2Do7fz2XA
+snn1Xj3SIwSDVtWPpCc2CeZEN1SD3lNckH3tu2RitC0bYUKxvDtCmbsD1mjEDwdO7HBGenAy7p3
n/aZaHkNhe6S7LSuP3gJ0YVxShAnHitwsgsiwpmpXPS7Rtb1/swVE72toT4KD0MdFnmhZclbTqRS
4FIJSCc40JKTnsoefmqf19lQDwIE3u1NfaKSvOU58yfTLje4rAQWz27k5vXnwoiebZcQ3DnDrWKD
PZ0a3WZHElRtic5gLiNXbgQNdxAAjLNhf/j7YSOyfB4KR4zqhCEfPDkRx5qHNTkTBPwLlMhaszt/
1TcgTBwP15Qz4oGgEOKwzJvJowkSpGVojl7RzGvwpQtSElxI0T69LqBLsCHLbgmo1TuOKnJjsNhH
L5myinhO/1+rTUlCLLFoKmgvDw6y/H0/BHHIc6no7g+F/1kD4EWZkQXe044WZ3+Y8vqFy2/UBEJQ
v9rHiHlQucTcgQMTSE4BpPeaILjj1Ru1pEe/yducGcSFHxk8rYfHhXSl8MXkMY+yIUbxkwV68a7J
m+C66cRB72sDZBTT49HG9mmkTay6c+xoco/5JfA1EueJE/cPgXtiNyQc61VzIUqlZW7SnmvkSSwg
RgY8bf1OrKsn2THVxTbXHdkFxK/cPTQFpEDe4F1ZZGzl0oAV9Ee6DjUS0wNqWgcLttD+i6OR5nib
ju/9eZadBsj4nddRxt9KPxKReF6O4LGIfDv4cEZkNQbKL/J0MzsY4v1Ji1ji9TZ9qQ2qPSQ8jNKs
RASTxaEIOQDfBiKzzBQ/6cXsyzA/bvt0+4A2ghQyOlPCAbnmPxU/Kpm5GPpvSmj3pqyZu2Wjbzn9
TGS/LBwvjsIpAAUS8AUpEXOr+9PaDc3obsAGm+91W+q0PPzfX74VoqVnwrrX3wMs+mgPAiot7Sus
33SeGDULL3pY3/p9gkBY40rC642Ah63zuFTL364dIkwh9ms5JPSyDrqdqvURqpj0hOlpB4kU7hq2
/NA5o6k+BzY2RxlpfwoAoPN79Fa2tqEN5LZiLc8SN8mKaZv5E2q7vwdnpjS1b+KNGBhvm3Po+hT7
n/NPPmlnfiiun/GmaZy7yKQ1od0bvtRumEzprQOdCQBbvhgtfRnOOu19Tkskdt/l0ib16aUA4N9F
SF0kg+6q44vu3r6l2inWAvyz3jHD4Un0aM2EkrcFsQ5t5Q6+kzv0fAfTrcz3nHNvjiwcVJj0Jhp2
xpL3Eg6ua9pdzt6e5GY0DruPaVsW1d+12d49Qgb+IetaNISKuZ/8P8K38V+oJK0A4ctPZaH25MZb
kagRbcWPslTR7eJi3//PA4cpBf/zZM/2UiizE9hxqpF3Eiy14BFyKbtXk1yD5z1elbhqhhz2zzJJ
YBK+Ov/dNREn8b2No/aFG0xyieADdM6kBX3MC9cH4ANM8207zZlv+QrKftjrOxKs1oMBEpZHiw74
dWzwtv92IUU2oy29kz86bcsI/yDzfSb8C0rJWHkb4TyQXdt8g+rEnO8HREnxTcuAjpCGdXnnfflu
DzH5uIHgHagNkVxSWH08AT2qvTL3/1HzuBm6hHmn/lrA52rJHK+XMAeahkOcROzg+YaiLZ8nde0Z
B4m0p+p78Py2XVe0BClJ0Tefe7GvmFM/Z/+FdCzl04QPXkmayksmGZlU0RGvYSO/ANHI34FnbqBB
TKTcHCwKOxRe+KYrwLtKM/tv8d38JhmGo6bS5zP3ATTboPAiVxSzzPPkZ6u8NwKNa4G2Jw1ysByr
W/mU5U4abzaV+FUV1mSsuUCK4rf2c2WLbLWKSItwL4IfABGsXrZhuu1TcgiiYpassUR1i1oXea+/
GOf11fJdhLhBHMXO2/zHmwrnY8N1sV+zZ/bIZvKILb1yekK5KG8JttSs+8jgJitLfTeOPCu0wvet
d0BcQNhrjE5hpPwxi1fARGcO9PNuEtnuuUwcT21JL0sR7XbKy0hdWUmrXNEtckLORoE+jij+ly4H
2X+IPc/dGx71OVMl7NPrtOiP2/K4uH03M3KGr0xga/x1t7sJEY35FhG26dSsflQdEjNGyDQXYObE
yFMMxBQ4RJzbRJ7Fs5yHBBeFnfJ+gY3jyC6wSDqrkuv8RKV1Oe9N9LfB7muSGb2+lCfVSz7p/0vu
iYl1RC1tZyNzzgVPU5KvWpcLoUXSkC9lxokHYLVOXoXSi4UEpzNjQW+aI5MDw5JMsaxgzoGv/EfT
8aQEnweXA+TwTyoWbLbWvOJbaLESAvqePxtNYZMU4DQldRPQLmHy7R/WJZFp3s4NfC0V+2F6clzz
QRPxBBHJExDTrOaja+Y/3+uplBc8qOIQHrnI/2a1qpPpkXPcAloh7YbWZ3Ej/DN9bXFiNmEL9les
2nmwNPEhCHTxulMvPbWxGjQ/IM2z00x6+pzgr/8Q6+ILKtihBF1Tv5pgtmOQiDIO15NfWi+9Quxf
6mVxX8eh9eDDn1YSxI8AmkFQsW3XUQP1UzgGg4qLLTsDqP/c28szHX6y9HyEZ1dbVqhdwsMhhGNS
hAgvQf+N6ABnIuv5OUTvVST3uwLyWAeC/hCnjV7FL3/0nJ7GBCHr+LlLczkiaMBimCjqB07cYmG8
cLvDVFJ4r4s5ZlsItmCBtGsixgJVnzinetQ95kZ8Hm/9fnU6GXFkLdDxAybopQR2LANbuqlIdUOr
5r7Qv2tlFweSc+s0jc5sQGW1z4jSIyDhSY0Q+LqyBJGicgfSQWOJoLloY/6ZOOHnejJtDpz+Ztg0
oI1JCin7WBxM9vfp4SUC+kWbXO8TsImTmdxJyqIcd1iDEIiAqLvKM2Ppeotme23ku5k0cIzIq0eP
jcs54ifSlt2sVDvU4fnVqljHvm0jNby7F8aOpG3JwBz7fmsC62EELIjNCREue0rcVV1DEBgyNYkG
CUIL66y8y9XUxcdIulJcDOo/XifkW6JrWSJpjb0TUa48KO1hq3XFTx+eCPMJ/71EIf9xm2HORnyf
Yn2ZPMfS1VSonexn+g2Zt/hxiJHPvH3W3YOhK68vNGZ5OLyrMQ5QjQDvcGMu1bA5TGPAstM/+sDC
4Ffjf4bDsZ/yZgztCu1MHNkGJOJo+WJ9biX0O1tqGeEiOIBUrSvGZDtxrkPEdEEjJIB9yvGOMxlT
yIysuEmqyFZbhFNvzPQFe//AOnA5fzmvApQepPNn9ye7dNHpoXlb7UE6UXWKkozKoQq4nS7OPQv4
RWKOXydcGg+qbq6Ck7PULJo/4AQj0E3wwIu1VmE20YTrDQaQMzejU5kqKXOO+o/8cx37wk/A2aD7
C6q+wKRjYPNN9LdSAtANDXq8UTTjUfJMood0w1WizgSJNvN9QKm/1avDcjcff0VjhT+sWzN78ePY
Mw9MACikizoGtMqhgyh0zliFiAO/yR/mL5X3j5lSuwDEgMbE08HB9ntnZgkmzkjjbO39z1Rgd1BM
vhaczn+5mwI5EmYcaNa6Yu4+xBeCbUQib5kXJ/BvZaIRk9Dmbh0LxxVCWF1j4XHmFf6p1ftLXPit
n/Y6VT9YruPJd1lMOX6TokmR/Rxwj5FeLTq5b/xsToVusCvxhUYnGw09wRaKpeSzUdNrnIEkwaOT
trtmRATl5sPoMcTRHDGclTGj0eHBelzDkRrjYooRJvGowdwEcNHZLUZ4doL4PA//OmuomCoyxMoN
RV39ILNAwj222u9ybn5P+NamIMsDN2pumulS3/JDiNbN4dNdNxX65GFobmNP0yxHKQVb8UNP5kya
3RTAgLGjgSQ2IDHvP+qDiCUncCmnfdKBHkG3B0ZfBI1hpJdgYNTclMjcVIhh4kI6UaAQGj1jaUA1
G2FJoZiTcfzIH/goe98ZbckPiWNxDIH3iOLngBV4KsBzzYLLgEMC5RFsWQUVU6FnHgnKy+uTbi3g
OVnvfx/QYbrp01Jk21U+v01agK5s3TEUj3nORmgXu0pXK+SA9WcPINwNwsy3BN310+VuhQ3s3e+Q
d5haFGEqLQErgtcdFCxeuEl4aBY0PZoKAGR0SDpp1iYNhJiYUPwZcPopQacIYJOb9yklWkjdsZLb
+6xkGEqvt6m8FWaT8EicVvLmrD6/3INxbXnHO+rHW5aZgk/kHj3xQGMzh+co6ApfgMl8hIBLEtUZ
UmJ2H72DiTD2zc1iltzJQrbR1lUPc/ZCx2qeADfIXltjjxDb4Gv6XZA6R9EQFM3eU5z1APdnPtqc
8q6Xnvmh4un0/HKlIgv0tvf+J8hWspz9gJT36E7JFhuUpVuFJeP59QiRrW977A6UIMMKhpgX+Cu5
dM0aC1LTyUq1D7VOGDUpGeF6OdgfDyvhbGCExWND101kl/i3hHS3cTXTfcDnMN4DX4VSUjl8w6Lm
SDh8eE35f2KP+ykGERf28tXG/u+L76wIR0iSklovy9b2svVoLAQYQ7iX0di5MF50n2LpuciFmpEx
dpMPKH+P3175AjxK8dEevK2AIFZRsPQt19DXy6CM2t+ofm9+EgJXVdwBKOndBkAo9q/NnoG1Vmx3
AQPgJGryBtxR0wPOpdwQdzHUrBgnCkTlzcYbYt3H2nJnKz/3GvsndpdT8JoGM47Zw0fZl+bflOQk
8JNHW3cOgAAtU4BVhfN17g2C/JU2iC45WsAnQU4w/iZ7J5hKyKMmuyOFkfJkWDL8Bc9fhTJMSs/l
5P6/SzZUnn8+zW7zohEai785RiazDpDmHztV+e1uGntE1uJ0JABn5UEpyv+1YWM54tv99uG51N96
uRNBNlnou1ybmeUwiHubM1/++QT5JIZ5QtPH3WVzPw43hlNxmtriL7I7CHLD6d0nXizpDML+x+SB
5ozH2SvhAiiQhyZwdk0OPureCEc7pYzYY6a/snysJn87PRaxvP8gvjTY+msuCv5nT4SbvNmxepjB
tG6+6zpmMOGSuDQsQnp4eAfLXrqPc2EyN6MH/fjDXKEPHW89IQeDQ3BNi35yBSbe/EmWKVuYRJ50
PWTRwIl82UOfSKquvA3zLcmnzKDPEz59dxvLOlCM93RikB6bcG2A6dWs1MdlJa8iB1pd749Hrna3
vr5MqCPKP8aB7Xol7PK37fzPDfI5upvy+/9/sVxCnArkilSVxwEYXBqkAn9ZiHbv2jnqvJfBqjRI
NVhKx25Dg9PaVJ31V3oi9z7/wrwbNRkJPZ8bLigooCQPVtvAWDX7MwpklFSho6n19tojnNS7ZHpj
sI7JS55LzcQK6Dm55P0Ccm+Nq95eRi7JkPcUOSUySVs53xZa/Xfsyu7zJXFfZ0xWnmKiPz5rT6rn
Yr68iq3gI+UYZBgxHGP4IAfAZKdbXqqEynLoW9rsNJwxjN/GVyYAGYwG/u1nD1F8wC/NGrxdHHEB
JLNGMWbAL+ItWuWv+p+iHcD21xTBO3V1rMZcbXk+OIf53oZJnZuuvaPvYos+sBG8j59cJ1OqSufT
3dwsUu/YRrImzBmfYWxWpl2xrnBJJodO67VsZ8drcm2Et6wp/rVzD3g0J/i9hbuuN+xfmWAoYRmT
0N3r/TcSHvtPLlLOo9xfSNWjv+Y4PaOnx3EGOAtqXXKSg8ZWXV/TcGfn0MwPBBnA538RfJyLuOwB
Jji3nZ1sRkoXJ4a9SfgoDZxR/UT5aSq2cqxtVCeOm4PNOiCLjuYc+wgTVlE7Vdp5+VZRPXHNORy1
x6RQ3JzGL842+HZ/lqhRt679V4sbWMYYVYxTOQBoH9n+Ubtd+bhxarYIeu/HC0+hspSnZiGsxDrf
VmCilZK/xYFFzAM1BLMY1FoMYfrqEO25PjIkR0+WIGyPW3qKQm0rkGaSWMIyjVTxeb6LlPI8BmOb
V2vW3a63DyYm5CXS3cu6SEkIdPYpzxrpbheMzFW8c56OidrLuVu2x396r89J+yg2CSeZmaxFc7pC
3i5yDFU0bgX3DV0R9364TAPygrANFUPaZNc5XPLx8mA86bj1tDKtLwSz7BGIhgRDkGJ5dsLe1hLB
r546S0UXYLLR3jgppNeIHY5YD8gb1uaEUVZ8a3llOTNYyP9YegmrSMOF1/nLDATZnjHCC15XjfoC
PnUhOKB1zXE27OnxQB7OCb55NHukQ04nmFkR0ZUmuDwhFl4aEeuQTZbj3mGlSdmny/lZdSF0fnDz
q2zkcM0qLemMLHhmNkhg1tUXs2ubl6EKwD21EPn+I0QSxUzDjJDV0ugG4wrtIxK2weSLuVy/pm8j
bp5ojL04vmcqA9f4fc5X/xqhcxokcesKzwZJJk4YW2/EFWsPGW+WkkDGg8ReEmBcwYVScypnEir7
DzeUA0bG2C0AQfjLgKZUdGmnPXLuptqSJnjhB40X4djg8cnL5oNNAPpqhhJQ1Wi3ik0y6jC3rhEv
x4yPR17c58cprFoRuGliwVxQUO4y08uz6uNMcUy+KRQlrUoW0+gVPCc5uq9RpK0UWASFShtkqxYU
9qdx0KNgchM91roQBbe29xDFrbJp8vGKNkdzBQ2I7OcKseF7KdfeaHWvv7RpIcZScUrYNtXnlnky
/TskICkSaTnyCRCcub2C3cNFrB0Tg+tm1y7oKPx0cEEGlLhZ2jqFQ/39kKGBrstd8CY0BgfIDaAP
3jSkcnn6jy1xDaBWIYsGb1ttz9tEDb50hOZh+7glM7SWLC0V0DrUSgA8HyrPPaElMmS0WGMZDDdh
10n35+WimC67En06Tir2eAVaaN8wOKrHNR7WiiVuEgAyB4KC8nohfhog4nng3u73n+YaQeTYUh0b
5lzRyk25FFb29Z/9Uh3r0YhH91QTomiftIzVIswBn3NrhdC+a3Kn+8qXyyL5x1fARGoAhnU2k4gF
hw2WJuTmwos43LlNLBk5LdlEAd3lbqrp0ZxbUPXLOdGZjkw04uFw7JP95kfQYY+qEdngGibbul8k
9fUPT1T9GH6kGiug9lVb22/A2tjtdpkGUpAhHorS4HHPgkd6lOAlz4kz0mFU3EHZZBhJtDFAcLtx
CeaqKNIwygx4rkj89ipxBZ3ABqAopSJTu41KuRlFtj5na9v5bgR90z9Ubbo7OfjmJlbdCyf5Wi+3
tq3Qn3YJ6PI8vZaaYW8t28pSrgxj5bxjv9mG/ube1v5Js0Zs61y1hDUbgphFIgFlAU5zrHigqOp+
bdw76gwp8fSKH01bAbjpoKYM/PyYxPuZWsIKirq8g3fvWeMafgZ4/VTldkJEsuxtCSKdEGyjEufQ
klfnVZUu8UYrYTTFqx1Imqr14diubXt7fFvinhb9AHfG4x8R+1CZfTikQ22TkHpZkjTivgc1UfPo
ogWpgnRoZq5hCHT7O8vk/6hb3ZA+wm1vDfR8CDTjL8t7GiI8hUcJKfIhTfqQy95+0F+Ym20jiSBV
iOZRoDHhhrctJ5H/HerdzjMXBSL4/oFFxLBOK7ydrVJt1Hr6HnpRlei5tudmT8qem3tFfWma5Lj7
DE/0AQFGANvSImQepLOWls1hJx2L2bfY+hRZ3pHdmOBME/92jbG6r/Z4ntTZTv6XLGV+CbqFu3ce
f1f+Nad1BT9kLLjG+sPFHz9eUZMzu5eFrPiBS7d1V5yy+xb46AqX67dcXjlpyiCMkjZI0Z8LKdLn
PeLkw/QrDyPpxd7DqR3Duojmj/wnsp0C340ZgvhGpSZK6PPaESASrYHzHyc5cgMcgBECpyCu+1eb
SQRg75xajbKZk2hKAzBkdUhQsEgc+R8cAkgLaM/pYBcwEcRtVXzPZDkygcd/9VBB3mTISk+toOK8
7UzstGbacbAVVzgSVvnvFQpvcxZZSPzJVf3paQoBJ2x1SypWWb77qGsviAH49Oipg1TGqa3sSwNp
dizOS5ChrOFVcxyL7MOSxxIvKzF4cyS1tOmVnNGKBF5Xl+HvZ7liM9a/jl1E7sNAYmP9F7pR3uIB
DdXZiDIDTDvbfMt/6kdl2tt3k8YcVDfaSctzwGhHjEg81RF65Skfvg3699nPGvolLAU2ut4icMAd
EBpaisYscR12A8T9uFrSLotmTEJ8Saud4Tr3NksXSm0VKr6SQl1EDuY3AScsi4XjCnNKI5I0ig6n
kJnMiGx7hmArkMsQ22ip2UAlSKtQks6JYOtl/MEGY/oVm508nSTvyseKx6fxCtJd3fbVfvs4VVQ2
FWsWyVT85ff+xkrRTYJ2Lp42zCZpWAQ5+Oui4qGQpufyVH6yu9354lcPb9cKCVCz8MIS+5MrJtAc
YxpaJMG3IBbYVNKcuObWtZcEBnQCVd2lxqazIQ3yvtkxbtaODz91mfI9hd949y4M4IFgtgNEoi1X
0kU14dgIN+mzgxs3NIr98n3axz2bhM9LUFFA0HI0fy5YOlDzFU2okeG3/Q5BernPTrXtKwDMp6I4
WBZ7vpgWbE47f1+SFdcSP/uKJSw/efpbstO/GTjr5lpHwu31LJ4RcEUY5VCTtCHQSSuuVaNnf+O+
q1lND1F/HjNFU255L8MG9BHk0RigCjnRQ/otazlnthANohdlMG3VDckdZNQ4jk4Air+QwtfnL35h
remkLTbVyNi8y+XWNwboKKPhamjn/DDxuXfcwWVMiuJ+3DrIIOAnoiwmXnV1UUXIlD7V8/vsfGYr
R59FRbk4ashdOkbI9FlplHAoEboPVs68Vh3vt80j+G9WaIvtoFrSukjTSX71wjh6J6RTAS5XBjb9
ysVwNtSHhlXo1WQxp1+jN4HkzPyhmogAVBonfjkmZcK08qEzJSMjdlPTaBfvSK6wXzRhQ/RkSJse
e3XVEVbKNS3iIksyXnXOyc0TkRttOBWc3AXgIxj7Wl1D3VvmmQ7e+SuqUwteUBIdPJefe9bG6kcm
idGyhWWlJdp7BR+uE8AM8XMzRDVXqDqWsfG+C0ceu7hzzQ8R6XvWB8eOeWLGFXTqZI9ZUhmSjOLU
u6VcpcLZZSeavBrU6T9MCvkMNaevuha+2mswEg7JbyI5YJn9PyFpc3XXQROqWEO5Ryd7Kw3z/WAj
plDGBUfI8SOO0s8g3eMiGKKV8IfJyy5kyht/Q9X87/KZqZrlbkvuYvCiYnEG1Jj0eZiy9JNokwgK
YU8iAHgEVI6tTPyLqGvnJ1hKn39oGadTIC/oHxyG30hCw30+Heco6DIDLiD/fteQ5dpV4HVgTafR
zRNQFR0CZcmJK2zUQPnDPGHvsXwg5+VQUbn+uVq67Ie3swd5y53WOTJhEEb7YGl3uEVUCrR0qeuw
uOZlOrRZRbTCsWcqVC4wD+3gVRumE+2SV7I0o66SGqFp8+MvcLlacv9qmwT21sWNnd5prinq9RA5
Bj0RKDj0MpcP5LSG2aBCieqwdP9HJ5Yo8YUnhKGLr0Jg2YGpmwOWMNYcBfvVCyVmsjd6xiUMbo0r
Azm7M3chTjWmsPySHOnnYG5298C/weGfa8Ni3rC98Vr/hzixIhyd6arla1/gfcuEln2hPHThcQEv
+5iZ1eRpsy4dU6/BHPq2002GZzVhMLfHBxPrjT04YQw1r/9TM1/VT1v3h4pCNH8xCUkymVmdefmX
UnL+HsxVSIn81VAeLjV02YFvl+hP0U3L2WUTWmAjpdqhVLcgsG75vBIOtgXRz5lIlS7fnkZLtuvK
/aKdBorrTawfJO+ZRqUgexMVPAanGpWYwe6ZNwMMmklOG6uJmC7CtyJ7Tf7DCTC1d1uuAj1pXEGc
uFIWHM3UK7hRYJyogDmLRycmU7beOAm+BaEvX7DW8u8fmJUmMrzwjajnv4WPaJzmF1OfQ7aHekTV
rvK+Y4LyyLFX3x2s3QiSrhykBV7b31uURM8i0ULLTowRv19exbU8xEeU30Z5kihUEb3kBqMvbsx6
FxNp8V4Acq8JOYUPTh/C3bs77G1It/tASMk9RwwZ11yN+FDdgNouQeiMKjDGR+RWBK5jOdv7cBH8
GXcwgIV1XlSiPbEP5eBuGJIm8qsexmRao2imWDgFJhmAaraUVCrGWp2cpHUa+0bhRMUTOVVCFFmV
2ryhNkGM9a3QnqaRWEnQx2q7PJ1Esp9eL8FOimbqg26idbsrBTN9/O5/blvNZhzeWwNgAyBKFi8b
dMy8bg2begeje35HMGQnmhH44J87z0Ie+I8LQYxLSKYA1mC0eDznkS6fBzRI3P+ze7Er9kmyijW4
H0o2pkPVPgbp0KAqIc6SA59XHV4Nkxw1XWdY8iqEhNbqU2MZIZMpzogKr6rIPNu2DT/+J8fb2/Hx
7NI6kcOeH82fjtbDvMJwOne09auJSZ21MXcolmQ5rSDxV3w8lykkiU1utSC4nuDEYWSOmwx6Xk7Z
o0+LojNC2vtx5cKjNwSQXhAXLFnaQArxJNxT2t/lWhthtmtH42rgMqapjzF/xmCoSkhttXkUrODX
sXCph8WJMEPzA+H0VkYwsVTBKGWs1BRivIQEIvatSLwDt1a00D1RUMPRFZrG80/ITFpEZl8ox7PL
TahCmHDu0HRx1UGFKISsas4dS2rtczAmxkt7hTrEjNErkABRmieAVlPtEZP8IXErbwsSx6rzBOp7
QAjUky91jDDTzpT1w/ahOpKIGMRz7yrhXSQC9HY75Y/LFNzfsPfF5Gkk9g4YsfJX8vTNDRKi2SaI
1z5nChiij7KTQ2iY17UkG2J8DySyV/InItaaeentiFJNALH2M87s7s6FbvZzapoOkGe4uYoZUK8g
9m6r+tuj0UzeKKKDp2CdOrUiXwemXKjjmXt79712w+TkrxBBP8jDoBX6lUOw+L1y7+mYsVS3tSol
c9TwziY/5PVUMid2JSBlJeIHLETUWPiLF5SJ6I5LMDuFM+kFNSnZXPpMEgoPorILdfbHiXfUvss+
Mc+OxTHJNyOEl1Y+hnbLXSCuZ4cQ9JqKFlTYe0t3ltzlaFtslQXXRdsiLkBisKsWO0RjDc41kCrN
S4ohrc7S8dMnOkbMNPupJP8v9Kh/Wp9XrcPZD8gznVyqavT2vRO3GW+uJhKzNadZALEjb+KJzEEF
XVW/l9eP0kFTvYNzIw16A7HiOKoFvcw5K29bFlNBALYehB6y+IelLuNFeTgej3vuY8Rrejn7W2q9
GZAchbJU8nHkb3YoZXrdgGw12oH81xe8jOCknzcgiQ/lAMm5wXR6xsVt16SNYq3+DgoHH+3TQaDU
+RTQspQYMoJnSy12ad4uB115CQcx8GGyncJfz0ZyVG4IPhjhSvN2J4QXFBiwHyOgsvu4VJ2uVPsi
A5DFsiv9tcTa9y+K791WQjucCVZEmTDzQ23kTS9dwwPMvHTKXu+TnbbiKHsxqmxV8gZMMUuqBZBU
89sfYcWuFE3Wfa1aXb7wXSnz7vIDdbN0lZMCp3KUbkHUKf8qHFTk+6ejxfFJSpFJpTqXlMc7+Ifl
HIsaL1l3NR00ZRbcIoNRoP6xH9qPbWqw2Stit/VZKiz95r/exX84YMQRL7etMHejsZmbW6WZUG4E
s+/DMkJCXplhvx70Ge6Icu/De1WqKxbtTZuGW9+L3qH7f0q/kUJjxNK4Dm+GE3fI0DqvANq6Uexk
U2jY+vFwoynmgeAP2cNfNhXQiN7LR+cjtTvXme/NEnQilsCFL6VI6rnRaRkomXJiBGU0pECbv/g0
r0BP0Rn1xj1fDxji+3x/P93QJ5f9qm3fOKh7xHJmjcarD+II+Br3ca/Wzm/w5lIkscEFMESJ3W7w
TdvSpIKreJg7kKSboGpR4csfJXq7PhnUrtUcz6/+eNE28vPlVW5k3aoY0PBRRBgi3aYOU31esDLx
RX2Tk3uNCVk7+6olEHW6zhnkHJEipKrjBaVkpNSg7zfUepHfMyS3YiwLlKg2WL2Ei5j8LfY5w3mp
nabfu283fpZnpQNjCvCi/Fe3YPPbGWOPo2OlyOAq+lSuH0eoPS0v52RyD1LJvAFjwNkUyc59F/W8
CYHCfThS+IfAFhTdh8ql6LvfqfUtu8N/ARsFr4k/bmx76TPTVcrKmDKMfGy+UofRWlV4r/Ru+QdP
Y/SMkIDUZ86q/E3DDEHtc0593n5zUOAQO/qI2jJPl7EShwJNobVR9sLLQMhsj3HukNWlz28uV0EW
qwnoEOhTqN2jEC3M0IYW/0tqS7RtWSa5bAo63I/eMYOsoCPDYCUhzlJ6H3BZzfK1trGRUgplhOAs
uLiW5xBflGg/ls0aGp7auY5vLyigQl5VryGDVavvWanNLeeMcAI8bQwDh+Vg8ZUzktAnSoclUWPn
WLynCju9Isz2+sxn9maRxt/G9OoQpaZGSVStz7Lc4pVcbg/6z5GiRDOCN4PcODW1n47RMevy3VUD
MGNfOHlm7WjyW9VqDxAV9H/dRVTohLG1m9A4Ioi8qb2vdkEys7P0zjqZ77qOfo79SVACENFQHsgT
s/5eSKvHq+l8vsZVHB5VpPna7fUFfVkkxWeBREujq7Iv1Uq2OrkrWU1dGvBTIvX1WbhFLzcMtpYk
1Jn/OU9N9gTk54gh9PHG//mLrDsCk9yXDEXdY1Y2cq5/ilL51dfj0LvlrI3MreuTxcnIKlV+GNi+
uweHZDL++mxlUNfqgDYTEO7KI9pEfKpwxMy6MQVD2FDmkeN9dswWSgANp22n3h38Gn5odRPm2Alz
Md02W2CJ0iz2Hcvv5T+3221NlgcQSvKkS6dILDMZvVbzFTcEZkGuRsi+Liv35tvoWFwzcDC2LzpS
Kq+a68Axd/hrTpftCtJ7Zw81EuJ7CHgbIY23kTHKQ7a5tWie1htLGNj96/+05nTu9eYYXllnuXRI
NbyrE1QcDN8Ns1gIqIWVm88xACXc2pxp3jIRtaWFpk2ehgKrLJ5hqD93ckmDw30KwopkBsOVAQ9H
Ay4fXDCfBeSlfr/I4X3mxfsj3VqMuOEvjqrHGIpv3JZw+t2K8O8gN/8Z4JOl4ScTEBSVQT+fNOXU
MQdGfoGaUzsxgrYJUwZdC7dUl0Max2bdOvAbDxwW/JZUILMlqNAW8q3Z3zHy6zT0HzOgUu9Gf/qZ
gR7hbY7aC4N2VOu835p0KNxz4pNUgkN5UpxmP9gpM7o1DclFwu6yKGRNb1Ulmz+mUJ6qzahilruC
yV/8Gr0+ryZrp3XZ/VC+i+6gHHVe4ThqeKXlXl9Cyir+HxBy1erRo9/GivCiYom3cwVFD/UuACK5
DLothdijKWdmum5CbSbTYlYW4dHDjrv7/rTPFt6SmyS3GDuQKGiGZY9I3cao+VXAxo72BjMu0lIl
5ShsWYKdvjcK7WV1QVR22KacyRndVj9WJRgRWXpj+7DBi3gOlsRWvsBeM3T4TckpHaTseOdqvz9L
yFCvV7kVrX4P9E0fIAVTmf8igvAES2Qx3dS7cx3gJNJYDttRI9Y2FIdy5TRzNPA9HIbv3LDh6a/F
0LK7l8072pvFE9qTQxyvzWUfV5QzRXT2Fs4edXk1ZttxxR/H0VZHyfRPHDIMH1RtSxKbBTSSJhU6
QKbdQogxJu42M0z0cFsxVub4BeL+vZCwQH0WnkZI8slIqKcSZFfnBhlooC/eMVJ5ZNr6fk0BylSX
c4zvX+zxYrqzdTw0929Ed9qAarBBqiwkdH6+17BLUlC9thQxbTjzlNFvH3zB9H/AHqNJfh81RR/4
pbgoQSQ+iue8lVkg/XZ+lZzouU1h+FY6yc9axCicH4ztmoyn5bBzlCjq2Ywm7MklxfALL1CrXRUT
880Sdap9DiTzFpIGTR7D6nv7+FlLS1BUr05enbowIJuBuJyipWvWqDjXQR3bN4BjNLibeR1l2CIu
uOvCE7UnL5xMbkFN6VNVLpAeeqfOwBf7T/VS6UQv3343sb+rzqFwXfbJcSI8Gd1LNWTsJFTAkmxw
/0200t4VxaewtuhRyPr+zf9gHTigX1W+uir1MrvEKoKzYNM1uczSzYR9zREF2dA6j/r7IwkKF5oH
QUX7NiLK7ynFs7YSg0UtDj1HtvloHdYVxgMk6AwK3U/RZEf8rLm4hMJXEYh25MgSWskTNQg6bNXs
QxsM5RENQuyN0oj5HSDDquZ3V7yxwZnfsua+3O5BMGhGgpa5rOZmq8apjatc6cLvzzevO1+m7rml
Qva/SlyvQ4CjIvUjjYkoS7oJSywNoRB2doh39bG7JsR8UgsAMDBhDt564wE6cexg6byA5ZHOjEtv
bgqJRQK7OORyZjMhN6k5GxYrKkIn+aVKTs3wyfvmq1axSIBvSWS6cK70zTYjUTa6YxrxBfhhpLnK
dzRHQf33uAgqAB5+BwNv1hoY0HEpm0u4gk/QN2sYeIG9ddVEZHUt1XNUVn7VjvfuGxACbvuBdn85
UIPjSFXjfWFSotE5fFEONEYDScvK5SbU5rHLdxxs8qR7XQR/H7WM9Pkh7f+mScEZXp0CDG9p/Tye
vyruMBStpJHXDZk4uWVZiZpdRP1PtDEak5bs5ZiD45VuHVD8gJ/tgm+S+RXJBN1A02pi/NNtwZqw
lvcOfbQle8nCnN0W3ft/qzvMgWCxsAr0PG0b3GiHQMYkLRJfOnvqCYlnMTfogDVt+XdiK3nmb6qL
6sn1m2vzkatSJmAGSyS7/fzbuvnqFgSgBFB57iv+URFlL3M47XpOdI8J29Rml+xSU6MfAXs/YipM
e9cylnVjJje093MU97m3G2GUgzAzkxN/SjakQ8pR7uI5MAy+VGFX8C6AO7FF30xg4NNpavcH5JnU
OIF6utF491BwzTGfrwe03OkNwq/Byh7pTEEJqcEkiQISfoLzUJhMstYIw0yfToKgVw7wqbWisH6h
Jck0+nZwFE4aZe+JpcKVvZBekFlq3f2BNyK9ykGqgl/c5o6IQcArM3K/5fQ3FRLtmJaERxf/MxZT
33LYw9WNAOasVCy4AqGz4+N1d9x0W9DyuqIRGO+LPFzzgVuJ+fqWGCZe5VC66PNAPFoTl7JcLQa9
1ypthTAWdika5lFrLou/pqVAxizqGV0cYpYKNl1ukQpUXNuUmcc5EAsoJbn4ZDDc9Yl9vb3U7Um1
LSKfmBYEAFQ8ARPHd+s+CNg4wEA3ah+lrdj999BurqWClJU1VaOy1DOhDoteE/RuWBJjBSBlmyzi
mab43k8mdhg8qvc5wxWpSYLXupLxaBdje5t9BExRd83iSrdFQlcEMpotoXuG6H6xIxFrU03uL3WQ
MH7dPn3YbIcw2ftCFtnRloLfxiY/IeK0GFd9n0GoMW3kDyN6Jy5B0euE9RMizRLjuwEJ3n+qHX1s
pzM7wxAkbVFVMTrRU7zM1T0JtShLElm57Ycx9n3N7nVc6qDRdvt5pKzyUDWkwoeZg2tU6VqrJLhC
IhhHr+QnZRmlt+5ThsrFnN9JlkAA59Z+Way+oUWp5rFnhKV7LPCd6tlFILh2QExGG4ew409LF4MO
Pahq9dFDgvXiQEG5RElqLmMudEpcFTU32rnWP43zCobg0WAvLIYsp4YfLs6rb6a2/gicW1Q6HfMz
OWPkVBv2zxI9Fh9JuUFYBBePh6By8ifHCEOViehRNwDP3VC92Twqa91ICXkWyvUsjZcmLQbac8y1
Ji4mEIgW9RpRbmZdmsS9fqmmkTPldZRdug7ZmXb30LkR3517eDqWqWFc1tb/plEKNh6SnLSBxG2P
ZT1Z6rZR/yFq8XxVlXlw1J53oYaHQvWXbBmsLtJ3opSQl3HASMRObh8nKZhfjz9UnvCrI6r5Y4MK
iWaxReO/RfalXZ8X/IiOZGQhetEqSY8X9pcZEARNi0Lpl4KtuAz1MYbcBfPeiBI2oPxQbN7qFh2I
vtDHqNphyx4uqcoSTSfbDMMr1HlgYdixFLo1+94dqcagU5NL/cFyX8zeAwTjAX8kmp3eoO1gfC+w
aW2n6PSeC7Nyp9mMs2KxPcote2qvZgHHbktLBZOqqBSFXyXMnge9hTcDDt3BJ0ldOBfmmG+XvL0I
QyAurdczBofeFBaYaFZxUm9WJ2/BRkEJuRo648bDma1VcM54viRyr/uWJ/rm/NQpqeWFCulMfeXZ
Is1mMRuI/MuypRFblGAg1Tpt0yglUuaV/u/JP1iUkSmuOFns5FHKlPN4gkWL+H/tvX7ZbTgK1DH1
XCDESdRxau26PiJauYazfTcB4YfDQzDf5IVs2ByVYpRlHHH/n0RsEEHukbXCb2gkaaQ3xtUDITj/
pVr6rCEoaN9b+SKbV2uXzEKDkRg/jbOvzgTUcfDeoY3R6uZKUviMgcn2g1wHT4cnbdPhqu8oX5Fn
OVcYb3+VmiAEbTqhvYEupwoT/ZF8say13owwJsCL3bwcjAzbk9iDZee/QiEPlSqPek64ZDU8LNoM
bSThG5Zrsk2FGd/wDFV7U4dyHQVFrS7HOYzKfPtJtCqvmxuPk5pc4aAsb1JlAD7hwfJSfyNr7mMi
WgTgvamObJMYiT6Mx4R9DsSIN5gGEkA5Aa+pon5PdKzN+wwZFDJ+PUACn44qkHNLq4llZv8tm/zH
WecNiH7HIpCEbnDgNeuasMJnaQ+TPze8mWP3C79SzIkNECaJaFkwr3JQ/HY1NTM0EgHCU/Rpc79v
B43D4QCaVVcbEN+vTDh+Dz90VweeAPpDo6gKTF4T062gfB8TrDLK2n+bInGy8HT+cUhwpMoWMpAr
/xJ9j1GrwfS7Hl/tNR6W6LfG/wbbvBIpoJIlqq3z4Xwp3eaF6KgxITXf3kBR9yskqf0M8Ai7daEA
Cs+e6XDZ71LvLfb53CQwI2J2nroCJrMH9Ld9tQonFFIoLJAR8hjzZa0I5TybWx8HJuEDly1aFYea
zLP7tsyBK/STBTLf1zyfOGl5BZZFlmaIhV5S37c5p7kOJJ+DxFFMmRiCou6cSHCMnj9UPBHAzt4A
7CIkP8lNICkiVJN+q+ah1ZJ5Ar2uzWVBzrQ9wcExczeu4S+uYW9A0cvlMFdoYGUpw4quqPvH/DC6
WKSBHAeUtAAOtde9DmT2iI3ibjD7Zq++XtiVBbn+Br7yDXKCT62JIG1DaFIDKpvxhh4drze8NQx4
3n/mwoGcLfySDtzEqaiyVI7r45tHz2em9A5FRjH03ArL/TYcBWfAcwAvJ5qaiEtLk4vxFx3h7eq5
gDO97J2qGE7PPD6umTh63Sy2eS8QNR64t6YBgEbPJ8tFJsRMuyag76dZ0PhhDcJDlmtiR1qVV2fe
0Ug6PWAnj/Sbf/E0uAv0YdO18r/CZO/hFIa8JKBv8e1lUdVrO+YRYbkGLzaWNJqS33SLjTV7Sz1+
ZHSPRgAAksNQeoLc79F9Yj4qUaaNLlBI8QjnacWtfdEf/Ai96C46W+qREVgiZGvoS12eUOVCpoBP
7EUd66wEJVd654zXsK+aEqW+0XpkUcfwvCorbw9xS5c+3q+b0peqyvwwjw0GMrpPpmQwSo4Ownpr
e8NgUecG/z07RsM+77ecumEJjoVEK62cGhnW56d8Ke4I1+zaS40rinuIXCweJ3Azkt3C2/b7E7uD
H3Uq2eq5Hd5pA0MXX/Qb9EB5Kytnv25IMfhyzl2fGX7gSq4QmJwGTVFeSS8GwfaCzrK0OfUa9vdu
9ovu+8dAugYBAKSQe3hYzaJRLw4gRGZhuDtR1p/p2eUx2ha9trkNaF5CtDC/gnk++Yn8C2f1WSFe
sGrfL04s64+b9g9esAbFNJo/KOdUFBbedrYh5TR0f5lYn+ARTprhL9AwFXF5UShOQi1Yxnq08QAL
cIpXTRGyGck5+2qSUl08eEj08OwI/+eUob65Z2/Yq8DXKhBUohYeZULttSJCSg5N1yKo8SaCLJro
+xoirertM3jmUqjPXAFfsAMsDfmgbui6r9/fHhtarFhxZrmOq3AQKHXSzlajK4TpcpP0ADX89mek
kwPI7epq/z6CRaE8M0Arfu8gz7P8XXKq5Kn7WzuG/1ImvjVOLNs00N+N/w48a4ZuoXQu6XfrKoY0
TDadjpHJKX5cPLSwikeB9dfsP1wKdZrHmA0N02+sQxt9C3QHT7lQFbDa/VZ3NzcEFlHRqUw9LE+5
KYdv86Hdq5Ya+fZCrfyXOKdIlE4k0DO4guGp6EHSj/Guy27VDs1pcUxKe+NtNTIHolFBIQd3vmLf
LYv37eSW+kbhbQDvLAPc5sKpamMpkCvAIq74sci+EWBZvK6PIRTCXACREh5OUbCldo5kNeaL0maQ
lrq37XkYhP0Uqv5OayqM7KBpyQZamQNbQHVM5UJ1JMQKO8V4711bMpiDUwt6d/6M4z9gx8lPb1K2
FFeebcHq7xHGDIJxw9gI3a72ulTInOK3o2Z1xkp2cEVWvaHbZ0U3KjIq+8eGX6YqySF7qQapyK09
V3fPNAzowJCk+w2Bg4MUMl6nrF9L3ExDnAwt6Q95Pv8HQNQTRypAP6mEvrzE2efZ8+n+VxB1JBgL
e0lH+75nwTVXYbzKaa9m4MxbeQjYvzKzBrW98MCyUs767PIRDGKsJPNAbWMDp7JmiVaV7fL+nZ6y
qw2rNnVrXZeFKRMuVYCoOBTIBbJ7UOpYNqElHp4UA13vDPN12T1HwAkHVTaeuNai2NQWQxJscTk3
OO+0KWF8TrrIr5cUtmdCSk19AJB0GqbDjnCEIBe+/rZsAsn46qfvDj82kWIPeMoMv7bqQYMPjvdF
9/CHNESibNCtIwB4iNoJAkL8w+DUJB9zZSooiWv6ylUuoHg5GF2/xa4V0L1VC6zh0qpFnwBdmQp1
jlwkMDeZvtNf9oy6YkzHO7GB17ptg/PXXEk3YIM5u65IbEozNmyUg/Owd2HH27DyQhKNVXdAtbNB
DxoMHkmizcEIpbY5W7gOZIsDeeWZSTCVhU5ZO5VIXvP1kPYIgfL8pmePRI+DzdORrL4YpizLLb+O
4fBIXKyL16lf6/swgCmqTFV8WoWQ/27Y2hF1jFSGJ4nBMLm+BHmo9iLXvAGXGfIaMWm2CcFiZxMR
m9zLE7FMXbVmjx7nq9guSwn0MvZkwsqTyJ7+mgch619p4K2e/mx3LKTcv9RECSo81GJgjausPFNF
LhjkkILpXORCeaok3KPtCFcWltspXf8h4g6SHyhvP6hf86k2wwUQYyXiU9x32ieHTJnk1u6sBtRe
e+Q4ayd+4tVVOQ+cdJoooAU3TIwNHKjDjejOmzGHKdMjlNDnXaaOTCVvDJe13/kr2nkuoAGUP/Vl
ovOZknkLVr1lcOzo4hrzg5k1HD1MSu1JbldEKpUdzn/DYQ3av9YhaJZTFg/swsRxOKxU+K3lWFVl
5gM9m1fdTXu0xKPbxSeFvNh+uGN+eky0EYsk0CCCr9Rgg7/FAiThNLRep8L9f/rsCmXu9qL+LtR3
zefuyNbkfFjioY/R7tA986HipK4HvygCTCaCtSUIgDd5Nru8KfPfBkm9zR57bod+geglHFyGWi3x
s9s3SSaS6qDq6kXEL9djKINw630+ZJSt6gI9G1MBmG+3rHq4ARop+sl3x6U8zXJHnNPX+HlWcQ5E
kNLYSgoL5LeNcLCd6CPt90vDKuhnNVF8gkMwwx3Pb5uCpzXiO8l3P/gQqQEuYJaaoaDLx5yrhS+a
o65pVN58w1SM2Ev3OWr9RDbWOodWrbi46fb3N1wTl4HGLFrvwJoXWoEI+U40AHoRYX3895pVh4tR
/KzYEWZfh0n1Z9DUNo4g9X8RZ7C0tgpGns33SEEbBGuUtdwjwffQZbfHnuZAGcN572ufQCDbkaIn
mM62roea/zT7Q3LeauQMCdyu8IwYFn9y7/KjkVbTUaviBqZszl9f6P6z/5WQudp59inMki9wSSNw
SPdrXv0WBZAf+T437Ftb+qOZW+Jt/o/7qCowZ/q3+UnbfJhYs53x2BwhZATtxJq0mTdj0WShzERf
CijJ4tqf3JeZuMiccrIJwZB20mx/zvq7q2z/ARdnJQcIL/EpWYEtBPgkrNTPdgat+thojq/Tn7Cp
l64xoKtcFeYsHa3rBapXhu4hg+RjAQT+i8aT7vpc6ljG3u/RGMaYUqk9Bcd0Hf9LHj2DWLXqDqFZ
1C4UT4tu1k3QyYEFBsmxu7xMgjs/oTHhqWDI/JuBsqRW07OPh6S72FWvvyZlI4ARWItZDjlfVWjh
Hwl+44HBraOhChGh3Hwh0Q9A7mwv47+jf6+0RScTC/h0OEUmJVKpXKGobo1KT/jEoCUb0oE/Pl9I
klIEQH1aRM774D/rOt3T8HDEgOPN854ij24ifR8NtzvUhdfB0Hcb+D/jkPJhEHC905DLcJRQ0oJ8
ffsag4VjLTo7M8zrQ0sDBapUsYNG8STl+PrwYC0FWwbpP6ATCxdpaI/eJPBaaCGXs/vYUsOIrG28
5JcLG12w1PBlNSsD4vpYBRaYBIt682xYBhzy/kXhoEM1+RZPS6DC81gfHeU2IeQ+hx3KJ4u2xmaK
0LqjMyd9dVpGd4xwy47xb3oN9vjpexTEIusycvuFhcPV1f2FxSuxxlS0bwUBfMEminSB+WPUf2Wb
CsYOOH1u0HhAuaZ3PE52Q3K748rUKvcyBb/v+j7E9PMGV+Uf0HBe1UPT740jQuFyhr4tsFAX0FJm
pjWRJ6/WKVngKRZVX5mG/gN2QY3cvvwDCgeSqfgttD/dJDPkI9Z3XHaWWX+9rcGStnmHlSSN5P/o
YFRZF4mUFK7hUfLMqYtDsN+XnlEAXj0iL9e9aHI83HWnUm8Ehe1JpPQJa+ICnlsMl/UKjTV2kCOG
GdmQ3C+whFQIRO+qPtQ0Ha5rZizplselRORAY5orDlX8sn37J+TOJkPdms7GHGNQAArvOUyQ9hoy
o350Gf/AImmnffW2QzrIPz3JXZ+3/87oc4ElnCVmnch5eAqzQBYC7VzPwGKJNmim4LuUO36MGcJR
NCtfSOsNdWoQToGrahP+EmEq1mZhL3H+o6XdYIAvgxY5knjzt49mkUdy5mSDnvi3nMXzZDSr2M8N
Dd9DsmW0IXAqMzN0CpU3YNEXDg5hCnBBo86lsBHMi24eGN6E0GNzrHETZlBlPOm1B7cHsiD6d4Lf
HIoVZD7DkEYegKxBhuaPzERQOavVTYFerNFDNitEwsdcGcDBqN2sFX7aEhR7uTJ3tPgT7g4Saba/
JGT/a4IOiVir81zKTfZWIkMlmEqI5WS303YikvMaAk/qS6La9dT+dAMa0gsJupue9FIBz3YEsJgA
Wnbhl10v6lPeApX4H34U8mGg+lNKdm/p/7IhXOK8iU8zlSDzlygahORuZk9jDmv1Hk89PiGQBE8K
oHdCAD324LMjc/28AAUGqKGqyMvB0Nb6qkqXU9pXdteBbGNUJq2vvn7jNN2YOFqNqkddWUJZGyPv
GLhbEpC5ivbz/Ju2yHc0fOHCGQLSbbMPm27PcH8ktDBz89rgKWvjIpfXpnaMjz63fl32KVDxgaD0
vw2oB24f3s59rSzdp6bp5zw2JTXyJbG/Gbm0RkxN0BEcbFGfcCYRmd7Qtu/eA1IjvmQ40Ky0m7z/
TjF4or9bW7w/EfWgTg+OBQ0OAYPom2vbnf4mhulUosCd3OiAvjaVAgYe8chpMZU8bLHiDIVusNYC
PGbEeE1dQVeGXCZR2xeAwu1U9pZrk4n/N2oow4okhJV2fl9OLlSKB3Oe9RPfIMf+7723YD63Jpwa
S94iwhM5b84uNro5qaXHzlj89t7BSyyiU2bitVst/d/C8u8kIDTbbzi6lY0K84wHpwp5FIFyOlKT
Xnmx/mjSYsPYxThUtnlxMnUgzMlxzJOdo7o+uE/njUr1ukwVnuB+Ex8r01jrl1UpW/CL9UDYvvIZ
kDWHnDLXhFgyvQ+zzQ1GKH2L260exwnn8vbJQrrpWTE5YCjA/Q2llsvK/Z7EkqtLiSPHx5u9qUBB
toLO9v0HPVuyjmk+dby2lEgqJ4O4jy4/MQshjshcL9yE+6Leu1D0R09ZF6jK6bhIoAWUoCiqBlYW
zqhNn0EAv6wLmRH4a70/NzL4x2De6ZFSnNjIgkJB3sdIHz6+Vt7cmEWk/rLY/KS76hPffXg0I/A1
IYAe3LLTQo/G9P1BItSL5ties91nnAJ2X6oIVzlYsd1yzowaUe2AKNB6VjblFTFHyxq91RKJroRC
2toivKmuK6f6vcTnIOgCpygF1OGJ8mR/9NrboAA5FQqJGYkr2zLTA+0BxWcDntsLzDC5RHnqpaO6
XdoZOP+rjaq2G/8qQFW2QdicDleyLp3HPhNFZMANeZYtD5AH+WptiuyLlWPC0hStTfPE/h8O8kGJ
rmluRcg3UhSYcljIPA6WAHSqy04EtNBm6Ld4mWDbcaG/QKk+dPI0uI+aYCUqDuIosFtPRbamVBp/
541m0QRmwmebLYmuQ59gLNgOLCNeyXP8tsxFvrLdhB53YUnsCXLQVkei90e8Zin808XM0c5fQHOW
QyzCXIEvWFVq6xWI3/jPMJwHvXttymUNBCAcmYgOlywNzmOytaDSduUd4faTvYwbE6QZqZJU0DAJ
gRZttB4ZjgTtv5TSqYp5S6acz5QOqAyM6yiEjw1/UbV49f30JPthcDC4EOVwdU/WvMuPc2zc/0q2
EnoZohDwr3xwj6EkARBP4oRaw8LJo2lBPv+RIzDLQHbgo3x/b7ZMEwMHuvLD4pUjPkohx63CeCvS
k9TzH75AHKqsU62pH96Lq0zQZJ+059h5O2rYjefAusT90gzE6fJfjb0ky1A2/kShO0TIu4gsQHAf
rF//hBHWwy5e9ASArW2WiIn0x/gsfDP6eZW3kkPQtZBRNRln1PyQXRR3G5q0NXgEjvjJC1k9VTrr
JrIOFYBUyf9gNfHPjUjmWUcvWJ6WTsko5XM4t+UdX3KBnisqA0ye1p1CLTapNq3Oh7uSArNySTwO
lXUqSu6ECZLqBxfz1wg7zuHD+bnzHLjTOaQtGEoiVF7RWbcVRXNEG5BmmfecSv4Dk18pQxdSllpg
xEMlaJG1sns2ndM83fy8GoowK+l1ZcMfz+wE0l55cVyepowZfJszuqCI8POnmeoHGNdlMwUIVofL
3oHC6taPM7cAHrfDSxByZXtBnVuHfGi2Me2ks6q4aa7Ss/vz1GPndqimfQSRbJkkUd1R+JLKKc/G
shD3Pj+mr/CtoNSeuYIXk/5BpaS2JT6LuBJ5NkKK6/SdJWrqOuriq0LA8/l27/4UL1T5WNPGx+GO
996i2Sz0C/8xTVabb0YxeoQm/sHJX+YIoJDvZdYMGgnZnGEWrcU+DUCkkeBgsj7JECNok+yAkPgT
uQdvCEl3F86GjKOh4zaHStaH8lv3qCcvlIo0uAyDSkZAk5toNsZzzWlUaZ2DnJt2c6DHVtJ74zU1
uG12+nzr3FJALwd/tIC1YJQDpqcvHYLXK+i2LHWatmEausWKA8KFZDmmSlimWIac0kmE7gKR/jL1
DnyOaQbuOjXgXgaB8T7SkTrl0AW0pS9um95k23HdSHNCSt7NiM+e/tpaO1h06rGnIxBBymWlfR4j
jaXlQdWv1gsdbWGxzZdHPPxwfpVUgxU9uCMlm/qiMdoThmG8e4lf/tkYfPuBXxBniP5BlX/yG8VG
w40gp7HTmGOuPw1bRtGgwV7x6DyAd/3mTIf00ZUxqAScqIZ/+5RY16WgVcec68IlBuXZ9y8PbuxU
d7utURSAoWXO2NbA939wjZ1J9+U21Vgl6KTA+AsMK8oevimz1EaM5OwBtiHFKEparh2J2j+lxVWZ
QYROosZswljspGflZwghTdl+zW3lJLPHJRI7RUIgB4RvZ32irTlyuEI15WN7hlxETZrVAVfREwdF
jeaxv4pwB45s0lT1Yf4FVW86j5Js8oU2SnNYU2bZhVOxF55bkm6DGByon+em76MjwqohQFfBDoDW
D7GWNwaUT3vee94o+H07EpnBQyHzZVfFmpd9JkCnqxNcSA94xaEtStilya9l33eglwIu01Fb8Dds
4jTfR+c94yQcGm8/GER65jzS7BFrwcVLRoV8ZuxVv+kXIk6uAGEetLe8EfD5V1ISpoUf7Z5UtOtr
k9gxYBeeokw6h7cw3XxI/1p12STluxvSLU+gJN95/OqZ3WRf5BvpqmWhakbutLkhhmlqlB8hGfZ8
4VEvsYHPCgzPnS6trrsO20wj58+dLksFaFPtdVJhXQEBQPG8uWuqqHdFkDOvog8FJb3cRjNu4ZSn
ELKOh8KIc29aWBB1VuaHK+WMThf2okTp9Jhd9E/FBT/Tp2zlWvb2wu+4ckJfDXFvmaKWwZ+Qfwjo
VJdHPudXUOcErCaW5OLeZa8yYkYFxbk1Je0oSMs6NnfYcUA+AkFIG4yCbuQYRKfnWuBmshfmOplK
cUEFmT45X6VNjZvPXGoiy91eMNOZ5XfA//FnArblY4WJfO9K974NKQ5+sKmJBUf4gf2GkWDDzUBE
/FQi96G7XTvE/mOBFBXuzViDUtCQ550NLgmQeUIG/2pAihlyhNfUUr0NugGEWxhORF0n7PX2Yzl/
O0f0NSOcXq6m07nI8+0ULZ2vE8r0uo+Z7a13ADtNH1C6E3jWmqUzVMmZOwgO4QVRG3VbNQ06G0Om
8OFqDHp3EmPvy2j1qqUuHg2bK5ktdZE0hN7+UOoUZBdFFlbdkThMiBot8Q09/nEgPkH+PVqx9ksN
GV9ypoUdw62s2ReDLdGkEBHyXHUEtBo4BBlv3KT8Dey3kT4rML4alwZCqWDP3xfcsb30Svmes15A
Lg1eK+0X/wdCqr+v8ilxwTP5anqCznZ4/xsHaB5L+NIPEIgLC1P65VXHqDE2NuB0bC6Ew0vYqn2L
r/xANUGG0x6P2jk5CK3QO7+ESFVsZ5Zk7pKRQSbwDILuSU+bwouQD9LNfM77pd0EFHe5LVTbahTw
PFJbgwy6/StpWlwji+FQnpAKBDQoZ50xYIk6ybrsj6ie27kXv8lSwLN6KHdyM7sCmmxZWMDD1ALO
ZuKEolzSppaqh9N14/Hj0rPvaG0ML0gG9K5LcteA2DJx8/WRnD4zi5AfKQSdaW0yasrqqE+VrHQs
Df6CIHYC90RyF+4jazpnI23CmFfCpETvC1EdDVvlooHfU/CGnF4gNi4bTH9NMsHw4fWePg21c+oF
8kdN+47fHlqjJqXs0XrPnv+uNLqyZozauuZP3p/cdJA476kF3DOJnh4KEU19nT238EaP7FRtPpeK
8YFNh7qk8cClRJ8GqSqyBBMK9nHYbd2JvjR+ZXCSsX/w1c17xUHI/cZVIc5ExGitkZ2S37YFzBn0
UcE5lMUu4amdACdKY2UxiyjoXLoYrthTwr9o3Evih8Z8D6/WyM8BzhKVApacCcNMAi8iP7/myAte
LwjUi/0WI3bHXhOLG3eGitlC81Q6ZG9JF5SFhRZU/kkrAUa00l0NmUoYKvh604btEMmThZSCzaD7
HlmpQ411hYMQ0ThuAr7MEHlsJwx8xUj0bTRiCXEj5hLmhQrEXccXf+QBMxqYxFQG2R8Sg+qpLpGX
uzvZB2Jbtf7RzTgSSVZ5NJiSCblaOJHSe873ySxT52iT3d9oje61psunsAPzZk4N7BnFJgfcquFc
gyYH+M7V56AF4zonZ/JlUjfoZSLQ5UGDWL70/yDvQoHRls/rqP1qd5QW5CF8hVSk4cnfqCCFpO8C
YdmPTCi1g/HiAB7/TZxNBrklth2VEwYLG6E4v4Dvpc8H2GQ9s9VXnv9iAxQjzDH7+CvHae6s6TlJ
8b7vdEylPnn5KjBqsQ07U2C+Sl4N6q5NaCiwMF4tUVi3/0pfv2qSb/TfBBWkwj/4UBN9BMFZfsax
y7CNy2V6ZeJgSiN6nsAGoinr+4A6Sb4imkkRb1udWbkm8R8YxpRwrWPZTXSsfZZdhd09RJlgrI80
P9m+BoFz3XElMDNmtYXeOqI0tG2IYL8j40sG3GZSTQigDuLHCbJoPsROYF9ApnFdkjC2IVx/4FoL
ywWN1UrivQ5EL8cfpCt9lDZLyFQzxfNu0Nmecv/u+Ispu67ufp1ND8paRp+3L+7iSXpDnpEL65TZ
hQPPQjRv0SRMWrk1asnThAdMVw8n+OuQ7M+U0q36j48gma1lKW5DW/BL3espID8ulB9R0HvKh4Wt
4+jlfAox4B5zUm6vRMo2WQcJrt+6CzNnlT23mZ1cpP8dQ3ZmBFxj92WwBFkeCDa48Q6DuQh9QOcN
X6rrPEgTDe52UNNlEDts9bi6PozsVb9vKtQ01u0Sud+Qgl3BcZUZNziZo7NAVxh/bS5yzfaBviYg
ztEoi5XtJpIBYBxgTAt9buCnqER9urheYhErYglKtc35cEpWD7VkslZi28iBqpI5S7w9RZn1R/q8
J08852i4IOStteu3dSgu8XLtrA5cJJRAESlYgFGLalWyAyO0iaEL5BKWPAwtPsk0nqieEp6pGENN
VLoePaOyY4gssimafbEh06/r214LTJJJojVadEMqV0/rZhvmw87aF8D02iN6fTHWj81NHaNF80pJ
jxwQ1O/5FgRiOUVXgQVXBmKTfPeqNjtxXuMMX+0klSQpI7r2RBB730//PJjQ+GPqFasQqPQoP6AE
L+I2mKi7JFrSNhwRfO60AtD+X9att4GRmKunLnABaBNa96k3IVXfma2AsClCcKHLKUiVI6nOYX0E
Zd7OCT8l4imNl4ZsgJMszjnApM8iB8sC5yE783vAxdFKYteHnLWttbQp+0nwjxA5o6mzD25vI2ad
75fwDIUrwFmd/nV9bwUe7Zbr+aK8WNMgn0PTVkKQgBdom0bkxXHbyEX5u3GDnNQLeOdUfbV3JHSw
18WXYvqxlGPTcPqfafHnAVEk9qGrluJLZ9QQWLTxqZdVNZrn4j4QK/onCURL7rIldb+j3kITtpIT
kz3Q6UwqlJaONaTr0EVA2v728AuINOFAZ09m1up+B60pvQZvz6AsDVBBZ3bcvIY8+5h35wCcDRI0
Y1SoDzdaS92RaxmqK+5W+WxytLEVOdPN5Ofju5WGhJd1VmzfDnZpuaAir/+G/v55NBhzjHtZT3BB
sNMpRuylWYzoV3Z7+3ufqoqTrPVPq1yRZlag5uRFjyNSEGTQvd+zRMeuMZYC4a9rD2W5RioXYO8B
Jjk33vkjwoo/o/GLtST7WcrXo03Tu7mLyiZEJEdkbDyPPE3lPQpJasTUz0jiU6iJrgTwpTRO1ZSt
eo9K8eB0lpeahs/MrJC7O2lZc9uISwPKj3uMO1m3jxYfRuwYeL3EOb3UKNJYNkaOiUz1OIZ7Z8ci
Q3aqdcDMAUH+319esZvkn8tdC5AQLoNzuMPMnPCtYKIe1LqkWzQ2EAyaJI+Q0fY1M6kL7b1zikeK
abYrWa3egLs9hZAz1tJUPEIv36SS9U8zHtXOtqk/UT0TYeWiOfvJXiYUHt+SMmMfUoVOfDxymHFf
ilraaR9kXAwjBNkBjhPbeFmIRs1pzFME08WXlMBFANbITUx4HxpCy3Rf9mkbdM0vpSgOXiNM57OV
/eAITrbBw0t3YnibsqhBbw/TW0/0UgGYVwfR0B+CKRedyqlqF1t/rh7bONb0QG19ApY4mBaCmkAb
NmOQtd6X0pjsgIUm3kpCkfthj1Qo8hA4A9NTfCrDgM5VnG13XfspJBQnv6tpU0/9t9PoLAecR+Xp
HM3eVDUCgA3yzoOuUS8luaidDnVIqSiP1nhhIYEiWnqlZjbKVxV8+yIBff+aoqHKkIxLKIXjjgFp
ZoxeCLVrogYvq9FZH2aI/hTfy/Mxi/lWcTuF/msr9tlvLQbtYMFTFBKtIobvvwxKw9WyjONy5S4f
hTts9YkX5do3tA1B/1UKlbaxM6jrbB2UxqthvMhA3VoSOt/fnVNit9cuWxj4Er3pc6TpbQe/23Ew
Rwe15FtpwNwIyC1zBNMPmthoWhgRarxI8bFTCaFfRQXzFYyRuFTZp+jqYKQc0+M2N6zEmej/dBgR
qASCYYNzMH1lNnQZmYAnL8Lsf2k4SPeLBcEbNlCZLKqmXPTu7xxqY8o4vZxUvqpfDdxeBXsZ8W7T
FBYBiZDSQ3/AiJ1A+xAwqXe4y2PKaL+BadcIr2y423QWuC6S2nrWrDCt1DBpkLy4/QPI7aFtDcMW
OH7okIABKOGk4z5kuGCAb1OuZWyajU6Y4CGzWzW0iN9opjwsQmgaHUj53jQHAulq0C+AYw7h9Gsa
7g5bQizDja4XvCJIOMp7SHDIZk0Fw4wBj0q/DH1GpGwBmf8UTGJd17rMGSMinZ830W7vR7k9x2Zx
njLZEIBetpZ6xcN9OTV8T8KIAUPPK01LWKurQFXeTT0XERrghI2YsNgTwfFxuaJhDzAx9hguNA59
hKEAHFGawbR/SAO32GRUEBBRSC7FE164RWk1+9hWofK17A9yJPveF18OCTBnISU9EPwL2RCeGVgg
wB9ufurz+H6SL5WAZD/o49Vt0QR+MY46J0ITwSXTBw5fLbnSWVgQNCqUmPJ94Tkxq0djgvKU2tEt
F7P96U083BH/iG0h+EC4Aorg2E2WlbidAyayrqmBKQq7YNq41UG1odLhtWmRqI1/CUlShJbMFGwW
ee1UOctm0OLQFB1Asc8oTiN9YIR8qQpngOCaC6INVW33iw/5Oy/Qtl7w6/1+9/HGNUNaXKVTiBRP
VJEdP/Y4ZzsaFhwVizwMAtsWsscQ7hK2VFLb3Vkk4+e89tZpdP8ii+xRarBl58on79yj6eAJUrg5
FzZ/AwIylXQZO8wgdY1nAViNJNoj3rJIoT7JwrVFtydDHEfbVTdey565y5tgOLPk5DEVxEelJnyM
4CBjhqcx1SH6Z3GY7GLvu30WaVW7y9dCmgCeidtmRLyGGlKn1q/f57M/DioiIXnTHV/uGEdFwyOH
B4gJT3vBeZvgSxKPevoQFc9xd2bbke/QkgRtyTW1sMUvU8KSsjeY8Lu8DR21Lu2l9sIMsUtKmkhq
kbEWv9RWBNMxaM3eJD8kcF78N9wUqquxOzOksE7xuMaGFXcavc09ctCIz9p2IlFi64afypFyJHVE
fxZ+5J+cn91JAv7k+p+BRRm0g8olRNBZ1gJE9abtrXbKtxUTkAmlEhCKo9zfdzaiYQQpYx9L1HZp
RI3zqKE8JKHjNZVclzLYkgzHFtu+FKTO7nPsdg4ybkZMuOBZ9U5J1CgBN3lxQ6xAN3rQsnxQMcyi
SZmAd1CG2sOv+Zhr3rpYHjE/zidmHONEmeKyfmMzmgdL1jlBka8KeaePv7d+nVrvz0XEm5udmW2v
2s1GUk+I3gsyLpOL6MoU7bx8I7BoOgg5WEtaQpBqeTjHYWfqKd90jfzSNXsvGJKzBB03At4VKVJ8
VsQES3f9gB+McYAfKeRwEvJcp7BMt6W1E2gM8UcDBguVvrMegMCBoo3D1RKfKdtJTCUgYRt+CgRw
1ClnBhrjAba8KjkQRFp1rw9jgaaMwXhzphZd76jZpINsSWXb/F5r6e0Kqb+w04LLk5oXbILU2uTk
0HH2vtqibxk/tvxZKfokdavJNWyMvKdehFLkRexnIIgxwxWEYS6chFIv9BEccaAiIB5EaxloPzSo
JfB5vrjv9rOiEOW+LEOTW/5RpF60/M0RoZ6/R8Yts39IKGBiF1E6sj1Kt6HyApReASDEi3PlTgj2
8XuYkQqXZKT4/gLzI7hBEe+ZC7RkJq7AYOMnB6cH6rWk/Wb50e312rWUV/iTFG2RRBHw0aU6ctHI
Qc08XxDymbXYUsxLhB7DKRIMb0zFxGH4GcH9YRMuy2GW22DYkUB/Zat372lVwvhRGUW/noGSWCV1
1rUgwys+1xiPbQH6UKSrIRer9VErAjUMWiw1HvWOrsVPnNv/HO1A4kdWgPeaHmvfyzqw2uXlZfP3
uR0DsD1roHE1oc6jTC6HPIg4pka+OJXpA7JwiutWR6pGwkiMPPNgrJ79a/sht0jZk0REaH4ajQJV
H1qOSxIBj1Iya6ak5DDDDm4EBpwck1aCKRrid5R4/0DK+RLauQ6isxcsyfFQ2ogDsND9mvFnST8C
DpIt0gnvsmy7+fUyQXXYDkCMW+KXfpOr8rwEs5qxrMfUp2kULwA1SXKDBfhqPKGFkFoLfHhvZG+o
GZ4LAbfXl9oVv1esZubRg9TMoZgUmGJFIJ4tggwDKW3tk+8OITZ/lFVpJ9O+Z+V//TGdj055Tv6c
0hJ37SiV2YSoqeQ71v/TwAuvHKFk8k4PUE0kMf0rucOdOZgYS5uldbSpIV0H+ZryRvhkDyot0yri
8g/r0N07RgalNTxhPJqX76qYJwpRH5snyyazc41G86KNmmykzafGFKN1VeZsb2APg+36PBhlgOuX
D9NonFqp2Vt2YnJZzHHY7TB3PrIKtGHsGLPz06IEloIL7y2nrntx4akvYt4nk2lqFp3n5jGxiS53
2YPdqj3zeWg3DjdNtUYpaHpg8ZrffWEEW33JHhhO1b3zTPQhBWzumlqkn2CInjwuEhrg5/vpnMi0
fE2u3D90dvTjYUrE/UYj2NHYV1ZEkC5NZvl97W9SIj7nj6S0QPJFSo67lmksTtLn43mpSfNPC6GF
6cJkDv21oFuxc6h7fP41blLLBgZIuFC6LdLVO5AFg5atj0w9Xh6c6p2wLLFCn3LzOqEdYtZOcT+f
uxcJ538NJdVzKft5aE6q0rxcsSIQ5qqXJMxoKPmWQondVHOy3LfQPu7G9lBXIyw2yZ1XXX3lEE6I
ckHSqmsDJas1OTMbz2mSTV9XsnY9UVsGrXZ3e9w8ncQ2TykYvhpXY0lKmhPHTZSHBptIgOQ6AxqD
aCI+KxstbeDl9y6pXSFLJWsZQyIf6cx1uGPERHguYdGss3isJuJ7ByI8alYefVwZ8huajkegprW+
a4wjThAW53nNDTX0ssgfq9ZXJ7ZCg9DCUhEv96q77/xoZYYo6ECjlmxQFfxxejUtQQkAPWL3j10O
Ony9HOoRSyQUBRIikUkMN4YBYm4sSjf4koIYbc4EdrcUM8cheYoXI/oUtkC4FXycAxfeHAzp09sh
EtdjQ8DWS6OxV6VnhAI7xPtCIdBacL8obZon9HtCs/QqzHJk+3fNf6AoXQOFwi/J/gkb3wsZSUtF
0Ptb5DmQ4KBXm6kCXhqM+9/eB4pMHZKUgkHRkSdKfEkiMQcnUC9bZJr0F9PzPxEMxkdOWI1aFdf5
Myu75jG3YLSPpdBilWTZPYzuYgBr+tljGY344wxdExmjnap+g+wy794jFyAaZqv5a5TDOmd4vcdt
c7k83SYm7u1UBJWblSx4KIxTFS797Tp75Rl1XSbbrutGeeR0Q+FzfgEAN5E/FZy2ULaBWQj+G4K/
zLIgaNNuxbbL8AVrdDYuOOKhBIicD5x5oVoFFeTSU5KE79bI/Co1rakwHaJyKaBOyCpm06LMP6zi
IAkA/4f5j7gUg2edykJfHPbsxMewdWOt5IT0wWASnXD/4qKj8bLkimT+bwown3Nka4iUuVwYkjWh
dmXXMO2ABM/pka9gGPeoTlllcpAcXYZrcFRVjuYlPOtu37GrVcYiS2xp16e+2466jk2CFV6GO6Ol
0mjpxHds0eHbUzAvd2CaNRruYgJ5j/UtcLlHyICPZoVuhODXhDl9QCJbrO0T0UR2VaDduiohjdMr
PwrlkHvKSaLuI+tdg3LrqvwYDRij5VsvHPpSV/IIfJMx1ZQ1KOwYoY+bY0KxugpGhWsxcUrZU1sf
4XXLLsAQux4xkxIfJmm6eI4zOjT0E65/yFGs7TNUpIFLrCEdZAYp4Cb4Ia78zY8yXTXhXhcuMLfh
TCTUij2zAMW/fhVO+It/GKNjcUsVytU5RnaR6y/q+wouo6X/vvg9iTrtvDgOx57lPV/+BQiOqJ3n
B/cw00bugm8SISDTmY0gyPG7VX4bVkTTzdmSKfLiS2ajvb1cloTYuOrTEZj5kUZNC4QuWtJy9JO6
5wucaAyfqfJfS3LgSYmKzY2UGKkd3DaA0vvwfa7I1Qyt3F4XKFJqKqKXSWb+3SBWU+sA0Hs8wsKs
F4hQqzWumsQPQXRCdJpSD5cc1/qNfD/QhjESzLi0ZiWEghT6LUwh32jxCe3rWM8yFDgeCyxraeGi
zWxzwIbz65wX3/2WQKaJio2xkxGSDcOnf7KlNtlWhUTO2fxQebHCbuUiEDGVlq0ocA5AJEGH3Q3d
uKqNtMbIuVAhGaC8CH95hhmzheYm1SNo9zlelWuGPBG5kri+mxB0L2RzdwhioTYmnSLAxU226X4B
WsKzTFPpmO6epTl7VsRTIJfXxPMtepqziaTElE5qvKDj4dlAgyTkI+UeWCknLahUee2BoPZt1QZh
yBweW0OZSpiwUOwF2kQtaoackNQGMtByRtKeK80Z6yd7wYL1X5FecwdxNzeswHS00v5l3Sh1Depq
wcJo2cO1GKsnq51z7t9kpbrDcwbu6Lo3jJr9cW7MB7u7Qv/hgKRq18WtjTUp6z1By1NfHeOxS36b
O5J9JoEPJENJZr4G6xwVeBJY5+eLAljavx1AWL1NF2XOdoprwExkUceH9lWvcy8qRIKC11D2P5ws
hlQmwvkydJtiM43mkAj5fGPuOYQe5gaKQS2k2hGyBwo2NSj8qWndVNzoAfKFPHt3cVOQq+MHDJT4
EbP83y7/V3z+Wi8pbtPcr4lZWQvtIvNiDl4k5Bk+nl6oWpBpxs/D8udKa90bN6m/RFWC911oDPXH
/cj85ZAoBoRvDXtrYsu/Mdpi5Er0McGE1X1ir4XNFdtaXiAUAR4g4Dtn9LDduRge+QIwmGMSpemu
KFw8pTasvwXI5vAn7jLb41Xj3DNOxQn34kSvjL4imfUN0XDAyZhY/ZxMXX52/5sbbHeqTm96DPJa
bWgtj7HWJ3HZzdiAWaoLZlLuWd48WzGvPH/ViVVdBgh96Rigj95tw+88Ks+cuQvgvCMOCqhcpeQZ
PnHTQwfXI9GV6q2magn0962KQgKPkxRz/ebl5bj4OzT408yX+Jl5rVk6rc1jjoew+h7HgcD1nklX
HM2l5g14jFiSwIKnUZmstnaxdKdK/ZxJ/9D96qzbWK6VqYjQ7XiGcZFMt7lTNxVy24cX5tvmOdTq
ro/9/qaWBb6Rq9EjPJ/9pyvK+/WFgF0Vwxx3a5ZDXC7MIStA5B+tQL6oCvTPB+47WmgfYcUzLJhH
p/0rUWE9aMtWb6kVfAyJgwT0AbAuno7KQ5IrtHatUvN/7Oivk6tKBkF1D3S9RV/H3e5UWMGtNk5q
jujM4s2RB8BqDVpAS3q6FhVjD/xOJT1AV3X9qyfu0jECzoLE/yVq7tH7rvxFSSBKoG89GaMlXEE8
o6RW+y747hFO0jQOPk8d0KHPilXEsSmDHAAt1yTOztdoo7bBPgkWrGpyuhuykXrCVKE6uoro8dhL
5kRlpitrIoUMs/4U57Wzjz+98ywFOJnvyAxE/KCLszeN5kfSNzk+NGAuXw+qobqUIJA5E/kQn25a
uOzVeqtG8v97pAF4oGOzb381nPUbBJAjQ8W7uYVOJBuxQfD4jnfnqzArCUMoLM8T/syX9ABdzl88
5FPCxiO1Q8c59TDRYK9tRR/CiG1C+CCTIgzqqPNjFIKfRco8fAqP+fKmTnEDXkQtNPSSqIAdoB7Q
XpMb89+8dH2JY29h/CS/G6gMXe6bUIq5PPpvOZOeHTjk3ceecv2nOam1/g6kRP97M53Sp2Ce8uOh
bwd4bx3JeJmbQvnBD7GpO/MfIUA++QsmGSUGCaxQHFD0DPJtIoDC0Ma7Rh1YTPZPDA5g6J1hUNis
px8RVNp8+flEYsn1TXV2BYuzkqdPjFis+fxxYFSYT5HBjxv5xodb4VVUO+6Er5OqeKK1sFKSMLDK
mHMxPnD6mcsGICwxIfFKLL2kzhnYggj0ZNNEB/m8kWgztxIrxJSfy6fEkdUKkktZN/yVihyR/oQ1
njIuYgbXHl1dhf5J4a3hMsvhSTqsIKWypNL/livh9F02AV/trTIZAcgiBTPndME+TV+SJjwP7wK/
Mkbvc8lXuaF+iS58uKe3vX/eqjVcGxGI9qYQbg8LbQMjNVU86py0F6EB3O6JJ6oXMgpWJMxWqAEI
lzpXa9qX+jLuh7wiyuM46LUbLhDrjFGY2a7PjBYl2VH/1Mcju9N7ZlkEX96BpSTJaK7YCgmPZrxm
Ps7BBt49WhmnGPOcPlmqAw5SOtiXewQe2t9z797admSpKYDBbzgLODdhd6RMOCxh0YVx3tJ7v4Ro
RSA0M6SWMru3KpjuGsmgkswfO/5pHlqnAgHglvvPsO2Lulf3FyTi9wG/uT5wuu3bqkRUciERj9vv
LUHdmVezbBjGONyBFNS6ezswcp9lcqnCYGOyOaUAUWHRj2tBsr0uEYfu+j74FofNTSoSLtmXW9W1
n0zMKtAJoMbSnQoXxrmZwFaa8PZ/fRaapkgqjh7Fftb0T0q818YM40P2fqSs66yugv0YMJhJBKSZ
4CcgRLHkaX+dZniGY60re7nmMrDakNd3Z/eBfKB3F58AFEfViIUJ3VnDB6Ii9RKuof/LzhQkYuo6
fD4S9P9LWrBq2qScn5luI3dZlWiZpilXCLbaYEa8JcBTySnOWlnYSz2VI8GVtsF1GtMOezoe6AcL
SOMArtraWxDmLzupfK82VlMSGLwIRaWOyorackQ3OMwCp3GL8yrgGh7PEmFTcYVbmT+N7YM8TUtR
llhiIwK/hgeEusJtT9yxcGspUGqEtdiCI52QzV/fGMF4cYYPA7sU5P1HMYsvgBkMvPnVMJu8sA3b
KK5b7BVR/aKvZLZagSVpLSf0/OaD8awITvAo1QklQXdDRte4a5IzuCTASlmNfXgBboZhvQjNDBtc
+t8OGSvBrFrYRNIRPrcB4n6gJ7Mw3RE3B4ssbf7OTZlEZuF5iW5TuQrGCHHxg6C/fR3ZAoqI4EfV
5SQha4DrOK534h/nX0fcvywJpdlzBKsGwj7no8DS6M3kflP8TUqiHlv3aKSE563EFkqATgkpIW3m
qWOKK3qD7lgk/R2lMcOAqtdm/cwUthRqnLLtbHZ3bUauuoNAQ7lDOIAS+dcrPFI4BgeN25Pva9yS
Mx+HuakIgAoPcTrbnNofWfmzp6/k7S2j3luJsb4Re8kaFejq4IgEIQSNSnNGokAWdhDbsQlS2tPJ
fN0mR5stbV/YNtv8lOym13u68HB4ZgN+aTBbx0klAhVNPEMx50hcw8jx8lnbLy9DyqsGXVdU89sy
iR6wk3qBeL1TQs1W9Zhj6lJz5yYDkotfLbmm+1sR6FnnKT6SE2HJegU0l5fQqbq1/Hl9Zqt5dbgf
2HinZP2X3rbJCDxar/BB3cKYWYK+plb4qChJdG0fKQJm+vClWt5SYkvQEYb0uiu0rsHQD9IZ7+6Y
IpEqE8u6ozylkXahpp2uWI5OZH+s+iOZFn40yZpPaIB3369qIzpsP36OOpPrrygDkBApVW8JJW3D
5Ajq4IwyK+aCuZgKThtR4fBXQVP3qpFWivnxsIbe3Vk24fztXoDjy979cfgTZfXx1zFgtE4IEZVh
a2bPsikZgTXCr0F/ILsg3FtxCoTG0b4x8SRBFWy+M8ovGnK/BXN3DeIJYSIFkHpftRXrhZM/+G55
YosBf94DaDEhfgofS/IfOsByaiL6+M+V1TVJ0DfihW/i29A3nBDoU+3/86kxUfGB0JRto+BfLn9h
CWXeLEZdNodhkoEcTplZvfAEfqlvjhtNUGJ8SfhrxFyQKvCMpUZt3ZwduyiAGWYbNOP4hSDzPMn/
2lJwOxjKCrtg2Xrr/PvCti74f93FASqplHGz8HU6xAQmdqNAkx14Gt7IgMJ7EdzXchcbjFC5Eqxc
QdfQRDUBhTccN/bwWns8L/WCWTz9gzB317ZrsSisNRxH3OAMPsyd8AQFPNIS7P2ftY5gIg3qfOqe
B+fcxdrONFt4lJ4fPuD9Y2pAnt1ti5W198aTNqghD/Yq5RWj6wanysUb7uLOktc0GpaYOZtJt0ls
l8fC3CjeYsSHyWwxiRRRKgAKtmFhyjj+gJZhNOKUC3Rj4svVOdwCCjfMn+fLFZ8Sju4kO6dvhMKB
x4sOd1K2/c7MB/7/2Xp/wuDil8BnWSPeRIXjFOY2VvCl6GkMlH1sdYKW7X/qp3FEC5yGDzJTPkph
cIeJ2Frav4g5VbEz45lskJYuogAPSoGEWBCEMAxVl2Vw862NdpE/F1DvO7Pw+jJsxDwvphR1fxYi
e7h62Tc3G338VsXi03TAI0GD4OSm896lgcvEVvxi1sBnIBRuWKU67tbhmgkSOEYJ/W4GiNmIzNnr
tvo5OMsLDnnCAKrRCBve1WMFQlFDwgd8kerJb6SCCX8i0vVyuq/Yg7bjRSxITfTfP6HlFexOAEns
861w+e2VsOoMLGD4fscmaGRlZcjXN5k6x33rRMm4kbGAx10XmouwskujxFsRZN1YKjJTSpT52FnA
OfhhDIion7H60KJfB7Xh3MvCdGoN3zha4M9En3pPftGgzMb68zFOFefccGu5ARdmp681m0Rpt0Un
xy5pzDBHDbMAdo4AXlAlqfPN6ZEr5pv/a4BhAzb0XzpX0y86Qs7IFVmEESNkCpB9FM4EKAJPYU10
4FblhSmwwb6h1JCgsk0Im3gmxj+A50gFRTKpCNPXz4fUETzxp+UTalKNygx3xGvec2ouHhqSTdiu
jIiGwSzQaYRjWseZn/Z402cEoNMtefemDZLGLOCftprgIgPsc7g7ZCk6+rM0HfNyzNnKDGEAY9dH
wb7fK473hgqw+R0tqSheDaFq8N3W/YTjOXIl9RTRkavzxNwQNKlRuUHXtsLNjqSb403I7a6/5Nis
Iinm+qQISWJUlRwVuUcFRxSJHHvkg3/Kayowl1hiMySXSdzfas6jSHrDpTWN7CXkhDr35t7gerNS
sx09/zWwqTqdk775sJ5ETzek6nI4wg7dBnvbSv3KNxkYGOtEUKmzjVdkdHsGouG+sZn4+amuJRxH
WXlj1iFr98SDF/xGeorNwmNbs/6ZXut9NOiOOwKE7jt2ic/y+xI25S2IkaL6Yua/6fT9cS2Penp+
y+AO3MPR20qho4sXD+/x6cw51sswrDCfXZ21LcbgK5o0OaTp9eovrDsEp3OuRnNdrqpSeLQJG06P
BqBARCaKSCXfcQb8so74Rxw2wdVorpYyxpqONWhCXF76kYZNyislnePJTlGA8pSyledkG5eoV4/g
sq6VVlHkzyF75iuajGK8v+fz72fWfQEfcmCMwLqFSKtMdWq6degrj/bbKEAN5oZlOeWKkqwhbevt
5ewzTh190zyB89BhSP4z+zaQ9rNfoFbnQ3TFz6rg8WzD7abprztsZVvluph4SPMQzA86cgBW9Lul
FnV5D/N+7X3CwXu2Zjq9Yy+RSOaYn+TRR3GZxVTwrOKQFruYkqMPd1Ox10izAzpHdVW+BfNsy+DH
h9LeftkI0vWcZi2y+Dct0t4zIfKBY3H2LRc2tI5bFKykolgo9WHjXHz48TFYVccoxHQqIqYd0ini
V++CKhJKYbMhfn2avKtCFDu9XtmSQw3bHmUHPFWgGfguycpC9ycJlCJIU878VKIMK2+K4x7w4TjF
LH6vBkV+KNmpgQ+XEva2Ki8YnEUZrhCurEvgwdPtR1OZwEdVmjqp5LZRKqtGkjrgWzYMaEbRFP4P
GdYCV4dDNdUqUuNWw0A8PlzicUUhwSXNsYomkdtlt2ieVAzSkRdc12jnv6AJPv42tiBhHABqr0vY
axofO8n+UhoqzdShDYQQHoXwB9n+4ldRB6RT92Ledrk1otnDgBXhXVTuinBQWT9HmY3WfKBeMTHP
AsYky6xl0ELGW2EDZ30IelCt824+gC1Gm8cF5C9gkE7qIFiFIOGvKz6iPQxkK37KFd2nob67S8TN
9G6QiDXsB0HGyGcpdjXO/n55QJRsvoIfTc5NcXtdcBFCynVLRh5Pc+4on5Y5bCWpS0b01ZHP3NcX
WTw1uSWXyIjfK4q8XLal4IE6WfH14TaJ7vjV6pnNHfQH2G5uYeHibSwmVlqGZgtb0+EK1oKXPu+D
hbxOkJF1gz6fqxdbcMalVUU+GddRWpk4VJBDWBYBv+UeG9TpCKR1lLNLIR7K/6eDCZJT9M1AWhqc
DoJJtVlpgmN9JuF4J1uWiDZvfmvs7wXizECIhPxv3mr5SvrNlddxq4mbsI17Br+/cIH2t1FGKFtp
Mi6ix5ZMs31EbnJhA1BWp4SQ0QGFs9kPMZpRvGBe2cYn6YurXlN30lwReZFUAicU/Stpil5eKSRd
UR5Eyxuv7r1MU8i2Zn8WRGzV5o3CLbVOsnnBhR8hCIXfhEUrdctUWHWQQo9n6UsKUZ/VZRx+wKKi
XoWfUI0UoS7ibzCw80lX4M3DkVk0A20xR5nja4SKXobrY11RORlAvCfT+vNwjLQ3COT3bnQ/a3vS
zgMtQ+vdjYZ4az1VnScRugHgf7T1viscbgp6uH71ctP+2MwcpCbAkb3WJG5VzUUodmOlXO8kvkFP
pHMIfCvoKfVskmQ4teieVvhZCTqlYmhuseRyN+L/kcEVuJqyPg/DLDwJ7aroy2utwZfYElp+Pqdl
OYoCkJt0gYXred/JpfTjqqU76B7pEpIFodXk42rv397a/GA3Fq/8N+YknqrSgdyT/PMyCVyjFSJS
jQSHIoVnPSU3P6nN+XUmdOnzSqRD9qXaleVBtHLnMslP8raAJluhtVf2C/Sk4kV31rcL+Auz6Txd
ASkm+5XgtjUf1UfXWk6ECB+ZwMyCd6Jnh3cv6K8khU11/YreparIlShQu9kbhi1aL+XYMNXM759N
UBabeHXWvA/wQGGPsmwvwMR0AeSC/em2k17ws/UeLxrvwctmxfptLOWXNoM0LmVKMGNTHwKr4XWv
bLEgq0mH6XcqybkDNneh52lwDHMMDQmnYjljVLRUB6giR9ApBjTJrMdbMd5+KDsDq1EMurPEO4OB
d33IGJozTDnQoJeUVUwlkEIIUQ5KKOU3BTkDaArdSLsLyUqCwxTMkTHdIjtL4kAx+5RSft+H39u3
pCtojj9wVmIgcoY/obDc7opKdwXVhnleiLUJmvhWObimuZ4mt7oIi/aXwwFlDtUJplI0e00c8HGX
EX0C7TrmFsjOUe+eYysq+kyTg8Gz1Nuq3uwN+Z+OkAcXsmDVDuQI0oBxoy5OCP0lWUJFXGD/dMuB
4EsUt87wh/+WME6tyR4O7YpN/fBNonAkjUwv32aymfBux5x1g2i2c7D/Ckfcz1XmXbbzWcXEtp7S
ZONPkDkx/kconu9To8xIvjAiEbAauLjcyD0d3mKLicqnFaTWQ3oXlPh9w4cXD/szmDCQeI2CQgST
3n/tzH3oENnx3txm0HFKXrn+QFlDHneWhe7ryH7I+jPkdgbTtzxU5rrJDWAS20Q2a1r1q8WxVZPk
9chCzHJT0beCo9qzDeG4VcLtXRo6wVBUDa8p4MLycTxTlbmodVZWMgdN3bQ2x5jsZ2DNp4s7WkDX
tzt233/KrnviWtDPKvg575Yz9PTaWhWUDRXzp6zNyaBSy7ar/baC5e5g5SvOIgG6ckVO9pPcKIQ3
O63AXwZgzbI3bNd6i7WK1Gu1ypkG1QgUoEPTiWXdpeBBl+OCCCxABVoWunQxLeWmL+IGxMN2UjAP
0+4SLsOUmaTFiodmkc3QCg3kyQGV4u/QEQNKRAteVxpLtbIKW5e36BFjZbkjlaZ/x5qhR5ot2aUU
FSpWRZsDROnFSJs5zVrDc1xEA7YM5WoxyNGpa3rr4HtGVEIt2oJGFP5UzmriHC/bzWdT7nt+TlVq
LXdXaFy3REeK9S6QZk9WtKV/z8pllSsATYcsSFTeJIGQLjR7fBCWla4S6QHNhcDwXd3O+f4r9VKK
q4k+govzzUltGWsyjX7Mv6gulCe4O/WeZ3UOQYbreJ4Ua1/n5ZhT1YpyooIbDBgpGNCP2yybXkgG
eHgsOSplNCrhUl0t9LK0l2AV1l2F7TbX1JXd6NKD6PpU/vsUvs4L/H0jp4L2zBGXgFTtbbJN054E
p/+tVo2fIExU2pFVQ9n3/ZAFkY7+h9rZIsASE9k9fD8i21QB3ojISoCCFWfdbMIr0lwJBS+475PK
b04e9MTRj0t1gb6k2I7wJYlokf/a5aH2MXZKTsUFNOawERWhvCSCzmBrVaqFQinatBiswMeImStA
KZNe7ibx+OvyyIudiXMCZ0Exg22R3HAd38df7sCak1fMYZc0D1xTWF/ote5Fb29rY4disch9owAl
QXyJmxNZ0vVF3plaJWAEKxL2mw6k3ne3qU9trMAAVf1//geVFWpvMztoHkTLCU5yD7CYFQvC60aI
oeH6ihUd2/hCDalKBZ9g7N7OX8ZaH63K5OwgLr8HmsqE8hEEtpxR8F8cuiBcHahqIOY73GBUungH
0CDx/zqhPqoFkLYj/uVtp6dZJ6vKG11tYXQ2Z3aWeoV2l3aNKykso75y6hGiRTWawLxmvOj7FSug
3XSbQXY6ACtMVpbUiBNktXZoPjC0KgdcibY5S8k5FspQsOr4cAUe8lXoz82FVuwc3xDB0JmFwD9J
wlQvJoxX4N84y08w8KTE39TDYK+heVIyidS4Dp6FpnxGexy/L636XDiN93NGZdGos6lpTLK+ARvH
CX2YOhYrKFkEYOpF0G9ulMCI2YqvsIOcplZhamvu9a1pklBdAcJpLKSNfLYnt5jWs0S5/rkjxdJF
GM9rstYEWs090PTOOqrFgPQzxZ9XVnMOsdRJm5ck/AwOnhxgZN1IDvd5+isBiuVLU6E6Klb0iC5+
E+4HPvEA8wZ7sRpKv84ytR0kT3bnQWMf0KcgKZM5PWiFzyBDnOWW5YEBiMS32htBUeWLMTRssp2p
pR3N7FEtGybUDhO/zH9Eo4EVD+GAzA5lLHngEzDrhrDbIQO/5vD0rYxYYbwK5wjtVycNT0eIbGUH
AX8AyTpxcYCLsTmu3hAkRbEt7QrX+6jjiX9jhIAdHP+F52Fo6iZu/rlm9HTSIERRSp9l80cFGemX
Pgyre/WAlhtTygopIp0pVPaAcNRhn9954qop7Rml+IeAmcK6OAwoV9bExZORhwq/vVAIdhVtmrKL
d+urBtjgH4LAJJHlOAQpG2Gpe78FllREiHykfhSgBC2Pq1gRxS6YiEmvreD5RAuiFO4rR0MWuK50
+xJUMT+3idiyWG4Vdk4ZJNzQQ/rM3o0J/vMa9xcrDNj+Br+2Uqvt8A+xZVrtSnNz/qYr7GhAVyZu
sewoKgTJPsOA4tDXzZtvXQH6pvsp7IcDE/HiOAh9zmkHgAg6MVNOcHTbBZbsEsDB3i6v069K9XKe
k3xGJrI7bWHE+VqzHLp3ypDm34bu/MmvwEbtmgUG036YfaZIW73uUG22MZzlOrI38wBIsEAkFlIx
Yd0VvN0RvAyZOH00dLJRKO43r/iCdkEPSrND6mWOn8rQ7P1+dZ62N9BFahKGPffPDpq9MSW+Ypmk
mZV/EoOje19Zh+J2CyU6HKfXJmFhzLK1f3t76owrvUCssW6MbY6GKd+jL8fwiuhBWQaa+5AUh3sS
KNuEH7OibYRySXxfAFmSpDsmmW4pOSaxoDQys+48VAr0tn1aoJPizhefJs+kIxjc0XGQDQCjoA5U
MqoIUGeZKtRbI5gk0Nlii9cAD2F41XGAVWkp7w1O1xKT+7z8VOYT4rpE5DtxNPb8hdpNbf7mkCsF
Ld3xG+ffdoSkM1Go0rHKpSK0y7yYaq8H4DMGxXB7zi3WAWtuzyAsaXiN6q+zr7m9dW4ASIeWYVFP
zwaKgtoijNeFwNhp52m1xv6A9YZwBwMzdtSrPqObrZiDiC7fCbp1sLlMu5m9zctv0IcMSuKEO5hS
2UcYmc5zXkMU3FaNp8k4JHfWsSIZNJXOGQT8nEHAiJttkItNzwJTc6Uyw/dEu0+MTBqtAx7QZzYr
7KnAwdQ6EAOPr6EGgaj9vr5jVnLvA5Eu3vmV9ngtPrq2QqsixoTO1EHRa3jAochrLo7LrYqq+VDf
N1EPRBpwHxtlWbUQ7502MQMaC5Z3h7zPC577cyFcbGiKMwf4CA0POUsE1BEpRYw7kvr2e4ncjGNl
rlWa7KOq59mUbKm/uCLwNsQhbPFN5c6llruFL3H98u6leX/KwlDV6UkNBoV7HqWimnuyyv3cwtwB
2hT/touAvkA3QgW4CP07tNqffIaOAYwcZfSTsspx8uveVxAeSvr/mOZGEDBPs8YLA3Ngb+XR30z5
/fGH5eynJNNPKR1DWaD5HzaGkxPExG994wmE6znD5Qsjd9ldsR6Ak2G8RDRxirdUPJx3tnPJDUyl
90pc87gqJU0U2WCWikH58nlReYZq/zGMGjXaXn4ytKcCJmIsSDMhsPd1gCWyl5lrFR4daYfax8kG
XsK2o17A0Dm10NXwiZL3XxifX4AFSz7ClrimxIQkb0AC684zVXby8r6zxWajyAqOGeTOqmw9Q+3Q
79MpL6Rbx04suDzv6wFR5VdiMoAcUbpLTC0D1cKHCMBojlwxadQESSKSUm+wvDKqQgFLD7gfmWWT
ncqV9uXXKt1afJj7+BWTvuLNWgXGjqcPGLXzCHjJffo5Kg6E4vfD7xfSqtl5XHT3k9n1QEwcS10o
pLpEM+uP1gAg2YWKQZbQTHfFotuKU9dzAkdTUNH3sbWG2MaIgGQ31L1+0AhLkv5n7yMoOpQ1odip
DV2nwt29nlQJ5W1q+4ebnMwGy5D0H2FYtas98+yFSAELIH1Kw+1gD/a3FLL3UKFCX6ticcV0+Tzc
g+WKt5m/TonRBoT4BILRZ2DhlrRnbSKpPX/+hzENhkqA9+JxoTRAWmFm0Qz8+tUrgIrNEX8rRKZJ
QGJBxA7jNrc6NxY8qp7VxglY2eBznQWvtD2gLdea+M3xOW8eczCx+xcTOYIwa9WOWWFty7EtnfUf
JX8H2uJG56j+d9Qb0iwfcgSCEop2mk7Q5avcCh3swq3mb3Yjy1IWNg3pTfna0IbMzZWxE3T7Auc8
yyn9B2n7WkHpZJ8HVH/F/4kk2t4jHKWnUmua2taqvYcXQoCr9ot96UUdchv6liEx7JqOVLykmhUm
aKkdNXNS9whDgHj6YAe3+83wO6lBb6WgKqhVpGCwOr2laQF4itxC9YmaRabOxEvONuPa1p/Q6w0Z
IrZnCKV9f4FhOQYtRR20IQj0apoQ9czEjP3anfeLXjOl/5lekVmFt2cSUVZbw24crgA6C8tOYIas
u7D2pCQGLSW4Pvv1SKuFA8WQLN+qQKouIYeseYWn+PvYKwgdO9wRUfzLdhTABbT4CqD90cODeAUw
dtcLT3Lhe+1/SqUT+34LXTUZa2Zil7pLknjMbRtTN6Dkaltmk/1AfyES3r1tLAtEXx8bf7iE3o7d
6ob3dnWyNGrzBBOF2fooxcFofBc+Hi+w+q37qEk8AMaR6LU4m3pTJTHD/D5hDEF5j07JK4wdJHnf
2BXNn8n3w+HQU+71Bii+xCWyaOuTQ3u36CtJEH0tf+A8DE2ge+gaiQIfS69Fx2gf5iuGyeBvNScB
NGAYTJIKcgUcgrGOYtmLMO+BzdSFWsGXDMwkqI3UtWh1Rd/nLHprsGTyY9pwJlNtDFDH6x6WRDx+
soE3e2xW+wVNocmnxg18G4enJQDmdb8dFLWI/UXtHWUeNyJMJDF9zv+lj5THtIMtaLwPTRdh/1I6
XgQmWvKf+lBTVPYaxPBsNKzVSZ/oFNg/QAaarkQfP7GJ+itn352ezWtmyGHNWQdvdf5aEKzIW5i6
g4mvgp5EgKXrVCEDl/sdy5hr13pXRd0znAQuGAKMr4yzp8T9aK24bo5RzVt9BzGD7+N9OBxqHWFv
VCxngVq2zKIv3Od9IT+GjkQzGDUv9tEldhUt3lyyUtdUw7MTy7GW9guaZKzwHeCWxHZgTXcXaaD4
RiSNpc3Kwd0PfOK07XyjbqzXDwPOK/xz2y8kA4fMhbN1BBZczVgYb9Ti2bLdkQAl8SkeK2HW+/hI
diVLryry89Ay3lO5ioguaM5tgj2sDzpsDPJE9ziZqoB1pzoul4+eLqlFlxM23RuzVBVKtbdYFz+O
hMfK2HO49UnsB7yPENMNW8Civ7Vt1drdQc5i+dASbLEb11YPoKd/yKkUUnJrF/tmWsCqEeCEe+T/
ov7gizg3a3iUJrBDtgSPHR6ApIhR3yaRCjEiCEcH6cV+gqWsUcb1pXGQb9OTjCJsigfzEH4PEWWC
ST+06ZsHJNHHWkzCbBYz4CDQmgEbTD/djL+q1roLKrPweoHKTDIenjehne27BvUR5xkocmHe9h1d
JngfVFqOuB5enlumrnhAYxsbMPI+i6zsKfjnJYUddeBF4hY6ED4vb4IqUWXU1owfP8YgjR/ve4w0
irK7W3i9JWg18cWypwA1rTXwANRZPY5+F/SQ1uSDKQ4D93bRRG0NuygG6pKiPznFc1A1j09De9v3
88e4Exscxvh6sJaAXG7RDAC30LlkL2lp9USp9gWDuRU2MQ5jxUpSSEWW7rWcY4BcS3trLqIJy4Y2
s0feAsOWD9MzTNY2sOrjsVYZYBtTetjix4gUW7UGtQx6283omQvSpoewrBhWWVZytvL2/XiFb545
VcmmnMtip8iVTBt9f5Zawi2Uo7LqJzHLmiltuupIW1kTd/Scy2j46zVR4cAmkHV7nJ+C8mT8hg+0
RUGF/7npMzBEIEexHSO0aufoDN/w6PzTZQc8bc5VFa+dPl1AaV+8GHqtHx6QFBa6HXwiKO3nJllL
cfbfq12j4Csj7FWRh5GnK5DcdEmP58jvbaG1AIV49XuQL81A1U9PK+578zTjMudWc9KtU/Hwcr8I
Ka7pp4VcWHf1++/u4s8LR0vot5uu1O+nmM8UbiP1U16Lpzjcabdyr495m46v7DHcKDrM+QUWPGXd
mi2f3tOmEW9HXYdJVYN0EyZYk74Qd0RmikOz31IBvE8jzpWsQm1aJ3GlNDv7k5Atb70N0hQLdP1D
PZeutI+p595bpRDGKqZIV8e0pcnwBKMJXr5sftxe+2mSxTdEe8PFD39ocnu4P9RjOahs+0tdOfMI
BJBBQiRT83TCg/uNOxjhbwXK+5DmUKNVhsjEOm9xnuCHX+Ca/NdtSkYRywttrhOUKoioMWhMXOZD
UtvZH6s5RIZDdejCquhwTHAuyz4VvGnyikaKMFLsHTd50iMJN8zOTKTfCmtXlSWEaI4XkYcBkO5/
LoIqVKVkBBqfRwZnuxYinJBkcbgtRtlJPe0KiN/KPWnCdRk2mW8JE6TYzJl2cQGfPohtAPH7UvX/
zSLigsm4fWs9CTSAsehqJFINozuNWMpAksF4u+fCX06P2sg+GsnShwVVW6sQiyrmdurAjuEWY8Me
Vhbi5LSAXAbOIGSyyRMlFugLyM11k7TZDdc5Ok9B/XyDhSFqYNHwmrV0ssdxFt72foq4Iwa3xrOS
DS4GVN7dEw7R1Mzs84j4aeYMuC02u+MBvif3G3c1eZUvvMPlS1v65ntZ+Gf2Xtrmapo8mc0amixs
1Lals+XOE6ztlEw5n/b8KrcGucUbwKhk10ppKZ/jqV0db1rh1oOLboRaNQgSe8TnlusabkqdPuBa
v3I+kUCwJWNnyzXCjhJ1m67PlnQNhTftkt300hOcXG3Vj5wcD8iDBcbNlVQgmieFRaZOexwiqkyE
BQQ8TGdATm1e7TpkJ8UHt0Q37koATEN5tajMul7v0lqtaoqRAsPDHGkRSLl9UCQs86gt6TAVv9/4
CKuzhI1KleRcG1iahg4Nk/n+Imo75dRjB27zkJMq0qqqVs2Vp7HgwCJpqo3+8A+Xyz4T0vUDOyC3
6XuU5I+UnSp+xykYjjZDTW/3/7SHP6Tbid9wdQkqcwLI5m1zhYv9rzz/rVA0DK6/OklGJ5fnLSmt
gPbUwEUFQLGtiM7bw1U4irbJRj4XdniRugcPB/1HN3zhp3FOxihy/EG+gg+JvngNpie471TYYV3o
WSbaScMA1Xl/OgXmUTkSgqsi3nbybcpLeQI02NIKG3iJ/2tqr5wF4kpE+sU08AYz06vZ8U0UX17o
DVuF8ejGtWP3RzXYyBMmepHUBboQh7R13CqhKG1pCXxBq7ZmeMwlpfmejCjlSwGeyBRHWRdrUq6+
gzYgRL8xfAedendK17mANkdq7LLiWGW5Buht9OHpe5sXZvU/Wx4jGuCpbRyNKTMHj6Jbyu7kic41
9ZEKczWJHTz1nCjEf4wt/QBxff2ZtaizgBhjnzW0mNq5eSxuyOemrztAXrLmrJGxRMJTtNV96gqB
EtBzCa+bJVOks0o6Kvp9pp8mv81CTs6Cvp+X9/BiHXlu+Ai7LkKzlphskJAht85JjDZ32/xNvTMO
2os5MwTyS9wJpgKS8aaWsbdU5suPIbAkM/iZBsP1MVtvUr+BssXptXcTh+A8vkXpGVUYQ072meQp
OQ6GzsO/bLW8slFnQyAyVfjdwDw9imhVJvSQWb4/1jJSjdcD5MJInuqgCf/we6HW1dLNsiTIjjod
sMv6si24DI2njcaofyaSa1iriVV44XUAtpdhDcoGX3JhD8FSs8fF1Tuvp/DvldbdRSAv1sPzNIvC
MmCix9MhOwPxbLQAY0mWrQ7z57XHa4oZBVB7yhQpZQQOxsZfN3/KyNE4zanpgLL2iMgGtNcCBU6P
cj8cp0PNX+FYsWh47KxbL+iAJ2UztLK4t9JBirNfXmYW4pC+I4ME5o56sL5BB/JeRi0GRSoPGHjJ
LIFcTjbh8XLVZqb5SBNI20Y2k+TtCyxM+tiidGgfuF3AZ7xCy1YpQbsJaSSKVR0xxL1Fpx/fChiT
CwAxRNZyhyf0Fp8EmQmtN87IiP+EPbXmWTMSzs/ahS7dE0aV/vpYM1OMqxy38pKtEI4AITJTSdu7
4GTzmbpmnNUF8aSM6QBfWGTBoomM/5h9Kyiqdzh9Zljb3kGGOB37E8q9v9hBy3QzEEtvVRNZxEnl
zjOlZ9cqT9U9fqxBPmQTJH2mH7YhdJW62a8Pjb+BqZSGR1tCFpCyDE7mZbTw5Mjd6U++KP3mGjbm
AzOKg9/6iNh0Ue2+WES/CFE09kJi4v1tJecVnxt2D+JhCRvLg08a8YsArwHbIV6OidNQhX2cSti0
li+0cpPPaDKYTyznFZq2Z/duxIRpOUMZEki7KF9FPxv+ufdDdBeAR7AHlFwHWtoYXL6NutVtaA9I
ZrGl56vFZdoBFOzY4JjaT87t6pcVPiJXgGvsdaJ8OPweVJ43vWD9d35wbg1wPop3KfP1aUJIBQ6B
jA6u+LhKlcvxGlFf9oAvCEyekFpuInMbg5zObTxZcxCSDRMINg6wn+rw6HdrOApCTHuFN9hvVknw
CsL9xN61d7PucPpa4D/eVmVpYKW/qBctgnnRAUGFT05wTPU3AUgoVCuabjTp2PnUdkNlq0T0kOfI
C+qOzFvgu2qt3nA2/r8WpDPdS6GWbCPbPqkvruRS5wISEPchDaosYp2z1xINZ8yHteXbixaTXZrg
7G6rD+fwCtYPEMYuvS2BykW+a9KFaxXWLtWUW+VuwGxUvPUuX+RP//nARrJ0QtDGXMnK0sDalpo3
P9J9FXzxGmof0Xi9VOYY7ceGb8OXOQxzp/T69VUA1b9F3+L/9F2bS5C/sqhHspz1mDNtkU7x8A1l
avI5GPOY4qOjfDNlkPJVL4TV/J/RU52Fk8ckV0Z2fBcubMXf4jJPsswXmkCKJiV2PdfsPA4jr9Px
B0WfyEkZO9UawABg9IawfVhy1FChCBqPwFjwjAPC/WnHrIw14gev7gB43oP0mhVMgd4Jw5KOGh6w
5IH0arVni4N3Swvber2SXdyCGKHcw8V2mTfGphVpBQeAtO5iKDItKvPgBdYYyg7YpY/VKTXqxdAd
eF+4VBs69+mu2LFTPvTO6H8vHtIvhQOGrVuOIL1lwpx5EW3pGwsll+MEnKWrPCMuzWEtojgDbOSj
9Gh5V34ck72S7dJty6DlRlaPO0CLSlJmhOyt3RjuEJJA2CelFEN4gmolV2oYpswG3Rq8WSRPnC4n
VwdHo4VuK1/Af8gw2C/csEoZ/eNUqEThRA/b/7vXWs0KHsmuGMxu0wBfr5a90vlWv3N29HY6p4cv
VUFmcWzx6ko+4sMkoFdjrftTvJE/a0pmTastOGBpSXffYX7MOopAwVlfwgON76K75h4/rIZowAY1
8nPdebOagVMXUeFK0EpVJISiZissUeHLXkClrp2m/yBU6ukqiCBBuQvftGvCJw6we5JNenOqbjYO
SRVwnZUsnxr5vPDgWR1qxxN7R7EmU5RD7ezW+4MhSQWBwX3KoG17ufqimJUG48/szpe9Mu1PPW6R
omQGlFGiGfKfLC/Jcn45joO5BVlateQuBfawEjugdkfzxomgMb69h/3cKcZVc+Tnujms3O9fN+pV
m2MYxCKv3lgPX+qjWIEfgecQeRsm7zh3gMMTU5SuHmC2LKgoB4ZL8RgH1UoLNvWuOFETVv0ady08
Ejtd6C3wSc1NKFZ/tBDcUyhG0rEboZ5MC0ZXzD4KKpKBdcNsJdDNv+iajuoEMQ6ac+2Hpog8ou9F
I4U7rshFxemtUDMcwl+neEsZRu7jdQtkUuOuYNgxpiWjuotR2leEQr1mlCyjeHP2RaEJ7fmFIyDi
q/GdD+JqeR58jQ7UUpMmlD/q1K87npssLCbMawlWEl5bJAHd8KIukR4UNT+xdMMymlL8UYL8f94L
DwDJ6rSXW4t591fjuO+/TUmXORPcXs6FXpIGil2qkqeNaK/mPsODQNidtbaAzIYF6eLN8VNCe9MV
0p2ZmB8Ks/2r2L9b3P0azCB+9ATXt0ZEPNPeFSjgvkAuO48t0qb5ucs6bu8g+gxZk2+v41U7xyxf
1wNce/NaejIO1/yc9i7lXVkO2HPWi8x1FJTYw6bKzw0Mgy22Mwz4SPif78yl3oWyDxBA8S31HBxi
InRmxLCoJQkS29NzqfN1VUYPBLeb5KFac+k8FuorjXsdKDiwRTLVXFbyVhuIzNFVTgqfvDuTWbFL
24/0DrabqVg31Zx9/hyrYajKjLvvc/i4k98emg5bYem0p1+dW0uG0eI/WK33cN8L3AiMJR/EA5XX
a/2aBoZpGUxYftynX0ppIGQfmNHsf/jmIgsZeztHgXzV07oclkskvtAh+jJCoQdpTbHwiW77zyJG
FcW9BwkPA++XDzKlKz58Tj4g0+ca/vJpuY+Dfh4dV6WIqxTuhmCykXWUNJDJrwpaICfblOp3o474
x6EbwbMw4lLZDKyhmavS08RAttcpb41lOZPo9PefrjG5mt+TU5tBQMYkO5Wn2H8mmtBORoNDahHz
DKHVMv62jZExAcNcieySReZqG0zjlkzha7d/HDaZP4KAYT2SGvoDnjyR7aD1pI1gFTyBxeSHlQZC
HvJrwmUsFPK7FezS7mEnxINH+C1iV94deBGgoYhtG5Bfi8nQcSkh3g4OBdJ/BY4B+jQ6bqjcgCAI
kdTUhy4z07gy6fzB8Vr8qVNcZiPS9UQjdnRAfeEhco+gT+2vap5baTYmcvWOzRD/Kc7YsXsG5d3v
V4Z7EQuosK14Zz6dfTmEothAWv3+0WzVtg3ktdKkSr41JjdUSUStyAAV5GXOrIR31LoTDr9ZwAQ/
jZ+TrR02R8Xm3hBfpGZCryWzZO+fG5oDxmJyxLVSBDD9SbifJX/W8PJkxxh2KEMxzzhOlQRYW2+4
QlnhI+GocZvBo9l5y8E8eQxSaZ7qYRBKF2Q73XitVetOy10FLkPsGZC7Il8QTma3te1PiHlTrR7c
gh4FYd3AvY2KlyqbwLRyG4TO1NI4dDtq7X5hhspEJvFKwPiR+b2eVbgdEWKzF0nIb7cncA9Es8wi
gPQWudrQcGozuP7qLBIHHKGBXYTlqdVvrCZP38QkkvqtWzssdNzPywg0csCQCuiJcCHsZufPAFgk
vy/WK+BFacLe9ltARLODNvYzDBXCbTtoV4/DdIgyMCWZ5YyslMI6ebmr4idCLlmZ6DuMma6DXYiL
X+KKL1GdFyZLK8mzGdKiz4lWYq4CbvpPSxAUx5/yrEU3gFXL0hgiQ5QdlbXMt3Nl+PfI7UxVJ5Xj
+I9YG7UpHq96nHrDJGYy5sStuaUw+ga2wwZRzby8vh/CL39p6W3ScjIkX0ZCDxt1rNrSZIh3O5Cz
Hby5d079/MOL237CMUydjQo3N8YJGXeiKIZjusOtCErH+SApq2R5ql0EnamIfZLY9S2Qxo9cRFRT
+EZyYKgzbjDOObAvb1iSMgEJmt80SqfxWrVfPd/+SyQnoKA0rUk0yMQO0S6hORpCrQat0MR3dvay
jqvsGGWT/fY2I6L+zKsrRQbSGBJYroEyvYZwaC1zIwxPTRzQM0iOEN6gdKnUBbAG0x4OBaxxU6zK
bsuTv11QvOz9RGixxUnJch62caf1DT7Pug5xb5iNxIj6XSqs6eRRxL9CNfxWFRaZ0AmUivRjohMA
8lGWxjW3KxFZAz2Pb9gSNETrTzVwmzdw0xSELLTx8asDkf9TH32zjS8N6aRITBmPAY6wM1S2hUBP
Pc4Bdm/6+MR6ju01LaShN+wb6D3bBCbDYgB840e992r5O8TPX7hR8XWaoBP9KoI/09C5lfRoQu1j
5o5xaFVUymANHfdT8c4CG413OjYqBIVn+U+lnz4RbD5ovMWWJQaTs8tUVT2lx+9Vz3mACkAbjb/V
Qv2vv9y3vC84IVgZCXK7m+Vv8ruGvxAG1xH7qf1c+iu2PiCTAx8lclPcovaOlqSsxSK+RZLrSlA1
9LZV8Qj4pO3uLqsEMAONr4N/JH849tSmXl/42kmaI3w+xjXERDpfVJtn3JmffleZF5zdbjYfHFFD
QmWBN6rKTER2aNEGSJ09UU1ciBdD2gGekLc8hegUgJzmI4RRLAGGOvmuZ7iwoVHCkLScgF3EQDE2
15aYWzdppt/dwmdfr7CAnv4Kn0HU8rilrPNkBbBD7bEVmmJoMWm2cdyVcR+Y0Y0oDTNy/izj1Ang
DQN6xxJR1ANX8K0scviYjftramU7kUHMFbj5Hbk+yH+tUp6+hGLnGhxIKM7psRKejD4g6wQ9QkVi
a7m7DjiAtoxr1MIi9VdMP9ZUKpo/aUJnbb0/suqS29LL/ULZaK2uXMESKHAQ808mfH6GBEf1I1rZ
NkHln0yiozQ9jt03l/l1G+ikOlyfu7da3ZdL3ElX9J4M9KCBCAy/PUc3MCzNuXZfDL/W7muEzdX3
44wJtf+Igou8RQD/w1eEUCSFre60wvnR1JmPbxDt8E9F7U3yaXWtI6vIJlvt4q/QfZ/o8QtXH1qp
N1eUz25QIuXqJ/g/cE+NT8r3KEpzYM9y7ay7BRNOrYRl5EPvrtkPk35PxGsOOn22S0RMaHA3JDqZ
VqKWKk4MtyLQnOo6Fqg3SvJO/aFfB1DDh/CtIr/CyZvoQKqEJAQw77WCcXuSbtKhbQG9e2/5ksQO
kFnqfPUSB47HEeuPqAgHs9KNOnXM/UqKHMhyiUrJcfU64YR8sVs7tCN+Ow6ZmhacYf90NlJXKDgv
gE0j4BsDiM6HGZS1ZLVku2thv6tpFryNxRQ99bsCJ1hsP28BM7f90ydiHlFisLeXBg73wefeyInh
igEdzl+tUT3w9/vFI7U3wTv9EV1m+y3NKxxFV464PmRv0zj06E9rhikKFDy1Jhbgj4MIXDaE1laU
JF62OLeezCeaa76tTJ+mboCsf6U7/kGkfKhduH0gZAQXEoNUDQksfeZFA30k9yoKY/lFWOz3+5I5
WLsqK4wEj5kwv3VpoqbHn3fSqZZXP7JOBKiCJQ+XSf+RWi0aE5+JoZFyZqGdu8jxgsui/XmgP1rJ
nuuMPO0JiqZDI2Gwn6n/FbxX0iuNIPyebC3bnSYfwfXx51mh1YIRhhAihxQkBsdtN+yICTFNsKCg
30KJAKesQ2z4G1oiN/0qsOSSDinvy3RrrWdEyXD63oMuH743m0Z0zvJx6fiZXlBfdYIgT2HNWwfm
DI0m8UPpnoToT/hPiRh4svhj84cpjU7kYLZf4KDYjVL0lUAoQCfapOTPBeSbfS5m56afdW6pK9wZ
GzbXB8nlECcZVJK8pSjdCB0U+7PeE2uDCf4MNT96PPNATD6xzkjuBRuv/zpkonk7z781a0TPUW5F
pSYuFYFzPmwbFE6pUypXg2MGTFD79Bo9k3I0GmaDmItAeiyEGhABfnz/olMTa0eSaotlJLNRIY8V
MCotq8HZ7X+XzyLZ8yhhVVphYQ0XWVJ4zKQSHisa7NibAFbMC6xQziuEHRZClPYRoiMkkkMY3VB+
HlWLu/XkVcOv7wNpCAVrx7BT32Oet3oQfaI+k3zAorPB7IAr9My0IdiBL30QB8Wzs36XhZ1Mm1wg
F73EotoWMuwDlrvpeF5SwGrzAFqHLzp5kapLZnCD1+aTywwro/VYqizO4afR5Bp7fvdGtUqQST+G
0YilkwHxYzSRVYLPX3skjEPPg2ZK05+8DZNBgiXfW4JK+SuDUBqGrFPAoykZt/WZtFRYufESDLxS
RmqCCvI5lHwV/bY9Ul3AZzQ/MFd1qMupXmrlkkXbo3k8np6u9SJCK+MM1k7uNke18y0mGO9sBJ1O
wDg6FLezpovu8Huh1H8V7Wd2IyICjNMC9UUg5UzdIcjAnoLOc9isYbkyaLLaRsQBvQu2WCgC1oSr
42Faz426w5SI4XQb2U9sp1QhA5G6ZnK8NlbsRBNulK+PHyq6HJlvqkXay6Id5hgGQLbXiCv0Yt0N
WsR5uCnI/xIpw4F+mqeO8TQnreAl+JYNkser67V2b/OUybVUmjPMa0RQuk8IhV/C85rqlMjoMb0E
0c3fOI3XSco+Luv7CXono+6AEOaORtNtmHV8qOljk200k0dn/ZFo6GbiTfKRJV6QX8gJqa63kC0A
20U6KnVyb+mcC802FITbkALnzCfDX5g/CQ0bNPmwhtciNVOkRItvui8GOIyBqlr1+TRHfL00u0v4
4XQn0/sh4lQQNRuoFDQ7XK2V8RMY/OX91wHS3vXp++UDdodNQq8vGMl3uQQnrKiNPJhjmoq2a9hi
B2qmTC6zB8ynA3bG9IfB9Ceb4hflMIuQJaD+G4vTuoAeHUfSybKyc5YYwebCKasY04jk+6m9aKXt
5p3IdEii+bqmdLpMA15QwSCKHxjw+sMOEGOT9s4v+SQs8XyXu4eA6S6NXEQMtFzolkcHM0rGKeDj
Tffr6JtCvujRHDX/M9ibvseSuI5FDzvNQOQjAalfzhfRLjHIiWklYCHpVaiceQPCO5bSTFzg8NbJ
/KbzBv33FQNreM1IGLPgTe0lhRsQqM4qRWMVl4GUnN43x/8CyRmD8L7bzI0llk9sDOEjZXR4sdDa
RlrNjzT0ASOmXrdpGWJv62lPKcDei19F7B6sOdlKATpOKrmZNyi9Cfw6ZOUzhE1vGys9fWLpHIRc
wytiVzfBRzCgTRUd9Po8d1DTYTV4469nFPdvlOvyAL8skFqzKsNQWvGmQBEwNjazloGHEU9V6WRU
aW9/iASbO+KElDz37JhlsSPofdzhPkMVuAUW5sYYLCmrDLaB1padEl8S4ht8m+YPjXq8piVYPlsC
Qt3NOX1Cxmk9RORXrbtrgF/YFpqmgdP8GDMgGlc/n/Fgk5AdT1mV4A6yMCnt24+A5L/eIZ1/cN7E
IydlU66/o6n5o7g/T2niwqLgMijZi+xYqu1JvjoPVg29O1tV9vzMKgwMCxcQLXHjU7lkh6YvZGt1
+nh+fE7SOA6q3Nu7dLZUhxB82jYdpq1bPoklbyKyCiT12mNA5wxbFjpjRzx10Zye5IWyYxOowjRf
CctGKtIKGg6uwsuR3hSI5IK4ooNZo/H+P8W+4GFAaHsFr0nIk0RXDGk4thkGoalOX649D/IzdZiX
zDencsBLG/WIwV8W7gczn/w5vSDb4/FBK+kmDbfAkPW+F7GPA7SZU3QeB5K+AaD7E6Wn6I7tyEVv
7qcwwj7PVdu+oEgOTCRRzaCouI9xZdlPuWqAPR7Q96eqYdyxIZtIQzctAQLio4KiTTEIXRvtUEmp
GKviwkEEPG9kG2IpaHf406eZHoPIjWxqz4NtAX/BsVNFtJCJk0sserIBg7+2WLRqZXPdBcmFzdVc
fqqHQ8cOj3QU4AtbsqLL664TqtEh+ij/CsnWRp+6DxKburf3Lf8PL53puJL671O4Tw3VUcll23Xe
mGc60ea6M7pRzHUHh0c1NTU3Iqbxecuclj0SIdMIrqOgOQnJdCwCFv5Vw1lMwaxfgxqDFoVEKbpK
pYf3R2bfmToyBElOot97ZytEz2XXauUr9DN8xScYfepfBN1WQaRZIvB7t76Q4aYySJVICOhrD4ta
I2vlADl9EhJrdeumy/0toI7yeOHk0u9YIBn+O3jCwyyhFRV13+t1E8FbGTn0xJxeTDY7F2FZjHsQ
KlcTqNQIOHzRB7eJpkfdIa54ZJjw3uQwWYgnpKLh4JYL6GtSV7hHTtdgn+ZEkfQyAYEH+5B5IDvO
rMzg2zJL0Zi+blxli8Vx8brO8S83iWaSBBirXaEFNHW31Q7i+Qq1nzzIh2HCahzA2e7qqFW7lwjD
IX9A2fneaSXrOk4WoKcW4saETxZYTBQJSIS6Kf+rBDleC72DCRle6e1tfuCJ2aiJHvrx8Xa2fBvj
LotyrcWWcJyLwmFLeyRbIL1tqr5WVBRmS9VQnDnrywOm8nIesh0bmqP9Zx1FE21xg7H1MIk4QlkY
mWKuDJbQz11QvV71BrCtqPAPkZ2/rTnyREIvUL/Pknd1r/n9zwIkfhGFSxTzi5f4r2UWX926R59v
+JnILKR+k54UcuuFw0FgKuLKUyXx8AJ2B612or0INrMdTveV2almwmOjpc4iIIpc8DyOseAsbSK2
OmAlCrqeMSHlbgcKSXKOkdIXhqeBcwiUvVnyo9T5S99iKurqNKaZxo0WkjkdHY+un7BUsuDT23cI
+QzofP5gwZY/rtWPzZaVDMcEPd7cf07aLXCY5xSgUJbVtHbr4y3Eiv8U3/D45reLnfll1nWPq8w2
mvq1PAH6F5oB1EtMYFkr0oOxKnDMc9IW4uCw7/0qDVB077vOppwEPxqOHcYeCK8Iac0dP11nnq33
1Ne9YIKbfy3jE74vaDzld1tgkDaY/QvdBSk+MbOc9NrQgVbWdl05FJCErcHo6jszzHCPLCtkS5ot
/HU8iyWDeCDZvFqZIPKjZUtbs9pHCPyMaYPF/xSom2GPy0nrhkOE1+zvYnEavWM4MqIJuoLo7iYQ
ErtKWhElManfm7PgapNPLVcCGaGn6LJ9RX6i+/UwyENefMXzqZK0w7LWm54gsBHrvjGKwzA+Lxj/
HRmMDNkX4z2CZ3zHJf5QOxF0qAxGNF/CCb3DHDhW1V2h0TauxUxEg2ots2IRwjN7E67GqNlIghoO
ZOyVf0QsAIfyga3mkSI4slpg60LcVEU12u2dtNKZqpC716obt37fYO/kd0gRO+O175+6VBx/pBCH
pRvtbD0qorpB0PT2PyelJWLNX/rHARZjYEiNRDUlCrrbM6gPU/5QZXDmqsPQz0aJlFMnr0XuhBTy
XZpQeC4zPM2QY6nV8F9mL0p1/aCIK+5YQT5xyH36tpHDiL6qxA5Stl7mLmENIeFcI0PjMGORjisP
3Z+vIlg4G3ityv+NjyPO2mGvLrlM3exjJRWh8OVfgf3yJDdWYzVcQJ8L9OvdgsVhvpE+7oICMMJi
HL0sM6RqoNCErV5G+kwBlvygLgh5j7wHbLbDsv4fQUO8dVxsUcpnQ5NEwFFUhlm811jwJ91iUZon
BQXkVVyE0/lMb86xVU1gb0C9QEb0so6/GpWmlSUoJM0lI5Oe9KvRxiAhpkT3Y6ZfM23vEDM5t3Ab
I0d/heHRQGlfVYhUUnZH2nCOiw+yqv5mX0oxi4lKG43/52WI/crEEGjCaPzPynUJS3NgSb8upQ/G
p81Dc03RWY/IbRhqBrzV7X9rMXrnbJqnuj+UF0Ja6DU1DaVfrefaw58IZhnyIjBJ7Nsqqx90TO1n
VC/dAviC3wvS6V/EzSC4CvEdo6dKDSB6ELYFHiMyh37+qC0/k+cAx4NihQv6EzCEhq3u8CrtLkRR
+UZ8LqNdjknvHrQj0OXP7/C7eiU7W+KlVh76CFmfjGAxVAUwY7sHxhtSKIxt3qq5F14Y8jJLl+qK
/M0Je353+t5WlIEsyYFkHYA2TUNdymXHDm4A9iTR3JD9CbwslxJB51NscCD6hA/+beady/I7ke6p
mGkSGBdJGUghQ4u5gWeO116qppdpiX1aFoSlFMKbCf64d2eyTmN4dCTZgcBZVTGfjg1O2Bq65eXY
jozFGY0UOz4Ed3KzdnjZLSVwVAEvnMU/1Fyggx2tpgG3LoT+31dIEmckEBc3e8HlC1TOK/DWzkX6
aDKPoKy2sPLxWygujqnSALQGhp3+K7qYzl/mBrwcPdMPCutiU7Xetsxwqfgs8FnF6TYP9R1gQMvE
aaKTkEmgY8jxG5Liy/qzouikAA82jquus3OXRqSnHTfQWUiq0vAecy17QTgiQbmj8b7NaPClM4QI
3Qtm6NI0EF/tIX946ti5PRezEc+Gbth06QTj8Lbx2xldZ046+MB3/m75bN3Y6/m5LBYWjxvLRKgB
fu+8T2pXqwxAu2UBFTM8Iw8CbFXtwz8BdDBj0qieBe1br1V+7vk4kXPWMa1zRPsBghFtyPJearC8
e8PhzAWmswVtykKCs5U8EGahH+P1eKqey2Hbad2cfG01WdwJYJ28MfXCeT61DDhVuyw3dZTojzQ8
eifkK7Vq8kSlujzauC8ZnN7o5NP6NdqDQQXYopBiVTwieVgk2FWBpHc8itVYhLeVZM9xumP1ikcR
fwwgdBOfVHgzK9f3aIUGG1P9TLhKJ0W7MPgw6aGqMC67R3If7FMQhFj5ekixSAsWyXIZ9S75XA+C
IgC4KHpd0VqanBNPF/r771kcMijzxDFKtTKXGD9c2cNDz+8KLfv5Yu5Fe7g+1yqYvVIa5qouwjtF
2DIFKYSOEdKudayV0tR3EUHka2DOz4TqBaaTW5OV9d5x9fTtxWWexbhaXBLA7vVfCFO81Nh9YggW
jslO/SsP/z4Z5CSrONOxyWTIw335jChgtYYH5LrRyIRh20GZSl1IdtSrsEnQw+AvtyxHN5Gm+H/L
2mxhE0ZGCt33HFwX1l/bVc3TgKlhFoPpv1fjWH5tFVHAu1UQzZRuYXYEJgQnlGCpzOgLOVT0E23n
gtnAS2tfzzL8uERT54pvlKkWg33aqH+FqO++efQVmErG0lad37ecywybDnxE7SCgSpE6x0Rmrgvv
/TNSeXMTwzuC00Y8hENp4mylzE3saXPi4YvQ/hvIsYbHWCwegB1p7CAA/kiRoINQ2QCKQavOmsG4
CHD381BKV7WStnbJvF8gXUHjA5/TU3HXiio2ImWby7gPTI36exfXb/WOnoKWDj3TjehLk8iS75ik
/WvE2Y1QUkFopajOWaFfRtq1Os9S7zVWR9g80oJtq0DMFBrbmcRDKGqCwGVcVyJvB2UrDUR9SLjV
jEZLluZVmnbRYIZaOCSa4X2i+uWAtSG4vwZ0GyLye7TghXpgqbC3tMIPmSfy4h9QdFaQRfRx+v66
CJJPsrEiIm0i8Kf6O5c0HSCnJjemd1UEB/TduxkRAnnafy5z8pDBnHwW4kpZiBQ11iKXo+mKmKbr
8Zlt1Z0Me+f3yvlUL4tccuHdeCKhdvncS8DVHBXNYf4QN7UTThnnfAqd3Z+Wu6Hxwo/4olghyfoR
s3myg3cVRW2grFJnneGJ7aoK0kGAJ15MUW4taQ5BtZqHjdpH+kxCQXxYNE8hhUpVp1S2sgKb/uSS
vBoAO+fj82yrHG9nu+te0flkl4sh/aY/dMpAznocm/QVcFVDVa1T6r/Lj9d7DBVdWc27lDYSMoI+
IFJeY+8X+Q9PlGliBGgjPbqgNroTdU9ThXgTlNWQHdFldKe0eVNugl7aYWWMh51ZNA2HMWeZkFee
mLWni+OhnHLcHbt7XWN4RA3rOy9/bVzMRJ45J3jDUU1RaPU/SgKYmY72ZZw6LWjAxWOZzprs0RVu
hlZqGPH8tIaoIVjfNTiMqmXj0Klg6+EkOjmo3+ypOt0Xwi+bnVpbKeTwz11kpjdFUXZTb6UGsMJu
OgAqI+0pRcq6LH7TquzmhIPjkyHtBkI8L4r1BtB/FvhHNBezvsjilIfQd99j4EmChEAki19oy5Gr
Y1sTghi4Tue6urg+EvYaJeDS5frxyZg36nWtZdogV0OT4+Ic7xhelklKvDM/k5PPl0456nlEaD+k
sItXrL5h/+lT6fz2/cKP41Ll/+0Qh/a6785gwq9LFWCmq2yebCdPugAwWtaCAbK77AOFkyletj/D
twxzEUE7bL/uEh/aVqm0AO/GFo7Vmcb3FN+v6JFSRbDjl2xmvhyBFw6bw145smYOMUYkg1f0OCGe
RS38pQRydCn2i3v8R7xpCZ7Qm08XSi0Tyhr8Mg62Lt0prKurcrRW1JKe77DUV4e1FNd18/BE81RD
OtpZhLOEPf5sew1HlYUyVwMenICT4yBJBKRJas5e6OwUZH/PkdWij5ZH3C3iguODtYyQ/4vr80qy
t/rK5ZR1MKfGBer7ibWeIYhjBSIqfDtc88H7wUUeG3FhMc/8R5vYYaxdvXV9o8lpgOUN9ebUHhrn
5RgckqMjPCOD8bP++4ts04938AUJIlI4XMv72UjCJsHTXY9vd+q3p48GJAzUbYm8reEn7sThp1zq
Sv8eA/AsNdVtwqxZX/pn0l3FsqL5NcoLPdKgZp0LSsUZ2YpJZPnhAVYbw1lmwe3bcOTrphSoCkbs
k6uA9HGL6If3+G1KGndeBkj/bfOM5qFv92SQIAWg6TUrIQgt96PfZ6h213Mufd1P76bnDVRBEmhd
LzK+ImmwjnQYg9xSsqqJq+H6peZghxo93dqVTobShbIoUHGqlbIqIewMfD2sAiR20zpPsAhHc+lC
ZPzE8ZJUzHcpV8xuBbA8J1M4AP+G4Jz3Ru8nO7Wqs+7T8TXdSIA7YjlFHiCTmAASqnNjvFwURq9O
wkvQCcSr/FG82mbCak4M2KEiFPHMbQzzNnXyfx1xt8y7wnsBhVk0D6apZPovC7DY4on4gFJxspEC
+XRuAu5DYu6i8qr7dnIM2UOOstA2TSGD2+RMv6PJy2StDVO1JytQpJiZ6ldqmfixhgZc0N3y0dwE
YPXmHdoX+tYtW7M6TRi81WP+2XOkMj3H6JZ1h+Q46+ek9Bn7HJh+lPx62Qy67Fl7oSiDZmrbvmAl
2IMEJSwPus4t3CTU1RbiZ5mZ7v+riBrWI851VIkQ0wg+oc+c9tx2kYEF5YcIGcit5iUOIkZbtbLR
YN44JDKFPKpsDYWq2ZqWWoEiD3/Lii4b6F6+UCYntsOaQz3rZhobZUkWLuOpn33PXzknRlA7PCbU
Eypcc9CPN41P4xEqEmtdEQRxSbOlJpK3i08vx5tOQ3aRUCd2LEad6oLeZqXYsk813nmDqevbNkrO
eR5zFdXdSN6iN/mtndj9ysTLm6IfVcuDP8nmubGKVZ80xDGQNRM6+Bib3wZUIDOWEL+c8Diwudbi
DUuPpeI0a0pHkQm2AswVWWc0k7BWwy2dv5K6LFC4vVE9gydlM30y/HuooaHgz/4yx3BZzGuKXOZf
ovTzhzBQCMhn8Lj2HmMLqp985RYqPC+/OvhT8oUzSlkJEgYPdWE6R65/gxofuNSLv+6UAT/sIyHo
fAUMNkS7LGevmb8y91pZq6aEvpEXmFIAu5ZK8sQ+6TWiIS7OSVO0qQCphRYAUKRQOYSU6rlKPDfk
I/x8uh9ryd9fPDrZTAIPmfBkIRT0rZbJqSlOF7yqqecPHqHIuETuByYKxG4/kSUIuOny49AcnkTt
ya7sgXn4xXX8reS/X9mY8dHPez5pHE1lE/IYDQKR/fDWETQFuIILlmFv6vnDBYXg0yoZSlY9zrBJ
1UGutRhJ3ua6V3nwTcCY6CNZ9fzAtjIZKQK5KwLFjNNVv3Tb4m8hjbxPDG8OT4Yf17uNXwzpcgz7
/m+qNyrJcn6CAW58MXaIrEvIzN7YuVYqLKkkaoZGSuXX+MNA4PyzYkqc1ShdtOsBorKKqBtOEO+E
dHXeq878vB5SPpu+E/kqR3UOwFCtnCd/deBSF60s8MQl4UsqI7vI7Mpf8URuE191Zuaiwbge9e6+
+P7bOinIlfYBitDF7nkHSTSOXbVN67DJAGFLvzP+SyA8aO7k9Ov3LqoEbmcOiBu7vVfErq5A7IoW
Zk3dVIgZZs5X2eWGZABsze+Jvp7Mfo+6whhLmKBNTD5td0rt9YJ3uBSXJZNZNUPcfOf7IsDpLP98
13UuPVIKF1VNjawonVjqhu+doPb5UqWIgNQBXuAX3CweuqwzfQEiGyUy3p4luwOtIkTe73e2a4Di
HT6Yq2+iJiKHF/f5Xy3Jq+jmqODjbPk6uol+OxWMPqzBSZROSwUcCFu9yx6Im+zWOE67fSyoaeJR
AAc4wnm6HY2c2TyCAdXLl4+42b4FfNf3qu7EPRBvUc6aYacBPf4pv4zVSptVZRvV0dgbEaM7sgII
mpa+nmFgaWhsBTazP5L3IdJ7Nvqow4YGFyXB6yLHgnmRrXmStKoh419frj36Iqlx+oNT0zHe5TCs
sLMKgI+sOTAfChY/lsWjZYd7UYOBgyMMJBbSOyVnBrOJA8881jW7AtCr1To6zP60KZH9rBitmb7N
aXh0BsDgnpehchn+nzmqHpIGk7QwR93dbjA6AQ4CYNfZiQpqjLHrdq7HTYKyCcScvTVpaqOKJaUS
ZKoInjIuVwTEVFTHIN2jSlzEXu5gMX1fp89IhLPoIEHiaDBgFUesuNrsoxPUig1+E6bZp5wn+yE8
yL6DH/t6SB+OUCXaep7MkwRygmguO+9CSBv1s+4882CVBu6PGBN59a4Mfz71RA6DABZLJvzuwn4a
uSdIGybUcecAiWuAp8e645P9lh4L65LYBFvurw0T5u1Polj6rL4JtFLVjWcpq7wMaPBmHJirsET1
IPEljasQBbpdesa5uOU0HKYWMHH7+UdiSIr9oVYa/2st/NVgHJ3+GhBEFxzBqOs4W1EOzzMxNYaq
dwD5rq8cbQlv7J5xm1CqqnZh6pMdztSifTbESnC6TsStiXrNl4C3kruBP5spkcsQg6vedAXuGfkx
K7GHbeKb5n1iwJknBnjwc7/jsYgqSbtc/3DmHueUH0sAQHjMhEPlzDS+OfGakRR+UqhKdYIOHyXb
FZFbaB9okCdxVXnXCG0QWrAQMbYR6IY5hrjK4g5pBifVB1R9UTN0Vt75GSJHcK8zIQfrdg+OkvWg
aBjMs0c0aMVFrG01LFFAqHUl7qeNTLYjqpvMHNeAStBtmy8IyJSzgPkW46VAsijVuign40cO7Vr0
nuGWofu9PX1nYCZz5bUG9vWDsblxJeIirTrwkKzMU3jmcgORBpGtdC15H8dzXKZ+kURtxE5tngpG
c2bEfV/YLA5t2xQ1PcSOx8b+fUK3i/xpTan0I41k9wv/eY7lAcQ4Df2sn5myPRnTLQgyKmhYKmhb
APRRkIr2z5n0Xp+UXdr1yOPqKYY1NgE48f2XhXYzgAWbXuHk0toQMUt8nNX7yZNDU5MbiOsjTCbe
RvRVASqieSQv6/fpkqkUlo/Nf6Yo76BzAZ5p65PcUiojmT8njcq9tTRa1UQYnLpPOITFzsJpxaRe
0iZa1GAaAPjSl1Ap17pk2LTqSFMYpwG7Ws9voHxHvmRu4u8IyqS2c8St3PVBuSalgnZYpB0upo2N
958oHpX4frbOcr0SLdkpSS+Ob2TbIi5HLTiN6rxHftUZ7m1NP5tNxpzM3OXlz7u3ol8WSvoDrToP
iKwp36+mwDhfgdW1be/QRgc0aWHwL24N3OEAXrJqw6fo+i4Dvlo5dDL/k9emNoR4cwYmJ5hKPnfE
+WPwOyfsszHPebs6LH97K4f+kezJQHrApxN2761ue4KCxk8NIYX20ezxDyW7F1mhuO+R5C9WbK7j
t5J5iXhSzm6E1TN9DC1+u75df5xTY/3g7u9XeEmjlGcAmGdKbBBHJ7PZsfd0CemdhREq/uQuvK96
BRUNhie5PfBV56FovFPn+PjEjsurujJElhm8hCx/QZxqJtkbmEMF7NulQ68rNexZHAqMifFWVYT8
Z+HIpsW0FAfG6C3Zlx+hl6HoHECCpO+qEd1zphkv4VfDrOgt99aiiu/DErq1nwWMMdCMHt1lB/Sk
y69S3eBhXemcI031laHOEFt8cHu0QJuU3dc6oAR+lEjdILYDOIgrbVxtst9C6hAI3dYFqlu2N2yC
MNunRYCzaZaos6LTlzwmKgl1Y+P7+YwucweFjmYIoUp1PjhFVHe0xKL947txw2P1yRrrMiLjN3Sk
3RE4mckr8zDHQQ+YNATiur7+YAcxXv5YkGRfidAvsK+ZuPub08A7KNOhylnIAwDnenWkoOx/rQJ1
AN2pPtzTAgLqKYuNtcIgq41KCuJwGFx8Y6BuX56QZ2BQpAybHkNX02k97phIFrs+11E3oL3ExJpc
4E65wgmV4sOL0JLudN17hXjW9L3T7Rk3hw9zBNkZrNrSiirg6PyLPMFkqrjAQRS1nr4Wb4mr75sf
MjbGRnyMk9khmbJmkoakg4PUkb73gUPjVpnbBd68fUtbR/H+AcT4y0j2QRDWmJMZND1jgPWrk0dR
wgYwTbYohGwSYgrkNg9sUBMeWxvSgicbaxHarHZGn3bHk//WT9AFDN4yLrZZIEIffZiN4oqzvUM8
6JziVfc2Vqa/75I7Jyx9+e0ydRV/PdVNdAJZtENezbg+m5SECSiymMw6PUz/lH3S2zH9FnUk44Yu
RsEMxqfQMyFKB4MTcwcx359mtOFDW7oBMtFTYMUOlrZafl8MZYiQD9msNI8onQePWpvygPwgGdA3
vXrwdbvA76DIERVsv5JXxIfJ9Rizxff7YhhktAJu1pT4f/ZrggHQqrby7rrjXk2HxMTEhNQqVIsj
6Z0napUKiJ16AowQkkipxVXZSO8YT8mlIUs0pIyNHV05tKrbmB3WSZf/NX+DmVJQRIQyUkMuCMez
tKoKmlEveJ1Yi27GZvRnZuPyPdo3NrCabeI5d3AhnPFzpRzLRQwOCmniw7MBDF2bX/wUHsGbFf+f
2xbFdpYpwXyhPENEyQ7oYbAik7KcQvnSAyKvDQ1wzMF3L62N75QnMXfMmwExksbq9oK+Hnr0P1wt
WUif/pmtwj4b+89i+Etw7QX38QNiiMmL8FC4VfSNcajdEgeG9wGhSrh4egSbM7BzhUjKRy3HGCY4
4kgj4Ms0r2qFbVZUiVvPQxYaXm3TCsq8LkXtBulVPvHdOTugn33pcVehw3wRU7Xf3Jza4AG77u7f
J+W8zyjUWBHyIDP7tAAIfOnLfOTmPN9A9UORi+nxyVz0IsmzMcsYFL40Wow96gMK/FfmIZOHxznd
s6Y2cHzWa+HZj6Oh1h0YvrJ2JgdRqNvc/ntTjqZ1oMkePABklVI5Dxl+eadvhhyP8fd37KZN7xy/
TzU/fg2sT74i/5pBwFZpALM4aV3krn0a0MWfE7q6SwjHFDGdTeZN9GynW+OtR/AG4X/byLly1sxA
TKv0gK1E4GxOuQuNEQgIiOlBT1xbMT7zle+swYjuk0E/8s3na+MkWx9o8+jDGFha3rkFVZSkX/te
QNyUZugpu/G0IL03l9IUrbCHEy6pUgOoxQZkoLDMAyL6vzzXgy4HFVm4waGE3MFXHaadmaBW5Dwi
HOa8Nz+F6B7+fB44hM6rpnLGa355uv70W8zzJMPlkhXElek9rHtTgnIow3AUkqJXsMlx/ubJDgAu
riF5qHDHowtO1wZgp2C32l8ILo4IZ18qgvBe+aVhOOd/ar5x+fUMkx3EaCznItWkeJ36Dm+npzzu
IN7NGx7Dow0+jEWOaMUcmjhFFhhQyQySxys6WO5hmrOEDAcF3LXB0DNSZfAPfAFDMCWLshQ6Ksdx
VMNFCC2KcAG5RStoWJEREPuWPxhpO3WrsZ9Ur9WujrjAs8+AbdiV+adkoneyxxVIfoxKkqc8NC8+
CKJljuPXCY6iKsUAUitquxj0sKYNOdm3ZVjP8f4cBCnJkGOFqB4WaxcF20kY948BtWo6X7p4qwol
SMQbwBxN7BYGzShBqTvLxYkolhk13Iam+WZGIYaq5tMPjaAxqlk8KvK2+yzg1gknnBRZrGg9smMQ
4PjZq4gT4gNoCph9+DdtFP10KnlUcCK+zMJDr34FdCMH569FErM/cd2/eH4o3sc3DI5u3U+FfZlX
Ew5AiokJzVDtinxDigDZsMne1P4lfm+NXNe4nI3ijCqVIy5PIEtPi7zhTA6mzU++yhMh3WpWFEsa
80U3+uI7A+WLe75pv73j+UZgIX0YFobjF6y6HMSR9aT+GaAXbm52g6S0jLA46ccxFuvWa/MoEsg4
H9m/J5FOtbQTvtwnaOr753bXn/afdMHCKnkwaCdrr6NI9rFwGWph6ZwxHuGj0BmjV7p/vjwfEYhw
rR1ngz5teAloM7fV6yz3WLkSu2McuVXA3xYP1JmNAQGvGpv7qx16uk+2pS6vvHzX2CFrA2YFmQyL
MBNB4TgX/pDLTk55eQIyqVWPH0dwwweGDLqX9Y4aM9+UYhaihw2REd7AI7srlg/9So36S3Lfg7eG
pR+wiHKHkI6adfQJV1ebtTWnECaOEBss33wMChssi4KUDKGwcaJUAUd/qtgf5vpLEfIBKN0TS+vN
6OJ0nKTmg5sd+AzyXNeToz3ansQd/JAT5Ouk9sl+g5GfC/pcZF9ZF2L5p9MhAz1+VNnUKdF7hKX2
IDvk8h/tZdxEcAOB9D+cCAwZBwtS4HCo5R25faFBHLgdmFt+tGPueX3Gg6P6e/aiT9VGlCyiPXxz
o5FfikGyGvx769+dkZa6rzpMGxyjbfP200NzuTuOZVI8bMrxWNJOi/D2PQBKIm4PTdG8tVhaEgn5
mE/W4HbuBk1APy+vS4ER37cKv+5lEKBLZHCLNjZVQWU1QOc4n5SeIX3pizmHUMPJtnpL8GSr6gTA
UVW05oA/7b+QoX0pauDFBIRhPivq/m3jmp7Z5ldCg1PCBBGsnLr0W5fWmpJd3oKYX4CBxcuyzlU/
J84q7HfXH5HKNbzdSmXJivT2XtIEFv/OPGl1vd87W8nDc2Mg2RKVcEfqqbeHUvEK/gHe4PViNIe7
UaZnw8UJs1ang+U3G+Zj7MW/AD2UTk0J04rx2jKRRyXfN3MzJG71pv8/cNocEel4R0O7zbFHHvsC
iN7UmTDcXmBD06r2EiVVHWBX0nZJywIYV3HnFCLv6IJXi0XxEAnzXcvQfTl77cRnlHj0wL9G+fXA
ibkMo8thz4S4GeBo/8d/gu9gLcJ9n6FoglwsaWyU1nQpdKFaa0O36jHqq1K0DAS7uJKXBl7URfIp
wMG7bpAryqxDgcEI4mthwSzkv+sjuEPvTUP67y8gQUGYYnaj82c6pet9ZYvS3z435iWphY8Rgtlo
ggFz1PO66byo3Z6WDenAVE6pZRQ6WSGsYmoT30KmYvTsIWc5iM/FOofpuefSxNbPaEtXQIzhbu8v
iln04fRpxlJp9LhTbnQGCfytlWcGaieu9RkcXVO53LQo+gDoTPuodWp4WKGYYoOwkcSu+RXp3GqZ
W/FsJG++6DFQAQDZurF0HaFn1psWF4F9uZ2W/Me2P/ZqjfCJWSF01xeFu4j551xUoaq/PGgKec2U
W/o+eEfC5n4pp+RoUpcxTCqZBcezYIAHBPkmy+la9VAplaW1GrXSC86/3Wqm5d6EccTq51n3Auh3
rruwvV1Bh/e3xK1tCun3neLbWlE1qkBMYvunDvgrhdd1j06T09+vHQdyIFsf/ziFVP2imk8n7Odb
iWwzkDOT1zsDXt1WEJ/d4V7CKFsyfSmATjLAW1bWD79+GaRNle30xJuwOT4tydYpnPEVVyrDtBrp
FrfVyOAn53bgq8xHxMV8nwwrNjoP1vwnwVKQw/QypqVEg8QmW72aCJBxUqzoSlaDIz8GmOWb2djk
RR2uzg1iDzmKnqrEbkpeTmFussx+q6leR6phR5nDnbHecYO42q2FWHWYe2VxuQabJlKapNlXgBF0
Pz0qj2Ae00FZXQnJAYM8MU9YkA7cq8yag+w9aLAzWR68Ukd0KkN6NbuDrLdNxOl3sJ3xzyGj1yie
sgDU95A75RIvH7NO6rBX0kK6sq/n8paGWWkNmhL1d4PjT875eqsHB1sU6modZskjkH1OQ+vUov6M
J2sf4Wh70mHMJK3ofENUQm3Vfg4iEU/nhTlO2Y7cXmy63i3ZV3zYqgrSQzZHZmKGxyBKKu9Th/14
ZqUjmZt5L4Oa7D/1lxj7q28xSijDafOKUzQ4bepZtXiIponnthz2OjOL2pmiFN8Uj8IleBQHjwb2
wXe7OsNCQwOywEAlsuDTvVBgbvEYE9GQ/RXeA6eSl+zoeY9STjob/53t5VGbCekv8vZvqLhTmOj9
6Oi5You5f21d10mnAdXYkjM5njphZUAfme9aiov6t+tMUHI+gwoSV7fEJ2QrJNVXIb9iEmL+40dd
+t8m6w67bSlTyhnkYdSa04WKly2O4fCY1wLw40LpFRoFjBu97OszY2zgTyZjm9up5uXIii4aT1Fu
u+yPilZU/STMG19AIwwjF/XgnHqtwOOLLDn3HL/KkoAedyfTCzV3gd1LDF5jlmFaFr7zAlT0KGWM
inpCSMK6KLgikt9ZqHYQrZmOxEI41h/vosPa5LcHrfTe8Atw5CCXV4NGy/cNxGhyis1pcRxGF5sA
i3Va+iYorl5TAbq8odch6D7Tqr/8mGgv6qLqIEA9J5In6tS0oJgOzOIajDyEgY2DqKWEp4v4ATpE
GR/pAB4RJHIghs6ysOGaxbRGMxc9yYKuRIV8kNLkuOKVfT3wkGcFDbtL65bi4+0rZeGqA7IWtq9y
f0GAsrENYK76y5jg1oux+raF269v0/vIx8eUHjbttiS1jYiys4ig0ZkhJbasMLJX1cNyRpJVg8Iv
c9B39StAFsoI+F0cTCzghNgRRKxGMZ5c98qSPd1W0bjZwQhVKtyRYMYUzH4U3Hm41pQURXfse8zj
4VwnUh/LPIZ7DXwFEH54hB6enV1bph/S3dN5YLtlToWSGIAP6moGVmzIurlsN31FCcSqrIHaFmIx
fuhDRC2bvCnmtlvHOPBk7MGjcyLrCnELkgMDRQideT2dewe+puSnyakWsjafy0NbSp5tGpUUq8Tm
bxft1GqLIwCBF11S87W2Oc3NMR80bizp3NWM4+N926OP5YlMFrwyOnfm/jNtgOyZQ4C+MZV9pY08
mfzqHRvTVV8ysFp5N45G5b7DAqIJI9J9r7CtFwHvLW4Zp8lTosHSz81Lp6D4ve0JX5TGB0ki4iY0
5bULQf33TAFucLav6VzE5ZQRXw8ziqgZx48TbCYM+/WiUjIEF9AGqzWeyafPDz/qRjER9OcSgBJD
CfH8qLc6Zqmh6/g9b8cQSnro4/BajsVbBB4fTaIr3o/hw343YzdVz5hFNWWMFh5nQzkcmho45zPG
EavxMeGLLsTnaKumA+ccik5UMhAhpazxFl/OtqjBMJrZZWUTxNuPsB1mNoQCo9XHMJxQwBZCt35D
FZBUHbsy7WsCLnyfpzfIRyFTa/7LP4ABnLTpjbqyvj8NlkXnaLbB8AoRUcoYDjCI0mZlCz0X4dta
haq90Bx9nQMFsETKZtSck2lefJZz3JMT3SqIo6FxAQ2JhGpSkIKHkWM3H+WDjDbhXnr7c//d2UmR
hX1WGHs4kcHb7vSsnctGnxRnIroLVN9evZMyfh6ywrtAEots2mJLLyB2osjLue9DD7Omvi1JKqXo
l90DS1wEsEXmJzTbC+01TXUU6tRMsywxAdqfhUvaOW4oMh4YZ6b+vsXpLcPZ/O81QCusqYau7ICx
AUg7nl7SKJk3+qWePcc0kzXDX//DuNv1GApTZ7BDTxmw7Yp3ksVA5+HC/icpM6br8RX8jKRV7zlH
t8WSiela0fmka41I7UsQsmquymfXDAwIAduSK6twtlPGdlJDrmh+Jxytm+QAEmLj01okOpc+IRof
4KzkoEsk2wNYcCM8aztj5j+819YBuvHJaCwC1SbDQ+oCkEX/XgH9wNY32rS0GpzAQbZQ0APNagD9
fyfLNE/4Fuek1FYG6qr8gv2QAUBma2opAZwYaz/t5RF0aKsi8+wYHN701hMmgz7Q/H9ZlRAtGO0E
BKNbAPlPPR8UAUTfiYk9BDVsyWN9vibMHxbLtcc66+U8hmpzG0aGEVIrbXss058ltQkjdYV6DtyA
MOwn/wKOQ9jne4WBIKXJTDuCjh0G29X91m67cCD/TRIw9pC16PCDAm2wO5WLYC0eTfiLzldwVaOS
rAMxE/VlV3tduMRgO+B7+wEweUFVg6Lh3bPJFv33ZF1Kc1Z1etkdMStXwxVMjbYFD4Fn/6EOgrLc
9yKbenf2suL7sw/XUk1DJrCqEv55iyRXFBlkD1yC1Jvjg+h2qE/krZo7aJYWzB7JNt1pWX6vf8p2
AeBfMpBsKj9WoxPFRFXC+9oGr75eGaAsJwQYMwTGREfK800kqlkFn44PFCh+Avy7fVmaSoRt2Gm0
Wy3bsSvw0m7V0wjX9geTIs3yHaDKb94YjGfyLqw5aVRcPWuaVyXsk0fARX1wvkkTQOlKZtEunr1d
itoiSLOhpxvsK4IWJHaR57mWbs/ayOMCgxgy6JuJfnS3dRRjgoBKF6/a91vb0gdyeEEASxFgWpn4
ZR9gkkOYoCTDj7K+JLLT2Ql5qoAz4GUfivhWIXSdLwntLY2oRCjBg8yulCC9Kd3kg0X5xozYGPoi
WiOYomzQ7FPdIqiGSsQD4n/w571TnsXqF1BI5CjAFRkaSoprNVSYPJ4FiPLPMt/STLnYoAyX+wBr
PNt8R42IQQP7H8KxFT1BFif5Z4E/FjArd/rrW+XRa4IhYWHN9Y+FkAGolRSRvAI/5Lyl5Gcs2d7g
UZLv93MZ1IweUESrt5P/NY67XT0rRCH7wr7dEZjD6NhHUSCqnbIqAoJTWQCR5DFisyjxnc7QjM++
ZZDDDz9JXJPN77AhZtNMWvzDO3Z2GJhEDnyvC0RXxAr0dZEyQ/vrjZH+u3XUcG0LoVqbOpT6Kt4F
yuiZ0qlRmhXO9tCdN0uTQanXbxfNE4CLGUXWI1LLhwZMuHuqTvq4GGDM3hP+N5TOuaKIU5YoO/0V
HarNzHd/ShRKRhiuPn0eF8gKhbnDZxErN9ZIUercXnJ+xTZTjB4wagDdEOnRqjjLKNp7CxxpszSs
u26PSX9aPP/RgI3ADKWECOvPV7r9EK1oiYvxb+kOjizL2SZsPYSx1a+w3yAh06aryJmKo50BifWA
u+WYyTiISvkH5e4X7OCHhK3OVv/gsIdimPXBUVoKPD6LFaQn7RLiAmSl0Fyx8iA6gh//3VnXfLAi
vvsfKHELCy63oEmiMjQP8g2i0x1JGiKzAOpTfa/I1AaFGhF6DzP8viMGcQYnNL4VJgGRaMcSNxKA
msNGjDCuuGu8h4Z/UFJejKOcOgqU9+zMsV2aFMQMBWl4uvlqbzdiF8Ul0LpJQkbDhkjv23vF1CeA
+9R4Cf/F5hOq8owVcJxcJqYafsZ7RZhp+8MbPyAyTVkL+EVDXJ4N6buVe4pyP/VtrL3bRYeDt4HP
aGmef9gOrwZJB5aOB57rHca90PCHPop3zeVIkCuV5HFX3yDtbrRrRV8h5TcI2uJW0T/gh7IICNG2
xWSnCTXErZcX0vZl1/ErKl2DpV655Tt1CaxKlEPNGoAKwX3TyLlIVxcW0dtuNiTsBc1zUozN6YoD
P5IFazop1tNVf7zuLOfo6GlCG1wMzJZGj6tatcoJL2D3/8v6b3IdjH05Vl8R88TORTUzpdxtyHD+
gaZ3/+RZkX7yQN/lTFpO3pTVtgTlojvznmp7gwnLB7KDsv6qLUg3iAiXpFBVkL3Alrcvu3R7k6kb
uY6Xu+ZoS2gcoV3OQ8wIy4W9tb7A3Dn5woNkX6n8T1qI9Ry/hTNCJpsuSy8gfn/3H+/cDlaJKXmg
nt3kIyIsdXDBqGuKemOxu6h/aEgbsf+/PXcN5Z3XvrQiN+NIStaNGEpvvrOLqVSviUrhXoPQA5mw
0nQ1JHcQBmmmMNtSguvbyr+G0uuXNzpNGMZ94EXEhCh33GVggk6KO/aOsctAaI6MXqJ//iW0ExWf
8NLU2Cp+qClDxu45+wtH8QFKpI0X9EK+dxEHeizFpLJrzF354hjleS2jctJSJKm9GFUQ/rAivKse
TI1OLreK9GxZkY50vDPH2feW29XoIbNzvoH0UuBpWV7NAjCC/uS6aOstIyJWoG+7kCvwamW28KEw
OUT91itkw2D+2DwuJTbw2QBIYqwALJLeePH3XFFRtGa786TmJ6aJoJrr7IXtP4CMReDKqnR46+KM
buapYJBhj79xTK6Cy0xCkgAP2Ttr2pyb/LMH0YdlKAXC6e4liqusBpAG0CjQGw31IPIDO+mvqYwd
SjaeajGzm7FTDN7uNpE2fvg+2lAy85FBKgtIoP+KbZoFc7o9HjjPbBw4vG63GdHYssvaWJ22W1ry
t+NkwHhccPBdWpIBP/R6TrTrYD3KUPmrGw7nHyOQbl7HyfHwg7mtNnanDv7bwZ8hj0HEtfAtGMkg
BWt5CcJpqLRYK3eoZ6EFQx8dMgAq0qA8pooPp+dBBei1K1dKX+u+nRyiFghRuXAPFog4aP8E3dVd
H6a675atWMhAu9w9FM4QOUV+LSHibYggklmchZ4Zq244wW8DfFayP6+YCt3O96iZ55VL9358EpFe
Gbhaskn4ZFU3ZyD1oz5WyxQ6qfoc2eo4wlj3/gCM0hWc0HUOJRq4qrWSslxyHMFMj+6E989j4EKi
D3SI757DglZ4JgsMBhJdUAyJDv+Z2Q5vlD1PB/0i/gdOc4LiTG7/7fVITafxWtEGVYZNJPNxWois
CCvFciS9tAbIlcPOfkK0OydzLXqWwKaDoc35ZbhpYpEBpD55lZS/6MYxVUsn7xi0FsFJzmaavYhJ
sq/sXAzrAiMJAFMFEDch4cruWmxISIJzUZ+vdRFoVoopJJQ2o61L/gaCDa6ZjA0sAH9QmEdbynIB
h90+UxpJuXcPqCfOnMe7Lde9LphNqwgpVoQGotepPMOXR+sNI3RCTLNdJ17c2ErqgxinhoCqmint
kivyUjV0hBMiCYlXEvUTiZ1ziJCKga8u1XWEgqOtWbskvquzVO/llgC7+RpxGjx45EHPYFQvRT+c
1QKV4GIs9qDist5HLT6221j4h0+i/LHAxks8z/OVusV3mXN2YID/Ayt+/Bn3R7rdC4vHcEZcAZKj
ytD+7kfij6hkhHSl1rQV4jOhAgyennYGOeIlX4VB3f1U1uviYH3yjAXR0FVd/ZLjZCfBeg9+V/Xs
uOk214ldg3WpbWB/dqcBqBFWG4HNGwGMItXKR3KfkoM30o57DpA7iBbntN3mPG59pA1EdUIVXZGq
dLT7PLSY2tbqMnouPsKV26HQddzWbD3NQCbO+PbpKj6k08QHkx3s6zYARgrbNbZYnhMrGouLRhAQ
nCI7a8VrJdIwnO500WuqvZBTKWxzFquU+BtFe41Q6BCgr9i86ktfi90cdXxwQ0Ei2F4MPhJbPX1c
8qrJJab0cWcWjAq4KVAgJEmYwNwO379MDFRGBuXujuawv12bbeqCsOUOc87c3Jr2RBZ8pNUXfJ1t
wyT2b+nhgSiOZtN+/zSM+C/MUqGagba+ukzvDj5qYm83ceSdnOrI5jk8qwiRP2p1MYXMwVBuTvwz
J4Oazh6rwH9NyPertLJMQGIqqQEyf3juwRwe2Q1QtdCizMGYvjddq7ue05GyTVbZEKV/wv6PTtkX
Amap+dvqddfyXMqfMrQrmn0d0uaDnp6OR3hDrTq0LvvlJpcZblwzEN1ZLg3T8I9VYVKDxsR/HjZk
dZll1ZvtinqWL+Fv/7hNe/KG3N9RYAA4q/bi9PVwg2Umy/L6VCx2uKozcmSfdo7T3zMHcfv5j95Y
7dhgjBHlaK0e0sgXwbl1pQE0Z3cq11GIagAm87EkY5pC4z6qwE0/pitU3Fle/POevxjIG1aft8ud
wlTpKwc99+Rmt+chj9Z1bPxjrlii2Qits3C/94WNF6KzHLbSatvmh5oLmtrx6W84+nm4cHv8CKwV
bgeWPTRbWrAE65x60iTSeyR1F7E6xcWatWxbdOVXVoWbPiX6eju1WXx4Ih/ydlMEmwAKZiO1/vj6
nz2XhhrKH6xGuPRd+YdBK7utHVVL7+/OQxQr5hBoPrKpoo88HnjTsiSGp+dNyNtqeSjoJKJEaliZ
uxvlK/O54yLuWfIXtsAMisOk7BZWU2usxkQ8WrMSh6/V4FUeG51+B5bZNX5431CeDW9JhCyo7o8C
Og5xEg4SiLCdDU9+Ul8qq/ZDudOGxxXvoZK0/JHn9zryBnLQQ3N/FE1GYvX1IlyI6snNy1jY4/6B
3L2rqVldtuaXHV9dfQsskMqtlp4iCjbqqdlfeaUnKQn+2A5Ahj/sLbW/l72/r7EkEP8brYoE+ofk
2vSbmamLaumAmDB9zNc04XaF6TbjEPTtpWCaygOEzLSy6zow3POn/+htT0LflwhRGC2YSRqBeqpg
+R6G3HmSYWqlKU8smEpsvPcThv4DrKRa7H9i+BT1O3moT+FiVztptE5wdrrwlVjJgzXTk8CP+hMQ
Vesl/WL78dM5x1/WBHgbXD03wpEMwc9QamUc74zfrVZqAvrkeBxDqtj0sWnE1f9jvdeOhnREdI+U
Z1v7D8pvdIO3VaMMbfzeQuQgcAsM6Q/pHsjNsEexjwpje5jcu8VZ50Y8tCwUw8IpAeP7jzzhuSCE
SJygREtqVFPCpN4ucmKelgjeGfUeqVeW2glU+buCuvnzuh7rL5Zbu3s5uEcY+rVnyq25o78NyTuy
EqvaYq+Eu/CdF9hH86/t944xX7aRqZTtM6y5g/U9jX6FHdNIWE0b6OkMUbcBnKL+YnyoElkf/HMh
KZ0y7hSJ7Td21PEbFoV1dHR64wmKrQew5hYiGSTeAmFvFK9HqZhTJ/JWiwAS63cHCRgHmEzqOsIx
29s0+mpwZRZ6dvReNfzSzfV+r36mjLnpR+XNWzW9uEv7HbvVsOyJJu1zHr34nIKCQ4ikd5zb86iB
m0z/+qxUnc0xbRVgnt18KolyTupR5ft/J1gS+e5I4RXJxj0lqrk2z5ZQ3YSrVoq9/Fjz1Hnr3Mp7
GHX1xT1E1ZnEPMAH9a7Vs1cUBqp0N2muwAFTcZC9mSiN2MBEVqAvLlFoUyOToCNxVerJDl22fV1R
a4xKg/2yyuF2FNAvBGiBeWFlUTJtFgf4dRuSjpYdezvVFHbuPE9yFRk8125ypCWIcOZzqLHBjzmC
53SwpSnT2FJQnfvkHoeFp0UAKBG5pj45GJGp3aurgDQpFmhnkLQWHTvdE5Ltt9RBR16KbUP6GQ8p
aWqAWffPLFrOj7+HfMehtBuLaHgJU6RdDO+0G6rtSYbr/dOuak62ouIjy8eWqy+hw5mLN+Hj4fa9
9wVnpR5y7yYGPJJ0KdKzGvHMSD5h7z6ghA3BUKWfEESNmWkuPRdamKar1e8Ol5Ct6sg/7h/7LVvO
DkKsUTBQd/GUHvdyljTNUJoJcPSniu3fC5wZniW4YG+dWtNLDf/ijvPDqqGQViqvSTkN054xiNgP
gQBJgaZzYXftmqnEkuSwiB1VRb9ftQvWsnhUoTBco+XqqOvq6jCLTSZAQwPeo31HjtIsRqhFRFbg
oWo70hVZSS6DQasXY7FLV9daPd9sn0CLYLJO65Md38DLwDCsEAb7aFl+LjGU4QmsQ7poZEcfeiQe
y8YhkB3IBh5dS4DG3zCYWT8KxHVvIYMLHMEuyCP3o7HSvanWcun73bHxa6/v6nuGHulh78GFPB8E
aBb0R2ktqX6TF/6WmCmgeRs5lhxDWOE6gIlwR6PsxqGRmsyEPzJy9AgyQf/6nKG0Ym3ca0O+BZyp
Na3qhgluVA0LRmIo81Ja3oxRlBd8dhNgEkOQ+kMVTjnxl+XCCVGCDia9u94S4uDiDO9ybmf4C+W4
kkMnjPWVwOix18u+FJ1Xb6uaIxcLf8AQntIts0ofnSF+f8wFZ+dtdivOaq+LvOheBNNvXQ+l4gGy
ndVPZ6CVEsbVlpjg9l5SI7VBXXyAiNwU0dHIgLYY9G92PZ9lUffRaugGS8Zwb9ufs3rgDDUHxsL7
VsRXdUnWKuUlnwXVDSvUIFu8HjkNaMt602YL9bL1eGAj3qxd6P7z2teLKmokaB/LvtCS62W1CGaL
1+QsiJs85Prc3HNTZsQvVcGO7XmGIQjX1CAvp5kTGcIDBFRsQgEzrPmH0QmByzcT1HDNZD+ePKUi
ddhprQuf9XaSJdZaQVPfazqVgVAWeQ9COQOKDtcVByw6kRd6+inJS18m04QFbBqUeo2uRHqte188
bsJNp40oQdyN7WKgS4iQ3pn9guo31GFgMttRSfaQ6saHEc8lKwcg1rfetV8QFSwYS6NmcfdjcJFu
qjIwRuG6mXFZqdknzSHDj65/906x6kLT+58Rwam4TdPyrnTVwHSO7B3eWqFE7mT0Rvse0ddnL9Co
g/OJ8KdQ1lOMlVcIaa4OAoXZUNHIDKO2oHoy8JIy64ENbS6JUe58Zrb7F8BuPpoqZYUc3hVFuNB9
4WLU0L1kPJ0vH61kVa8Gwv2N3FO/KQ28CcWSTO3P0AYxJ1PnXrWI8DySukccHZAkTFxGGaROq/td
Vd/z2x4O0bQQ3ZN9dVsQ6lawl6mW9lRB5/SwV6fJy1NgpU5wrU1GYKcsG7FcS+V6vywVWlDmxfhp
B8goy0ZIsoGXvoaYR2VO4NgWQUri2x5FdGUfrtevN2J7VFpOlPsCzghGdYHQfAVCc8BdzNwSqya0
nKlGgvnk9E0LI2Giu81V63KRK2yTGdXze2/S9iBPCPNXiwYgc5OuBPdbdqO7eltxEisWtPeJpkt8
7On72N7vBDy8V3BRLt1H2cQwSzprOlF50wXWJB1ROPHVuQU19/8qdlDyBMjnN1EPocp03YcTgRTx
mVTCkDMxy2faAzVwrxXp0pdzc1R3ZgANd71aatEMqpIcgMzzdn4l+/eo1MFHJYCSHqAdwnRhW8Cj
cJk7UYVhGa1SVoWMuSNwQOLJV8EI4dEpFqHLhEGIXftd35hA3a7/QUrckBVCAerYAxhidkUYznUJ
VOd3mmTmk5XVZtiwwWxqDn/3Ge7FhHG4KpJh/rq1Y6GkbYuzh1KdI/3RgYUSAtlwp2UgxTwTswuq
rAYX4kUKoez4y+7VVFJnAjRrdfXaOzkuhsdZ8giInH6b7H4c4T16+uVgiXzq/C75nNnnY4G3HJA2
pu3rYkcxNhV02BoJrsFoXRnbjw6myFBy/8h2SrIbPZxspXN8KSpHsQEHD28obxB/Z8GXh6DIzjnn
8iJhGFAjObzP3DwshstM0HNY3gP4drUHrpqZLEfRIa72Oovo5LwYTGw/cYkxmQwd6+l+VKcVV9Dm
cwP3POU7ksZVJdInyfqGGDZiqEXCTcnG9eea/MzfIDc5lJDsN+aQ8czsNBnNi2f6ll5lRgZoiNOi
Gx1WFZ991ARVIjEwopCoECr7VCZcri1RsR7yGVkrmLYK5V38wRFwInxK2q7tqI2DyG9B1Ximnfv7
+jFRxgcqy/6evmouQq2bzvV8jkXHY0AWvgxEJoGAfdiP5Gds3CsOlNJz82Nh8t+E4Q42x8lyjD/p
zPKwS+r0GvFwaTpD2f/JqDDq9adm0paFD3pzgTQUvlJG4Ci6RrcrZjQH9ryXme9dERA/NEQS/nIE
ychxD6c9eGfWaPG2eMAAUhiHCjuAZY8aai1LLMAR4TRsa6RcQN2VIKB0B30Mk0QYZlXjbFuRNiHr
lhLXRR+7cj4+xRm8IE6O6/hbCy7HzOCBSED+9TlFgExV3hDoyXctcByNFW8OHEm48CYvqVBGOMGD
ncgcvEAZBEjCIoZeV+i8NuCH5froya1s/BnHVXhKfRMeSGjBzZmDgU8YAVU0fQZG3utup96BZpor
dc4HW+gXOTUrIbtU5qCW+mx5ZdVZi5NtuJalVbVkKhQo/X77hS7EUPnwfOaZnOz3COio3pBBcaYI
qZAHzRXQuZV2gB+LEiUgSczhBXa08a/LQxjbIU4I1LQ5AiwRkwVl34ojO88BZZiuwQSl2LC4Lj+O
5NqmojKLt5N7m4W8RbwHKFXli5x/ktD92SKY+dDA599pfM3BkoYmvEn0A5Q5iPyr+B/pKxW73I6r
sOLb3AADcdPYjDa0thBU2T8z0fW5BSaOnfkkqHzNaeSocQ7PuFbsmMiCoIsZ4ykRR2Lzm4xy9zr/
VaEpQqh754B4dLysRDMM9yO2E4mL2uAIdWX04MBZ7Ld5+UvF44PGYoBZHtv7XTpeM9FMWXfSD9aK
7cVwp0a06T5lRs0QxUbgTW3+yXE6KKOeM4m/h0sVFRTA2mrEBi0yxatB5w3hIwyNlOK8/YDwXLCE
OJpd56f1E/VjN0/UHedjSBW+uoig+ZWfNAevcVzr4kqrmUvZYCIG/Mt5QCLINoL6kOsKL9K4cfXU
DRVaNI3ar7J3CLd6QMf60XzGDkG4p3rZvgZXQS4VwuHlcJ/eaUiaxoBlASn14zbKPVv7h/SNdF2R
1/oz87sP5p0f/rRZeUCGn5ZWNNRkA6Vor9OrpqNKKUF1PxmCgZvtbV8qqTXXWFFhDzxsRGOePKs/
sRQY4T4kxdhIf9Nafwl6SAzbhMvR41ebhlt6jIriFpnweMx2fwX5IyJYg76vpptch2TjKPDXkhRc
6ZmkABJiTw3fB8/XZ3tUIF0NYSOuXqkXYHI/l3aSG5Bem4aFKSm8wvzaprTtLgSGIMGzmLUiSmD+
Pj/F2vxSUGyjSzEt0j9o0nvrTf4vfIqIlBmE6IrQ2WwIFV1/xwlYnuwzZvM5ImU1WJUb6WoNWuIt
02ozWkyMHaqB4ofapt8zbamN/4B7xQB/1pKDOJo0E5j6HosFl+DeKSqjDHADvTdfuRmIw8pxKIcf
wr7ZHvtlXhyESy0PUlrQ0FURHDZd9gxUsNOa8lgyVScwxONgINrUpZNoSU+scQsxdeY4ocpkYHmb
8afI2ltpUicBRNlmyvCOrmZRtuei8HeFwou4xhezGI26ZcH0+kcslS8ycWLQVklYCRyPDrFdlzYm
Vyw67X/9QrUVB6Srqgbre11xCMtlgfMi7aa6OZkQqe9mybt5VKlqhYSeY0LZ11/xDHUsnxesKusb
k691IN/lGL42+MgT5hPZVVG/AFCOOHMPuR7yPVTkyfd1nIF1oLG45pxbyXpHZlf0SJGTe+g/b4gV
OCNNjm2S2WO4+Oos0jcnWnZagyZxhZ1ERS2UHhCBigkGHGy5UaOtrI0bno4RE9fDH7KU1iH40QrG
gv1oKSBs+Uh2Tkbp/2KOwkTnRsFCgKBguRkvBxw9dM6mBtMmiQVxkM3C3sczhQJjNrXk974BmS2e
kabxOI5VkbX6MQGDjfx2jtN4olQBh1lGNEQEoBTkIEuszVMpF+5CNNvWZIJbhs0FmD0Rd5PL1Tz8
rPnzX4WGUOv/Hq9I2PlHPsTvYtxa+Jow0OSUgqp62FBBc3EmyqkoQcaSTQWYWIz+TDN+wQhVR3OE
Q3EgFp7M1yYVllPzMAtNbNMtJwNnnJ+/MhRHTmS6AFK9AhNpOCaMuPaANWQn97JRhQANJor4BxCL
uIHkWEnt1/A5o29Iw+IdJvV8KSha2OFF6SThA7WCi5f/OAMGf9pnWgu3QXaYiB9eu+M/ipgQjbrr
/aFN4Q4lUHNb4//HxuLCBpdyIJE8PfguX6H54wDXq4jbM/Un6A+f5JesotK2RoT8A8cXOxP148Ec
boFPArwufGp1HT63WizRZ1A7+BWCBjtLRVsSjyXynV8UmxTtAZQVRqd/BXU+ohDL/qhQujUTq/bD
jAR8BoOlP0794MSi32b4Ru1KSIWSan+SGIY4MuIOK7uM6W+gznY4Us8DuwnTvMKNWEnPxXPNbNPZ
TcUF+007YAi6Km4D8Tu18DAm0gkaXR7l2G2ZptdBD8GiYrweZxX4jEfzywUWpTdpdU+ymU8jsIIY
t7/COEBJZQU59R0tVDKJLAZXRlPy0wGMMeZRSf7vZEC+29+qtQyJr4WHBkr2dKJM5jZqPCEI77MH
OEAgMnTe6HC+WIKuOQ0OHJJo4hBzJNbu01upWSULRqu+DYN6SvHYDYl5VMX0DIJc1zhuXkU8Vnzj
ZOjLtOh0rHOQXMvdJGdvOMQ09TgZdJ7cb5prOzU3I8ttMBi/lzjV5NsSND/pBkZCX8IWDs0EJG2/
7Kkym8Ua3+9Q/Dz5aE8v9hY80QCsUtj4W0grb/HOprgxFT6eRnW8txpTfyV5cdKzREkXl1nfhMiK
YdhA/B0m4Z3ZWR9InVS1QcA/4EvAnet9Aw2+Lqv0bARmXiTkParDiy1Ca0GTaZJeRI1porp8Nf+k
SVCHC+nlqLJ/w2TyejYvHCUb7t0mdQ1cI8C7lQZnaY7UldEAdU2lIcDzLcE6N6sIxgFcIvpqXCCA
tA36eZTx0iGf+VEEkvbcL1QspIyk5Fif44ICE1AIdTsXVeD2Q653M9RRzXEmRzGvd9VxDfn4Iycx
mu01IokNzkGZtLOa/aqVc8H8fhj9ZA72XnAq44KcbNjCJ2V40pGVz+o1d++3sQIGcy14JHdyWmAC
ECnOKM8+hYSzM/p+B31IJ6P5hPxIdZrkoRDnTZWUJAqzBhOkgA9NWAqqV9PyFR6H8zD6GWf9UIV6
e2cljs6PjoUZS4e+iiq9EMIz58IcZTv0rtQXJqJtE9kOvcOHSU5W78UiSFLtPqhw/Z5Vqodt9rf2
r2SvOLWvodHN7JpwsXKYIL/Q7znRCHMsFLLQclnozbiEwbc+Er6zlyDzPC4OtmOQpMDaJlWVVFDi
PvFfqPOI7ZbLHxvqBAhhI9cStBV2j61C306Q0PCDKv2QrK7oqCvFzwBBUlWpCysjzPWThtVhREnN
yHcA5W8FdBhAa5aklDSkAKq4ETLWXlEA2Ef/d7xq0nY6cHuz/xK6jnzuJ0CcSQJsi/6JWwaIx4Jo
VHSQmwDjPhe0hxIU1CH+7kPlmOb/MyLcT1q2/PIj1PMbbCuuPJkIWk8qAfjJIsnDbKwL0UYvKGmj
c8Jtw9TbHUoZwJRAxrfulurbmCjiyAqai9b+iFaAmEVhUSjxmhWWHJnikjhFhW5Gzf8eRBHjYq84
FOyw5M7TBXDaRLV+E7sXXbTL4jn+xG+XiOThKGxkZT/qS3kAexxSfqZumlCoX9Pj538jYyGGmAyC
nRaVnwcPEyueJqWktrEdkMPAN3sYVNW3ro7scOI622bUlOr2Qq5n7Tpq66KqI38ESDtcKMqMVvfy
qgEr9763BL38BIkFmAcglSU4ViJzYSJxu/WC7S7mOFLquj74Pj6o4zrXKeLuYQMhEwIdKB75TWyu
cnfkYe4y4hdR7v2Erx34l6x6o/3yhIWj6tdOYSvsuzRb2Uwx0LqRqZzpy8cdut71Hf43Mkg8SWn2
lzDW7WtHV5rKE1nC+QTxRKgJTN9x81eqtJIvc58d5ZBT7ftgePJCq9W5wQIbjN0HLzYx6TYOkXs0
ImD/oi74O5BNJ9mDbYEOdQWL+sM0PdWpUsDKe9f5a/PBBSKbuArzc1NOoNYNaEy2tPo9fYNCjbv0
m1qsH5NvT8lLcaMJ1r3zxu9uS28aAXU/WUfWMPn1UgYv85TgQyUC6qdw8LmcTel5MSq2gEkmd65Y
LdR16vmIAJgi7v8o+t+f00XU2eyuRPpeOIjDT/iCd0uU2k4nJFuJ1ZM9sX6Bh+ShD5qbitYkCmTP
B6DQjKpeXR8zTJlaaVhBrvAAjBe3TlfMJKclW6Q396PcB4NtwDcoYao2HuIIjhHb/mvFt0FUtFRb
5Gsj3VaqGunzjlGG1JBPcVvI8BZa87VUwPAb8lKA5QUGN8fPT3Aw5DD3d95KCt8/3RWw1UaWvhEN
93qVLzWyJedyPLrlGs4/t5AaApvkTPZ2Zr71Gtj6C3X4XXAICXlpiGahR56sbwdZx2KRqI3g0ncs
U6ZnFf1yov3zPEe5BjSHUK9zOVylPick+WvOTAD2QpfBLZeEiWmrinqccHvid2pC5InuJMLSkvBJ
ey+yH624Gy3ErZ8tm91OyFFB3pxeQi3hllzLi1qaBElupJEYjSomS6F928O67by9I9Eo7280vXYc
6Do+tN/u/Q1TV5Wu6Cekyq/N6Vow0ej4JXbovH9+xc5m9pAGLDIsJMCe9c9bV02SOp6groS+815x
8I4Xq/Q6ssYS0Sy/LVY/4SzHurZSxuSSQtXYdNmkruESyhlyQyK5kuWWivQfBi9rWvOqX7gitP/w
hLBz2VPMViz3vS2BLO6eiFTuugHFXbYpwv7C6xC5C1J1lvEj0io++zUZPp9bo4tt77BvpY4gDnQM
CZxohLsBvdmn6DfX4Rh37uG+Zw2eKYQCftjFfShzAGhh+F6eYitu3GmrKeQe3JyEB61WmD9MeJbe
2P3ccgqDqqXWP9NbBlt2fLYK2cvQbehji7D7nGVcUoh9gWIMy0UAGKiKw0RnDcaboCctHEA/q4L4
NbUymHFj7Wvm2yhcq7vaJ/dSzfAcenuBgt5nbaqx2v1FreqCAUjIFstE3FRipavE6HE9Ggqa+JHd
R/Xq2jGhffcgVIAb0Cw82zRrDFd13kO4GEbYTqptdQmElJPm3q2egZLxpZ1e5PKIIrJ4sWttO9Ot
3dZec1kHuEzZ/DnIYY9RR1iZ3K4YZ8KVnXEV3+vMNWDTMQYTe/XLKjzw1zH9skEdFPmslvNazHtT
EazXL8AgohXn5vwrr7MHvuiNnALEeC0pqldBng98r4K/OzX+RcqML78BU1XhT3SeX5TjYU01u491
uONubIkA0X5RQ/wWaOZIoLKTsC5O/kW/UwEkYU+Oyjr740HuNlKpafO/maLICataFR3hlp67ilUv
oOBtYR1A8i2Fn3XY9+XNQJK2eU/apw72dZqUKTeguFT77VR0CGWXDxARzJrvUlIo4e4sX7unczl1
7iL7NIMYzdgF8/L76CPZJ8ENA02BRt0EpTvn4mLIxYGWi9v+/q+o9pBkpi805uKVXFwAw93gJ58G
4EeKk4aVHUtSmdLPvsA/Yy9kydQb6d1CySOo/uBwH90RH9FS8sRtvM5uanL9F9VXzu4f+9VRFvvC
qHl6NmYD3CoRRYDtWSAWI2nyZBJRCy1dQ1d0FtC3P5N9UxBPIYzXgYaP2hzmNNmZi6Kbc6lDhJ8D
uPzMsD48XuNsRR7EBcdE1akp74idq/1f63OMlyhxpXTlkF+1ULfTooQjn60vIx+ggspgTD1uPsBx
ggURls6dITT208SRuiENIBPSxfg1ri2X8lsZxwmGH7BWL+dZ5p0Yid5INKr7n1DHgnhfY6025mZV
oxA8GEOCWJXBJYpHrghzIWuhZcsrkugQR4QubW163wV5wUMS/uiUQioxWWiWZtDGx9BMKKbEoTP/
9MmC6JAM8cBo0ZzCsK6tM7im83J2/TcA43rWl2Riy0ccEKh/Y75NiL3SjbrRlEMOZqegES9JMI/W
FW1yDRllc+9gqIhcqTCPRC5/GKdJzkDyGAu7puo0JsXJKxz+faJd6amS0fFOrw1Ynd0ge9EbMxB0
ESzHCtdwqmMfH6alpGcf042hSEulTe5f9KHVq6PhJXuoTntEAmgy8w2EHTOFZWqZBKy2Pds9exZ/
7seUxKK97t0WCKK1ON3oNBg8wKm0CPdRVUYRkXueExupPJpcpijk2f1q8FHIh5YE7133eNkxS0W4
9CpAzhQMezLFdK8K/1OufTjfl9ei3J8EbAN0yddQDDH9D6AqbpISUUr5+MPj9YWpImfjh9p9BmOX
oKqIN26s7rF+opor4Uc8DrUeAMtdEfUScWaIOENRLvnWQKN2VpIEaMlIJFCeQ03kdMgXv/RMagbK
d9UCmrfb8+QFD6EhW70CQ+c1L8T1O405AFMuIG8Ep77COqrQ5uuuuOmZ6oHnZVLAh9ipvGZCQbXG
eB0lcrtmiXMm00QbGCLmuEFUHGB43YiuBm+GomUNkdF6HM/Iw6PQrBdmVhrLBaMvt5Yu9yTTt9Uh
fxTYqa54AXSGsZGs5FMMpolVvfqAe5155tbJS88d1QxcOo8vbqtjXpRBKVLweAukA9J+VSdxb8Xc
LPbL3rfNx086HebRUSshQHwqCD0kBH5T/uI+ra+tIFYJ29YlOTUIW6YAK5xADJ8/QiQt+OkoqmTx
xWxQ55zlYwUHiL123KMtT+IFDtlRd9IAxGyAYeWSGx+9qxyhn17eO1y+ZJpDzVcHbygtV/FerBq/
KY3+z55WhSTEmlptCEsmJZybDC8+ePZkaenH3HHGjuTLUxobdvzRoI9P+P9wq5hG/pCPHWF1Lzkg
7mxIKgbLGa9sNMkRou1VHaHaixLwO/9VBLSE3qiQlIGHMwCHcWjy6sm2wboo0TRl52v/de1NTYb1
jfj4385W1rkkVE2xBOkOahlQHFW5ZBWEAYEF+8+Aj7uRXz4eZzaWrKOtLZwkFbuMP1Ddt5iNeBpV
rBVEWlCl58fm8poAVtRzgOSr1hbhVipWzT9YFU8mdhWmmetVPsdMrNMg4LYKP9eFKHv0IcX6uhCq
YojABYtJSAiAfOXiLmuKgsE+XuryIm62vvxmxeQurKnF2j1EVGixIIfEXamkFbqitiTph5n9PzGH
Yih5T8ErBTc84Bm+qT3NxTvGQ+reIzMbnKvJvfLgsBX6CvEuLZc4tqJGLx91U7ZF8HhAIngunbsR
DZx7Nk83zlh2QE/8j+ah1A242RzXUebSr8LsqXA9eqaMVDBU0pDCksxVF8pjsW3zWE/UR/6R8kM5
V7qTaTCp3ey+TGXHq4ocOKI+hwvknYzvDDWE2Q6wQ5t2NAQK6tFif+RM5LILHu/JQf+4DvGofWE9
YRnXVZhyhk4UEvah9aQ8PpRcZKx9BGyC6xBDk65PjP6IchLWGLXB+NggjfYqclA+RwBG7mQKWHzY
VokE643ndNlsGDQVndIdfQ50IayPxdd3v5iFQok/r2l82x+/+JaE4YsM6Q28hwNscbKHQ9FTwFro
XMDz2M9jfPSe0+aUr1R3XdyXXDRNeU2pYu+7+y4RS4WKv62YDL1LXEW85Aaj4RnRFU1oUzebU7OM
0bTRxEldjzeNKh0R6iWO6yJm+YAUQyMxvhBSJP1Ndyu2Z7cF6FvQndq4Jg0fLGGOWTADwiWRlrhp
kPnr+dnuaRREI1yXLE78U+IbZE+C2dhoc+fsS2e8mUpaavycvGQbu5fN/d7JX5m9mQTKVKP+D0P7
gncZ1mEIJcyZ4uVg9Fao+pw6QTR+KFXipRf094c7R/JyRJi5hkm4owIzFcjgX6cjYQ5gnkw/hl/L
mBsaZAgkYh2PHmC0Aaig0/P+4NCzikcgAhy7bhpnh2lOJo7mPk0wHlLYqaNgMBxgZjuCcfBn2EQ8
fZVpAQbKmz1k0Xl1PvYI7DZMC+odj7N8WwgNgVeQ3+XQt/IMUzy0CI67wsgIvHnFzCUuFOXGYBTs
Qn78L+d6q+oBoFH5H3SA6xMw+gb503to9C32x1wvLCgyeAIVQJYg6vOZKGwguuvKueOsN6HsXyj0
EOW0E7hIHCPUpn6EhP5zRbexxw/Sl4/WDKxZXc2IMcFyhjdDMYi99q4G71MAKSwQzE8hKlP/LFZu
E7qm4v3VtfL4T3LOhBv2Cv26PnkTf8Qp7FlIBerp6lz2SkrVc1I5q92hl6iyPLIZHESr5yhumCXE
J6bvllTt4AlLteZqsysWvUUvF5aYHEDfraDVdYlR2wAEhgFsyRbFEfGmGQoW60DMT2OtyMNXg3Lq
bImdn4ghsR0RgOHPm86ByujJbxHGMYplPRS1eO9xiAV9F5J7HLIuymm1Ea+q8Bc2ZyRjFvOSPHuX
J8wI+Th3UAvVTS8zGagVyXzKMYBjopnBg1rQHVVcCFvZo3eE7jGkusI+DC5ztglqS5cN9Rpq0K7a
2Hz6UeApqaLPtud1zZUKVjeJXRkB/cZDrH0Rh7FNrfNAM2DFUbh2/E4fxiyl8Di8gb5dtplkl7QI
3UScNJ4VPjkWIgIDz94mKR2qPTTw7xs3dTf7H5kakZufi8rvVD3p55vTQ8Of2VTwDIlmF0o1Y0QV
LyDa3BEht5KShHOPl8sGZh6o/N94FTHrNbGUDbDcaZRpyGwmXU5hOp0rsN3q7TK73RngEdU1ljxt
Jr+Pj8sH9Aksc4gRJKDejs0FYTdGKXePWNVC9nhNp9EFes3aMgfP4Y/g7jxeJLCrjXbbYDPb/KES
n7iZtxjnMNMlgZc+Z4nrwLbl6RRY8Ym6LWKJ9ONCC9l6DKlHMO48sThrFLSje5fVGU6+P6CaKyZ1
1zQqIQtp5SyYEBVAUT6OlmlJbjYNNNIdLXBBt4uPi5QW0JeltjTYxV8iKiJjdDMGR2bAXH8I7Dx4
1CCmkz3ecmAKByXvXWubn5yKo/LHyVxacijKij+pASxKBCEDUQVfou4t1VvhKlrhS12U+vuyzv4t
w+AeEUsfsVygul6iMmQQ3oRz+/hX0mzVZRE9AQSYIjvBZ84UWj0VDU+pc9vEO+8scBpun0g6NLyg
ou+FyMZXL5mlvXByTodipW2R8cuUoCobxRJf2pLsSiWudErpX2CA3SOutmEqs2ClvfzP72UG1AXi
aRVGZfB8WnO9LGKw3KQZ6sac05jVD0Ysqevfrefvxt9k0owgnLcKVYoClPB/Ul6puMgjSmiL2GVi
wmBVthOALBnCfp8hZquYpi2YLpfI6mi+GFTOUmTvSbZ+AVnvcubrx2xVrFn7GT50EoMYsr6cmh9/
9jPEOCjmbRuZi9QtVc1k4I9n4BuMCPla+fx+y4WWvGD4aTcWTUJV2lbRUEQ4KJjMPgLX2KWfmqWO
Uet7NtmTCehDu3AU258JTIFYXhPFt1Farq10B/yjQKefAtJpDBQqwAIItESDsie7DSBr4mf6KoSN
xJiQjMA4Ubz0yQZzKw5rjLPW5lallJFutXeZ57KmrzUmWNNieYu7aRdDJ33frsOe8ko1ESkuYKNa
Vje8no0GFivc/JjnikYRt276oQNb0k7CpH3a2xojhRI0GHcMrNSfrnI8wZ89ahWwsppVNsZaui0q
Clyvpw4l4z+DQIU1Hcf10V1TodUp2Z7VUyuDzzAEFjNh6FzqJ751zX/svFg29NoDkPfO29mEtog8
o9BTL14Hsr8v6ofR18E3rBbiiR4xi3Us1QBZtfbYaDKkJM8S6Osxx5jxtVswAsiP3yZ0t8CnV41M
EOtdzQ4ALAN/3jFAeMV46VzSAt6tqVQ60eA+s7UNK5D0XHU9I/ZdvEq6rFF6m7L7c44/qMhrKi4p
Iw+LeWfUYUav4HagyIC3xmWfhxrDDQlDlK3RRkkggT7jE2DHJgWxhN+gly+sP7HKL2oGlvz651Ga
GbV10iihAwAtsPE2eD9p2biHiOvK2usUV9WfPFmwm7dxr4BXnxJ/LpuIx9Xc3wYVO7eIh0vMw8MF
pHFBgF4/VU9q1GpVOGT+aNwdXCxwvHL+Mnkd3+w15EFb4o/6gjoRaY/Y9yoD+DnsX0ZO9LrMkeRN
MAEGWDnHDvgiYk4NaBYQ1HkfGCVPiYxKtmHK/5DTkfO7L4osWJM6lXCKK1m6VAQxCn8Wfi1RY7K3
H/ZDkqk6f9W1bA5pvdTcMRS2iwdc/jF+nAn583h7NsdSwueWfy4X0kTfOrR6sr0ewsyJxJa/djOZ
vG05EkgG63fOdQhi4gbjhgJ89Z0276teKBhhXB43KypWYfm8jikjdo36YYhkaK4cEXhBnRGF4bov
qRrYmxw75R/oITt+LV2tiRJ3aO+7aDIdWtHtyZ2SYKXUBg3+0x6igtJNvx+hzAHBfynMXvd1BWZR
7NZMersyzcOnKr8A8WgA0exJ5uLO10fS5NgC87B1mPXKxUcF0QuHYQLZBmUXvgWebrqPvwVBG3cP
WAEv2rv7kdPBy7DXui41hspCXqWJAuyCySVj3XTBnOlXCuZg6H3gxJH4owJS0HfVVlsfNLSeKzI3
XSffJnrTk8MWc8a1nQdxDkaXsNGJ0wb1CtL+xNsPD4PxyCUelR+/vbn8E5hvWYvUFQyzuh6V+G9K
FzBkrDbu+bC7Cr1E6QrvKBx0rYbPB91x9wuZcmAbgpSB4+S1tqc0avs1yK6yGtFCrpIXCaM6fEDh
sPDnc9pJp4nvESU+4YzOtwRSgCUa0xSER2iw8gxv7+b1bhO3rOMOdmy+8ZzhecxbRDcOKWuJqSg/
OK0T62fsEpHnyL8Hw1Yic7+knL91UVffluODuSxMXyFhT9bxm4yRQ16amK+ss2DfNn2xk7A73TUG
jdGmlIA5LIWzmLOS/Jtx6l3PdZp9Y08oG/nwMw+GNd8MWHRkKYjEKbTudhbEc9X8/rbxswzufI8i
a5RE5lgQlTZveAWA/VFUg5giBFTguftf+kruSAaJnar+J1M7tRFy8Nhobnr/7RAeER3RS0J7OA5A
e8V2t/P6ioxQlbKvTYrAcb4OeNYzJSIZxBdAQ5ipJhogg9lRQYwvxilJvBZoE+hwU6uU6XPLZuxN
N75XT6MZ0ISjBY0bsQn1EvtUa3mNQz02aY4b3XdBb8H9tNeXriUpda4BGI1v9uB/Wm65FlP21VZi
5NQ+49OzmHNBSs5LTcD4473+kBarW5CShXDem557XVBtSRT8y3cethxL/rVhM8icezChEnAzBsmc
qkhx2NHETCpfk32xwbn4TERpImBU9cDspbtCLwHIBl5nW2/dHDZVzQ9DXAqA9AQ5cvW/KX7grTQS
EuFBPLWNnpz4GWAGoeAeDsvq7g2aAEwFRJiT5pjgQuHWW8f947Mi8kPqItJbX+r/osVmY2SCM2L6
SzERPCCxc7wSmm7O2+NNjgbXpnxY9AuwAWc3tSH8whU1DWwsL1cglOqjyOTaVqUMt49gBhbN+baw
pm4a3a0IsIoDg7yGeQGhPELfEORPKOHfMVSkX/shS5FwQk6v7RigGMxN56sscTko1o5d/NNcTdmD
wzZ/49TQWNCgKOasHrlnyrGIiHz3gkgx2nMzUbsadhn1eEjZWNNqRoJXC8GYwgaVIS09s4y7Vxzm
JiWFKOAqNM9co2dV49gxknCguuHdbVbelSvoYjpbC5fv5XJJ4v3Rmv6BgE0Ae2BHs0v37x36BXcM
WKT+NkL3+nJDq1YLXfid95UaKYYj+n32WKrKuEzEfEHRxo9/SM+iX6wwOKJrMYSPD0C8FC3WIWmu
2gPsKWecFpY+9AkOqghmtlYUtFSftaeT+WBOjCxDxXsg8IwYByRVSpnAMauCsQIyBmKX3eZGaLOy
V17RVZqge9V1aHK3WHSxeJgMwhYz1eoJST8EM6j46lGpGFxSPwzsbBoneqIiqZkBTAepd+/Kgh1e
4kbZ37qvmepdA3PoSWtX8vd6xG3hPd5ypXdg/93vTPEgZA+klVt/5coZfG0rz38I3a+GGmsbT2Bf
5b8bxBzVnq2Ys0mILSjka7ZrDGm/qrwZX/gHLdiDHprooKUDOLD1S6iep206yWiKStJT0s8KXm06
UZl7Bb+Tpg63gfbpf7rRjrNqXyqAEVYHs+518SrdXRH0K5oieW1CboIgtaU9tGelCfvM5xq3+M0L
b/eRpO58p+tX9HFVfLWanet9aId2OSIUQg2Y5RWhaP5lxLGHCSvqLEc1EpVkNLaz9iTnqA2lARgA
CL4G+1cnwywhCo60iqzyoti9/03mWqruJmnp6UG4ZCCyj5X4KSfIsJYoewEEHj2of8MX+y+cxWFQ
YfoGHbu/NZSXwgQAHSfxrGG7cIELxZb+2FsfbPhHFh3OiVbpWN78iqORioqZa2gCLOs+Xa4zBeyf
8I4N8ubaMl9nYRkoRpZ8eKSY94UZ83Taa5Zi60w4lO1J39+Kis2j/Dz98o1tmKODOei2mrVwl+h0
UWxl4PwFoMEZFXzDMfAOAWtzjVW7ApqY5u3roxtEA7i8YtaflKev6Q2CmR9UwdAjHWPaJr1KAVYC
3EYevZEvsvuosAnt/Ej7KtLD9XOjmHsiKWovoZj7ShQCMX9svp8co0OCFBqqa3fQ1RmzDwjjaxzY
e5W2I/2JNJ+LcCroApYhuwSErKJJIZwH/mgdXGYntv7dFQfM4D47FYrvJRFu+n5hq17WXQXT/5qx
v4jLb2OOEhOUhH1VoUKqUY0T2GJMQi5vG6fJ7oOwKvjnbNQLl/UbkUbxBTdVS9LekkSLRHRxkqm3
Zy6M58jyDrJdqmiwucYoXiRxt5HBgGCjARkHxlaY1QWKEUbye27FH9Tw96My4RDxF0lO08Kdsjrg
HZmNCoR1j4KljQ3HBkYlIUKvYl6Nn4VmccwtThNzJCQDhGy9MQGhdvWfKXSGcUC3QCHZEeKQR3hX
Qxp2avZNbnRxGrKOY/bZ4OXu9VaAWw4EYUkopyf7vxPzGzk1/e92TywGty0/VzPa4o2IwSaWBXJM
VdXqOqvQVjmacKsGZ4WbJ3mA2KBBhdXIo/WFCdaecGnlawP6CeV1vQLOA/JNjL8mQ7vI1mMOMI8m
EwE/1SddKmbV53OH4rGLgbosb9RfwbxDShSr7hRvE46kgJudHH/rz//V2wpSXu0x8/ZDhqbJeUuK
niZEfMjzPJpJ8OXjLH1NYkmfP8vk0wouJuE82EpouAzFOFmXyI+NyS/EpjMr5KWIiWzes/YAq/eR
+ssZZJER2LC9Na0/OL5S0hs1bWApx7vTlWw1Lx0harf+UeWuVNCGnwu6ZzO7hCijxKE/zMzOK40+
u4wcEkLmKn49E0gGLOSrIcF9bSWFK69JE5vI9SeCl9v3LVjvI2k56lN/DDr1TsDFWDaj7AwEHWp9
Raj4nrcNMuW9cDxpLE43lArgo2lDBSXsf6heDfGp4U2LHUq85quvP67OjLnx2TjhziCrI0c11Re3
MYlCukXVI5dU9MZNty22ZpH7r9IL4GG9w+qAOwJdAMY4s9Xj/6pJXg4UgK2zWk+CdrsbD00PqhzD
kjGTPfEHls8OIIPQrlaJd4Wpokz05yrG//OTda9Xe0TMSarclTg1VHV2VvKDZcAKvJem1Ka1B+5r
u4Mzhfdanmk+NEhgtriOitoeby2RGvcv5xbLF9XARlaMFmI+8GJs1Ck08DMBSqnQgHm9C0w5GXRZ
gDTPunPvLknHgFKvs/HjGJJsNEZ28niT9la5wfNsqCNwSHgrW45SAvGyu03noiqma6Xog2L5Jo8T
Gont2XHoVbu+wNNZ32BeRdFe/tFvFf9sbLwrS79PfAH094LEaJohWcALS1h8U3RMdKnQVqEfQ69u
RXtZOU7F46ri/fiBIvxyhQOMKmHc1ivOE5O6RpOUXFz8zh7g3dSrueun8VFOAXFnoseGVAe5PLvC
wnZrIjo/8l0hgZaZ/itNnLgeayj5oTBomZ3n5zd8dh9J/BE/zRoDHvgVn7kgUDpwicLfI6CMxWXh
BezHvhEm8d98aMMSLebaSvTe4V8JveNzP/FBeP/mmHBjCTjBZcPgdi6gcShPNYTWKReL7AmvtB5g
bOyONV4prf5PnhBLnLELG46nFEVMRXkAECrYDFe4RXNCYfIqfqOj+YRXZ9Vbbe62bsV2ZoVUwlQM
L15aO0/AublX1Kq2QFK9KuWrIyXwvzxTpeEtGMszhnlebjG3cj/nWOyFanIZUyeDijferjnh/k5m
DzJoiuGMwBrdulNP7MwCKlE73j6G1XJeATxtCHRd3mKl1sQNtsyASpv6iNCSkqLPW9b3BLE57e8V
y8LZ3QcCNLsfd9U6hVuLgA0EXva6A322iyRIHysM49pCR4vwkm6c+2VGETBbLL3J5ECcIb7cNjAc
vy6vVScaAgQZZ926LG3AmhQJTdLfGdua5gqMQ4A9XvUj+JgMY3Ol+ln+BgtKKYxrWur8H6m9/vfu
Djw1IxMKSqCzI0AlOjGMQ+fHeT4bH9wDKN69jePmIzO0cvv9L7T6P2Xwcxp6yQDXgaSlDZT7PqRo
rz5q/3dWtM7tV1RCO5AfEWf6U83XqATq4HqNjnqqRV2/qoLIkT6YR7goeNDd9blyrC8U6huMX4la
LnuDcSNd7E20sbDHOAa1B84nHw5oPBSkZKrgXCiEm+r4t32wdG35Kzx3RfjGF7gndDZmI9Dg5F8z
QSlSCf3NJx0kMTTbIu2KXNB02ry8WCAa2/dGkXhU1XpY4wFHEKPpC4tIiv77H6y1jMIJBnuOeiBG
f7PpTz+YO1SydE6TAM/vjytSo8b18QcNANZJn0NuFrjxnKOKqyog+2UjAvHd2Txmo9Ha3o6zwoTh
Z7CuQJycECLCm8snRNLEzGQWzasFrNZcGjTeKmkBc2Tnvbm8psgX6doyQQkkhdkreXLppa5V7Vkp
Igf4AShoOkAor5yVs51NJ8piDb22NWFP5KYNcDMJ/ptmz7ajaiCL6ZUmYTIhN8ImJFL6P4og9nlz
tcotciZHyfOBma4LJ79+jLxCv2dY5b/KdXQBmpp5zyJAg1PzNucHdWN2FpgPJJKJU3vCa6Fwr1h6
TRy8EtMZ/U2V4gtB6rF+XJy6UMNNU+1dafKFplgiGw2OhDkfKFErxd7xQX9GHgaJFUYB8MYoVC3v
NK8TetqlBYP/Odenxiv920/O2aTVDEX7FL3E5xm/vpp8dhg4Myw68kOUu46r0l4C3MH89toeHG5H
eZpfSeSerBfJMcAAbPnLjllJcJ7CEPnmsCgf78vu83rfnkaXH4RvafmtVCxNty8Fj9L85kAjkyyP
kAinCGcCpqN0d3gkQIYPuZH0D5VjtDG7QZRYHNcECWlRdrshYuR9co9Mt4S3Zn9mkDIm2nt8CnNI
mJsjT2L2lNfWZAA8hyKzF/4riWkGGTEP/jiuX23SVHjIVO0CIz4FF2NyUx5vgVucVOgvRhNVHpdR
icCzoMZ+7fe5OmjksPH6zr9kshE0mbKkXhWXR9Blk46EKUYt9o8hcBZ9yTRsrOrCiXA/HFiWsY1k
Fa5Rb8zk6TgFAMHsRaGNJjmlzNcuipbE1AuSGZmeIxmkFTw0+nYmggXKKuVCvYaA97YUfvAEOP2D
+p5cjMIcZBjr3M36O3pSQXKood2Cj8Es9XPgOKufSweYiwLFCO70wRzHY05t0txIEgQy3nozhbY8
k5ARwEcSunqDCJ3Lsgas6cdVidQ4tZiz4ZPXcTYMp5SB+j/cF6xSgQzQRh9U1DTConal/2xQBSo1
RnvUtnMWLzbMYAvputfGL58foMEbrbdOiXLcwcIB2ZE5vICw1c7aYzosgpD6T68J+0Q/yvUuXi/U
fLSkt8bH3c+7n1YD0iw1KG6L2VmHS2gZsvfbx5xLVxXI3kHvn1oZrxsvp4UXzGTDRDDhf/BtmFX0
rBPwrrhwxrlmrGg/z07XwTIVkhLaXmXZfrjJIpBR/hfHm77knkOisXg4xBbhI2J1Tg5oU00P4ubu
chCalnMRvqz0cs9LkE/oaqhpiuws5VORlRfmHSJhmtEZf1LcUPaokEL7hFjmCAIIT32Jfw70i6sX
PnlAJ8wrRFtbSPavrFeV88HfymtJB9RD9Hj61XAYj9mcQi0CPIkVud2huKt4yK2+AYpEPs9VUrMA
ky+AuVaidREx5BcsGCIshSGNB4uIedGiYjPm3gOVGIqk3Y10oNlAd4X2jtWkle8YNQG6Dsy1gQPE
dVgiaqIvd7wqoSRNsKhGo8QqF1vvB3tTWjWY/itndt+liZW3X3RkxLJrxa3CjTM6WZsN5AUXdDeD
IPajRxJpjAWGFSbMIUsIOH/jy7atDzxocLUxqEnyITJAalX5Z1JCzO0xMN/fR7g4fLV8dNGGRd4/
U19/I5iFkHNZnP+6gF31CTVBJP4kxvZ7MVmrA+ozAwWJf+DrUgnq7wPfIzDLIGXn7I1ctCUz3Y2Y
HgwjGSRjbaVkuVU8kvLv/6BYbfz31QGwACdltBcikoP+ora+1yi34BhUm3/Nn79zKDHQ6JfwWLQ9
OuoJ4yxBeNTTll7mYx84A0jP6FRPK+kY6KdqL885CrVHzVRUx9d/ymglqdQtGdiWR/iEIIgByUme
awGRlBwuYbYELqDPUMORCsDOnagx/KtSXzGD1Y+aJl2A0O27AYtCCoEg9TUtB9Nz8q4zgsg6QPyt
raV+6x57VaLK/+ur7FwdKquWfq5tTxoU1FFx2wROVwoGLZuWgobwPbIpnpVyuMIlec3a0L4jONau
ht4LQmZ2IgcFtE9OddhOTuIdtkqFJZcHPysDx7bX8jXZ/jpYP+lFG4jTn9rGTFGbDLCOBGJZ1xvA
TvVEbsctT8TXiuKZiXnH7Sh7b2Al61hL3+lKKwOD3hiNn+2yjhpDAwwM8RKpY22ewqHF7prdlnsL
XhIjQwXE1PooL6Ee6vG7xTGa0zfEMsjKDrNTtB/suZdT6PGwA5UVVQdq1HjgQbRUpio23KjPiVxF
WpHYr6W0p9AeXvcfco1U46AiG0JvqoCigTCX6TmjeiXeXSjNHvZDmmhKC/ZypxDsZ9ZPyR264jLA
OoF0Tx74o4y4JfHf6KnsflSo8CirgLrTVQ1PD2xMLdHANnwdJjewRoSkHw2yRUtUdpEi/KddlxEy
8luxha8DxvBzQu88x6nB4+NYKFx9pzGoXV+e9LatnOxTb6gRfuhZuUIiUTDhE6B5IF5lqPFA+I6s
L3TiDE1i1SA58O2sx2tdqj8zKkYC1LnTKLZ99t6MvzrG9eozn+qrckgbhBoi49e8/C0gq4jCHjkR
Jho0UmnG8/W8dCw7kCzcKb2g9viaJNBSsz9yLkNxegouXYI7uk9yrqlMirmvSFtZt2fMOuneLcIV
lrcPA52slcPjbIq1u1TIu2RdHbjuWuEFZi0Qx7kspBmJ7/2GMSjzhkDpDzcpnymvu0rbh85MEMKR
mYrVCyq1TYSdXTCTwHXIbBpEkRVv6ZmkB5iL1B6jqHVwHIW9mMYVbuFQBRJzWhEIHVXcB/I1PXM2
+brZlrp5nV8w3CBWvM1W2/65tQ6oNNWYuTO9xwMJrKxngWwO64Qe2sDXsFZ+nRqSa7a8PB/JTLwC
m69KczyeUYY99E1bn+5n7hNTdrbNKqpRFOcWQjENxSgGINirXV8CxBuQwJNrqaKUj9Lg+OPCf7Xo
4dx3a88X+TGBhYkd3mk54HULg5tqF3ys4ME8GE+Kq1FS43i24Hfg1SzgGBvPtxnjYo01mP7JlEfK
X1xUyCjYxuc9V4GP1FF/TfzWe2KjAOlT+jBi8oKJG4mxfV7bVya9ChoQWle806kyKJkImxR2U4tn
J/uOtC63UqixfJsN25ckf1Lmyx9de8WePisoPJ0NktG2bQzYUErVDe6HGAGa15aqOwBMEoB1Bh0C
joxo+im6QWKakeYe/x2IrzSaucolUanD2SYeEK/ktMfehhHWNoeVS1/5/0R98PL2uf/XnbmUKtpS
DUGd+xgTPxJEDcgSR+702tM5Yv3zo2x6dTQsMHe+PJ1elD9QqdF+BeJHRpgo9N01ScU1QyoGr+hc
0yaEm2LNGL+oNDKVRFoGIIHSwHbsxOWDE27Lj1TPSuOZZiWLKDS+APU07micaCkUYkJ0Ku3CFIRo
wxiKrBRiHzGMJC1dzGKCVHw8HD9snRi6rNp+maTO4ULYW1dJX3Z/U88rckIfgrxuO6WBPapqhQ68
FqLe9GSDt/XSQeAVlZXjJ0Sld0eilmATd382h+KsKreBWgnYWIO+oTqDtiXmFfVQ72ilA1CW+M+j
L/SW0c5A3TzO/oEDLK+n1zsuQ0RWwJvo06imsAXo4Nzyp7w2SFAEduEsCH24poaoFyUwDJFtjkaO
AMBSJc4iadip/LaxIv5JHUBfyKiJ4p7uwyRo+rLMpuTM81uKlsRoYDfLqZZrte5C/cFkfj+zSoiz
5oTPAQwafvZ6CoP99HNk++b2Ccm+wmsGoC4OHbYIUMG8cctW6RzoUaTNutwDGihNR8NNnfz2OLGY
UV95CSMhpvLfarGBJqDw4MLFtmVGFvUBYJr9CURlI17We3JaWypJr/krijZCwBBah+NhRjzIy+br
QaVCjiSNPMOhL06e9NjVC0KTRU/9CnSX7EXH+QLBwNtWaCeXm2I98pyA3i25gXrQcEpk3Lz/qkAA
cVUz7KOupXGSwKEW1DCQcDzmPk6HtLSVvwYT1wzsPev319UXGS29+3L+mLsKbaJw5FHRKSZToHHC
c6FOf8iyhILX7jX861tuP4c6d1Jvw2+aBj9wxRgocv2SUtzIpiLLoU9lDDY0hCU3/XRDHLpiHZZt
ZJT80+GBQznbVekflJirOQ7k3pBQ87AcUgz3uBXCw+QHkOybnUUm2FCHb+E83MA50uDrt4Y7Sgnm
DSEl84M1ZmJGicTDpAfbE1jjpo8mDVy7eoUIeW2xgx8Ua0x2y/2ifWTe9qZY5V4TG+0MJ0LC6mNC
ox2zDshtH4hbe20P8VJQSHTVp702wYwtzlQkJj/rtZ2ow50OO1cpG3R7VoHeq/dyMpstZHNBA2+F
nm/xIIB3Uyvl7Lc/KQrsgxrz50f7U6aP0DKdxAlz6VuG+R/280XKp+tHxkieArU5OldKjSuZq4d6
DQQ0JBzFBTldSg5Q1dQiRAnSY0950PfOZ70XC9GSqWy1Gwk1xH8gprk15X48qQ9FJb698huYp4E1
xna+9sttKhCHFCiIgxwalN4wPV0YdJ/LjpMF7hDukTL/EH0dXyNSECwTPk1ELrv4ediXKmwhll6p
7CvEoY0L+DIZEYpIvTfDFVTtTiznA1qO9UjKD72eTMJ6DvWI65I3oEYTydx5ExMHni41Tb9q1cU7
p3swfjvRqopsp/ibZhpP3ktUaiIUyyQQvUcQLvLEDVgKfECqnjFRpbS5DBvreICxsgnBWMlNRzLo
4Wcw5Ctw42Y7/So14TjgdSHsA9cn38zHs8MeBJjw5SO0oWgso5+2C4r+1VWi2M26j+1cz31Po6KN
JNZBpOuzW6QcDSh33O8dmE6vb+2PGgQJeN+ax0dGIVFj27JZ6KZO58Hx63Kkog+BZAgUqx3xsJXf
NY6vmGGE2nqZclVKu0ltd47+l1JNBH3XNiAmLH8RCQTo4VxUjA3lxDm5h32gDdvR4u+uZ/ArYQPw
y/pT1Dr0UKu3FXCapMmoXq9Jg5utpfnfQlHt+2aG13+BvmSKSNPptYXI45rnMiNS5cuDmmsa4zpM
Ua04OjM7vdujxN9lF2RnfjLw6mPwzH3hLlwlBjIYAUdOpW7kx08nABVPeyR4ZIOBQ8TOc4uKx+sr
NCNa8mYcqO9xysWZc4Qf2+ERuNF5pneQhs9DHKLGtkrV/4MuAGG8ulde1w5f1zFtWrOA0uCVIjo9
RAN1hILjtUhCvIhwtXBWhGCc8YnX6jpbDaVmzfcoYxKQC0z8TyWVJkslBMNo2F1BYAk8GR9tT1lY
baSJ4W6w8ei2caE1ug+BALWmxOdyWrFHIMa9X8PLF0HhgwGNKzyqGUgMZi1Wp7BFyqUyN+pRgmSi
y7wqTTLqNdR6rY5D+GpeGaFafU3wznew+/t/W9c+0hMLM0Z5//xQEdIOma7G2KcbzM230LQoGXw4
omqs9G18NtJ5IvOmArDPioiC9UAnIqyRXlQ4y4720FHRCjnBEQHJ6VM1kB8N/VqIK6o+fc+g3H/P
ZKXKmRqAfL57Yp1c9VXsoN3RYFsxG2YTSPBwrtFxK07tNpGebxU81gTAd0bWG5/AwD7I1YcwPoTl
2LbjFuZmulfYCm60ERgS/n8MKVgWIKq6pEcqUPmsgVozaTvrFDYyhNIef7Y6QB0tGhd1TJ902CEr
EA423QHDQW7W91SOf/4YDGtFJXIti2Rev2BkY/qkrgWGsFdSeejWPFEecf+xathE3KPMYkvUeCWf
mSCY2X+Fg/trk7rT00TpCI5WTBEaIj9CDmk28Wxyo6rkmzdGs5l0dq4XbpknGAyGGd7DHvrD/9k7
fuMtWRG47gjwooFS4yic3ClNcMaUcscF6EFiALvcu5J4Wvfe+3FWy8m0q3XxeiTrzz34V1wtsgLy
15vpqcNaOCp6Q3LE7cn3JlPxEot6s3uAaQafzJf7Y/Q/Xj70SIaKdPBE4RfXUKQXf7ob76SaIHIe
rZ/72VKXbwUuw7jmKbSPlOkAo64VAiVk0uHb/L6fPdnvS8hcYPItQU+PNOJRlAYdH3EUvp7/hNih
DRH1muGK1qkpsdd4fJ7uzd3A5RtTc6oJ4kmr9VMcL1yU4UfRy3l88G92oNbNLS+/aSMrtUdHwoFx
O9AaoTMzQ6Q4KrNYrRi29QXqAG1wAJm6avJOmDNqk4Az8EVJk2V3fB281TXX4SEkLAjS1RfhNpBJ
pQWQroNkilRKsr9RAYHrkmn/bp/LAeOOgyyHYcWpOJpzyimLaW/SwdV/5nHvN/oMgsKpr6/lA3Ou
4ctJbK+c+JVNXsOpbndPGXLmQ8NJh7XthlwQK6qvZ1qfGpf+Sg3ha0RGMdOgWlXa4TLBJpe6spT6
mFIdD6t8ritsmYJ4mhBK5ER7vvCHPH+M+ot3rtG2jzS7JzcvY/+VuMRyWYsG4VuxYRAIptj5qwfO
KHmjnrDwxJwLJHjSRCY+7gEdmrya8cOawssOlkkwzp67CQXR+nD+LNFPkhXoJB33YX1Le922aEeD
JkUjleVQJ8bgeEyv0n4m7y9KMuL1ZfBZeEHduQv8gnWv9ePXI1vneDRoKYS8m1hsQdX8vEEyXSyT
fCxqdamE496pldF4hqn7nbWKT8d4YWDjB+PkSR6/91tEH4aCOhjHUQSdqBj509WVRsJHb4t9RTlU
MXiGxahF8CiZbFgeV95ZzSomJkspez0JZspFEDRKpOm87qOOEh8ixcdSToSPCOBCR5HrnVhE249C
6jzKa2Ov0S7+1awiP2tYBuQDTLWtdROEZWJG7vblnzAUYrdHpmdSnlYuH85pqyqzWYrfIPGtcq+R
UVREainayyR31Ewi2ahUc4uL3a29AnlfKUisSZ2mgqMpIfTC35tGTRh2JsZh8EPfpksH0qw6GBAR
gM2PW1xL4HwAHFoR8m57VHcY2rNPWPU/ldxYZrmDqbkPUAgfTb3YiPy3W4KOMIGXDvjVZvopXV6e
uin+GJRbqrn19oEKZWd6L3FUOx5THIWCwT0Fu0z41A42nBNGGcprfZga6WEMPFc9BZ3R/vuT9Vwz
o5QUL/c5jg1E1sb+S9xs94wIFyqafqXeG8JmF3t84yH2tA1Pr9tFwKe6hRT8VU8yPNFhYdgv/Y0O
g7hgqlWWImgWObR/LZAT07ik8yycD0sDd/86f4MthUUBmuEgdddluWmnOjUxj2jv6711AJ0nsoRR
s2QNYoDaSZWW2s5ivFCVRA2bVGG3GsVFZrVFRRsULrwH6c+I0osnrvOoaw4pWkEf6uwKV2qBEWXU
PpnNS6vi/YWpLlViDu/NQOgyH+q/h/vcfDwa7jxsPv/kB9wAZOMo6JHHVDaA288o7GRUCFPQzxmF
rlDgtLGSqv8xHUCMncJHL5JXNaP7/0rNkm8/gRwzAK6zZ59KeWL5HYFxCooTZ+59bZGSZvKeKDmB
uU/TjSxbpzEnN79LNkTkUjYDQThoBuG6TGS4PeesEgN+BieHdNSrwH6JZquUeXzr4FGfFPzivbrs
sxzNqacwUz2Kj/L4wfZMxgPV03C6tBjDeca/zXaIBBQJ83s3ulXWhoDiVyijJEFRrvw0XZ/1COHV
h6K3TPfEgNEoZtDeQFTbdpcpKuGpBVWTmJVFHoW2uF9fl7PNHDxkIZtnwKdtFM1tT7BTqFLp2+Ra
7yFe2gHh6pQvXKomt2d4mLXaqhkW06NuPV4DRnBmN581M8YeCDa0+jvZ7/9hpX36GToLrNd5p/Es
ZuILT5Aqlx7KWg8S7KhwahLSraAy2/wEEghg7yoSecnDEAhnzwo9YfPz70gvFZs1zgVVmHwJWaeE
qMLRMrUgNffyb7H/8vh4XidYQxZQcOwbPguhVS5GKP2R7ajRRTg2Bxw/QoZ1WDXU2oPC91N1LHK8
lueCbzCE7RqCRRgK3iB+AIsHtyL4dwP9qWQv8NkSy0CDz6L2ou38cza3EuQR2Vxr4u2hbhT6g7S2
29nFsDcpte9995O53BJC438BCF3fp2Fhz3mFRdtmXWYcN3rekHnHQryi4nPb6A1M1X5oka/w9D1s
xGks85tsIhU2X6ip2HoyYCxrtW53lEfbrAz7c/2yzoOsPYv7LmocfzXccc1TMWZp7roJ7l+YFyLs
xPPztVi4LWilZ4VcwP+MzziGMhJW3Of7Rl/MZqLORFd+dB9RniwiDoLi9a7Gz8jDtd6mxXHhDjU5
0iZKnyZ/GoNfm1t/hHeuClkLZWyQQA9QOtIsqwmx1ZXnb52Pv8aZVrvKkjkxvKtck6jKMwzLJ2CO
ABefoJpAx+qoAneS+vOHLWXEOO062LneLmaqZwUfy7Th/nIHFDCnIzO53VpgNSnsWjgG4G46vqjg
8oH/zactrLrFgHyhGCz60RZdrmRWSHeB4h3Q3MfLnjFWT9ued821Oq1zrFSsGkHE4WvmJEAgyh9G
zR7M8Tqaw0Itgt09EHAd8gd2/dShNi3Xts58mfAce05oaHsB3bBt9uoEr/XpFBK9c2128sPZ6ekC
l6DpxGfXUjG9tLiVzWDPlHK0e9n+hRTvZ2/iq6CiQnaCno65Rio43KdBMLUI4RXnGJ9F4jRh7VPc
VyfZm6J4pzENKQrcfU9W4BYOt+QvZTy6HtG2V7Jv1jhmvucRp25U3zgPvG+UX55mGfAD1S1urJRl
DdcdelYskUxXc/0RN/pWSfAxu8+P/07ra51bn97+7rDNn6ySqb5BtU4EIrAF6HN7+HAbtGz20V9o
Zjgsq9Kc+Jz6r94hFUqRz4w2jsFkDuGro10WYesuCQuAymaDGQvmFsVXVKnHCxfsOAuzl1ecBOmY
4lF6+jWj4kLT/a8M99tx6DRi/5I7qEp1+DtHhBuvNRlfBqYjiIdDxFADEMNSdGYCCHxDoJwkU6Dg
/v7VHcuBj1jMDIBVAttEnoeqpbHOQzWhZaWi+gWRp+sNXkgaqF7K9taSahltMBsAQUgTV1y8DdNk
6gjeJzrulkhAlKYezV0zObS3TDzd4S+5o5ovGuZsPRCervYZWgwKtIepYDD6/gPV3H9OoHbSscf8
UebeTBhtko1c27qzWLKknZblKqJNG1Fh6vHF/HIIlRUshwQ33r42ctdKIiauhIXeVHulHlqBWsr+
Hyw42iTSHMEYjzmGSmVtnGpSZjLIkEaPiBAuKyj0YXwltijKz/ia7dW7qhXAth0xdQYKaqObJ6+g
iRRc7eU16Bc7+1tn6y4wNxkGYQfGAhbks6LMYRS+B7SPvri/ZPFrwxuOK0aqgbA16wfZ8iq0I2+F
ChPmcEgtletq8bfw+rkRPq9jB2f/tfsUsuOCR3GMcnTGoy+wQKsNXbMt67PtKn9xzSodvraHvuHs
ssvjTEDMFN4k0iGVpEv/ypxf+6edkOtgAV4GWkAlQGxMiY9nN2/WFyDCv10LbNZoZY14Qv3bblMb
lCAesb69V8iJBI2Spr3znKfjezRUS4/v8xY3M5WRyDEpoiHyTUSjVEMsSWhSAeyLG675i7XKZxjp
Qnvh2TINMm5cgei/GHv1QGaD3Amz5vw2dr7P6dPCr7HQzCH88z4vXtdfXGDERxrBsC7fvCqix9VF
JrfttENbi1eJo2eRCqMmNxznuqNPenufHWEBqXyfhzRlsTRL92KfnWvD4X2sMxnbiEetCNnmEsNp
PPBV9jcCL8c3agWYPw1LZv7ypPq6qSRyj699PJYdS3SpZU4dnqaGTtgYO+4JW7lW9gJ4Yy+p/G9v
5cFCc5FnRJKPzagIhgVQUqtii1ZORdC56LLkJIPX4debm3Lz6Fqb1mZkvArVMsOq3IQK5fdhamG6
BkBC9LyTYphRuTweN6B2TZyCp0DH9Z/zjUOPCyftSBDprRWmliJAGtplQ1SfRVwOdoWBzRhjZK0G
+MMhMk/MiQWdp1iGDF7hqYe/dj0abUxwCi/4z/cnod9HH+7peqvoRSnDSjLw9bDZ0FZOOhSPfKkb
Ghc55DH+8zE7eVoFfFHBwZmtExUUWTu1kZ2C+JqGRz3N45mdz4X9YXQkSYzkCqHJSgznKZjkBYpI
DS/6RfDs5UN8nEYWphfR1l+hhnmw21NRxYYFJNYTI7wt/mYL0pZb+gyJ0F9V+e1ATTirtQl5XWKS
aHAkFL2tvGW61+VsysqyPJXuLONgFmh+YfqGhSS+1gcUdqWjE3afINMSFlf+PTAgmgXJoh7ohtX3
RTnCC0TaBkFoTUf5B7dkpUOZ4wn0VIB/EgcmkvQfRVrYJwh2Kli753K+4Gigdx+thkm3A711bi/E
v48pyiisfZgAY2nWpdcr8VRBjacTinxSsDe9HBoqH84p09x/9/yeWga1FjjdHCwXHB6OhrdpJ9oh
pXU1L3ROo1dVF0doU63MrC9bQ+NMUsbmraUQvdrxSTKzuEEhFZeAX0dSzgljUwazdL+tgObfio9I
33IysXB4aV875qFJKM65YWNj9bz0DAaYSKI2qKy73gCajjvIw8JBlclaw7+neo28qViWQxcO2j3a
acvKbvw9YC2i2uz/mO+bI/CMNT2cFT8sCP2Mbcx15ZiUH3VhmzfXbco+sGA1xLgPgalpsREYSidE
bXeslFtOlayCN5hvdBFWlHuIQOqtpQEFOdAp+LngzIU4z+jDFHMrPYYGWlEUtqSyXWT3ROkeWGe6
o2JlfB2DPVE3t38MhLMWCxzUDu/kSu9MCqvp5Su7u3Krz3KsTqAfIwQ5jdCJP1fey7pz5Gox2MUX
xTmYW+5j8V55I/VNVc23PDq03NCvIQ38pkfL+epJdoy5xIxc+K8ESq601uYejqGdXnACuCZ6GJ6V
XtScpqwp80HoZCUVJ5UaXpb0msMa2yg5naVIYFB5wPNnM3Bpl6dPxcpGl/KWb+w5X4j7ml+3xqzC
+ExRggNbC3QZxiemWTLvO2AyC99qrYecpVrweJCXoJMKpfeOKWgSW/BM2GmTKDPFFn+o1OzlVz2K
jgK1dn6J1wX6qy1HMOHA2+MlenfHjibO1BJlyy8M0fFfUhLlDpEEJIDnggERgxQB+tJQsBHO+AIG
D2IT1Jl3eutVRdHwQYqYA0XlIrbgZ3f3Aju2auDPGfWYljowV1A7K9hW+3DYcAfrGPyFGyEYwA1H
N0I53jpS+JNk/x2xvPLtpenjv+hvRQ6Dqar2Hj8p3BqguCc9Z7AhRiCLAAmBmfD24rXbfqvcHXGf
76BIFQ7ux27Ts1D4pFHSrUTLoF0wVUfr0HuKbV/U9yLx0bKVwU4/+j+rcihLGYvxO6+VsGWEBPFZ
PZ5T0RP4wd3tKABk9NNslBY83C6u+sHEM8nHk5pO/22+Fujue3n1yhEQwuSmrENREuk7sLk6nVf8
WHM9H2JkYkbtEW9WJV/bUBpc9OsBk2VlhNHr9df2sT2q1lWICfQxGdx7rE8dlCKuNkMOjGK7A3Ts
QgmrshPmDyz+sa4/3Oao5brU/N+ynhvJ+ncWD7bp5TW3IycRnY6a/S3XEd0mP5MWChKdx+QZIkfY
DcKwYD9M5mEojJJXUM/t0sBafzgKgH6MuIE5fWQY0Jkly2UFlEt3FaNk+tTDWC0/ubTA3Nz5bqXe
UUZ0gM11G49HVgfTVk9KqRWZr/VYiRnqdzOquqVkepyEAtLCL4XZMTyL12dmDwW+jhVNHF0jOY1W
o0z/ixDmjtpShgSCF5Z6VQ4M/VBX+rddh6lK+8qtgGp6AObuFBRqnxJlQnSwNfls6DHXzEim/N+H
JN5yJoaP9JrHxDwUVE8KweVeinSxcvmlJEkonKulJKtILaJtpTP322rSD1PeJKRnxzqne6DyFMa3
qvNW00rEtrTOSCIgDekZFcVS7Rloo33fCAli2Oo6g9EOBS84HALbBH6b/4gN0y1oAXRtfcfrnU79
ttDOKZseMvBN+25vqE4vi3KXiloExTaXJJX9BjkJEXuQyXXefedkmxRQ5DxJPyNzLXmxPzU4ZU9z
0e7J3hohrv88XgEtya6hxJklnFMD/cfld6PA3q05AOwGibij1wA6PEuoY2tvbvny6YOt7FtCVJEK
DLPBrsm2WqKB7JWKQ12EVRMu3l4gQfkAzy6GWjtLC1NEJBoq73LKdvK0IkS6DBUKKGJrRE0bKtCR
ZYGt410+dQIUGYBUPYYoEikS/DmSKbkGcNVKFN1JloK4/lsTGOvrRNoYXEMoeIi0MbswO3ZulMRn
VHqKOdJ0QeZVsmdMLICSeVkDi5jTu5kI846fj6L9OpQJ3H3e8a1YclFLPtrnYrssCmg6Uecj/b2Q
TjbGAbvTlxtFhwQCrWLQ6g7y5NtRwqdi7PpY5ySd4OcwxRN0VDyxHWWAlZtm8Xpkrb5/a/1uPu3Y
hE8BcDjg/ZmsvdN+QacZe9dJCHA9e8URfZm967Ku0OHHvUCCRV8ey4rHVs6ikL45kDDCIS3fvKF+
4ogpDVUTz4gZK/J7Y89dvYBXnpf4/Fn32Wg+ufn7g527/dX/6mtXo73pU1DpcsjAwtzxWLHptJI0
XKlSKsbX1goW+GnsTFvLVyTOfPyrSHaFaD27Np1k52UyZ8vZEDek4nR2TiDxdTB0IzYwR/uIb6HI
JROBpT/AaVwnhjOSotwpQJ+KSyObzpt1b9ReCUZSEYQtYGrsLsV1VVg4PveQTFdn+TuP23uBwDiK
erGLKc+MJUp5O+ny9lPI3L8Yq8ReOvBdu6/zhfc8wnGVw854VQVL12gR9u8pEXT/KihI9LXwpTec
562SOW/60rOQOOUTNmGztJp+akU/5rnakLKnaCnqCobpdJox4zoq8XxSQUyJlhviG0xkiHDpn+wJ
YZhc+nNz2JbiSeZOZzAYBVge6SLqjjSAZllPKenJAF24xNriNxKUfwjXuRJISM5MK6F3EQyOD6Km
9oWMng/KTjlBbaJ5wW9bHxocGD6Nudqq401t7SLUqm7aXCic19r49A4GuFu3BEzU0j/c4RgSsUmv
wWXCbioaNl2l/OwLk47TqzRYGNU/5jlHTl2HqxTGN1gi1jpM4NaciKJYPb6ujqdDH9q0sDfkp7Ho
ACEyIa5UZkKer+bQAqho+IbRwrvW9ijyceHRGs9ZXmbbGsn7jGLDK08ToPFTyIv8iWQtdwHMnhlI
CpbzdsgO5dygecLLEW9H7Alf4MajQxp773oHFiYZHw66hmVZBw+mbBNRKUQDShH8CjRicqB9Z5YV
i/sLlzna+h1bkJGlyzAYZJoJEOPRh2/S52eeMoUjna6nabcq2/oeBRGTVj3qYRLnN3af0wZDNqoI
Z8GgD+b+sbMZSFRvXE6wInKMRYqfnEkmzhuDsXSkjgCwaB0yAx7Oxqp3Xn4+JXGjEsImTIKmH+SJ
cypOTC/t9fo6cA6gMO6/NirtUyvY4oFUBifORjJ1Swws6KUVDNZgcS9F6VInZgb/9ftKana8GqNo
wLX5stbmVeKtJPEThG139ISw3Cn3OW7nnCpZnHIhCdhlNZRE1E7goY6Cyr/sDg5HWVCRj5OYGHcI
TTbduK8gsgC8x6qJ57oBt9E6NxEoXoirzimVLjOEHe3Epek9Y9WSddQiycmFzqDmsJMIEIVWhewL
XuD1O9s6sMY0Tuzzv8KutLXMq2F4KausK0/1BtPa6cVVJy2/iVbfqpQNFVQDFbMsYZGkP6QLi/bG
Jq0yw9wKNUn/6rPnBpfj0uh9zp5GYOPdYRT07lqaAwcfPvYSpkKUCvdlUcTDalbRi53PliMj0JEq
lUMOqb5tLU0rQkDvNTW6MtnXRv8HYgq7/kq1efDrkxctsztUOwxeJKU/90rKTFkP+qGk76mbXPd7
qLPzin2eSLNy9LN36lCkHp4un69vBhrnNhnB7uCfHj8TqvXpiRGKZ1P+v40b10kNWhv3AzEq7XI5
rzUf33DIKmyC2NlpcEICS893e+r2FwOgzXnKk4cGg+/zjVmK8z2L+YEbFy5mkgANQwwiODPfH7Hs
KXU9UZVmj5Unhgfay1meGKRQ2saBA/RiR2aXMvzaP7ZadDFWcgTkgWBKCzZiB6IzP2uuBShYLPN2
1WS++cEjEzsPeoWpAd9wFDstFXcug2/mXzTWNjVoxR/JSbBkKfmFhCIwtiw/YEYzdJPuzzq6slqn
9sfdJV2ujQ1jS8MkDrTaweNs9otCJsiYHxuzymzDsOxM3do1X3jjXSoKY4cx4xa/aGrLuClGVfrT
JiT+QumqbyA8dNQGkjt9JqKNFi9LGC9pAjaPrauQwYHalvtASV9uX1VZXUdYlJ+kWLrcZn1qqbdz
5Jsa2if94PzwwClvUNMi/GUbSOJRvJAVYJC0be7ATpA+K2hwQoDPsCyAVZ+4ikFi6u3cU3amKslJ
0L5GOOTIJ3pa6aCF/rqKX0kEX+96C7ra8WaWayThk9kAzk5g4C9elcH5iiMbpzi6QLsHEIkIXfOK
0oZNcGK8j00kUu/8+PJoBixKhhdIeQ08Us79Q002hHhGBCtQk2JBvg33AxzXyTmPBBPzbsdF4H4V
nJy5HSwQZlnDoS4N+NoXZxr1uM3Oce2cv1TmAw9LuTy2TdNwbd95mIvVyPsgbkPkGS/ixkezv643
iK+j9WR1q2SpLBobcCnVEOGXAznzWx2uin3oGsiFJat97Vc6dvRhY6zgCdN+/xzGN+ffZtCut+6T
YKuhhdquyx9fjBA70sk8ujp/3vv2oGFG+qonu8yEUj6PJiD2km53Vj6RtMY7fg8fP35IaCXGlXYF
oWB5PfuZuRpJiLqCD6nk/m0SMvnUl19igptBsLXkBk9bM2xVxUy9AiBKHGLJ8Y5kqP4m4CcDybu8
UI0AeAts9KqTw+K7drBzgbW2JW7UH6fweAOIf0ifJSVUVqkI7rxEWwGF2fmHqwLtILxyuNylXDSR
ZnaVxpz94knDxZCVPSJsYJrDquEQx/+R78gixs3hSdfTs69EN3geiedLHAWP+v+GzCuQahpre8CK
dhIRs8NNh7gzTuI6+moUf1nlD+KiXURqKU+ubQnVE2fpivDsB7D3Jiq2hUALOPze8O2QU+ySHysP
jyBjJN1a+uYSL/5TcJPPzaAeGXO9U9EVQOo98lw4jtCKvKs01RTfO9T5WqKjsP3aZkEUA8wKQ9NP
+4ZnmA0TI14fNt58vAaQWAccpfDMNS6BWBeFa/Zru+WWhfj/ZjWH6y1gqj+qC7kSNvrVOzlb4CdZ
AKuNbfTfpGaGJ7er67iHc3f+mF5vbEj2HjkAZcu/pARM6BpWKff6RPgfgVJtQ4sSbYLMIut3n/2v
uEeVW+BdLbB/xJwszbEnDb29Gfu4gHV4Rx2aaA1GRfw9xAZ0XmnoKbEqpD/mpLBKLd3YLyQUmRQd
JpYK0A94C+a/4KwuVsimKAQcma3OR0TOyd2Dk/IDfQU6jloPLm624wKOG/G7F+/95Um+OdIvpXKY
sw6B+S7IfybFvdLt7LK8EO5/ji25Ec0CQv0aUcnnMJ3LgBMQB/I6b2dfICAjHte86ZsecrukWPu3
rdZfDSOzHVnkuB1amoJiqiRp16b4XXht+dgm3fsriYbOZjL8yaCFi3iBBGWKr9IkWG701/+v4iWq
eU8nqPy+i3dWzTygta8rACphLf7Clb6sMHkOt2NxfY9/2BpymiFOaXMwAcR20l8V4IhhCr+bB+wi
VmduKkd1mcvTSLgscE6TypX/TCbFfXSRkzHGmfE81YKeZAILgI+yZ6gq1QIxzVcHswQJoVrf1VYK
C/pXrzp8w8msMT/4cwPsUnxdTc9Wvc7VHrJRMYRptgvOTAdFcF/QsAUBATTt6SAZEfQnSmtb8A/y
/6RTe5tAucn/XL7XuTkVFSHXaKaE8+eDgoAnb9RIFdew2oA7UlhHpHLIswqqbUstbvaSOY4SKNnL
qnmXnWASqteu5yDqrFXZb5PiHRS0mKrx0GeHYNDZYEOrGKgWbvkWBvbo6B7slH2OsNNoiy5CenmO
myc7bG7CUUiemB2evQa+2z6XFxSDeAdTyySo0ZaXrEn1BCIeEEf+jCXoyCqVE2htJZwzntR+cQMp
qVu7v6vtp7K7hZl+t5A1MX6pmbCfCUgKFCUN1bMH3aRXoN6Wv5wakV5GsYQsGSKIZvFKfjaGx/G9
F97fk1zEUr9tlFlNyPXDdKh1f7D7YvpLTE1fk/UNRpYHWYnq1qL1yMM1O5uD+IlCqy6rX9YBEgnj
S120bKZ2OFdKT/bwN5ggkJF3QT6FwH1edbzP8oKmZqt97uOsB0NDhxq7ZaXQRCCQqqdGdoIFpBum
Oc2L/Gt+Ji7mqB/yCiJS1OPaeLV1roTaHmIDhtBVz+KOG0G48PumejdfDOibU1SepZ0WTBc7Uo/P
9hUqVjePqjv32vhEMi4ZzOkWxvyw1y5eucUoAaihtc9mbeDA3Qtd8trt3eVGub+GYfxMUDW6L12A
gt0/cH1SPofLESlVbyTtwOh7kYJ5Jl9LiDHNAyvWyt3s6O983olKtdDGgV3ldq0atKAzeXBQtsLU
Qhbk+dTsox/JHLTpTtMyd98G7a67vmaQaObVp/8Oc86YAIaTORxwfz0sUzboaHKg9m8C04B2+s6r
KLLygthsbf1O9ojm9nndS0ZVMLKJvJP7AtkOCuqluXtYPMcS4jSFCLSifUm9I2v1dMbQXYTj5uFR
WfCDXUNFaFsvGxFjm01uooCtGLjRrGvqpdnvk1+ouG/cmQ35qppsI9UW2y0/LcbEg0zLgDHQYEjU
90cZ/Fi+TmYBjXI2dnedTb/314bPTRxoQ9eujISx6PEYKIMizYkayH3Qcn1UyUYtCdZ5JfNKBcPX
OTTbhKNXbgzRKgG9UZWzjCObXfyD7lSfEPWZibUsxRMCcc4Qkhq8Dyw57mGO9BDkm+hcspq8RNYd
pRyE9eS+S85NmEiafTA0U9M1Pjb4QxAXH45bpMsNs+QLas3WaZl3RtgLXqlNneEkGUsAV42QFeJp
EKwGYyQzS9BXnjnc20HrlrEf5vRhli2at738Q4BzKlqvoUv3lghSWLmQKNIplDPh68GRu8jPgGnM
B0n/JtWgkhCnqKboJAUafWu8AhGfJrd0/NIW5R7fyj11HPWakca3B3jIGKBqbVDU6SCu0OXttwTz
o7Afel2XRBIqkTqxsfqss9EE7deeFmTFueN+98QRR82RKd/h8EqmwogSsHwE+muaE1+GlWzb3vgL
BST9V+SBi5Tyg1t7Rcsdk3eRWw+bvVb/25sPeklFFRULxO/8zakg3pAfnpHqVH/pknqSkt1uVm+B
r2OGPS0ythNRoFRmWDA6kAdDy4gs1eteyDlJ6HYzTrfI4EcKlXi8ABUzapC7rZZQCJkR3VynAe8E
MGBa+UDA3x+e/h5xcL0tD2qycPah5Kow2nXNIvvMBafA0ILmlLuhSAg3k5d/EkHUr/DOBB4FhJis
uUO2adyQvaYRIMp1umonD7T17K1D5pC8Me37Zj+Exb5YFgEQDRwWkGUU1rwBbm7B1j58/Rf/ltIj
uF8Q59hqJAc5QY63dYz9K4B7HA1MZULMt/kq11WIlByiB0ZDbJcC5vk7bjFqRo8HORzSUL0eoX+5
emT7C9gq5FruYzksSXhwu1znfZ6TVpJCJuRed+QAl1YHM0HobHr3GOXg2pGi7MAXSMevHN26UeHT
iw+ncQHprhlHMt1Jt1jrFaCNxmK1Y1kX9ycxZAraexOqzOmOdLCCCcTcFYdf+A633Mw0jGpVxXL/
7SPRQZe6P6aHvMaf/V2c+SanICtqrTMrtEyHjLj3GS3TBDJCUkvejKPM9bhy+a/9sfXat5aQr+3H
lc1IMIXKSFG2kCpEP+EObMgaf5S0BpM9j6NhxGaBmPDHYBK34ewSJ4oPX4ZA+jk9w1c2cByMTd1g
8p9wr651s4u9S/GvIJY66CJf7GneMASh//kxtQZ7pujHAkH6IpsA4SLw6DoUA+IKGj1dqN3mRb7T
F7AQ2oqrtRuIl3wG2bW0QHXgqQmO+cdm3PdQIHYZgM05Q4IkYlkChf1LFeBRFW/zwiZHJ0E+oTe/
x/RYCGGE3FdLWUuXbs9s5l2s/bkI88qPvWQ362KxfyPK16ObPRg43svWLDbW9HRmKi8FIciX/+pY
DiOT9oufN/mO0DDUdYvOwBiWwEMwKHFy4bi4wZjYeItgEyen5CrvCDFCAYhBngNzONH7Kw5SDh/O
5ITYmqz9EMaOxjmR3AtRpgDWEamyJj5hIvkd5qsY4dEYOs6LSTcneYRGE/TStehl4vcIAtgMSVpk
uETt8ndsk6+hFylxvaPFxPKVNOYQK6vGT2qsATWHX2tA/EH/41loF8C9fWWp0x2XCZgVxnraVSLY
JCRKm+RqNUwyDdLR7ehdKx/Jzcp+7xTDvFRu6wVeHrGf5VZpPerYXwho/HNng3qswBuF3hUylQlU
fv5yJYmAWIs5Zp3noMV9k27JpPeLoEpcPllvsLaMBWvwKj4y6S6Hyurqnm14IRjSeLzKajj6Dlss
bdKB42UrcGIQhOhcFpDr7v6t02d3SMnQmYKLx1OV90desWSiafGm0JVV+vjE+ZC2P/ZFT0q7UEn7
AL+t0u/LaohX2WZ8CSe/nYIlKva4DHnmlPXYBI17zV2ZYDMZk14YBBcrj+LRXmk0sFREMj/bmHTC
p586l6R+n7vQSN/Wez0P8NeurtaA34/WZUGBMg+TDCpL0mAEPVL740FtvSehTT+tVTAUUjGg+kDI
PQnGuzjdzcM+1jNbGaJ+1ANXAOyWc2lzA9RWzYSP6V/oDk6mgaJqaDLxyqfh5QQbaocTyUjtbEDj
8DBj0F2ZVep8VBqWolR99ST4uUdtW/B4xHZWAZQJXhzOAYDx8JOx8AacKAUAcHXY7bEKCflRV0hE
ry+eMHshl4LHm2ga3+iQZs57xnsqWcHbAvcYQk8fQlTx3zME59NhBBrEx3DH79aVc+VabxylTcgm
9walMn+i+aNFOFygjfKGDlNITvAH3RpaEkPTA3JduVrntfmSxIW3GTwpaYu5xYUXVXtPYLEbmrmG
TXtAc+fdu98XWQnDAKXn9GY0AvxYe+yeH204ujf+K4TfE6QUsxppxMKWgBoYC81vCWO3eSZDp53Y
MQITTLkgHUNX/znO5gvZ79NNUeoHCiXsG3LFuYLU5KQrlHHzkFi0q1a++y5wQECy5JQzYOR4qcy+
ESHO43046Gw3+jGZtZfHNfIVMlaqpS2tm/NRwV2RW0KfW6OPL08F5h8yGn3/MGBataNkjb0VBdn1
gOrBzhxDUoFEX4ee/RVmFjbpITObFb+IMR5iLhyyfwkA/pb6Kxk3tWtZfXq2kLGI4z05c3G3SGyB
TZE6/twcH326RhheEL+EFLbIdAl7VaEOD/Q6zVAbqu/RUKkkTVrS4SuCuwmmXegaLcFbJtMTYhSR
RJ8IVFJnpRnZS/ElUlFdR/sl8JMFq6NLNBbKZ8JybkwGIJMXRG0ionFTt9loQFZtClSKCFSP2OCn
+/VxVsNSTRM06XHVAN4eBoePFaXKCSthmJzg3IkTg72QlmcfmO6xN9txdP5+STHxIaPMD4XVRpBD
Po1+2pQpokca7S8zaBZZSfw3yEdR30/YRTv78lfjgNQANqnwt5LaKRE+FSG4CvChI0vH4f69xnJx
6Iq9j8Akoo2wYgsrjlpR2KZ0mYBsDEeZ9mLb9h1EsGg9ntdREEUfWP2ufOuIziPRDcgasW4tbFAT
VmsmgMPzgyxXdwrKNloJmUC3xGajsfHeT+zuN6XWlCx328WMOMxDap6dW2nqnqWFCIQJ6De7EKlV
hTuII0XjYt8mqE2xIBhShgqbcWBinFZN49Joy3E5JkHlQ0rXlzvNxSV5vfpUjrxCALjIa5ZJLarw
8xmgEFXFImMQ3N2Iu/ZSBlsx7GkVPGOA8El9nhFWDjlvqnyS7rOV9B0DgafkcQUZFzZsfuLdWZJQ
cKwIN84nqPLDtm2FQ6lUU6Nnz8UgtpeWPPzq5KHiQXo6SxOqbOC2ou7kHVoLr/VaEMNA8uCCDAxA
tIfXkO3Rj7DFrXO0wYKlQcP1CzMaNJ5bBKHsfM4RBNDPE1IcTQvE9+5fNgkQgfHSPBvziSptq+XW
iPybt5wXhmJJnOBMXqrIc8CSxESl2lIqDPqDXh8x0resnde4XuMFRtOdd3Rr5tGIrPefJ1oi5c4e
6CTEyqWOnH627IBbheLJzsZ8q2d1wM1DKXpKxLM2ShE1NwPUORcL0yoklFdGakbp9U79IWw82KB0
/elc72+rESVVcsuUg7q3dyykoiNXt0u1+nZr+Txz5lzhmeMCnpLwzvKxATvM8fKvJoWar0GWWpyU
NMhSTc75FWhUAFcYqdvqdSiSc0Qp12AaPGPoaM7rJ81ZDB+8hGmUl0M1rHmhgTWgJh/9oUpPTAjw
fZT6XocbCU4UVsR/a5dOu4kWdIuiuBwxf0JXa3K49F7Ecj3dMEj493fbUIPrSp49tb5xU75TUELr
zOF6fIr5gkMRR5t9lnKnY51dO1Hxt5HLUyVbLNoiO3xpkMOV7IMuRHWEKqKSFYt0EN/TZPw2Nytd
BSH9Gj/gOxS43iYqYc7dmwMj6Ap8PlpmCmf+tdlgzTYkdUVEN+lo9QfBALmc5mBzLPBLydkFgdAn
G3AduI6rQnt7C8azBMuizCOiDJ73Mm4ZnUY5vH05pvEhUqhdbgHY2Nv6ViwBaRfJ1VczKEiIj1DO
gislIR29EV+GsvABmiyKRPcaddO5mUqFWkUIV6o+uS9Tth2Rs07gwdTZdvpGOzZQCSRLLIYO1Hwl
Pmso1IzpA7WDtkQmmvY52bZ53I2voQntFI3Szv7YMYXsVtl4XtytuTNs3cRdWLsPGPzV+B7gMVxD
aIya0RgBrvnnMdpB8znFDQ+SXAXIHxnKZWJ9GpK/yTHiuLojhXYBBMZ7TiEyNltnsudUVSNbX095
AWpeix59ATGxgJFiScrI7EChxk0kkbqv64GsRCj417HZnIl6IkMhAztqM4304zYD2tK23QiRSoLe
F8KsLNl0/CcskpALp8nJnnMjAy/YjrL698voONe2rd+oWJpzE3TovZPwJHezUE4Od4Dzx5LGzkaT
OZzSgJTfn/3s1lOOKxgHrM2A4WUxJhIIIkdYr/j1ex2ira4vP8l88u3osScyq0AuhpJkIC7g0Kqm
zNPf4jxV7mtnasx1qGIIr7bj51f+xmZ4sRRNR4igMGUbWHL8R0ewzTf1zf6xsz6bkRc6frEEp99p
J45z+/oaa/jYQNCzxzs9S54XDsEr6GMitjvLNZvtWDgODN/Jel8XiqpC0C/paSWAzF4wlLmSErEn
OaQneMrSSCIdCwpkBHkXX6TWnppS97uiZMSmujF/+zW6hztgIJStgKV+Ek3hdNh34oEELlF5cDTr
osk4yZ8v2YFz7kaKrwqqmDwmLi0+JV8gyiX7ntiEKjh3zM6kavg+q4QrxG7Bw2NtxDgJni6+rCw5
zqfx5n4EVUXqcuaAIZSOQfezAKpvahKjJLrHLfexA2BZH0KIrlvi9jv07axCDaKDacHP0MOk1J/s
GjuCmkfuxUMTzbPQzAXm8TmsNvQ9WOe4B5+WK7HkKXz6z63soyAbKLnH1hU6gLW8oOl134fHqwst
Ob5rSOKtXRFD8iKFj+Nj7e0kFHw30FCVdd+2JsDexRAdqw1ZG4L+GLG1lGRPxVDCb/z0H9a5yhL1
e+lnILjnQHvZRSLvJODCCJfo+suUrVh58uX/ZLQFFK/Avtuhx3Jlg0nG8tEclyAapmBYY6YETBnw
4JcESnSKpirSniuSuiG6eIQsaYDgTm8LhSjvMPcCPdsZ4FQbgV5WsFxnCgFDx+GK74fC4Ar9cvKj
++CKPMUhh3PHf1zUPhj3TIDhqSqkhbcGxqeA5674V7atIJVihgzg8E+xMhI9+1psY/1n0xNst1Q7
wJhOml7AYD8TTVwQ8jZAGG0Wk53qMG+eClN2gXcEm/mHb8+4RXbLcA8av7FcmJ1HI6iywaGF5h43
2I1uThG94z0Zzykco6qMyQKx5/XgMeU+zi33MRhXsyz3TK0L3QGgfozLSitoNbYfNeKUkQs1hCMb
U73q2AXXiqspZxOrIwQ4tPGXBa54avWb4Hr+/SK56cz40GI/pFnWH+FFEimDnte4zt+EQTRxfaho
vMD/tNKXPwJfRvda1ll+LgbTep0N19mZe4OiueQTDGKUuFlrfchwxw3oE5d/zReriaE92vIMSqJ1
2eJz3TLyJf0ZvDjCcDUP8e4tUMQzbphIXNUbc3toWt7f0FR0AkO8g3yHhctbG0+xeFYybu0nMN5j
3pN76kYvj1B5vfPhyTIk8Wz1gYJs8+Gs7hQroAJOnZUJs9YTIO53+FH73ntVXEYRSnRKoB3EIMb3
uwPuz+Q43zRu1x/qITcjlYJ91y6WehMJZLM2JQ6AJ798PUlWOlFsWJSwHMuL7IcUg0ry0ea4QYIj
NpJ5J9IPzWEJgkTjp5h/rKvlnk6mA1x2IAztTqwxyd5xgMYTGH6nR0iapugmLL0Pjbeg9oIR3OD2
HAW+5x7UauH+akQu0Ag5D41mAglkmpq0TX93ACd8KQB9adI/FlUc44ydp8nv+hjP2L3KYtXaKVTb
JSXdNaRuY3O99JeIkfR1Y7KYIaUR9GkOB2HQG+j6fqxVj375Y3Jr+pZhhINoPUgJlwmQP4UIwXVW
ksr3hZQEAQz14n/IJUd6ApxoIKZeparf/pu11ZW8fSk3Z0BUVPMEwS1ZM1W/Smd17D/DLBnEenM8
DgGG4nCxwwqtCRDYdq+uwxYMIF7jHdgYg+hvJcTdThx8ratEsx1pB6duuoE0U686XahXB8YgoWo5
Pz1OJ0mj2X1ypI+M4QzLFotZHYegxzzhUEE3K3rGGaJNJLvft5Fq5vl2RCsjk7BrwrHp2aBof8ku
M14tAkpsWNrALnCOrQLwQv+lYfSdKeMVo53YQszDwY+ZB5IEdNntv0QQo2FSVakE7n4NK9Y9zVsq
zd/2whzXAGMmOO4P8DL4dXCrpvYKjcBsQnqIFuhHsUB8wFVnhEGSzgEBSWFduVggagZLG2FnZDMS
0QNm8kl5pF+AInmYs3zx1cCEG12x50GsKRi67g7CTuTfHJVgwBFi/653dtHkaBo2piGS48BqYtRU
edZe7//6mLXTgKecaeazZ4CUMXvUFIk09lUo0WhJiTjipG4RJs0Dd9B3Tw8JXqiTkg+N/V9F4Z4E
23yr8GFcUnVUL3iaFKgtb7IPUAIF939yac+Hd/xetj8G6ATJeShwUQG0e/SUL5Z5HYQVT1enaewv
QWP9THOp66Mgv3jd+34h6j1Z6EO/F12LrVDTF3EmK7abfs9/9ASioBfFUntiGvPJJP87xvr6AzFE
SL08AERMTG4Igj4DF2Q4nzskXQkbum51IFWnw40Mme8mgxL489nDuOMh1nuqUtYsL6fDRtVuI5ta
SanMd4P8sXjHYI9Be5DvCd1jGQZP2MMgDsO1SDnG0KsHUJPU4JzoSwJxMrEZuDZBjMoDLuKFQdTE
at4BmQehFXYf889Oi4MO/AuLOX+ae3INJckcu1v6YwBdOaJf/6LMGl8naqyZAyaJImCfJqoiCcY6
Rfj4BqBGXYKX65boGPfC0I4pzQkgmCeJlLfiJHZiBJDmgvckdba/qrleBJ30wGnvP4BgZ72otYOz
8fom4k/JteDgGF0neMQrydj+hPsxexVnm8dwUiS++9A2Ph1iJX25ixdPMY4AwYS/Vgyl8ikCiPOi
8sdFqBB71xV1FfG72ZBLgPVJXRQtGbM7eGn81sQb8fgXGtHhkPxDV1VzNCa8r2smkM190fs+yVxl
1n9A3b6ecqhoy/2iPStrRE5GZd4DlrhWA3Hh7k8rxRQUIe3oC5iV12VWIsC/+ljvHjpvvsDA7BeK
Zyn60lipf7VAKGFBMwRj8r2uwaPssfHQUiMrNgfGm4ry6QBd/W9+ouaZVFijs2vCI3vJnGBlq6xk
b470UskZecRijkLozWSpFEUQR9cy1ly0+LBpumc8P8mjBazXOL9iYuD3iuhFoLy5QFhvAribrDJc
4ohZzK6fqXGRw32ygk6tf/UcNu0szbDmqHm/ArDW5qLcDfp85PW6sivMJADEuYdewVxlkXlsVgBp
Lbz9WgjPTVh710dqwFnniNXVygANxQBIMjM3nUohfIxxv9Osvm6nXOqYEnunQcSh5Ezvwa9xpWCb
U89sxssPpi/YBrgpE+G9mA8VVqALucQ/ixhF+2TVp7w7p+B91sxOygVrDaadGLjSg9c0q2osZGcI
0b7iImj94+TW/8XiufOQLu5QJBooyaqe7D2pRm4ZLj6rVkhzFv0Ao/LGWHifUJIgXXfbZg2qRZZQ
/dvR+ynZKWwBAKtQvGJaGcuDmbSN3ylszO+36osCCkxal7NSjAEAdHF1wCk/pFUTw8TGsSzdjqZj
T3sD5LeEHfxQs/etE7NNPx4K3PEIE/H01RL5I3XCVRuUNMO9q3+pTiRmrHQId2mFHr20DN37TWHN
y5vvkHzwUhU+BfRAwgqCuX+eoLu3sXMW0ruWf+qDfKkOn/63I/tmSw12Cwfm5w0N7UJ+ilJNmmEF
HzizfVX3XlbG45bjDTlpwKsvDI7duyjqaWmZc7Zu4odEBbUjC/snKU80H3elPU6RnDWH0ktxIBmJ
5gmrSfJMUGhQF5syjCY8mPVwDVANYYBhUGTu7Kf7OJ4jusJG887r9f9uFiwRwOxwoSOUSVJSBmW6
gy9NpuyNpXuEGKv01TnUHu5mhL8ZCeFtqeXMgM7otZfz2y+VcJnNl+KJcxdkX4D+muLj22MbQ/Nt
fW4z1UYt4vBm/FRP8YH9AlV4qr6mfDncZqvGCrtno4kP2k7fvZalhVi972iRgkfpursNO6aclDl+
Z14bVQaUGSPuTFibf7iC0FHzI5YY1rsmrpH5+eUszKJCjK12FB18F0noYRgY+XD1dV22aEmMZwlt
2pYMWp5m14T0vhGV5NCH+fjDk2rFJGNCnKcRSJaMXoMsaIV0/lpgx8EnkMW/vx2C08AlLJUr8jaN
aeF4qsxCcTtyyy3zQlR/w5Kg4VNtXaguNYCWzN7hZY3oMK9FdEyrwpLG2L7Cuo3NbD/uyDBQqabn
XD5HR5eB/CU5z19Mp6+tctHZDdK74PQ3Y/6HufBUb3McmzndNQQiV5wEPXxBNWU93iQVjS8ql892
LymAiawKT/HjNCJxxHmqSZcFnv1YTaz7iL9SSCg13KCfbtY7mH6Npgecnv+31cXYcdbfyHvxMc+a
pqA8v/E+TMcDUquduuvoVqswmUj/qBid1zE2Beq5oVHHFeJKy8/7C3vA3qUOJGCA5Fh/KF95LNsT
b2huJ5QlNTysH3Af9pSA3CIsmB7UBiC+HSH9Adq4R6lP5mACyapppgfQtJ7I2lO6XcDwB89uAm5d
zWmQA36sIqQiNYlNr2pP3dhcgXNOOXhKo8h8xY58f9/Atq+jGuVSXrExn1c7Gm2njzfHds29nyxI
qbISF1OrvqJWVcwYg8jAdh7hyudYQomq+MKHycTgIqDleZTUzoMtHcQyx0LeceapTs4zEy7bWKTa
5ir7yhsCFXmWXen7jkKtMCBKhYRQUrd64TwhgzwOTEakp/TqVPlE0rIeqdupfwXTiEljrq92IgOH
PFZb9RsPQjHtN0W1/sWHOjNt6jnAFM+3/o/B0PN929uMAa01zZChwdi3pnHDdtojxD73OT6/fBnC
X+SJah60ZVkMTJ/fgKkCWwteFPPg+oZz2qGbg88d1r2McbXCH7S2CUOFgbMsptbJxTmq3O9ngYyy
aOfirvWmmT60Xs0GzFQUTIKcCc2lX3foGCQK/6Ygw5VMzTLrzVGOZWZbUMZ2NAI/7d88SNvbfEb+
5YqRZCa2SBi1+s2KZ9BoCwXwXOTFrVr5kTxrIAFAj6cAGnMA6F5DMAYz0MmcYGQ1kk060MlmMhmI
kR0OPg3oHQmD8h17PvdYmwD/DyR+u8S/cy+zQcbC2KBP1lTBlqTqAQrfY5JiWGdjPefqeOS04LKV
lbYfo35uXsGX+xbveku1NLFODahc0CDnREPxSEGXRgpwum/1Gp/qcrwh1bzVmRcMRaosQyDSV1KY
dt2+Zbabp3ekGg4BTQdBHPXzgcBo72mqybmbgpWGb5lze78yKV3GVs6lCxpQbPn3Yk6xaZTK3Vwx
habAfsACN9/0faztWroV21WrXIlNKyLstcoGBkRwRVyZdVd51RGcxz7Fs009lDZ/RdjO6FOkmhtQ
OS7n7FDvfVNL7wzxvX5x3GOn8uRk/DlHz+g66lPgzCxMdQcQuFGmq4KVHzreDxdM+d6KoD+JNgI0
evAPAuAAXMoU/o0BP5Ae5t5OZg8dWP2ZPJgQdXwyIHk2LxCjxujTeWZIGNiFqjaptmXZ1jzZqmi4
V3xKttxZMS+qgJCtvxF1NbAZG+tC9hyF5JqPlQALpCLyLeIR6lOQnp9zzHUaVycWC89QHPVLGlqm
NjFtGbYH9LR72ih8wgnlsdqnecjt3yUo+X5m+zXqLTjjGvlfGMmZvNfcnCQg8wz533pFngwVWWzN
Lxm0dhpBfvhNOGNnAu4+UxrKowfAW89Y1J3Wx31elHh2YRMmCVwTnu0FmheGz4+8CgPYwNssTuLB
DFCSU5BOyQBkaj/yw+QcuJjl/UgxbNdTWFC+ZspYgeCqjOIEKCNCvefQrYsHOvaSaJuFosb+pvnb
JH8O/xFDbCPsJ5cABbPTvSnklBjeBu4a1t+WbUIqMIzxXCAhVCQYi5O0IW3VWHHmkPYComQCQumN
pUin5Fe3mYJ2a/AYqdjXVlF7SanWjj0wpjM6yAubedM8Bv5edjm4K9o2ladTcMMu7HFwtXzXWRBv
X395DAzrbFavGo8tlZKBIYHssr+z9F0pRQQ60tQRjERXz9csYWg1Js7FAySdDYhP/jwvo4+e0fET
QW3lPxkrDdAtJmkLsaP4Vf6P7nw8a0MpphoxtSeM1mwhTNTDvpLs1cvXxnS3rrkpaSO6z1I49b7n
/o+4fFOqUwknJ0Ec+3jjup8Ux7gzuGmneBSdX8vLILUy+wsUC7Wy392TkpacTU1J2qvOC+wKiqzT
bRNI6e+VXRnOfEp5KQGOg8a9gOw3w9o+3qP+POx7baTUgrcQssnnDhvF4xPoyDZfQFsm72agBy/C
NzEfDxQFwHwiGvfPOb5sWjBm6F/nNy4BjZIIlAcCEVm8x+lpQ2HnLNNc8jp+DfvnOo6snVC5Xxys
qMCfEfZdExFHWpB++ecD9HD7E7DmiV/11soxNl1oy1ACjnAOTGPInAxV5PXi9y+hGl6p8b2tbufD
VDiQ+vCJh4LrsKDgWS/+kOTQ6XD02LKdqx7eLg1rORr52MDqMuyNKeFO5CiA9Wmz9dh/K6ZHCP7n
G8AgaNePEohowoGlaopwD3BJ/ZCrzvWe2zBGfbt9gnRVebfULmI3Z95OMm8gL5czLZH3bJUYRV9a
aZADdWv10QtSzkhNE34NcnG7tP9Q0rIejyGMJcg7H8hZmvhfKovP2tSofUejqDqwLBlNsVIqMuD7
Tv6bS3zXbWRWmwLNwmuEzXp/1N3wWYAhYDs6apxlq8UkZr+xoCz0TaASOONA6fcZ/2DbuXc0vWkC
WgtoaBKL2b7+jTiGGAn8pXYSgKDx2Hzx/c4gIdJZH2PSKDFfVYf1g0Wgm5vY683xxI1nWZLYgtpr
DnFX64cMfAe3HsJfHtNMAmlqgkveGl7a3jgM1S7/65eLO8WtFrvhXIIS3FMt1aNkkWd80faC7Y2W
WXIn2YordlwL1b7slY1PzYqCwmes9SJh1TqJQNwLJND5v+J6OUM0/L1bPG2e1wc8M3ViLF3UMxU9
3A8vpIPBSZcpvbJsJtjKBJ07b4hI8qkecmZCRWSDqsHmG6YXAA9xiRx6WiIvE9eDW1E7tf87t1KO
pMUZndKBxGXa3AtjLzyTdWqFDhsVHwgM8AabURw0o6kQTJ5k/95BIZ0JM4hZcK9SyHwGnXrbPyvM
Clovh/gMcjHn6UxArq2u7F4rMOHVsQQkKom1Sv18JVA//fENhs+l95NmXiGyR3H+8VRsc4V3Kvvd
BAVcg+kZkCZZyFNCBAppW1gAaJBdc9oqxIQqFM/7Z4eQjU6EuevpPGqjRxQvqxQOpxOjpLpgZxZC
vbqVoZ2aDUFeP1fTvQpHN3Y9jl8/z3fAiwblyH9/ankFbOQsYQL19nbHsqpDUHRm4h6s1Wr837uN
VlNaSLbbBPTAy2wCbYTlkwYbN6owyIfa8M2xwktUzMaNSusPz8OpTOsF+j5zClnacAbKK56yaBVg
yRb3+k1LdNhQPtDDFX1f3PSx/SZ4EgQpo2opYxDxDNTXOm0LofB5ipq4D3+4xgf4KE5+vK9CtRJf
/Pdv/L18AZSJ4qMzyoxMgnIqqBn/Z4O/cZ4N5ulNVDNLOLObXEOP8Hbxe1bFnu0TZ1Mxwx5ZQvBD
b15hqlH5ql3TCPhzIjH94rVKDeUpYFcrAz4otHxskaROGynrXZybFtb+Ie0EILnZPcFRA4MCxC6S
ylw/TsDVPVHMtCMNr+1LBvflcy6na84Rc07ROm3Mv5ThsKa5Or5fEowxRD/HIor18uwZypFPOIVu
M0LgQu6PynZ58855UhbdfeZQ9lMRFeoJ9BmMqkKZQjP5ehxo7CI1DRRimzuH9yIYW2S+K1TjmcO3
+76jcE07V90Ez00BmJiQW8PBE4fdE3Oh2BuPIqH2wdxhiHrJJnFuxsNeGkn52tBrRqpYW972Akl1
7M06dEIqFXQzQEvMeEoOeBPCvI3lzx7n6Zkci9d/Yy9VoRRr+HofnA1aRY6qcrr1u9CD6pOasjL+
Q/yiiyWGpModWiexQ3de7H+wRQPed9qopOZMX3eM6Mtc7QeYUMr/ZB5e5YT7Qj0d9lhnNVUTy8m3
My6opL7zFTN4LqZDmF4vh6SQ/7/nfiziZT3gtLlSnmGg9I3nsGMRdh3BkYfMD1ajJbDoJO98Cwpd
2Qeeh/+6f+IbvAxuq58CYTwcd+m4tj0mDHkiQXypcq0hTdxv1s3UNYT3MZfhSHFocu1IaaJ7MxiV
+3WY2fcN+D73bOWTSc3pXYpGKuMQ5TnbuacmwibgIuo5dTq04ZPKisO9y62lyKg224GN7ffOchNy
cLz25J0lR3yRJPPS2xhUt426JnByj/Z03zZ++/Ydd2ucMbXRD75RUXKMgobhA9ZY1xyrKd6ujwk0
YXeVk/f1noWfqH9oTAaWRndT2WN5Si30G89YvSaweRJoxXXhEt56/iu5FejIJHpxfn0Bz1aoeH13
JHncyVnqfKl4Wz7lf+AzrdEmqqQQUEfj7yJb6YEDzEnO+KIyIkAOMbQXyNLpMngBFExGgZpok0zQ
ibWYk/mGn+HTik51fRkPbpw9SHBESMjpw6jwryL6yqNIKhC69udEOZZVAV7ijeVOpG3Du1fjNTPw
WDbTmjb1tvlRoKJ+Ta7ih+kafIJCDaPnC82wCgCVyc9E7IzwEXceNJG8/hMb4l4izd2CWsIQCtyT
GsbwcgRPvwCO6iWiNXR/Z3Kc8b+eESO0WcXHt/ZsEObA11n4YZhGyBQSA5Eu21MFVjfwE03Zr638
FcpIttFTBg7qT7GPH2yoxWXCuP8uNjZibKSN5hh4CX1BOSvRkCK+XyeWumKhnr5zsY5rW7xrdGsk
xMmzPe6pi8ZK00IDg0kiWRsEsIkvP9Vnsha4MppcxZTHiktV+DOdFdZVjEyB1wxcQkTYEBrbp5qr
PXk3o3knM56qEVQv/Jg+PorGdz6ngIB+9ch1jJfx1MnRacqt2LBO6DB3aXB9uABlF5NPSPUKnoZo
Er+8gQs7NiHeyZ1nEa1Pnl+SUx6B/v5zJJlNcpsGLDzP56JnUU35vFNstyJJDeg1irsGreLTFYKg
jaU/SDxKeqr5LrG7qYwwHlTFrpuEk4v9PFq+pr3FLLcJKfkOJiB/kIi8x2y2NmvbTQK/9FzwWWbz
AkfNqSahNSRJCETK3hjIg3r+MJG9GU2y6Vd8hQXl7xlYCS5HW1xaF1X9AzNSebh8IUV9keR8WEC1
2s0qJEiWNcp0wv2rmvSzSQ+A9HR2t33ygCc0XkaE0cFXUIO3sXY89YQo8PmeZaCC77nRfKX0cd9O
4aVRuz8Mz5jovAmD3ZzbcVso19CVIe/GYR3cac01b1ROswR2nrO90rWUpBxBZdgLRf8EruiQKds6
ouDahvfq9qKuX5+lQ1NJa6ucAgPBQruEDTEQcEhmbg4Fip6GWAzYhgtIhkXnHLXyDsukrxjP7io4
XCYgEnVcuf8jFut4GFZhz9uRY/UofbGjIjFBkjFuyoCKLXQCUbZXTf96NfWO4NhKU+pL2o2joyxr
w2xfIPyuBE35IJ+B95PTWQXeBVavdplGEICRdXt9LVH+DuJQWlZQF8IxkHm09CWEcWozmE7S5grD
A2J8vMnkWA5HJjEwismTYeXIxvcLxHY/GWgZ7tdA3UFvKMt74x5THU10M+6s5mSw21uGKBkbSgNS
W/uOaSkWB7lKP1teoRUlGBrik7Ihy17jdoeGRDS9GZs9e0+OX57RvgqoDfAUvXCUuC7n+6fgrHrf
/WJbvAiJmyaQBfdLjxJvsnfuFU4SBkk2biJo7qLNOnwZU2/+ErezdP67ivWGzYKsoVjlGC0mWLjV
MJmvJvmzRShMgL97trv3M2u/YPH+Ykp80pUSMjnK2WdVuUOnh+ZRFtvVfDdjZEppfgio0I5pHwOo
6jmzBMq6rGLURgz8aJ6lVRTfCpomJVeSrrJiErYk8KtqoDVe3Eul4O6yhv/o9D8rKgb8KnOIBQRD
tzPULY4G1kOFaIeX5PYwxv99XwCWk49GqE/0XoZgi9W804uK21YIRvQVKhKxL1HkjBnaL3EL0+8Q
CIrAF8JWMKArQ5D+meIkHI22DPw+0nvVb1n7BKTQneVxDZBNed+JfxzASv17LT3IkOeFEKz1OyQ2
sHOfvekuYZFROnLLd0OL+jzEKDcUdn+n+z0pALhgEoh7AeXMC+lzqkhzE+h+9kfF1y2ZX7zls5b+
3z4xxWGo01Uy+7+z3pXZ2OdRgh6DtnGFA3gNKvh4iOGXkX3IcyTf/5AckZYW34QZ3o59TWLb1uTZ
2hKhFEByIoW7vUDQGtUM02HXX70+7J9vVTozzIrQjY6Ca/XGzsYv/JGDcbqhRAeCeDM6KrBbrbBq
QL2L8hf+zOaSX1tpWvDW5k3q943GAu8beQWLk0CG3pw41UAvJoo+zO6Bv8VfEZYRM0wAtju/Y3is
OP0X9EwswrDGnutAhdRz4wsnrt91jS7yuSFOb2e6ivTzPn+B4WvcQGMkEeXb17kt4m0umc50rF3M
QfZ1Ksj+f5qCCA1Q3gVH3ewS3/o8eLI7ErXqYYcAZpalYlBXtWYT7F2tzkHw+89WuRhuCfOx3dZQ
FEmZKfBflXtZ+Yo5oqElGYr0j924QlxwFuz4mc6kMczpQm4tGEnJSKZ4LlEYo+Cwmq5gDbGcamgm
dQLXhY6imkRuGMdCABQkbkfeGSahc5i7fkntmwKNUdRTZaLc0yY00B9Od0VkLqu8PETz9Y/6koX0
Z+YF7AtNFXpLE0m7uvdCWtbGhmTxAluHbaVDbf6z4AefThk1A8XV+Ib0pl6HffATDaOurps4FkEG
oZoHnd6rwLbKHtwjkiB0uOWOSkyHNCCsnsPYca1PHhCDzIvhEn2MoYoHysH2RW8aN33aXQyk0Uxt
IwiJAoX6pdD7pZ2cdLYEuBieX/0BAbqlr1i1Ob+BwCFGZtjimWrLIWUAxJTWAICsR4S8eMpPrT2G
6VNK/A6eeqFOPXJygOHs04IOerZ76mZEGV6aBpPhRW6kj1bB2KcVEEmb9IqDpXXSm+i8tPI8yB13
I9ckKzgnv5kJJEEhdojy2kOtoMOv+fQg5P2tQk9sjC56fnjFdGBYHygA52qLOnWWJ5leBEfLSUMk
kbyWrGlxd6UkizFaChO6rKahSYQTVQUZk29U8VFaljjY0siFxQABYqTYvSQAYRYBVV9HlyIONx0x
aKaKJq+hCMBArui911FW4Eu1h+R7LBGfFJtkVX2vJk30FlaGAisFRb5ogK0BhkkQiXJNNJxmFwb0
KauS0DBoLR/bpsUwthqSjUNZ+a6oDjcvFW1of4xC3mIoE/WauCAlo8OIf6UnfhfWHdQB6/dPYNMi
jc4RFT/eRTlhCeFjyYRZWw21jijDTf3BbEwF8HSS29SXusYoUk7oYWpWojy3V6+eejvpQoLdFe5h
6SUDkOF5vRiZKjBVA5Jeaq/1evZlLj4ysE4O52RGChax+EZUO1bXK2FNv5/D3FTg4zVBofCqMcpq
+utvgNWT+oCRKaugdRKMaPCalJRGEI+n/h6SAd6EjsRqsr+Uh9nazgRUjp/NdAN+JrLMfLLjAiZS
8B4263h1CtUGBGsqXZ6g2WYAExuY5lUEjNE0yGxwbxDs1w+MO6P2PN0jSi24lypzVQpXLiz6EP4w
BSsj0XrhfjgyJnIRLRyNoyy2dMlbOON5A9ykGnDF+h5WxSQz0WbBrgMx0gJlciFJpcQouI2o24jw
GFldo//mZ5f37fkZIBNqW9vyMvMQRSdknIps1r28bfaRRaS3V9f3nlswmsr2EquFTEIzBKhl9Yz3
PWggBApg2k7FPzNYFyp7DUT4WeXEPVotN7bepEIetexoA3EJNxS6glZg+6n7GiTZk6ZQr0ybmRQv
t04Du8SEgPKFfXABLBnIZWLRtYMv017BnN2tjt5CzD6xeGMEO/SyoEQg3w826c4wInB+Ifdrb8CY
u2kNKoVb94eIbKzWppxpbw4/yK9Q8zLDdPzxM4ckiLXqayW+WPMqdi0qBtdrldQFGKEuGeFtygYQ
IhcObuywOJJvUjHs+FuEgS+5nFT8VM6hCaLxJ8DnGmvQ2Ek1+cR0x9nN62q6oxIuji9YBmSxsMfv
3DG09A127U3pZAKS7PoVLwkHxE+oVjGqz4C4WOCj+9EW0+OtTMriWMNQNYV+Iv9XleoRjEWZKaoR
1fVc2zxYAAsgN8XP+GegluoRQHwhpn1lozoRQbQ4Idcb56vhmhkDls2w3tPjH6GLP7efvV1HdJ8r
CVkRtnP0UXENlwVK+FZnw8HkYA79UpuUYJtj08tQpUXeO5/s8cdNvAIEfYcPquWf0y+0MXF6gr2D
SirwS7e25dw0U0IcfhHPAlP+8BZsr1qDEWidbfOktHpbBIH5f6P+rALv3M/y4er36UmGx/rK5vBu
ifj+OGoeFWQ/PMFH0ijhW3fV0Dz10RnkYxGxpBV27JXDZtuxopPPVXn6YlBwygqn9w3u9Sbt7LZs
fJl4YFdLaCgZJ2vvv3VyvEKarvoCi8fN8sQxjACtNiq1PR5jktBWjlxu9FR6sJqFQ1YOJlaE2cao
+khyc+w7SypeT0BXfuAUxH8hoa8c8hTT84UAWEW6HFnhQMk7QT3VZ81CbbIizui1JOy7Eyx4bZVZ
ghbG4Ta4ikTX6kTxhN4Sh9Yn/0F7negFSd+BBPVHU0kEuiHT6S8XRcWtXK/4SxFNh4mV/jmghxCy
GEThKyvlxQvhhu8zsggCuPlUNt9h/njXCmeYfAI/NQPe67yNSQ6VV0cwJZk8P/VH0rfbS97fR7S2
Vuc8qbe56qosjthvB+sHJao7Kypf6gLfL49M28dQOCfIy8/4C30B/iq5PNcSIWmHWycKp/QUlIZR
xExb2httzG4moV8hxfFNw+lqi7hUYgD1MqRp1BOiRn//kUALJqdSkdzevOYa8O6jyJmNWkB2hUgq
4p4VCiKuTwXBwxfnZ5RfB1sZnMhdqepG8KbIsQK3V/zJNnJT+AKtucCrxROazxJcXkZMgRX0E61y
IXu3P7zClAS0X4SwxiZ8u/p/eQRa0an/9pzDoTnWeQZyHk6TDwHMZflpXyXMLQs8kDX2JtkR1tPW
kdUdF4+Ioou/zthDXjOV5ykvEl18YtnG3Y0FP7qUE+9qZJiAL+Z1VrrffZv9k5v06zaUq2vbL3Ui
m5nZ2SeJE3gFnUVOHj2U+vs2UmGb5Gzvbnfn7LMvovpSdrsDnp21oH35ndNcvjryvq0Dc9qFJxqx
d3GVkCqsf+gzULnmKEK6YtsmwCUsT6ra3pAceEBXFzd5kzQ59rrrB4T4AZEI7V4iZpKgdUueRmV9
EznGeMrc9FATkYUqubyjg8y4B1zJ8qgRcx/dFYhUiKTAYiuhr8fR+wBylDP7lUSJwHFNgTg9GjyQ
naC5rCwi1TlF+3KeNIxYzZzGnOVWaSVpK8Je2xPvTyNjShbs/GA71VSbmangqomkwWx8Zgw8M6Bj
uew3x9pzZ20V8WatkME32s32cGfFDxtA6yImvGcseWCSwHGdQvjPku1+kRm5BzSBJcN6gX2CNQHA
Yj5YeTZvs4Itp7O3F/38HEhL4Ketrkx8YX1d029e5DvWAOFMDRcIQ2FjUWai91DmvvSsBRfS/zDN
E7VRdVhdzVU1N/TV2eB54QykxtUBa1hXcL3w+50ZUehvZs7BR5QnAwSgMKDW+6YdDey5uZHv3REH
e+h7hjqOBWkb5XZLaWVXWQlLbB1ygjZg8vihqd/DFn9x8jO7O7onIolHNjfiV3ujIeOrR1ZMM/WE
rpoBH1MIixdH6BFnwjiaaL0+LzX5YUJ47sS9g+bGTOJMn8cH1x8+Jly1oOCnJqNPdy16R+QfX5E5
dD4aOFwO1fHPSadmfzXnsZPEVqjiAh1oJtzPdweX0b9v88YoTyHztbRxB/gwEft2UiVTMYsIh5m+
f9LQSOexSRkkh1/srhzVN3mscXFQLj9dQJ5Q6UdEL2i7TNnwyvoxPzyx1Ju0XgbZMqPDRjoIX3RD
RwU0i8k+Q9GmQdEmfTuCvjsqlC11OcGIKgDZ6zBKuqLAKEKILelWDm42UUdvh1PwUPa/SIp/W1L1
RNTVT4kYIEaAxpVJ5Jb7d7AcVLgCWNXONkajN1Jdxte5NR2LhcN2hcWKUt6TzDVWbCCy4iwYKblv
ygHxvoXt/v09I/40xGuUQy+6LF7XL2aketNRaaJaOoKoSrQahPX/9walMEb0PH/PjDWMxN3rK5oY
qtD5PcGl19asBJ+bEO6XG0L3SCn6hiqIFUcgPAj0BLqdqutl2JtCUur56tVlLYBM1S4MjZ8OrhdU
hGLO5E/YIZdkw8cD1VordTgIR7sfmN/ma+QmXsiE0JV+Kh1QVHGfZh+ChHceYQdIrptmyq7EZZfu
O3Ig2m6C+Yr8sjYffkcRFpnUbcWBgBl4ydHk/aHNkqXXRM8NRTgnLFY431lp/2fCGeTbobKoUJND
1Np3SKEP75x5SsC80BWYS31OgcZ/grm6OT6xN+qA2CugcovZ2NGyG8zmO2IZUw4L0CHxTmTW8pbm
AQMNAG/5TgMkTJfXhJ6bz47CQ98rMGk5OBCPwOBXAi3DCV4KeGt8lenPm8noW7eVC7SOAeg48BMc
XjGnUnWyAPTmC2ZBS7V8kwIjEchZvbTCKK5S1LRvK/0dVAz0b63zBCMycUyB06aomeU38NBh+ndo
0JNYKG7ltPSyfzWsP/BP0qMvRzK2GXdbb/KUz0Z1Rcccd6mtZfR33vIwU9DNUgG4XsKKHTNXxISn
YNDb/1eT6ZcWUvRh4zZtcvlb4jRDsFexHUHGYt9DLkhBwuanszwpUi5gxl6DwbOxXOFWrslfCqfU
KRekZx8uSv8MwI/gaShbyQk2n+MKPAQ9ZvdDDZsqXXl8BdRVfBuu0kDKMuwwhBCiIXVqGCEB1HMc
TGJKrMKS5uaGdQePotzY84v1R/qQfL8NmBqIf8rZDGESByGhSUlmlWlNayQ2un1jTiaqvQEcKC8T
vCmyaDKvKnpEpGu650u8pyYPhl1VwG/9MRBSU1O+l3+Y+y2VO4D9pZjTN8k09jlNbPD5wAZQlXWv
tE4Vf27SF6kRoTF38q3HBg8TyMbVihJJNq6hQzKg1DIeT70Xwjw+R0UYk8fu25o8BgKPMmPKRVZr
1IGB4YYLEysJxGzRsPt+8yijUuRbl8TF/Kjh7W13z8or+bLz56TFU8CAcxmjleouiMtS6h1O2KAo
iVxyXqu0gNHMcX6DgN0E/9SZKnWX2miAsG4p53M/XJPU24Ty8dxX9oDr9yRrLyDbnZe7atTa+8BW
cSxKwpwA2DDlqsPbHEEnOBNJZHPrf4k5Xy/gDPby5L2r1eW4e3C/dro0PDsNJaqLJ8w+CsZKiEOI
vc6q7wJwYhEST+6c1q0DfR9z/Fc6kT78HnxXbBj8yTPlpMlkLOK97IW0/GR9mevFQ0FlaNsUqxH1
Vl/JqAZaznL/rHCNEF5Wnz/Eet3SiglPo+LqoIMTlwcOqD2B3RhgP1c8wkl5bQ/x2SimBYqG6Cs9
wtDJiW8x7zPjJpeIkeDf77jrkKY6I4kJhnoLj3Pa4jvO82ditGwslrSUtMXkw39FExWzKLNQHb9C
RDAW+DNWhOpaNi2ndsuoRu2FAk4uS28FdALigy/kmr5KUIi98n1iNxTopyDW/I+YvxUhMYWI6rsN
A9cBk5lIyTrlxKICPEtnQM7DUVAZvwhO3SahzUONoOPnmNZsbsFjckhc8deTEQymxSmLC5ImkeVj
ZLppQ1Ho1DRF9d5ydn9a+jpqT+EHthS5ATPFvLHVm04lCBAbpBfgIJqfU9j4ZxuXpP9jWF6M6YG9
Fvh5PMI3D9rphvAr/uqhcYV2QQqr/o5HnxL3kYHmZYUfe7Ryzi8gTGgG4A+usincwG7Qzb36UNIA
eGW+mvrmQFpDLcImj+dINPd/0TB3NUEEkfVqKpy+f/8penkG8vdJx/MaIYsBk3z3J3OLQ1EK9oNC
sLC4HUMxIUkYIUwBdB9TdELW5y7NcMcv0vVJZpuwZjoiMdVed1St49LMB3TNZpBNprJZP8kjSQuC
snc4Rav2rM5kSbGOG4Pjy+nW3bMY/E57JT6CPwuRZSrFtz9mOr3yFYRWQMLx/K2+KMdkk50jIdo8
qViLOUrNmQcD6wwb4X5VG24HFb/yjmSaERYeWJdOwPBLHZzaYLhqMrKgNvcIdm2lQtGf1MwRjot7
Z71gq4ZTxMahHB+4+Qr/3rWLjwTjodvkd+xDhcsWopny1gUtmWsTb4wXZxZ7pd51Iy8iBSCnn0nh
VWnx1y9oB9QBLjPvaybjmQCKiTQdWrjoLprv/DeecfRAqY+DLkx9D88KwdpTk+0p/EVyP41Dkw4i
1cCwNI3TqeeuQu58HuD8KM5DFV5UZ5N5Gg4Y5IxFIUbdzG6nPh6sooTPXXTd/8E50hf1OVsmhaBP
LR+LXGS1ugx3yHDFklQA4KaGTkoxpJuBKDc0nCfWpWakHtW7gtr26ijHDF6oBuLlDkFfGiXD35VH
GVtnoJzakUhAyXUzFrdvBmU0pQyI2aNv5jFW5WU4/Hce1bN/s6hgU/c+P3DGZeleTBAeJ9ckVP2y
IaLVuovj6Uo1ctBsG1vHlKaPKv7PSrZoRmQvVeyoXwA7lOisztr9aDfE8i4GQtkvYa00b2Htp8Sn
fLvnE8DeNcNyHCxI8pK3bf822XMrhRZG0P9q0QGWjNmSrhutS/46ScIfbSSeO24mWIfLueIQRiKl
MVAg0QsSWOgkPYExrScWFUASpmHtrAWMpfWqBXbtqDYajJ0srF7ZU9DX11xctv6neBAlY1G42qK+
8Ls4czqc5ZgwdUPGgf/6+PSEC6FVHXEiaIILeV3f5iY+i8Cf9YsVojzAFQ1BNMeaaIRdg8zYkCXA
O7IcVhLZhVCLvvjiusb2arSgkr/Kiid9OyKVSTVVlC0RmACqFbHE/kRyH9pxJlbPseef60TnmwRW
RioNd7+ke1ZMwr3H1Up3kcZCTlfZ52XUMVDIYG7zwwWSmkIDGiNx52AFmK8Fgh5Mm/1lUng/WzHe
hOPcI7Arb99hV2WeNW9zM0QI3Hu4NLtdY7TJSzId0MBS0Y6zDygB//WjxErVqZ1YRh1ocAOME4ol
jnDi66PsXazryoAwNKtrzoZmSA1EwLbgnMeckb1DWd88iifjQl7GYvX8dzGHHWMb87rjKHifds0E
9nbev8KjLPds/Mdep+NUXwXv0vRCs0CThZ5ozScHJ57iSkrJbiuAckhCDNWpadi8PaVb+Fm2hx5b
WkeDrtRKJsSMMR61qn62V1OgvNImI13e2jEmWBTMFHo5sfP/dm/tAO7kYCINQp6OApWnh7VDjdwP
3IJeMmiRpmWqIQbZZJ4Wv6k7oGVbb8m7JUEBjT5rzLIwkHcxwHDl//haInjWixnaoS+HetiL7l7s
7q4VfNbDyLUlAUy5WBGsgKRA1d/5TgLIN38mReMucBANQreUlrEIFY9Yjslk8aPJ5gzp5ZkQRFUe
nuFRlprR5xPsvwyYANrNJIgHN6k+H7fDfHinls6MV9C5QCbpBOG6T9qigfPWZj7eGm3Ak4rteNgx
0+Oa/N+MN5wecz6PKlb+2oAnk1i11WwacfjayrRXG8txxRGB39V7YYv91VKuBPFAFTQ2zzBaf2HH
htWjQcNjT7UdOyyXs850ZNNAYPjE/7YHpLBAjOsKOAgBlx0eOvJknGVPQ9IOSebJ4Mg0v2jW8PoA
4WfVGDlK1iSH/GBp63ztJZfM4fr7zHI9UJshqDrGebx5yA4S8K7aowToQ2ZFc8+ze2C98XfQAWkV
kTZ15yfiCCxHeTOAzg/LzgWW6XXIYS6jHln5n5cBibU07AAhR2vIHJsBzR1hE/7jJchJZ4MJO+BT
V36zMvIEeYA0wdokLCZak1hQok5gOh+ylsPl/zmYKvzeOzeVden81PF7Dlb7MtJEK6hhUuGVDOTX
nPnfF63T1os9LoD4xxuBIvAaqygkRW/lcpP6VJnMslY8S7IET+8z0im510r32OSn2SM97hAXjxzP
2cXtxe4FpwMW599hhveiWbSiOy1l9SmKYQREDyot55hdAICVAJbX8s+3NfCRiSfvpZklAsCuwMTb
6mE2YogeXjeGLNS/O9N3xNrcTs1hZJu3IHaunXss2B6ihTsqhFubLK6AAV+PPI5MKBacq/2WBDr3
7yWvptLYIrXZejdIV02gDdJn+DDyYeffbECI0iqS/RaNnpjk03e4ORD2yrWMg4SG0SItG+yW2PsU
SDgpVOKw0EEQbcVfl/D+0OyOU1S9EykF7Ambw0HejXHQ6fVHQnq0w028S9lYVfejFF2dY+l6wVpm
807MONNiwcDktWHK+SnyjKoKUsFuI2zpk1OmkyhIiaA33Nx7wc/XEzwkGrOiPw3tk/+/o+DMP9y+
V5lP7co9Gf3p9PZyqdj4iz+BBY6njhLfRpvxGD52i4LCxEnGVb1b8lLyg1YZQergzq2/LfY0AKut
8ing/x3Vaiue4rzZm9dE1buEkGzi9+hNXnZgZPlVLpqPANfuTNyTEBPeC3DcVY4JXmhzhFM7CDOs
MR1JshVTaUM4QwDItm02K0bRA7ZXqV8MMTIMI72GXkpBs5255BcSPNK1S+0l/ZETeI7S7zKCL/5o
+ZjNmeEuPKQpsZbwd2H/ryL9FG+FJedY8VejX9ZYS0JlraldB7/WsWcq44qV2kxENWHEu/IgASrp
HyM11qwVA16rMvGmQueuq27bllJhLfJTE3+9KWrWi2wONXawaMa5LuJvRGTTqSharm8GBDpm4aOU
/Rg0A5Pa02pl6gyFlwUlr/zUQEd2v0LRxige5ZSv1SDPoRacTDcl2xnqBa16B5dedF0jWffcoXOE
/fN6gnEjvjgd6S5QoOphKYOsANSyBiHUXWVdymj2PUQVeBWc6kjT3hMOEPgDFzFE1a5z0yG88ZVu
iFaGgpQxqJ2jVSoGwxZlFME7WehibzqxmzZzfWvgesawH3jMNydLmsrceCZdgcwE8kevpr4a9mXI
2CGVW9YA+r0fL6xlLLVepfCSCTxCcyt2ZTJSAt04l/cZ06iSRI0y9m3AJIIKiiqEWLgxvsxs8ijZ
ioZSa+FKoZuU5jmq+ZePzoiDsrtx5/IveXtMg/MJEIciFi6V/hvQpqXd9jMEdbWVD0TLcFtjA32e
9keFrY/IQLcCafMvp5jajl/YJjRz6QtGDIdVbNnLARDRP9egjPMdoUaTGG/bfjX7XqxtDh4vhWIJ
3X9akjVT7/gfnV15lF4dz5ZpsKnLG9NC38LP6kRhyEYW0lviUMkOoS49MxplkMmYEv39Kveetu5+
NfZPDTvnbb519XMekUSiCNUM4hNRhZjrJaCM3zlTGD3mM3WiNs6DdpIe20DJCgUlcnubPFUsUOvZ
AGZMEaB+pS3C44iIL5Z6ZD+FSZKvG/eHiyiZLhnRqQgnXpJhO8wRpa3A+fQYK+VGTXtj7DdHoWYJ
9rd1JJOv3CmVUkZ0/HS6sloNtWH+NOLdyKXwwepSbgbchVIpgoYs2/WqH+xsoGrq+FcpmcgpmPqf
1mNgpoNFHcaEQYNjk4wloLsqlrCaGBEXPDG9gIQRstkWcBr2PCGkbdJs44BOFIcaAhTBjkV9yhy7
/NBXRxECf1vA9vxgR5cj0V8SOsjHmLa5w8wAKovrup04A+y3pvQDHP+leM8qrIB9M3iWf2INQbLK
mz/uDssKfk77pe/MW7ZEeLxYKpnyqoXZdRhIcXa/lr7lndp/BDvg8Q99TFZXO8H7OjjkM1zm8veo
Dn8VI962/Dg8BVUSNDWQmJyfMeh83lBF43/FlFntqFCEww8UeDodKkMk5/HIhHPngUjhaabWJCMH
Ag9NZR3QUjtvTz1p6dVrijZ39XT7IvNdtF6mpScD0ynlDb7o9L/yCKYh4SSqVGD/GPDtVl8rLJW4
Q8QbHjYwxiMXX1Nqb5LEopdrscbCSKpHAgXWxoFn16hjCHkljfK9TgYGbdkrxsNoWFosGKFqsDhC
dyBorBlsSpF93q3czENip0QGJfhlmbrsR2ldJKMssz0Wle42KVfb77yKGid4pr11AGDvclWDlLxg
GToJqVa28Q88Apjm7TChjiwLurXnieyB+tcywoEREGqXw9kTBsP/w4Rrv0D9nWKobqCHHRvF5iyL
6wtJaIVqQJG9t72uC4l/9prbTPxDyYChzTgT9G+EyjD+vL9vYBub/DUy5Wse4+5FzKRqx7UWf0Bc
0E80A1xR7chnpcGJodk3MiKJK+1uBsOqdhTkueQbi37yGVQCk5tqYCgMY+v5WD0TQ+PUItF3s6Ur
3/H/Y4AeztT7lOmitKa44YG1/xNnIm0elxXfdinNYihpJF4fq+CkNPriyDwudSJcSz340EAxVZe+
Tip+tOqBvnJTubq63SGN0IJr1b1WsU0wJCPLYAw6UBErU7mpgig5Hqi9w+vN/oQCNwOJfJh7JbSk
e1y2bQHhLADEIwlUkMQD/EEjI2m7CBI6iT/a1Yk67lJ+A9NWJGpW2mUoyGox1k2jsXKWgAosUPoo
7uKzV4Qq+zoI3cA0RLgxZIIsMx67foy0MZGjHTCoLcdnzyyhnbaydtphS+Tu2f8Fe30/WW357JFf
VG8B3pk9whvZ416dbdUF1HbLbZwVODJCLFaNY7ku9TwFy460KlRzq2Rm01/FcRufQshjPJmSQyVQ
4U9WXDW/R5fjPxI68yqDKc2WKx/L6rc+H+Df5IHGlHbOYAGC7pLorRBeQqTUE48e0J/d2ocVrNso
2auoufuyTD/s5uA8q5firpyWP4TvpXzR5aXO/QJK6Qm3KtqgG9MAMpb34CfOTtypha9fhSNc+gfB
/46XVaPWTwlu/wljTdzbmUA9gcZLzUvaCbM6ZUEuSS0J6DqaANrdN3QA1dGzM26pmAsIlSjqixGI
TIB8iTLzt4h2Iy20zfh85KZ4KvL/kYwrVYkB8fV8vvT96QfzF4HXaHep6QuTw4QiY/tSL4OHfKOg
dFDv7t9VHTTrEiXVl6zZDteYRex6g8gUVCwUmF+fJGZYa/5T6LZBlN2rrWHtHoKD/KsJ6s1bhU4j
+Dlcst/h76V5tuF5wP5qr6sJT1FtVZwWI3XdsJse9Saln3U9awPqs0A/ODvpN8oBI3Mmid72PBRX
RQ5REI2/yAOAXXKDMiHhS55+P5a7tVf1RqjTa5PMxGpU0Aq5VpNg8zM3Du8qABx/3ZBHxl+bLqnK
Yj18+HSgfpdfqtNNNjrdajw/g2q9HCgVitxqYhj7Z/eYED/gf3F8PWJr7K+FMm6Ivvkv72WrmWtB
FGTX0+COXKhCxI3a/1e6scOaVB95otPRabPXvNVHvwXbsdhAmI4XL6Yacs5vcljfzHv6w1yhjIXQ
SkiMovWcpU+GDyWofqS8KAdvON+3/FdUfWx5R/DwucjmBfU2utkrQxJaNq/GpduBQRjIHlTZEUb1
2yHnQI/AIEg9xrzo+8juOoGksfbB5E6DsiqbQUEXyCChRNFBvPuQ+7vTR0r71yWs91FwEnwh1MeM
zXfcOK1ut35lYyJ1RbwoJ2qzuJfIkvf4frLoPSyHaeFVlCwfPD4yw5QlnXsqDuWjv3CxTGXU0nRc
VIASiEw5WetCte0JSxsf7tq+HyfctLXKaXLxadsXBuuXVzOUngHWr/3yTsmF+UvqJ6zWkp/XUTcY
l7CDuI8EidWcNjpx1ApOb2SE5gI4ITx2MyB5ORZApnhF+W/QPKjorCXN4p4NQ91x7PHA5MaSM/aE
E+cE4ULAIQO1qKc84CHZ33BmMgOzBk3g8oNYs4tVn2kt3Vx88N7gAHAjcv7DfkeA7jfpvoIGP7YM
NmfpQNhF+DAtljyt+jD2QJlEbq9M5i0WwkT07r9C7BU9I+bZv5/IZJkEVfaGC77yy3l0Mge7UbGg
796OLr2RLuvD67QXLKLAfK+yk9z4C+yZQnxI6YyYzIX6XDDLv2jIUGrgc/SHB6IIxpKgPicg37ag
5K+JJXWpPZ8T7Fv0VI0QX+smkuYpCTBL9IdcE+TXH1kvnurp527KW2xqYSq9sXg7J9zWEc7gvYua
CoWpdmE8mUbCDHCRsoOqWf8Khr4l1UxqigIqCd6/L/6UYlExLV3QlOuTDRQFtJ5lqv81Z7lX6Y9k
0OkR1CBOHxX83NDaMjbkQ4BKqbEtOmuzoy9u3fiXu2GGIlitLhH3MzAOvBBQneQaLNYIUmCp30nU
uwv2AuPGwQKuYc9uW19FbuqHJtvS2Nvu4nbcFzOb59KeVeZEDEUVCaC9IBBUX3amHzLfuAOh1IC/
9RoYM8kZthnogHB/C2g0vmAXvsdhwQFiDhvkeldiTn5ClTaHaQsPPFe+o4yMwf+Xi9ME3XX8NI+N
BGFZC+mjPKJnJg822mE9AmzxO1RUL0KhxS+cy06cVejv3rOsA6yncNzfEWKFxuXfLF6x+UVe1q7h
UAULhKs4IYed/RYNmJJzrkEzv+BZNSWCcV/lsdiJQHaKILOC1uWCbhCRdMcfeV7isWVxaK27I73e
2AfGKyKqlW/PWmCEKS8sBfdtPxx/nem/ISLrNiySKKopbGKVywF8tQsT/RpEWQdva3H2Uc8MvSKG
DyIPC5LrVoqWXD4BM6nca2q4xbNg5felvttVSM7u7NYin4Q5rhEAl3cAV2s7iLLUk9x9aLpPXb7T
WI54eRzS8PzIFFX5A4HhoHwbcmtOTpeyLvxQq28jhvwOnyLiVX+QaBBvFnI4aHTZo3RoUZFM7/qr
3eyMmsIWva+DbD3mULEqhIShL4j4MNQiksqAIas78MEbvNBT82/tc6IeretjCeY4KAIYjqVP7Gb7
r0LRylADlXtVcXpNPPDjdEalg+9aAWx+efKc66vW5StlInHo9a+vZVytBrudPXjOxn2AhbAAaS8/
B5w2d4h0EUiaROAAa6WDRA9PxEqjht8SqkQ3ZcuKUWahzAbAgbse8tBHg1G/dXE4ngSRkiOiNbGt
RXfjFRTKr769VeR88LktsLgh7mqZ3H1PpEcHrv7W3U5f28D2awhydq03PsA1Kust2ed98pqmXaIR
SZ5+nEYEzhcoMJTIOtvVbkUMKOEr/X6JvMH1wfjzyL6UP3KTdI9ax41s0icmaiET9K3CEU59rit2
kr82ZKi2ALegx/7I5Du9A16yg/fQZ+6c4xZN+VSj3UPY2FxLif/1W+oZKUYGh8sV1WXkPeS5E33b
/85JxmX5SZcaqJzM1PAv54ub5ueqiB2tXOar67nzrjI1mSXnZrfev4Rsl632oNRfUXaxAOz2tiQZ
Pm8le/Cn3IAWPPLKkxattH5VxEUQ+yoTjjo6vCW3z3rr4Y/+4Fj60sRihF0IEH3HFtqn8n8SMVEz
WfBKoqKveZ1wQYKPG7HcO52oNY/EXjpGZKKFW5pkqZrKQ8/5WhuVPRGdOG8mwsrUCIjENNtns+Mb
fFy1wNhSXzKImvu35i1vXPjGafCLgQcG/MBJKENIU612GmGCeA24RfK8Woz53AE7yMOwqsjUTjji
7Vkdq9GXTTVWQFP/eS7lgefKdiPqMGyGVSPeX+OBz70YkY8ra7ybpdKPkGsBZz1KKX6tjSRmV842
hhL0qJ+yY9VfC7sOHT6XndFlhI8fPyZVDSYkYLRJdgtxgOY6NV4n0AMfKI2QWoSRNU450Xx/eTNj
YNfWffkLQzY3plmI5uSTdnS2dQX+/iDzF9I+mB0v5mCZ19k5FoNYKY4kUuobLuZd5ZVA0S0PV5+d
0497uwGyDeYhBuWmvBmD1+k4WfWKSfSeVnIUBzTmqU8QdKxCf1FpBMb3rMwSic3a5KrhWhiD20Gq
MsSgqcM4FDXeiB1Min6lC1ESgMewhj1/4rYqmxag7QyAX84wZFLqkp4+lNgESgTGMTxTb/EsZbQE
HKbZHaAwaW6SuKyxo0hv7s+ML7HuCx44Q5W6QLJeVOkaIL43LvUoJLWPuG9ORszcIWt3vABFhEB5
RQBjksu1hSIo0K9RUGNR8gbfSilj0T4CQQqiOYN+iheDqrWtBD9fxnvR17//02ZMnqdY1qaESTPk
qRZlsztYSR65h2JSK8a/L/ty2/VAZmcUPgpRXRog5ikZmCTPQrO4ojqEBGHMNcV9PGi1Yv6enVeb
cAI4brM1Av8m+a2cq8OaTa8o9vrM4ZeitfaAqL2EH2noE48MJSFOH5UHbMiIxeirllOYBRAaNarP
K83YbEAmLxgensr8wVg3tm+aRFCvv1Qzmrv8sqIxq6bSA4vsr+/DPo8vNaWtKU6jTCKghUFFYf71
qntsU3NxcLPZ/c+RH8IJFnErudiuYD7vH48uW+GzIx9zh6FFz89Hx3rh2wc3tFWvIb+dZpoTtNTz
ZQFO0PCmKMncLYllXwevV/KhntV3uDuRR/5L94stzTFO6tHrLpKkx1gD67dmA3L+gPUl1p64xKLr
7LO84BYHTGawm2tdEEth9F8smk0QI9m4FPEQDZAazqNH8ZaUI7/p+TYJtMS6f2+zikvq8uCroNuo
R8zGnwkcGx+yhcpRmO9BaBkkISow9IlNpK+9Ag+TuV97jR8NImzkKXpg8HUSO+CxW9Kt78hksCMx
dfdnsMW8CotPsuTX1ZI+SjeKEvl+papWjc2DP1+MkrwUBrrB7LKLG9YKmBtuZTC6+XvOoaGhgWbz
V0UCkKqLCChfaNkFJbdHB5r3L0rdVBt98mwjBmMD17c+ScFtpwvflqWGkZapusT3L3TrD9cvXB/R
8LdxBhV5vPNUwYIFv/OvNUPdEfNfsUd1Lp94uC7pEM+eaAJSmtD9XuXimpkmdzXCcRlg3XlJdF23
6z97QcK5bglW1xxC9lmGPwn+TPNoscWgawANdmZSkaWrbBhowztURPPC16CDPBLklsCsaqXyV7yR
dz2RNWsUu4T2Qj/Zr1fwGQZKQFJk7aKB+2a/YpwlkZhxZ4BntgCZr/dvsFkIAos5p4WYh8I6t63g
NqcVv81qprchTAhulcBlOeO9bYH2f3qbPs6547RsOBg9WSjGykboqDYxQrQn4l1YZ4WBZcmv33xj
uAPyL15ftqVVy/6W+NMo9UGpeeCdHwo2vh5hFQQFW0ohCUSupjNLZGn9cceO/tc2fdgv/3vm9XtN
8V2W5iQXASwS/GImsTTRwlHqTJQPZiWBazSqnLf0AO7n1APq1KpCyKgDJHGn7JeaCPxdm8kCvBMX
k/8p6CfWGUMUUB9k/hcC+0aYIRQffkx/7IWx/4zlnEY1cvc/MexU8edGfSTv+qbCUNSwZw8B3L1z
ELtyk8kUFpG2hWzCxSaZo4Rbf4soHl5bT3epUTn0v8s+5+yUMV7VRqpFOzWp6g0b5A1gIFkmmB2R
XmzexTX2pwIKyQQ+oel3Uvx/O5nHf5u3Mqkzm+UsKaoZNssNGoaa6CwQ8Rd342F6Wf3FdtDteHqI
xCPj2fOxzqS84u3XrQRgtVDY0oXQRlfhNC7ej2GuQy4jyXh3QFUwzSzAT/Ctf5SJje3EqhwrnHeS
nIU/CVFrOOeaGW1fi5QINy4PVGJSEULGbBosu8bc2/dcFy6wiB+r4fn6RHNabW8HAYkxW/F4tShP
QT805pQhckwDXmS37Hz1zPYUOUzabHiVpjcl9feYUaz4Tieej7Gz5DADLslc9Avlt441VQMp5+v/
dblpXqp9qLIFfSDbZiZHemGDN8WIxIXGGCDN3t0F2KitKDBm4RWbmjatMj6MtCHbkuLRpbDXgmzq
FiwzEDs9w33iPzIdw56yW/iGN3O7pBCMkQWnMSYGhqZgHFBjOUgEh+IEBhLGC/so+adX+a+VKH/i
nDQ0A68Urkk/mE9hsMzX8Kn5HGKWJtNbBXMVBLlxSWKIdsb3Cij4InAlmyMHsMy+447j3lNL+RPd
AXOBQMdfe5iBJt7N3IrGUXSYQH/mUbDGFgyQNlaJEclcvsxZOZSFhkt4FC2k5UzSKARpqV8OX5Mw
8/JrzLScFkAJ+ddPyKfJKLLYCyPaa4nL/gqfCOEjl+dJ0e5WWHT4uT0KSNImiu7Rv0v6KlYKXXgh
iSsAKYK4L+AsGtrCwKuA0OrEGzIdPXxDnx2QARw+O2DLvbHKiUPr1tEIUGJ6Gx5QIL1iy1Yh9RFa
RhWny7iDlPfoi+ajBkSpLmutSfN1wkCjVzL8uPZXcxdHY69qfYR5JOZafo6y1NG4hu+SEDqu49JO
HdhVZhms3t6eaMD8xoqIv9ktrlaTt3IuCKG6lKcbjm+oQUf98kikyb40JDRB3EXVowqZAi6mp80u
LY+qKHw5hTeNVaPwxdkDIK1Fggb26FRRo6IF0mXSTH4e05fEvJX+KuD65nzdPnwEaFsR0lflDHgO
IYTxBItv5KncwCtezCDb5EWQAy8bsSUxZqFb8kqu81GJY9dE3ywzJ+7CSNz4wBsIgJsy1M7501+I
q4xz96yuNZTAzvY3nFIh6mtn7pGNzXyJ0Zb9poI0wENHKHa99P2YDq8n5erPWeq8O6VPNXza32Jn
WuovTn41/s84h/wRG2PSCcfdfrGYXWb4QTeb0+3oh+yCOCnEjB3XC8QAYZY+Nt1lpGvy//kipV26
OzYaU0MsNXc2SIKnQNCIAFJ1b4FN2X91Id0/Wk9vX/0xRBg3in+ThLTgNOYFiA9F7/XhAGuUonma
/oRbsKj9JWICbCu0Ky7kaN67rRO+axmCjOebjeE883q6345eAmwJsJwHFLXyJk1s34SOoDdTzaAF
pP3gJAc09+GRZx4whmYBwxXQl8rTAgL9y+7zGYic19PPNm7IBAF/Ac4foxbJbmqc+eLumIBGGK4Q
Z4TTvAODDkzD89TrhqMLlcJn8kkbsclI94CKJt0kYVt0SuNe9waJxH5MJNUjIowgrjw/o5pvDg5b
I7nmwgdhbUPe2O6MMyPwrXATINkCtUguZlKeWkN8X/mhQLx5gccTd9YbHW3z825vPFvuYOgxKb2T
jdriHypij0aC2rvcRFiEH9h4Y9CHsOEh6uGb0sGyj7psIymHF5o5+alddsDAHsC4Mpt2gzItZwV0
NOkzJ+wXvzX0R+mTAHWR6Tzuouml3y1JdtFzQ9vzTRKTcjI9RgLcPlmtG/aolGTBY0ez4nwFO8Ma
DEFyNelbugcJpTXUi/dKdC1QS/MAic/yoeFLlSzHxQTxs35cbcFUZQcH/n+BtCvJLjEncIgbader
76TmYLSRvvrgOTqvSO2cRa0IdDdjgEzkMMA/sj5NrNCicUdsPyRC98JRNcqT7lIpZfREUNBrPupK
n0CkyGygnzRp0arpKHwHu7mlYaxy/exOvG3Du+fwEzlFY5fqmT4EELsiJ1itt8y1KnMscjjZAfG1
HNSKeXTWhfgmkT6dSZuHtBY7uo0tcpqu6IjtDGWMpSRBJDkbAcY8yYtAVYA66qI89bQsWIF31XAP
SQoF6bAS1FzcQG3ow/kOg04JqKwrNx7PW0Y5+91P/4itPAsRJzx1EjRNGTHToNLBzKJ6a0NmmFsy
mhqeo4spWv9ZFiEp99StZ7SNjTSSJh6SkiQ6RLnfJ9IVvy9vgdSPTUWUMqSv4VUoPAumXvRiQy4Q
KX0IQ81LnPbLczHsHl9/frHl/Sqn/HJ9msvInJkTSt7X3kD7QbqO94pRxbEfWV5KEcHHp7oU/NZ8
eydafLQ2TVNqUPmxbQP4nG3l+0pUhQqJSNqASXbH55RDYhkZi6EybwTt5SJanNJTe71941UQAxGn
IRLQgevl2jKQT6dTpucz4Tln56y35YaQgaP1L+6Hq1FG/ycbf4lDWzII93uDLPd+SS7TE1a3Kk1Q
KANYfx0qFQZNUXFp+BN+Q6aYeIvEPTY0SVIOp1DpNxb2M/j4hk4kCGKFPEVOODjPQtnw203ltA4s
aasIrMVGvHedfQosK+b5rXeU6jeDunWxvhk5Rx9X8a5siSQSUZN8a7YW1Qde5OXDR61GGRmMhm8C
Xkr9OiE/ol18vwiiyy75Hhzbs8QSobhhx+EpYIMiKfELceC57T55LF5uYNwrM3y0fK5pRmrKlWkG
YAnc/34TofOT34CQgz4Cf0Z+6HB6+KQzUR+dPvlxa10eLqddorbQext6yRKJF4Geipp7KiijVu/4
2C2b5b8cklOOuX30dNlg/LEl32VHdOS4PfIhKyMNjn0XgB9X6RDx8q68cL6OVvKcdEGi8kCRm583
/nS9KvMzajKvR/beFVZmtvRlt12On7w3MCasdfAwpnCnN0Cm5kbGY3LAaI0/2cJBUpTdQouQjAEM
LBrFMM7kXtI9JzvWPst2JYBkb4kbPSxydEKQxpOJJ9ToaIzVfhGE0Ne35st24YNc+66XbMbqTSwu
fU+t5tNLI0S6zl6FVWVoUwSOAcZ6iWfMHVzx3fCrCF3hPKmw+5gEDpaI7RJiR4+/kCDAJ1pFHug8
/mf/EfphbReBCHvETCZ69baWIe1tQheWEK31uIZ8oJYBGvp7sWhx3Q2AcOjLHgiiti+ktFypYk+/
Vz4JRcbY9Ff8lh/B6mZIFT7d3bi7UciM1bic8LKxy9NmRu65OOhzD0qbe1/0Gii6TMnhn69W3B8T
PKlotYuE7BgAeIi70O3f4MQNPRaJaQtM9NGX8Wf8Ad47UcMv3Z4eQ3mHlmmd68gAY0Nvlr85X3/R
s0hWx1VI4ND1K2Dk2uDYzKk59I9CWZyCz3frJ0bHne+/bCMnYveVg21Nvt5posHxD1UsqZehOU8t
9pOU3JdqjGcSwJP7j0TzIPTwE2ep11D4c5l7KlCHlJ4GLGJNow75f4yGf2CfRjSNXEkpoegqNCd+
6ZKY0dsVTyNGN+XI1VijNb0mpYoBusfPjolpb0d/StFvRP6UWS4TH6gM5SyYRDLT1xfSr88y9hhK
BIcuGO9DaCC/UY9OynNLIdMWW2TxGOapMlCSDkEBqEZt6EGCTQVYUbdrdDxj1HEefKDv/WYF0gTq
lsivhuhLA6wnSAbyTQJ6nEaPBXw25RHzA9EFlkjTB8txEAjgPKX1zWPe7pQ0GAIPbQSdhMQsJFZl
1ztbIX15DelY0oF9Gn09wr5paborl/RM56MQiquo2x4mlqFCBUQBwUHX3B3dLTyKeL1aNjv+ck+v
eQkHxwg9J+tgOPdsOFfEkqgGeF29XPEA+uka80/slHrA7U3SW0dDTXTAAh2gdlR8jo6ikkTSYs4q
nI6hw1VsTWLAn+JJWDqSUuikXV6cJkuN0puYhX+9/761muLsmyjXM9xdDB8AeQFNfJMcrZOIV0CI
jV+DAppQS1z3DqnbixitUgZxlAxOSYEyvFPqTMsc8M5KWXrsoqBcFlptYV+aHVbTJItvpOGXKb81
GPYm+MtNNJYD5Pl5MPuyrcdtxLl/wwUqFgGHxsGJrIINckYsfNXigHfSFT/nk/mhm8V639L3ID2b
LdqVslGAHhZLmx9RGOEQawXJzYDCrrm45s2z6qgVPDpBaZ2evGWXAfyHqIRE4n8bP+fzncdpO8V2
xSbpUlNWge1rXbw/9Y3jYYdKoNc+jdu2ZLWvZbiqPCqlMh/OhrCZyT6sV8OoOhukHRNVnjps9Qo0
4bpPZj51r/lLs14LQ+5piYygIB7p0LEZtnnaHJ4Y7HdTXzFKwO6lyVtndbQyae/wmuKMvqsqiIGU
PvWWgpXbdXKDtpE6CmkQELaqt9Xpk2RUlIb+S4689Q15k6UGYc7x5tJAvzkMLIglR8t0ViMHXIS5
F//3oOKS/UhRdC/MV55wqr40KYT7yEvmmIvstKLInr481SOpyf747uPNVVNxmu91ZjlrC2lUBzmM
Df5Mdj1XWACCyznkgTsYpQDW/rXvbhMYNdoNUeomk9u2Wcv9eumrTudjba4kDgCUPVPbs87TDqjd
CUQO21x5u1Ex0PxeZWxoM4iveW0ReL+DoYN2koi2wDMnjaTtmtRYo2TJ9IkvToVWGSEZ3MVBiilt
hQxk+XFMXbOrAxQXTuZ11RcXSWrgQt+fLySpJHoA4HcMSNQhXGo3lS3nEqPIbVGy/tgzNNkKG7Zf
xH2XAZ/qcGfQ+1t04DMoxUWYYWgdIpTMoQj0afx2M3AWYaE/dPv5zmV/oYuoNBwvcAEegQpkA9d9
bACKE8MnR9108ePF0lyaWiAptYvwZA40y2fFDAnMZnSTJ7Zpwza0+fHdn/bjv7D6OJN+qbajCv37
akTA3MUnMTyrK5NcczH4+8rBSkKsyLzQHy2bCe65ZwV5YlA17aNQprfYQNPiS8vMLaP4X8XOk4BM
tWrqRVPmRQsX7dLtYcAe5s/urdW6YANervcR3DKBT41NocSuTucNG4BaHKQv2XH1M8bgF0/fRGen
lAGixaVvIq7gnCEoQwTKFHBcweXVqRL49ftlZrJiCSHo/mVx/otA3YCWNReJGTV+/gxJ3OScX7YJ
J7dZgcv1J6d0PSlkl6VRWV9lDpVRsGOLB8I2C5Sg96E0v6KjOEESLCtEY4TLuIWS/i5p7bv3ZkIF
A5Z8AWJjp+4Gd4CaT75lwrj0hHRicuHhsFvjTh0WMAPyCGbnpTdWYLTQNZWBqxqBkQXGlWC0xHwb
GdFP/HbCoRV8eQ0WK6s6cuLU6N3Tw4CTGKYzsQXigVMbBxG7qlHDSfiUqxpmiT9HOTYVziguUf3I
qQnIFgQpOWyQ6dZDC/+v9qTVZSxtp9useXIou6NA0j/3zyaIZpmzkkbWFKawP3RM23Qmg0xj2ljd
iPu70VqDRTxcwkh3z//wIV6FYbd2tLTlqMsPek4dK8qOnaP3NgkfesfSdDFevEdSSUY/8CLGG4Z8
cZ44UuUqH0IOuuEdeOY37vek4MJ0qqsLm5Q5L8jiVyveA+hhgMzzQLPtW1+4kicNe4c27DMoA3z2
xzTJZl5GVt8KlkqH2tmhW6aiS7Ys4f1Pnt4sEvds8La26njqCUVAk+ySd8ztrvKPFjRoWFA9rTCe
vERUR1ibDnO/53rrCDKqxwNTaFl+Vy7xnapN5pH4Kqs+eO9alOFjXD6WlkBXp2huF4VFN31+Mcxs
q4YfsaCzaxPdR+Cp5Rg2oyQRNim/vteOTQAuMyAWYm16PbS0THjBkeB+W7DI1yrWYQnxE+WeCnOK
267whDwmxKmitWMm1e4vJg4SnrNQJjVr++8vTKKEPgC/FfWHZCPg/MGTlQe4x55J+3TJirGEsgzQ
3EGXIOxfv8b+jfMmLwJLoC7k/8eFNUyuGwzGZrfXNJIt/HOgBVPrKkRRXYjeEdAtq4axBVl+8jop
Und0qDzty+/tnr9ZT5X+ZKgDoqXWtxYCLm4RvJRxVhYvKTjfA9aCovAbeEPst+pjhoCnRyk5ZUA8
vq1bk1Sywbbf8maym5CPCt4VeXwFW7Da9ngBiU+ag2pSgh/XAhMH8bSNEDZSd6g4i8p/jGm3YOdU
fxnuuraRqYHmZ0iDrBcQoD9oVxC1Ba0wMi3uE98s5NmPLFAK6Ver7hnVg7MoU/lb6D45UxVN5raL
YW/N3GINH7XuzJ7syrvaC/YEYT3z+myzbdPLSHEdASkmvsTY4+9xmdNUA1RaUDPf3sVWwCuJDGPQ
TbsMRYQrZlNlNyFYdc+2WG32TxQEwlyRwcK7NyW6CoZGJtC2l2AC0sZUqiZ7XEAeXaW7xR4rtgfO
XXpkV9xlNG7tM5wFlIZbk7o2DFwEHl0NihNTpRfX9syHwqUs77fqxbkDLWJME9qNGRBjWyodia3Z
HWEMEGeA1mV9lb7TTlrGp+6mNzfvH/6jTk1IMWuCjdSXqYRSly7lZvnQTq3wEGA0Et2PnHk/LuiZ
9Bvh0ocGV1yBSaYtmXkIPhq35oJNuPi/n2Mj2lXro2/eDHXBaQUDVxgfbTWX2tWLm481aqTMyXR5
UxzQFOOnaMxljXxR7FyZs+GPcoc0m/xrSUUlQURukZVe8OYXJVi5Bc6vZXr4F6K2iGYQM63K8JT8
Wcy5+pgkd8T+4jkNguXzsF+a6xqM/tN/qUYyNhHSqzsUSSxga2QvwZb1KkuoKDA4Iw5NDHS9F8wa
hI3c/bnSwYy8T+GtpQADFt0nGkVT9q9wPtRKJ9/JCxgMj5Svsks/gZn10lPjQIJuLvmteM3TmQAj
NrpFb12Ub1wt8GGaECD7ORYHZ7ET7zvMF4UGF0qypBU3e3QgbEoHqitRUpM/sgQtx2EFvta2ac/K
kx9xPQe6uKz4vP9JR8s6Th75541ZU37h8xLAu+eAVoJWncF2zXo6Su1VdRel2d2SJPyTMU1H/tQL
vqLEgMcEp/xWXWlu2DUxAn0poapsuhXhQj41VV3nOXzRMCFbw/K9cgC51tuBoUwDW1HHOUWggZrf
ZTaoiQs5tpgcCC1PtSNBv5/YoT2mElN3fSLTosyQqvRSzVdNSHhUs+A4XvJshAEcmWEpfn6vxuXT
tmMIC8gQ85Cmz1rIIZ8vxcRl/X48CZdjwE6H0Cv88bB+CQ93fDjjz/Mlk9yBvb5ZgCO227X08ZWx
JZmGO3+ZSneDPHcIcV4jZNWY3iOXiXNbeNsJaj+zQjQ6lvz53exi5VQFhIjjPgzLfArm2g8Te2VU
WHrAxcFIqrW1gFpRHgIZsgjDyUfBbgd9bEDnnerx2IKPMyqR6/kw3Qef2drrXE1NXU/bQ5x3MzXX
wAiehiaF4WyVv4BEaxXwmmp52/9z8Bj8ao/rfCIAsMaIRvll4v5TqHzkrZIWq2/MkjyILFlQM2MU
spzNp8YbztjAb/lhHf8PhCrO5iyGo49l05HUiANMf6oDgkzkERJ18H7Je4++uQfRMl4hVve9XO5Z
3XbN1KP+Zh5pgENkUj2VazdetoPbVrIhKnnhkvypmcfpN7lOkrGYXy9okDzj8Z5CYhmMbfzQM1+w
PoGdMa+AofO8dw1JrmDK9JPWCXANpOvCG2vm8y3TYRVZROr1XBy8tDdn8h+s1ayuoowmtRjMd0fm
HpuTJuw4+HQWQElhV9c3+Fj0KMhGViJny6u2nBeav0C2E5QHaNxLYbMLfnjzY/JUWdKTXO4HzvbI
bnHLJvUe6WDkNfOZhozbGQrqs4WXB+hrQix7Jk0RumTU4jaEtYwBldNTGr0wYsF/jJl9GKXFLDlP
bu58EUAzyJSciUrVzQ6h0Zegr5mD2fsUPbJuRGFJlbEJ2fHl8QtWMLwfsMSyAQ04yedKHNEVUx+M
oQARN3SAEtxow4vWbEfWIGzOdj7x9dBpMm3p4aVdCx76hB8yS5O+APWXi0vhYxutB/lrhtsKfEWM
FPctU/GM7xYplxDYIMjutVDumHsVJRsUnfr8gZ6fH0jX6YpsfDUj6Q9kWecWEQGYGfeemPP1rHeA
E5Kcb9FJxmISG0A/+4bnuj+AOTi//5ciOYIQcfXqYk0dWHcm6lWIRNLaGvDDVIcnGz3U57cMtZeN
exfVZAsecWbdC/vGVSo9cYJgClpeh0iGAlh+sBeSA08s3rNsWW9SSreTdFX3WEv/d/0Mp8VbHmM4
yXY2zdq8CoY7ujkPhKp9YAaPEmRbFZdTxvVQ+/XJkqepYDx6EhJ3StSRs6rgdGwYgzOGZGYXV39V
16PSZia0/WOS3FPJRYPfGJrJtKVPhnwkC2dzn/dOQr1uN/abYPxEEiiRKBBBGrIf9KaDXX+H26m6
axqhp+jnSDX75AIh2eAyC/qb0FamlmUtzu7IjZw8+gFKNhEPe0uAUSJBDBUgKlzH0K5i6W1pt+f0
KpDzX8q53Qbfqo5RthPe26p3sbZnBoOm+97VVfptFY0ylf/BePaBZY3XOIUrLBgxv5MNCnFj+QH4
4/70palbQv9OoHvI6GNfWGdnHhLKVkUHGbmZkd/AfkkqvpvgkpuyxrlZIHmPQUSAOk5ONIp1FDQR
K7WLdldltKmUQkNUCirpgVp70lnSOh+2lEOaxRfWNNHMvMulr4Kmf86fc+DdRCoNOSXEN0YXRXf9
HctO3Re+L++5/46UvTxnRCsEsmzVkX87Y0wrYRN0rH08gkZdP9a1/UodXmluvcxcNiLO9PEszfcP
mU7GI1+g84JJBD34GtvoWcIZHJ25rNf0MelbTKCZsE0ha8KGZrmefs6SJHejx58vHWIHnGDdkkWA
Y2RW7rzc9vvmQnEhdW8SeSOYDx/hquDReEoViTccSgpBZandTQCRg7vJIUlKKBwJgP0bgEZbSp4M
ukuSLC7IYLSBIsgtsk5dH+IrpgE9F3jUL36FwuCFDNWTrbdq89O7Nts87qaNY8mmlDH1ocqZTSP8
haJIJbDrBQNeSCndgNz6H2FYPXLnmJzI+/JjnVLtLQavMpFYvocHlFGI+0KNj3IuyPBlKN3eQ4U3
zjJhMEgNsJhmNUvXcSMbTfKbawG8GgW6tLO0sHWRgCCy+ijNUL7p6g6BiWLdPL+7Dob6i6fxZVQ+
Lu+jGfkpRd0NpKD7zf3tbHmJtKNPR/NJ1jQInAdcqEIVIoaF7c84v+jyDPsZc3hIs8+tMARoI2y7
7ApwyqkjK03zI10hJS4eCsJEH9ObFs1so2abGdHH0epCEhe4E2ksbvHpc44pa2w35rXl5UQv347y
uteVi9XlsHuTUnba7RNCpQy9hZP24LkY61+kleM7ZBBtiqFF8Qio4l4VUihIe1DGfRpjew6Z6u+r
qEXNTubacjC3tkD+QFA7Kj4xO5eJeGzsJ+XZ5s89FA1hBBujR3k4J1iLKS3D4rwV/OzzVrpEsPVi
cY1dZXilML20UAYuZgahaBQHyT86vu4P+c7lM7kIgfaV6bX9JTnnzysdItjH5PetjTTRTs+Ue/tP
BJ9YfP4zDptiW49Bk/p1jI3QPhg3WQsxA82+Nzn2Cm0qQJDdEqPtJXLQZSlgqvJlmwuC58CtuN7I
Dol69W+Pp7Zp1lhaLWeNSaYbmFSkfXeZ6uR/I4A1jQKUFcw3Pmsiqvb/Ut5Cha/gqdjd9rpnW/Ix
mVVdnrbkpJ6Gt8weeBnI6RcxxpQfh2Mxva2+GIeNHoPhJt8oG8s28TadUsuPALI5FEgQWLRRjtRK
sJJ9R6k2HwxCtmINm1mPr8VEs7TwbGtG2qx8Ff9v2OMVF9MloBjWG417JAJ2mklVKEXEBBb4mwso
SNVTVOwJ5FCDIWt5flo4IZ6e9UFacxgRgDtBlaRwVZlTOQpVxcz+sS6pr7tpFW+mHg81N8YASD6S
hNLCMH8EzjO/X/dYuEkcGjypwwJvJrt/4md4R4SvzI25mAerE7vRv9o1mk5uZCVckF+UrfhhyUkl
+RfwbPnJ0izb8VO8BQ3oSRVaVcvBOKKBnBrYqe8V8npxghFKGtu4xDdRl0ea1/EbX0SdIMnydzB+
PmEm6fv5qiOGqf1L8+HsAreMYXoDd4HdYb4cQrSCXCvrtTbfjQby5jDIPbuVVZ2lSUfo1lZf27NU
0xodkOIeM/iuAk67FhmjdLaVvnAqHhB08f2JXxZK/YMeMYrDmSrYhI2/Ldxc/7Be2TZtekoN6uf4
Q1xKYAO/OLnzMBBUnnf+WltH57T1taYaLrkP6Hpqz6QU6a39X2fHpUEcBeW2Qe6iZjvCGDO/przi
IW96fotYnF5GH2YoV5AFf5OmoewfkYy0ptiIaxxU7Zxb+nDMDAyU03HWonJAyg2qmVsqIrUpXHIM
QxU9qfXtnEbZ1yvOUfmI5cjJe4BlPougOGtUE8+6XWct3Mkx73qWLVT5S/C+4psDjOWgGAS1epd5
TAfsSdXtnnJqh+eoQcNOfFogWdiGHQaX39zBJysz0lLZxZSxkf+DhFylmm9L9CSHCUVyucxYOwhA
lx/+JSwuc8AxwHKGNvnVqQyj3k67guoWPYQjBN7cBoi8hnhjRc8dLIm7n7/VZD9aco/XVe6hIgMH
6pPgDT0qjXNpxaaJewbNhIbB1CvEd0jaZ88gpkJZbu7RoeKmDwtt/W1Hhdm58u+rxD96CqxhFo6q
8NVfK6uRElmT2rtOAxyygnqG2rpA06Rzu56bAhfobHUwkkX5tcVOsFVbqe3AiAMPXaSB2LQ3s/UB
c/gErHzMwNNZeRcni92jQ4DXCEOcwLGPg66yhWi+xZLQ+/+4D3rXFkBSw5DmvtSwp5ertz9wHNld
KaP2d4GStoygF+grtKWZDRBfUmyw7E0bt+89g+PRQjR6e/AR4G0ZrqCbiI2djk/UqP0K2xFKae+T
gHDLCYSw4eJEZpttDZZqmtVwHa/ZxV0Ab9HXBApAAtoqesbsj6uVLLbaeMO0cGsEFN5KvqDHnXxd
DtYrTmHa/B6ZA9Y0er9awqDyTi2PZHyowt/2ceKVsYaz2i+Sprdim4Y/MHg3T6h25oBI3cX3WcgH
Lqi78PZ3Y6CBk74PU36vBheVVTIhU/AsKaGlL7n2vix189ichIueCMIORNQEySQOrQM3o8q51Qmy
ezK0owbV0xhcujfheLPCx/0FxkmkDQglnhGyE/D/+QtWqTIq8IYcHTxrU+vtssze8b28DFYYueDn
8GAYROJgoeMxs/vmX9g7IosHQEL6an8bC3Shzr3R7jhBo8m2ex1ufK71GtL0M1QvyKZLF7YsVjXE
CzYxzIiqG6HDXLriaXplUphPYKGTe9tmCLTwLz9D4Hdd13DHn65K346lJvOiHDFE0yigHKOpbeUU
eIFqkt9dgtqHyiFNvxF1KvvFdgNWSVLcBiyg7iljS/rZUdW+6cHOww/Z51hd0CdR0DyG3w08FdrF
eToji5gnvob1ESxUms6fQ56vdiktU7zIajwuwDQ0EJYyHEOArjvAGBFWfN3CVNRjhjxA69mZpjfa
Up49lLZYNbYRgZSaURYTPbQvGW4lND6M6nGs+/oPWDYlNvD2iBlCt/Hnz7Fqfyi4YIBPWfzg+3QU
Fq/sX1rPQMhpjLoNDayrY6HzBX2pzyI0Co+5OuJRiJOskDKxEZSsTfwS8B067ar1TWWFmnbsup0k
LajkgDm3lJOw7PtCEW8Pm6PrbBhkXFX+62dWEuxTiEQ1joY59Kt3wWYOOQy2PcD5v3BW4Q7L7Bw8
6v5GIaTIjnEb0fzwiITmZGom5tftR7gunE8hZB8KfwqNGbWTfwIfAb1zR6z6/lNvMhyzHUA3n/fJ
F8XBllpHBr/4GGTStV9SnKcPDNGwmuVKeempNToQziHt8+gVZcsSImw91a5tKyiQf3K3oPvlbh3a
5gOhWGADn03o08+zjarkCIzyiLOysCkM/HB9XAG9evLgvBIAa2XzNPaCA6XyCeeXMZmwBCdUHL/I
JCbpLvqtOrz9Xe+ta+EIIu1RixNquztG3a04nXw5avM1HcaQJtRHkKaquo4PBuaX1twR+57APjlX
alMM5/MYgQ2ZQf97Q28WjKbe+lvIJ5vYF9Vm99ozsrjNi84F0E4rtqC5OG6IGVC055QlHpN275yE
GWOvIC6PMz1zBp7Q62IqgN1XXFwduMjmiYSAE2rSfulSVp+mkVMI8xrLUCbxNSGlSMNUU/1HtMt0
4Mte/M0Sdd7+cKdSzHCNCJPpSHfHDVjJ3a2ZUyGdtqreuRF6eXlt6q+fLhuu7JOs9e5ovhQj6q4k
0hXJNIZcS3FlC9W7n/v4JDor02GrGyfABI100JFowLpMtmKwX+qXkdaS1w+0xShK5RoP1t8Ufwqy
MAbVVWoO/Bk7JvwLzrezkc89y+LLFicwmnxb5YHksddjIi6MkhiZrdHeJK/t1oeNJU8I8836X+2/
pzbkirvk4n83Z79gWFbx9e+WGXkh6blINZtzgL4CVp5xXTt6xH2mctRmIvwxdpJO3zo8Qt3F5UX5
nGiCXe1A/PIgCH0njZrKi78dbVB+W9SVBGA7OUU+x8mwiPBrTfRGz8eDNg8/2xTUuEtcety9r32r
sdd+TjZNbZgU26swKWSKaoHfV+AcvbraLpyoCoiDcS42Zvvok9JFXleN3rIzAo8LHe5X84DuF8En
leUpn8kEpzTglaalmPNpBjAbkRFk4hDFxNFmzUds+z5VicG+aC6ANt2lh50WzoOU990ntchc0rQp
NcHB3Ef6Gh5ogw6HNRrPxXi2bkbSVvHcXNzqKT58PK+L3W5YBR7ghslKr4o4v1B3uXny4oEcueAX
to+6EbN+t9AHhK9/QIU7P6XeLVhBw+LECtwxkblTe9NYbt/aoUz+JDRCh0YcNrD8/AWyjfXrOQHs
qUVhw8Mjm2S7ltkWH7cEsxYXArZTitpo+86jmTR/xZK1RUIN/32DctAeG7CArsH1FJoq1MH/1Pr0
tLQgz6qvG7FHIKlESuxc4eUIZdOLBm644qUFzUBjLo+BFXD2oUDTxp769mTtJ+08VlBdE38apKXw
eWtMVOVZFZlc1S8Xhswes1s9O4Wcrq/UVd/NVSpq9yedwh1jrxEs0mXuCo91e71/PAuWJjErjG9i
XODnGj4njLwmhmpjg56aadZc/QboZT/YQ7cB096gLbtgPluiPFY6Kv45OtjbUSS9sRPM88iCEHaH
ltFZudoIeYYG6wn+nKYaPWsaFDGUk+Nt6ffFA29zH74lpLW6hf7lz1XaAlfYGe+Ig07XA6qMswAB
sHroMuf7OBFYNm53oBSYONMac2MVGvwb5TmSbN/XlkEI1qvM1625UfUzAO5O0v43kHEqDYce34Za
+9utlRAf0iyJ4tzmapEutgHps6riZt1ve88yGMvrw5fvjY7t8jhTjfaN9nSWNjPw1G/TPH82Pxjp
9WMSMij3ESwYnYMF6lVoEVOQCgjEnMGB1gW12/L1keyTodMPiLOvVLcQMywpgH86dE5Moirot1ja
71laqZJSkUexRlkFlDrc7fW3vh0MEHoI73cHXB60L7y+22GQSbFWBIHmAL87/S9YSHNxPYawVhzy
jxkg3QHE+Dtjed0eCEi5GIIIVDSntV06XMBuS4nFTO3zIxPXPfYQpm4QEufyRP+Lmtd+HMZdFeLs
5cEMxNvreGb995FalecKIVsucni8KhaQueau9tectuXry0wYwTM7+hqQtXlapwIDWYWyix89rxeT
VBbVqJX2xQiWh13inW8vh/bkj9ByIXJSHcmPOK9lsR2jR7YEE0yucH7/A0TS3dIL+xlghTZl2JTj
f6ZHir10X5NqxxtTqI4RA2fEHQORdmB64E0vYc6MBrTaxnfFptiSPTJj24vjfo/nACTHUxEU8tQH
TaUkv6zta9lHP5MwHgQhfekITFZ2+9kaicM2qHZNuFJcVNTfVPDbFRclMpbT1oihinWobMbO+Vr7
D+rWwrljMLEkrKqMMatFnZoG3oUpuuFQNGl4blGDuIh2QEhO3IXT988ErbQiwrvPr//mjGT9ZcOs
Epq0swEEX5hma6KitpE0fFYCr8XljZxewDY6+dWHeHl1tEH3x+6r7mDrEfR765ASg1T2wH/BbsCq
9G7xzSUfqwyEycf01t0cJccm6qisdZPLh0Q5/4hdjL/8yFOJHRLK0Ik9nwPQYOYlGyP/VXPttevh
FPeH+hEm08KvSM8Y1pedeQC0ElrtkpRP7BvUHC7bBWMqA+kxn1jXSspaSpMGhqXEmNJ+SgHooVmk
LvHSAqOUZSuFGRkvJ+6CBqN5J9WJiscwBICdjNI/hjyiNB+CSdXWiZzzXxeFQciZHaHX/ywzGS/k
MvyVBYkZoeJzgJRt47SUGOn0B1v205VliKqPAbjIounvqepEesCBiXOnL/SXhcSWrheXuBngpaiT
IBBDTlJS6BMG4t/6dYseD4mxiXKv32Aa0F3iPedqMo1aup0NBzjgtZn7aGlZE7W5ogjrvAq0lwcw
+76KDbXTof8LaDsHqwYjFJ0YNJ9yujIl+O4t1+EMhg16yEkylwwKpmldQ93W0Xhq3y7bUGPUipYH
mJxW/9sO6xPUrxD1a/YCfOJHXUc6jmF6MOHNaVkAqieIuV60a3OHWHXnz677MU4nzaTcWnW3Doy6
ISZymBgJi8eIbi0PO7Af5kN0tLjmDP08P4dervDwcfel78Hy1Awn2bBnIImKcWbKS+Yfgg/28wsg
PFF6p/UVNoCWGu8kDGt202PhC83xIUqA8boV7esnCVuAhtuVpWwDOkotxaLU6I4L3VQyMO5FZXUx
NVBfGvqwi46+vMVEYu1VhoIiPHrqXdclb0Q51yU4WUrI+VVF01x0yhSdRBcpZIMIoPJevGBd+Nsp
rkJ7EgETrkJ62uN8XzLsp0dNJcp6ZKvLfYZrk/E9YMBuLVR7bAoCjUgU/8AVfZ9xOLg52KnL9sO2
NW5MlgMnN85JPPAT6vNrVU9yI+gq6AJ7CZt115g8o0VsUpCPMelX9W7+5cAedLVPfzOPtY3sD7fW
Ichmf/ohCjAjyCfXiX0UgBwPxjjT6tuafjbxr/D/mVuYnS4FLRLQXKuvQrSf6Oy0WLstg8l1hlZQ
hlS5AgP2YlrWNfqdftbsVu6YK/nV/poj6Ur0LLPLY2euxnqn0lR/hUdZ6JBH4sedgniPluXbRczn
Ae+x5Nvn7qIED66Xq4ROxYibSmn+cZrOf7WRgB4uacFZqQRiRBAUnAVBCQEwxMpBe+/FoysNg4Rn
E3YxOY7YRLffBqedDVfjhYQ66QbfMdnVLikaI6oNb08ERPuw90vyVmDnK/vBfKkKODe8G0oOXqKO
HM8SwF9ZM5O+tWDxvVWrR+oXQndp/iVEcrdU87Y4C6KGRb+cAtR+TxDiVAo8eNDGORCLyNPtwkik
mbHdyOw+2ldKSApInPATU4TVbQBJw/nGHvWKgRM6q1gMcR8YXCt1MjP/wJyVR5o462PKQrB1I4v0
j4Geoi7u8h7ur29LyinTG9qDKf5obFNIN6XFlKGZqplk22UF+puJQ5IsPH10Ou00K3R/aivn9Pud
l89zY8Eful6ssMpM2O7TRuXCQWIbTtcHOSa0pWQbTBeVUETqxtWPRgFmlBkow/bPwyIAQs8AIUKk
ZDlcR3wd3BWN7L91S8H1BNOlzfQC8jkXdN1pz9OeQzYq/vv4lJ0OvooPf5d+eGUk9RZ2KYHyGgkz
aR4EsGTv256bmhSdqZ9wzbumvgz6Z5vywzYpfM3TzMnk7tiT1TeNtulZlsSsT65U+4Y8hAKX/YCk
sQmt5DRzzUxukjdiZpcKwUiytXtXF55ITItqaUjPQynHdZn3iJyYxTDvWpjgfeRb7aUMGw0V30it
btYwtznpGgxazn4qJv2dG1LsKyTd9DBwEQ9ZazLxaEUj73AAmnpfiAMcRCuyPjYBEZb3NXm13s+R
XqIXAfIpMaspIO6Tgb2zdTtkqonh+81z4ydW/dVArxyUc2BgKa/ks1/0kEo+jgdWQJo7khtLPwUO
mur8+EvcT5m1u1dcr9K6yzIoDi74fBNrl1+p0KlLUejSaok8Y83gaRAZ9lFjMT4HwjZM62thonZk
WAvW2x8M7KaLSrCYHiZiGBjEhujPgyuSftYwBepE0QiA7L7EhXHhK81jNryLEbltNjh1rZCxnfz/
C+Zyu8jawO//btGiYJlssKRIf2TK7+wXEgVXh4J87ZO0y51c2CALJUueap86qIhv5S21yvYnMas4
IbFvzBzuDYLnerdt3JFfJu6w8SCrJHcQ2Pv0YYhWRoBE6uv6MS22sTPNxusDXbr2xv+bkWrpRxyl
EqPXAUbR3L3vE/IsNvzMMYVGCxJ8UiQXqZMH/TLQPmKLEZzJI5uqTxl3b4jJHFZUHiVl6EIyWcuR
GWSNjcrvYLmb72SsEtFTa+I+WZQwTtbAsIP0pRtFz8IsTUvasErc+Wi8QOJeAFK85xzV8cM2QG7N
RXeezOMB7SR4bK/ZF+9Hhr9Ydyrbxt2875/6Fk1KpkDGtPEulk2eHTK2GSeRpjMYk1yRgwqTHEKA
c9rcH8/lh0xXX5A3VCvkJAatzoANO3+Hu0Bys37QwvhXJsJ33+WsiSG3klV2TkqlHITgnCmq1QkW
lhdipj9PlSXM9DZMnkkyyOLmf1yDsEpRYHwRfesk2tk0K71W7m02dIhC5tfqnZ78sMO5xZCqCrRa
9b2GDHmPBHzx0Fuk9Tqu9wD7DiINGdlakPUngVBgRPqFmcXPRLEjqGaQBGDbNRDpLdDrIQSqqQdF
MN8JVbxmqBUQ29IxE8r31NmiWNaSqBwW4Zb6rY18NX1SOd6d1NpYa8EboVa/ZgMOoeP/QbHvOs62
2qA1Ltspy9ebOnQBARyasKPu1KSc7FdUSvB1DcyQDUG6H/gg83WWobjYhuuXSL6SIE5drFmDuXaI
q2nrbl3xdcq6f9EgWTlKOcWE2xj2Vnduxys2vxSLCu9rXEyB93DMGBHjUkqlBvxP9ppP7XYjzXBy
Mq7ndpl0VELNT1L3qFLRCdVSBPpMCPrKkc84Yx1ZH9PcIPk0NO93zeXJpBMBXeOIopNAi7NS5/Xx
5wXAAvbjrP8KtOJEArLtPuwunkSOK3ZOI7cNBnx+BCucJi0Jzl0VmwPV4KfqSnQyKYWGH55jGjCO
9AjI/C8yDdTAvrdTv6gal2AN42U9uRBbTwRqsAWVol3bmLYviFXuyOBtsgIZwUr1cLYy0e0HsZdd
tCH6+xL5lh2GqREFqIJIHXn28Ti2Z66Yw2zpRWV5mHIkYNQGOgzDmKGzWoLxKt2/tIad4YtD6QlV
ce4AJdixwoRrBCPH2X+rtJjzLC0q/1rczdGsxNM0myMdXZKgmM0O0W2tQGk2FuARk33RmbOEglt2
hpve7OegHYr8Uh4l6ItBRGpmlPaB5nGyt/4/Wm2+ZsiJCOtq94ysIap10Mewpcj8A2aOWvy0LiPx
TjKNp8/oLtda0L8chgsYy3dujeLGzfO0alcKXiYObMioHFobwzShbaChYYhr72wHPL//O8kw2/ZT
1qwMO5m4Ew4oGYqMRr0r4TJeZatNwRs3i7otHUfK3KZ7LbDlg+VYnGpacQ1MOr9WuQYOlC77whGe
R96MzJ+QiHb1no9D1wn62BPaQpnSs8nip6bvJm6pXuEQJJuVjG4cYxaF24HoDfUIHUUEaOXGU2sK
oYyfIOOF8Pqlv4QlSuz1mJBFlOM1p1xFd3xvKEx2gr5EtN1yW6FrpQl3ZKJXtMVlrB682BiJ0aZe
wBPHZdykLpBYmMsFHagijFVW7z7/xjhNoZ1uNhvFJPfY3aGSxhITjkelUAfDkt9/KyWUPDHNszes
92uYco/ZFTjd5kfOLkXyqMVWUnnTQkbrOHaYzp25/UcAcEXRRDxNyNDhE76DL9XA0O2/5eznDCzv
BIAx0reoSPRZuMMZQkBw0GeFGcRKFTpXzERGBT6jlpYX4CWdp3Wvf6Z60cTlebVP7zgEAV21W6Pe
BVK2BVBPPPSkbaoCRXV96e6mV74CUs+4ZXNijdBJ1PmZh66JNAWLQaNHJSHZuubv9gX2QErEH+/4
BimGyB6Gh1HEdvxduNDkU8HAb8PIRW3JUmVucjF3M286Z4c2jyyy9CPiYgE7UPyzpVM/NN78FxeR
d1GqWKpjit7KXIGZSH27tVjlr5kiGJVYsBYYGEe6Fw1OuBxvSqPgiphYo0UpyGwCyWW8nZGT+WWa
RP7FvcgnNMfF8rpMgaf/7vGmLkzZABuY+PunOYMWMMSXE7lFB1PHUdEpgNqx73513ezo4zh8AgUU
H5Yl3l0IXX15682c9nDEYXv7czuBXnY3Vq1TXJcZzGxg7nHPbhRbnYRq/d8q0oDeNMl1Glo0yHgS
3CxRPXNtRRimH6TrbUNSHWAwHZXtU9JLN0hIvR96BzSvbc1xnlBJLJ+FYuZWR7hBaivW66jRYZtm
IDWltLqXMRAmNqmxGUW45Y2TFjPcGRZpLFuUnFWyoaGd35ULCqV8r/3KjcSH8Knj6wxbMVVTFnMR
phKRjXklkU410lv0MtPU5lp3tELTyw1fQvshmDP4t6Rily7dnxzmL9u388hlfB1/yBjZj03WZQIr
VmYoknGcw0oBMeaO0ungVSxwaHcAu5E128Q4DNhn4mmzUI5vAuAVq/w9ik6U3FElbZWZ43jWwnkd
Ox2SM/JR9+riOd/BtTXlVfZLFvJfrXVGN8OhefyBvZ6pzHNjnUbtraCpmnR4wVlA4f+CLF9aVE0j
SsFUHg48qmeF8hMUp/rq70PB+Ww53o5PP7BvohlixbrcSx2yFdJWMm4TkJu+hapMYw/govz2BR/0
t1IEEYeNpQer46my8MS1QyjL2SKSMyTxYZbyHySucIg1pyK9SYw6k/EvE+ItZenmQCT/kj6EIPZV
yaKJamJeQtALHr8EkNXgN9I0zEOIAx2L9CUJC4JS4zIgrKwxi1D8QsC4p8+iUdmcVTPPQhOXGi6s
goivHE6hQgUjrcY0wEhZpTOywYtDDYJDoi6lZAmvmU80WlH8zAKxvRRs/+X/Swm+i59o75gkg3l0
xuNg2n58jeMOyCYo8Dbzh6lCahhkKIuuYxrCOBxBqnsE/KBTfdk1YMNMdr8rkSmLq04U23pYo+XJ
eJkULjxJpaccgWIhL7BtZikIq2eF4t67saJrEssr3GVlMWGCtpX2u1QEyw/ys6Xzan58WKHDSrZ5
Ze5Gz7pNUfj8fmWpaCEd6LaCLD/n20oHbbwT3PaL1OdH5fGNNXK8UDAA7yrHzP9N7nvoPY9jGiM1
29ejWaRSUNHJw/iIsqYSTXVBKQlbb0oldtE7gY2f0lHfT9n34R0B85TRqh4y8vKiPRRRBO8JSvey
HG3v1dC4AZIlfAPHcDYheF+b3W1tT4SqUpTIwm3qU113qAX6sCj5C8T1Ic6z0NGfjD5MWMhJLmvL
hEd8I5grrmCqJkH7YTxl7fELHW8xHTMHTDPg81JZjaxsDI9kLPc4FMYFLXmuXp+xxfIZRw8XEbkK
IJpUHkypMZpM9d2YcxRXPWpkf3DicmsTgTQyoH4h0+O5j9ok2B1kU5S0st5q/OnR+NELzDeDCFWx
GrZEGU3OKQPY4KJ+h18krkz/D3vdRijDJkBoaHUbN12m9Y8xzedPGdlEQWu+L1VeWTfgXS2238aT
IlY2mGG1u6fCW7CjENdoWS/ey6nJ0f+4MgR2VDYxJFwgXqfZDP3QxNlRPvQvxq5f9GuRv6rc75E8
r1/4SF+Bb6HoVvHJycSNRVrsPVi/3T9e+CgqiK7chJC35TvLbuWTaefxIjJM+7TL4tBXwCSigkXK
yYll9/1T+TwIRf66sJmmgDWVqBgNUPNn4aU0x1y2UhJnpclJ3hWeG72AJUJbnaSl6R5G4X4PTmO6
9/i/LwDVSEcYE9EY4Qx5j0qEMGXDfLm9NB4qcdP0x1ceoN/CTwn92jP65i7e9EAZLvowiKEVy9jC
5xXXmj8vj3O9OKSWKK1V9/VO7XEvAiGA5nIlRyZyx6ZT93RwWnP76wiPffxBwvrk2KawIMeZu27z
ZuYcIcv+HB/7eLskfGfbbcR0wJZHrw1f3NL4v1lMSxJdwuapiQK0yGOE11ioiXoez+uCVrUrrgWC
k6bnMZ5lVirokTt0XjKz3KkWT2HY0ve0WzlMg0Dh0KCeDd0RfexeZDhruEipXM1BRc5XkYrU3Pik
hxHUGn8c2pfJvCmdLzLYzlPpv7QzVUV07DBuJb6BHSnGBUNiqop7TdMgQSqPziQHAfG/U7Wv/Lo+
P3+88ccNCaTboKxHbI06typW2DQXzrGAsEyIXok9qy364MZ6lOjM180NDivTlvTouT1aCNe5wWpv
9K17JjNOYv1PFzDNQLwakPufMN77kIJUiIV3wMGcS2yRcbMjFWEi4VctqU9QntzBMAhh9unLt2/3
W6PSBKD3Jq+ikQ/7fC+YmKx3xuhBMgdklFNKw5y1BJPoG54rVp+JQmNWGYRDzOirs1hYa9y3Cgtd
HdeeM73QBQExsAy6ry9m6JyOQgQVEb0+XXDnqd+bnM7ynotxBU5Q6MQuy2VR5W/W+eRJX11wrRyW
+6mdl06Bcf2nqL9rxKHt6IXvKFeBKbNpojAnu6+i1fntHuCvcDq1aj2JsHwpJGzPM9eKnM5b17Sx
NGv+L2+f2+L7E1tyCElOjLZyrHPAZzazzrwlYIBxN2K6jupPeyH6LmleZjv6gWvK/TXr64gZjwhe
DWh4RRRXu22W1VfHOntSTewDrO/hBOYBQBtYdhpvyxmci43yTfJ0TsK+wHMb2iMW8PZ5anB00gdb
B20iT3R3Rhexf05LGMfkbbwDQkt0zZgf5224B3N7Gbxejw6r+Zgpt0LCAhHgWVrZO1ZwsD1CbznI
G2fO6oYuaoCucF1kN1aM/JJzvzYCiboKL8gLAt319Ue9lexuamQwop27W3+SnDe2S1u3dELH2Hg+
X7L1ZK+Okn1n7QJbLmCVbZiBixVUfoz26Cj4OSELEBzLuDVE1rfxxkL/pPnwEsCObp4wfPpW1+SE
nlQv0KI0dj+s0/sNo2XwsAwJqFiPuIA2TupqG4cRWZiT5RkSTMII8r5+bu55P2GKhgAuu8Jwyj14
r340L3+jkd+ikJLfjPLrte2r6xItcU/ghraPQBeovclJhD9O7UWBAV4kZrm1LeaQOSV9RsTlcpAL
Gm5uwVJKnuZFH0hFZnjM3r0NWcxzLBllpwF0XWleNN1rKzHCRVkdy34coodqXJ9CKMmj4pZsiXZR
01V/626XMbSA0p1/5DNtdw/HbJWKpme2LIY/Z9Qa53TM6GiLV5rQ05SDv3U11JBv10WVgmSHRoFY
05owtxDbka8KS+2n00IWwC2Qbu9zSwkFdDqe6ejT+swP3Do02d6jY+5QgMfASFOxamxneMx5uZzx
nOpFMTYyeeCLJy0A+OKYYFN9syOifDltnu+T27CT5eJSL7IMi61sd2aCHyKjrD6I9WXYBIQ5IHZv
uu1/hzZneLazPwVtkBNuDifl9KAuHTbjq/V2r16Vmr4BMMVF1BFxgIPU46AZ8S52wbfQ3bUkNwOT
wm50f2avSSVh3xjH9TdrhPohqHbDJcQJcquBy8fMwochvxTPC5hnmLO0KCflXhMxrSUNVPVNtnYy
E6d8MyyAuHH6hlmENd+Gmo6lvy5QkhtC+PkilTaxCNb/oZzq1RaHaQV2XHTWPRZjMNyqUg+Qc3MF
DdjfilvcmrN6ilGkv80eeHrF6MN7IAI0NDy0syIz2+Z2ZjCNzot7787Y5Futa5fKtjIFDIjT6QMJ
en/nPsWDqRN0WyVyN8n+oCClLUCFCUXcHRzU/E/R0CN5RZfjS+Bs46Eod4aUyVBVrdh8alxKGVsE
Qf7q0CFSctaiZCx4qwP/e+lLi0PwPwDmLXtk8hgjesA0jvCijPT7PThMTQCAPf+S5GDkH3BbHXFf
hhqigi9Zgi/2HHOyZk7AvUS+rGXyJ7nvbM3Fvsp+JXHpBtUZpBbyW1MRu5fpiiuCKUGAJZUJ78fV
AeiF4PmUlmCg8KvzcOHHSWd27uovwLkoOUcnkiR2TxjYnnCUgisMgBwF/VJxuK/nImkbOvfMwZ9H
EZRpANEWbOwBEGCCtUft16wp4gR9sDwfDgAnisi5R36r4Vg33yCchxEnimnONXpqXgc/95BBD1hk
M7EJLEiyYaTAGNGrtZXk7y4PVSZXvOpep4t3vQNMbEnJvYW+H45IrjNaMPiupQNiEUAMA4FLwYK1
MyQYr0tcIDk0DtRn+5NfC3KDUd4V3nztH0b14gowzjGJ4cBiEHVEicqjfsrvsIplc45CyLfZCwZ5
g/9iMvzOumcs6PuIZOYecsolmHQqV3kd91U0P/Q7WxQjGwYbZBfgz1kDU7ersz6Q/8FsRodaLC8X
Tt6IKVXQUGOPuX4DNLMqnaKtL2QCvWW2Xda+lMg+TffVwPiIp5LHg7+SwMZU6Tjh9UlGmBP/8V0C
n9ibwZPwaxu6EDOiKLHvvrngURdWVjmHLstsLHGGQGWGCCMgCBcfhaVWpNTLbCOHuqSlt1fleHEt
H6Lsb0szkqDx/A1k32Xq4+2n6I/eUqe1bjGmBcnYlbc3ANiKSAZo2XbJT4mm3eEUbOtqevkW//ti
IDlPcFQGpLV2mAxFMwQmEX6NaQpKBS4Ge7V1qp7ATsET4tkd7kwVhXCHe3wQFHKhQNxX4re+6brl
MMdF57VBHNpQzTvsg5OQoE7d6VyMyIKqu/uTT8gdKLfmxhDq2+lGMwR0UTvhN48PsHpFb8BLfVTW
ukyCW6L9QJti2Xnb8kuqtdjca51/VtY4T01XcUqVjQrcrEmOypHd56q1b/nTCCQGaazv1+Ftkpx1
aQvgOlwwWRA4fxZzVEF/zb2q6chRQran51ENdCs8vTUbrZnM2YgshLwHbLFxgrqdbJiK6ZS04jN9
rNoNA0/Ec+okc5MAlXycaXdXAFtpu+xFXpOvW3/eSR0cWN3+j/nhFQ6KbmPpiw/NuRJT9DPGJIeW
CCOJsiX8abatsl9cpwNMJec1n879UpDObXdParo2jlm7h8+IKnKUihHRNDAu0FXHwd/piq7VMIWx
uBloieOh8nSrJG7DUPNepYBOslYNcYkxHI6JBwa86JKXJ/3dnRgzkAPEixafmATGdIZJAezdkqpc
u2Fd7pcsBywpqcAf7WZ/7VwiQyNcAo9k0qaYntsCc1QPI/EDS1egnT5RTni1mGlfDDj/qclnoWtq
kncJZ2vjefgsXKnW3aAX5qJb/eZySxunhyZCHqLOqS5O5E48XU+X8krgnHTwIq8to3dUSzn8lfpJ
nznCNZxq1FSaW6h/otV9I2i7boWMQl/6w/LQWtCq2tURG6raBBDQHko/IY7tbDLyRh3sqvE3feiQ
gleTFQqyFq/L6DWbhd+9bbDe6Lkb0zXkakApzmw7SI00SRG4L7zSbJwrVM/wmNOFp9VJMQ6A6GDI
5mQkTxASQiiv2y+xOee7JTK2MNGx5SXbKXBLdP9WLPGxgGEaO/E8nc7NYuiSnBEwDsO/RzQzGSvv
PZvLlqWCwy8DPBLN8VRv9GwNwfzuSyVEvZF8UVyi7D06EPZz9CK/8C96ga0IriYH9yEdSYUvvzsu
NRbGXZgbC2bnJ9Fgf2bO4yOhGhf3PLkyb8r1dT1O+hmh/RHpxXCwirU41E9sXd9LnVw2A9gj3r2P
putKONXs8WxXR64+ZJ5WTXk0Xc3ance7iKQNuotiUeM0g/TMlX5ckcW+INrL8Ix7Ekoo4akYv6jm
Wi0bMcBc9S5MYZAlOKnVtfIgOHUutdIVviUozqlQe/V908WImuwKyTzFO3xDI40HGSqqhxhoaVG0
yzPmE8CWbv0FZ+o/9c+EBIG/knFa81qdsZz8xjBX6+zunoAH+IKY23KlhaPMs7Udz6oZxWxa3Kf5
z2+1mWAHxA/6KY4/nNVXmlKNYNSblc52nUXLlUQXnKqDybv+G78Yo631WI9mB4h9KnESn5eARHcS
F3nJEUNtSwVYUL/DiA8JJr5cbLBRXE1bpMXTYkXd4yCsipBN8M6Cz7WS0mf4l1D1S3K2Ifh+zwAw
YV3DSPwH2R45kr6IYEJq+6ChDToPjFaRnr/x5iNM5UZq2aDrNqJBhfNXwFTfEezK1PgOXub1aRjA
cd5tb5k78oJG9dq0KqHE8wvH0LDN4CXE8dFHVOJ/Yn/NBDj11gHks6GtOg6wZ7w0riES+pmMRH1z
ZSykBWF9iDNpAR8RC276egKtmFGOh0c0+2F00XxULmLyQzFqkvzESWsGAAeMBriBlfy2pngVgG6Z
fakJJIXSS4Pmzp6ulotit6jFD19h9CxnAjZJSZvxzLoBzDvrtIKawhiUHbUztOLFIU/ndwStWR60
y6tw6/QAPgZ0KqxQC88452BO+4sB4LU2xXs+idf2xsvjLylIXQDK/Ik90viRrfXbIqYnm3M6Tukm
z8EsURg4M5Ipl214My6UMlGrjYKNCGpMTWAgkok4aqrgSqn27UXYuFdjyrekPzDR+OJjNe/exm9y
gxcz+np1iPyVeQtHxWd1gE4asjtn5ZcWWEuSVDRyHmTYbzOYVwvknsuMDOudSK8Kza5MJpaJSkz2
k4bR6sjD3oUMvPJDKOdsiC1DvD231QymizEC2TFUuaNI4MKM2I6Z/4GcRO5BXfG1vIBffwW6oXH5
ceF9udt6+HaBrPFVvABsL3k2vISxOMrflDBV4xoZoGUAo/8VRE/uD0k8l37uOgDYWWIhYbV5wjUD
gOFNW1SlavbBFFjTlhXk1SNz5sVWlKpkO4dgrj8SAS80rW66on7rVxaQerNTI6eENxVkS4CRb0FS
3e8yYqhb7lWOOXRDYqS/Zha9QjFqQsppdXvHusGVPJrz32Z/LZORyr0oowCpEWFVUkCHpOkiuCzn
nMTANpeAB2gBJ2pu4iHPoZyBcyawQGtM2dyqLqhbaF6AYqPmBbnNQzDHI2vZ1BNzH8rx/ODaxmxQ
Zazk9Lw6ppuXnUiQRKWWuFnFr487T1xMiLZ5gLkunE1X1p6a3lwu/NTsa4SIx8po8hJk3B7ld0Zi
4mLwpJxvT7W4QjSuEgp+R0IkYkvGwEjBG9Rrz0t1Fjf8KKFxwvyjTLgWvWL8FJmvsgW2moyGfvSN
mksrEDOaG9tCfi7pwChnuQvzVkHjjRj1XqJ26US540POJJEQuT1UzMPdlVt0EBJBDTimPlk6E4IF
E3VdmKmlzntC8pMhn5AB0NDe4FBtX+2FAZDxDBPS9vsFfAAQ3fB4oNpSIoAILkld2IB6i0M0LpZF
eXN3foRJmnfCXXNN1xb81Yxb0pYMYiizaywCibyl/fu/+71IvrqPVY2aVIDW+FIIQUTnm1cGtY7v
zVD/FDtTHl6lE+dOFRZWvluK1O4nYopGP+24updWzHTOAelZG+uozfzd2+ZfNZnQLTPDnRv/58Vf
fV9BfTqq44bfhxmfm1wi5wlsMD2ikAaU9kokbt60KINA5uq14pjwTQs7qLiDWN1WUS4ZSLaIR8Td
Bs4CA3iNIynF8bz8BhrL3EdxpNhdZcAxRDuQmtUh12R6AyVBD/8x4XWsHwkvT+S+E5UjZ6+uFQdO
EKtK0aaEa+iCTFy1V+Tq5OWwmTZV/7WoNoFoqG6B8x84NyhA1REclaxGr4s7lYuOLCNIiz57jCyU
yxmZfWPqQ+ySoobGhnUOi0Xg5RHzZt+VDjyoEg/Z5hUbPKPfbEqUdzBhZa1Hq57oCWYiyX1tWwBc
Jtj1inaSwgdpckp/pMLWKG/P0LPkNwMMSdC1fPMUQ8qL10ixGUBfDvY+Ubiw3AVTmQ9G2slVHd8+
6oNkZdTBh2KCXDRQSH9dVJE0ntUPTBuI78LfC/fnQ7q10bJ0StIkgurQ5wnlJrXw6RuMRZOK60Qj
PT8mH7+xu8CJn4jllD8s6ApT8QTbhb7SSP2/ll5UnGoa/9lVK8PZXWCqmureWNsI1LbDY5puotCg
k9EjpSeIfHvan8YmiqE1CPCcajpxBVqZyxUgS+HqmlMb86jIR5SP4yX0patNqwjoGkvb3QCtEQKs
/w74X26i6aFKyA3BzesBN3iXbsefjoB6BIzovji1OSEsLXtAUJi00atX0dK1rrK0BF0SoYSd1nak
Sve+8OMLcFtKG8cymvXrhykPUUvt6H4lmmWtbWrs7NdFcY9mMJ5NFaWtIFFQMVYaE79G+eiiJnKD
RA0bVw3eCdWvX/OliwN2wM8FsflivYtbw3xtNANnZs6F2Go5J/JZVWFLcT89pbv99WNNcgoSZ/nZ
vljASwsPvXJ5XqHITG05MyJdtNtR4cEIQ3m3rZIlqM5H4TYZhDJXeNhVKdJWyZLJNN/UUidYEURC
ItMLYagsqBFaroTocjkHTCULtRYqv6vN1EOXaZCFOWYNAnS5zGBZizRN2WO/FTpYPa6qHeIpYPK1
5GKoe0e8EmmXOXf0mhiRgk6C5dX/WLCW1VxQGbCkqKzxgo71Oo43hqB4wu588OFnDzNA6/FjQIgo
RpJdc7ARC8LWQspoT45wBr1ajnSoktg3OmHdOt9DBXR08LvZ/g/VzwSP7MUIMNmTzgrpvKtUqIK+
6FH+7zPevkhfei37kijL8bW0tyaxMM51RzSuLDdd6WzEtGPteysBiaZjXBVWxJFwafaIh8RCU7PA
TjKgZIueO69bMk+alV2qy7qEBrI2dtT1U7F4zpdgEf4P1hu1ZWcbp+LFRU/cqDoRWK0ceM6Ajgjo
ELOOodfbg0tQ5zSgrTcSU9QAu7ItaYFOU45bErQ9rrphxE7i9oeuQ06jSKOkVGTjYGs8UohtNGci
mYwPLWwF9/NupaNT4u04z7wVup07bFYkpzTGzYI1pXeKoi2AvoJWbu5GPOwCT8cr4T/WBigavz95
GdRVX0/2XjJlA/NrmZCfDUZIPY9Is7KeL36tGeKvUo6z1Qgzd8xkn5jphUWu5byF6nzE6zZlY9CL
ARWXsQX1qmrhWb5JAfdps/1iW866Dlr/YLPoBCycCUE9SdhydKLZTzfIGdP1e/1Ce02wrIcDq7uv
PFYsEObx6wgMJH7Lcafdm6W3tpsqdwUm1KH27BfxR65oJNFtvMMYY7Qa9bzhYzLBruh3tQ0s0/5m
n3zoepfjLiMunjY4f6LyR2X/Nreiafz2O9qSNk6A3RW9Nh3WC3MfTd6+3hGDZ2K1ELmR7CEH1eW3
q4kzyoh5Hgnc43tHRSUvHFISoPhU2cVBMp4jy+Fp4tLtoMXSgh7CnVZspQhrgogK2/U3kw6JLYUH
VOIlnlasDYiqPYMfrD4efzHqYXHRL3qVth+0xB9eSYFWAmiDn1PwJR6vTjRIgFUzUK/t1E1+oHUt
1l0LpM4glMs0Jp4hRZUxT8zxtHZB3a5dPVbsrXJyh3F2smJaCvz5T2n96e7/ozSRAtp+l9JpGJJz
UtbEYDMvg1tYUdG/Eqa1zF9/lrPNGSbB0qIZS+EA8nvajW1lDXMz7wnlyVl9YnzFUEjWCdTohx8T
cXw9RNdNbP2kRrSbxBupyv098d6Xwl34OknoA5sDumv8BPwkJgnAJ5fvaazE8XnzTvNDwj8d/8O6
+MKrZBBCjEM/oUO3ehr46Orp8Pjd1+39+dk1HBjk3Db8H81JrFaFFoqOYqIYgingo3jJcbuTi3oL
4/cONQomBM12MFiabcvj5EWVEBQSy7JZVFtyZ2H53UsrT2bxcNc069fH5jr1idjTFYxVZb7P1Qco
TyvYF1PYITGKkBpVvtdcmp5+O+M5ZrrvVyGpzYyFAdom7HeYd+hf7M3JDrqt2fvx/KQU1pT+4ay8
EaQ6tmeBM1wesuF4Fb0vLqyLHZoML5owGZFvOHX1OAFBT9ouK36Ls3bOFscTW/N9kNSGJxiPt4Un
p9HVNXBE77qNpRYAcILbb773TbaFuPUFLI6OyR0G2xH5pjl+KcoXGQlO0Z0W62ao2M3+QrmMG+55
D+OBv248qluJsEXWKagw/PLq/jlISFFh56w2HoA0KdyiDqFOnAeKi3yqPjQLE/84ppJDoCeitW36
g6NPT8o+JZYrn9nMT/J3HVY4Eu45Uly1rv+lPZpoHFr05n7aSkKvS1dAN5kyHxj2p/BkNy9ja4p/
nxg7TdyBmNMKkvc+2LAFVg5Sp3hGR+MDH/ofu2O38AksuphFlqZdLCRooefw3TVcUpXHxfcnULkS
Em1cTBOCBsFYzUAot26M2NpatguuBmwG6QiSzfU3ToAYQRuaX5qhD3QsvjG+l7+WI9MGu8V3bXg7
w6B9NqSrX8KnwZ/m+MkkvC5gb0lPwGwQ2DBTFUz615EyRsHMZHjsjSkUMkrnNV3XGLRm7T+8Ijwn
sjBZ2OTpY0a5EoiyhVl/P9SqF3MuARKCS0uPbOUMUBUe2523hrYpaLZpfK85dME+eTzpin8ig2aw
In6WKGg5AoGw8/vJu/39t4l684fAGCS+x79yh4aEBwOWa4NZSI6cpSy5g10cuEPW+N+N4zd2my+M
lCzeZjxJuuPlUdngX4wGgxP00lxF6J67XvMyAe11RP670d59QsqJnATnWw/nwjQKcgl8zgbJjDO2
8gOOomb6o9p/S4TyZl3mZu762n/Mu2r6aawzJGObQVn5GQB8Eu2LkiNqKcjNF6leOVikNgzpQ6UX
PLC3M/Kx8d8Q1mNrqOpVAc4HXMqSLUf/1QwG3ZBSlgvRc9mbscgdkUfm7RKsb9Rippd/1VenVCjy
2UAOUN5yzLNxBrJbRIqeB2jml8WJz4V0GySSVgAVIDxoSDXrHR0TwKdYMixN/x/XDrfE+Qy9Povy
tqzd25+pnj4u/8Out9/1CS10PfF1ChRekN6ibmyxgTMg0/xMOGJ+SR3X8DZMaiSpWoJ9eZeWobxv
tQxQejui5NOqvqbRlvBFvqkyAArfaw+bm+EGH88RRtLvF4yRs5asGS8w28qIHwUCAJVzjxT4gAUY
b6BljtsRQM67HMfI/R7iZXAYck12XZZ/KTrHgKvUa4ClfBif1ZfW63a847x5L4Hu6O+ZG30+3000
5/ookpLXalr3fL0m1ao1nQ4a8U2BTgIBljb+KiSQX3JNs7a7cIoQIh0kCWQF64t2VT35u1GnSFcd
3vk+qMZGFjKUDCzTfw5t0kd28Zc+4X7bOY7UarbqBtV4nB/UDasdqv4P5KJxPVDhQm/ZzZXIIihL
tSaGVwHcObCQRaBvn9jNA3B3ZTRNixOViXPMhKFtdVjx3apdxwcqPfFvvdUHVYnnV572jt4lpc9D
4vPhvREY9ZApRCFn81NWTFk7MHekfl/xkuRUfryQ9VR0oFnOEPPd+dN6KQ4grypIpV6Qk5KsMiEm
+Oo0F47AP2u+OV5sKTucytJBn/1Vb3qcs6VsKeoWbFAeQg0pjLqUwgW/9+r+2oUlUERsZzYY0OTA
U5nRW2C7pKNsMZf/jgVk9zAzKNiqLhy30kU4hrQDItMzrZjsWo85fEC70gt/gXag4pinDQQOn461
+wiCwoy2vmhCIdOfeo/B46joT7iLy/orsmLgpslzIinCcZ3TyPefKPwGVlQKDct0w8IFpplWrIQ4
UgoQhHogWFqpHs+M+wLSikU3pH0iYzFy17O+QMeLAG7ewArpbHDnGO2NQ96m3mEa+Qd9VrF2IVRH
kA++Yhpde0oYireHLsqEluhBCzPqw6s76ZdsUGi9wbzmX5jcaa31q+6zYoPVrQ6h7BMHlRU5uD1w
4m/S7TkAeYqtig7j8l9H/EcF7Ydx1Qim291ZxmMZ1RMeVPVVfCbaEjYG5YnSrbeRjIXwa2sHPBS5
EAnPxqDYDe725qsiUHwIYzR2ZnAuDMgIEXNzsxVEitGyhq7E8Uu5nKAhRtRMn5Tafa9WRC98MaG6
Ury3918d4k1rzWnLS06FTmCrJAxKoak1y8fpBlm8UH54dJc31nDD8Co2rsYVXF/zCJCdUy2Db5Kd
5lkG9KjVMOZ/c75isfSLtZsWsqIF6Rj6jbFT0CQe0AxOBFjOFYIyOylmk/dx0lojY2RNXacocZ8X
U6o42Is/BJW0riYRI16Yyp6uQ/6MJpkTt0N0hP+AQOIxtO05KwJopTf/aE+yGH0EHmXJ+3a/5Vwb
+OYZegUrZ/SgNF8mVRgQ0YY2uA2DGLZGdUHKlrXY27SZdRbC6xy1qENeyf1BeY8i7TJBtzUhT8Kz
zzec9qwAq/2Ul9P5udB40EjVgisRLej+uabvlhf4EBp8/DPu60zuO8H3AH3exFAJNdhW0Psg/fn2
2qhA7mWP0joZllvpgiX/91FBJWkKgH94m/jjLFv55VnZfcZh+gfF6rytpmnFEHUCazxll25ucKB0
w3M+c/MFLbHd8bqC3jnL7AkZhIidi9V6QDPdF5GcjL9cm9b0hUdTcpmJGPtE9+cY4AShMN2f+3VL
CD0B8AerWWYR7Mvey80wcKNllVmO6J0vnhzs3oWgsiTP60mjiTYobSk1M4c7LvSxCNy7ISXntanZ
pe0H0wgc7a5le6YLtp7pougoF0m4s3XeNCK4LDVYdXZ27dxLkeC3lCbn+TjsyrAA9TB0PWfWcLfs
eJDKi+wjG9VI8XuUMJhcmKz0yBShOmeSbRuiJg6kUI7iJWsPUXQmSfbptfkVmiT8tnMzPsrEAZxu
QyCoIQvzi2aTGFzRu2c7aWoRqF1y03j9FlIo10Q2o4RVZLHsMaQrVVUcMis/PEjoAuNg3TNvpTlc
TD5E0sklV5BNnES7nO+77i5KdRUoE5q8tGqyoHJOmgKxM6gbjdhv2Sk4tBBREdhKiVvcG/S4eR8E
dZ5p+kmSypzv4O5oW4aIfc125GyEYlNkmUu0wej46UVEmSzIBRYuIu69DnI9ihQaYEwXDoAkckpB
ec549Rg3d8FzdgBGOqL6GAiibIOPQb8QnGKtHG74AbO8zEuHamnm4ad2oZg2El/nIuzLJKUx5CdD
Oy5P5Wgi5dsU6USNizXH2YoXIpqT+HcZGAVKfk1qOTiB7t+dNSChFqW8mrW6v0wujChOEoJmQmh9
PB/atMDZot1BFYDk5+U3DDt+J72dvKirIRo9WOMJ4dsLfaG3wCdRE9Bfkj4oFAFzg2WYo01x/Iic
NJW68MXCmH7pTUJ5+LIaBNFCouT5lTXbYtOPVKvVE0535c1ARlp/FOcR7yzSYs5Ck7vG5/qz4geG
Dr2lCXEpnuqje3eys0uWqoid0INg9gE+psgS9w0z3GdxFQLDh8mjaMaRjHGEQ/khaIx7PQzbVtHT
Pxhoffb9K7WIyAJMdhI31tG/utfaB3eShDNouoNJk1ASqk/YBiYNRi0h2pJH5cuIUP91FRlY9Byu
2BzTvYaWjjavsshvKZNdJm/SG0WISatSEUMqEA+l6eBZgzc3xe/6VXBMgBTNMStvX2tTPvYSlDbI
J6IPCibGol7vxK6a/Eqp1knHW4rWwg+X7DNfh06O+sLfaKdolcVf9ZUuDhjq0ms8o4lOMkUeW06A
SfbDjiaoVj6o5/tsPn9DTwBkI8E4gKNVx7xXJMyweUwoZIxfU9ZVC934BfPT0f9PvCytC+CGYBT3
BJySznxn8Cc4cIIJ0h6bJdysOxKane+zCyTSTmsyZZC6/zTYtbjosqpCmTtyJzFdb6xbnPSlaCJ1
oL02sM8VabI5FBZ8TboBXotkbbp0+VRELZAKHDv3vq9HHkBuiDZuLBU42Ceubb93Xc0pmER1D0is
NBwJYNMkMiG+12lD6XKwyU2IWJShHinj3OIWkintM4L91WC/pifQV4dIP3qPoSR+T3rEimXcAW/C
IIEKE4hdgzJMYIRk1jARYpVHjwXhPeuNu67H281OtH2HbzX366UBxoMh4rMiemp1BwEvj8pKXk50
Xxz3wkjkJx+pc9Zw3ea2+1R6rqFoWekLgdQELfydDnWpznbdBr1eHAve0Gwm7cVf6xuhKs6TYp0x
BaPCC/FCbuEwRqSqkF11QCBuyKh2tR4gvHq16lJ1kjRoKCCS44NTYNIrSfacIalM7DhIACbYKqb7
VCa4s+XL+pL6xY0NXaFmpacMOu/5yCCsDoivjC+FH4vB6m7xOBWny1sW55uiYuRTb/wm+vrSCz1g
QjPKgyTTc7/XqjFhpDcwDxD6ciaBAD0Or2PGBJCEH0xPpvg/qGdb6oX9BhGrpPTknDRGbqrAAHwF
hwSj9R0f/kclVdYpBhSZdfVxcb3xYwxpp7QA67RWcJis/agweYDyIJsR3LGq1BMl3DeyM+k454q3
VfpC+uJf3HHzdKfBoErGtGSS/YYvJRUwW8ZbciI2jJ7B01fYHnhQW4JHa2Hndp7NuBM4HFAX29qy
JHPVIcM196MoaZ0bcxgjkGRNpUCMermUKOUKKZfI53UDkOVRrccXzrUJJyK2TW8cGw45yUv/Eqyh
svp13rdMvgBo8OBN+6jCDr8tCOqViuuoEfUhd0LItCVB4lzhE1sHl7MnKecIwPKRfLCBgRhHyz7x
PvKEBby7eyNDfRiXdIREG+5V7ivpSvOMCujpHXqGTP/rG37zmCbvhcl7tWB+JP+IbTLMqUad8Ktq
mkKJPF4pk5TYv7ycsXOx/8MMVe/xuf9piqCPdaoeSI+psGGQ/otc7EO9N63GUlWMxS9WXdE7ndOJ
WTcbbqhvhKuPyND7P+mhBQKnb2ZY09ybNVCl23QkE8jNHs5fnE+b9dp+fzCLOHAymQyxs4iAKJOr
fgNAD/n1/sR0V4j7uEwaKGpuchr6y1B7gZWKw4iqdr6njCqsRVsS6u969RTKrEGWMxOr8dl8oelM
OGiHI5BAYA58QYAyDEVURioJEArLucigzwLwVIKaZSXP1Dz5Cmz7TBxdrF9pL2WlJILG9GxpHiHo
UfAHtiBEZSC/NtObhIyS0YIKrtzEdiyjzPhPlrWAz7d/ha3v/Kj229+4njDpLL3RCK1jjNr0MNkf
jEnbnlXYbhXH4fzy1Dtv/1JFDGW90+Ms4WLYHOGllpfpenNr4rVXPQW6k/DON7VzEAz2p6psppEw
uuqDcqwKsWkJNxhEKZOjgenY88WhZCP8BQ5ipQmljun5pL9tZv2r0EBL/SUt93T52zHpd6VeixNV
Aotbpvzqvw0NEAKolmFXUvdjj7OXjuGXo58qykfTlnIdFk9ghr58lsbiBMxunNpmNGDzINQTc6n6
p5lcWmTXmpa7bNmBhZTZUEmm16X37O+kfnjoHJHY7O9R/o33I+neOCFMgQSPxeDOCdOX60yP2Low
vl4YTK26DOYG61h4xB0X8VWLOr496vozgn1WbsR/N9uIofNk3k8ETx/lixgVKjRmLrcPsiiaHO0c
vX9mJadvRMolLjyFB+EaMUAD/SPIg2toc/rpcP+/WyqaEkw0Nc2Ywc2BKUI9JalN0QK7JDfDiNsY
9WKKwJomV2MUOHz+/HIIkZtY/xZcXqwpMYz6+qUO1yQm5AVhnvxr2fZTVIwVuMLG6vFHoG7LUjpx
B1HdHJekMt2+tYUU+ZL5BftwgKs52POqMpU4X/p7ChPxv/KGycf2PDiPeM1uKkZtnO9j4PqYAccT
g/IjAIgQ4Lq3wy8fGto62gJlOiZVrSVj38yQ5a/S+3DZhuPm63Q6Rjplq32ebB8bM26PoCjjSBkK
A3iTGxK6LdsTjvqcidU5nn7pQXDH0He1DMO8Jc/R7YJZTBD7ye/vLVTLCtoGki5kdKrVKR4Dfl3S
UlU98SWNVHqh25Nj0RSq6d0YiCO+/cLwPOs0Y7GWVo8+nQl8W6CaokfKLHScp9kpoFwU8wS4sU58
M9+Ce64h1LNgpwhUycDcX5F8E74irvC0fiUOkoHEe10njoQkblrVwtXvKOIDQCLqtP6aj88NM3Uh
GlRxqj8VdIU0HzUm+vR3Sp6HK8ZXTl/ozHNAETvXmTP/mWqIglP58FD/Gt8VnZDxLl/VShJIddRP
VYyrF42trVoVdoCTtWpYrnEIdPpnWwICjOfgx8Aaghy1VDE/eHE5Um355gMtM2vij2SPrbIs9M20
hx/p9bQRBHd6pGIDMAL04tqTLVTJ2Zm0Ff94O2seax5xQmPe4XiEje5TTceB+tpiVhZKIXmykh8R
oOXYwl137Zc0ptIDrUXfNJRmnEi10r3g5USmDQhAfTLOdaQu7yZ+dGVDdXJOtdQnlZB9IQADB8ST
teuCM77+k4+ACatAHWmVQJY64iq/OyOTIvw3TYLH3uXSK1Q4lwt4AzTQTRazMTIWQ0CH+VAfqaF6
yugIFunmBMyuE3XRhwurKlBBbGQ7/xx+sLkdAoIHKelupVaqc1NPTRbpoguyeVafygaGe9HdhRHY
XEYBpSXhRkif7aR9QcXIiE4ojeFTHHf0PJJxivLE0iZSbCUA3vlP5+h6+sKfcq4jDLcsmj8qgNlg
rrAy89VriG2LcPK0mxgoj6uMSK+DU6+uwt5Oq07QZ/YkWyISb1uKntsXCVJ0rfeFJ/eJbZDPJIXP
/pOTsWWPaMrIGNwgt1eh7mMWg5iQjNbH69sawHybA+FoTeRHfO+A0u3EqxRNfqf1m5bH7fGtpDEP
VmP4gEaT4glK05rx5Ns+1tstQppiltA5EQUFYPQxew2Sj+dQaisY9yAWS8VU+Efc5AXDJAt+5OpX
E1KVIU8yVjDCycHh7tJhlf6DDGRz2BSfeQTSk/rJbKolhlpgELEQ33ltkIe4szhgvIX6L2kdpiNF
RG4ms75Zh5Z/hBaDsHAi52PYF8mY8PCnuAqG+dcGk6BHIVJ4t2eAfq1Z+g6VSibAhoR2tru+qYSd
D7GsPalYOAO89R3HDtZU7F0iAp9evXaiBs3cnKbzP7yjiKR60WPLMYtNFyBB+DKrTsomRfR1TLcs
l6jY7+Kg1tN3ROWLApadKvFdrCWbWEbAs1LBTUSE/2Sp6YPFxCyDexUoS2uHi1RfIclKTn/6Dfdv
6GJewwVcJ/TlTRV2HCDKIeUxtPa7imkbHc3mZCCwX+JAZzV+nlYESydgtzJ+mXIyWqFANi3TD55Y
oxBQw3JrVjsyq7agBPN9HgrozZfUHyZKFhLtdAA22B+gPY2wkR0DC0+zUeEHIxqmawG/ew7OOQ5o
iydgnhuT4+bfVxCqG/l1BCymeefqva7r5JwfBr6mZDCAOOuOYjkHcEwa6/Ax9XgK0caX/YFq+zR8
EOnTDOzHXXclKC1UwQlNpkJHtNhzIwIv/K4anoBlpFzUTbxZt7fX1tA70fsULPG2G3Vp/waT/QTA
IhcBsQeaXAUPNb8l6Yxkx7kcO0NkcHcLrGM7BfkVM4KPyzy1dt84DNAXcW5C1Kr9A0HB7b7atD2/
4ajQQHnGVdAWbe05yGlhwOn/AHKI8b/nq3CoDB3T+BN1P+rsTGWlBnf5j5TQvsxxQP5ax9ZpMFSF
prwAGPcfxiGI5lh/CBrMNmqrxoLnUJ4XoXuA2751kwM/Det8Uft7K4Teix+pPAStF97kgsoSs8A8
P2sRyiSz5nq4ERnoctN5/NSSefApjZkGEVUBWhGvBKA80GHwO4c+yuy+m4i9T5d4r+qVzC69hxkh
eKCKQm+n3p0s9nDlNfI7MN5Z6OZ+DPrNvw1mTkW+WNcyHgdxBDLIsLgH9TKVf9XjDS9kvojFER7D
BwzpfEOh6EgOmlepkcA5bkvuAdHtVRtJ7/64pCxjj3R+EFzwFQ59Br5FjjIJMFs+51Dtiqwd6Got
/tciXbLUSv1+hy1vG9Ww5xVeXLbbOH2PogQYno/hH9c1apWEqvOQuTt5i18xxqqqZ0N9LwXcm6He
TmQLQBu7VMbK/WdC+F3nr21aLscAejr/969J5zI8VJf3jzvRCabUKIo54i6RMojN7gCRfK1o9ZuA
F9kbhqD5LtDpV/3YEYkOfjNn9Guo8zHCWxlLVeliyA54zhBPfgWg674/jjWxANdRspfnYq952yvT
/kdlfslWrPTiHoXrzIEnGkkettvhhZsLKmvDaFNcSxzyD26yyuw6ovYuJfupxsUrz0PcNRcvgGqx
WlP8fnTWHXcAHI8FZzm+86M0mJOgyrcIK80V27HmZUuRrSy5u9ctMBfV/iaeAvyJLdCJq+zCESO6
xksyYQJP7pQAQAfqdBrwEtvI/QLfWTi15rq0qkJBH1WhSbSgBsj/QlWgRx9xPbxdcK7Y31jnjVaN
HcJA24+CJLhNY6jhCfeBTsAOdpcphRuoVulEWxf1lc7kCqYmCRgpeTs7aLfojs6DzXs6wzc7XeXB
0cUrnYUoCXdHT1mjLbarEcHiVIg6sCNzWFNwopIBfA+xmTrMVMwnPHwmIJE8dK3DhOEbrZTKHCCb
mQvZOKlhUjvgVoi3wfHUYmefNjL8bQ+C7aa+Lh4vEjTSaH03kZyAykHjaxytPpwKvzc9yXm+Pykd
HO2J/BUsP18ynVAPmjzIgzgyMJ1MxoF02QEapAme0I0dmQPVZCUEKMyVxNJ9fDOhMucfotldxC/y
hCRCe1YvYoN5YJy3b8d4JjTHCvifs3xGv8gNTq+JF5BVGZNZWhKkRPtX1yuNoxf8hn4blZ+6EuI6
mhPMI65h0cdNJr8YE1mDkkCe8qGiICOc6sexh8oEDNrBms/NTZdQH0mJm3k4KsYQdTr8bnzf3I8n
R9dRBiTEQILS2UUcbJEPn0wqEIfCS6KsdgcpIdGcCe+xX6PJP+B1RSCYmhSDCyRGGh/ZOGVIatVg
qtZq7ciWCcFNny1VMRRSdsNyt8ivzCahTc1npakswJnqkZSlTpaxVziUYhHDv/ujJgkJ2KSp+zzy
wLIkzGUET7m+RdFxFiwQFDjdr/b4o5yT2e/cTCu7QSwkkOO1BC76DxWx88+j4nHsZ603j/KgSQii
DPYRCaaTExGO0kOwO6JxMoYiNBVaP/9UYyMC/t1Z/e8vPRnL6/d3a340iJjwA7aev0iDtNcdGzFu
3C0VOJ1W1hGtVXffutjEjB1JxhksVeZF/g/ZcM3r1hKjScPzCduoOuU3doZCeGibFR7DtD8MmoJY
WclCuti2oogFFyd1alPYxp+IWkRn6Ef2XWGB6GEaKVGoCp3eTbJ3wd6eqfA3HM80je0kLbBeAlkq
6ix8mPfsRv+CukbknNMlhB69DoWKXMCZ14WKBfKTfETWQPoKG6khu680irJ6OEJ9PowGkJsm2x3Z
4fXo9Vt1x8IwpyFHHqcaoJivvtGc2IYu74Uk20APBYoK4REBh35c5R82spl2pIJHxn5Q+1u9y5DF
ap/RNmlVZFDXrE8ZUELaUlRIgAY9QMvYXsj6AcuXDbbIjVmDulUFSyi2/uCPWi6dYLVoc0RqTlYo
Ips2Dc8zRZ8NXZRWsVf/KIK0pXAuc0QWGAx+sN7Tx6cp2iierfhwC3kvCnID2XZHgWFVw1/daw0U
Ir1MG2G4O2DiR/fudfDacNTQdOIRmZ0292M2dcWYnAjH6LMuYc2F1L1hyF3nXtXHJxkGWY5eLKpi
8SDUdJNoxjUOYy+5emYOU4iPKgBfjvtsubOJLYSEsn5T/r5ejp8/p80EdIdldsG9l4/l6C6pOSVm
QIwy/lc9KIOQisC0r9fvEz38pVnOvv/no614eJjktRDIQMMoWw7xREmagVQnPVA5K5xytrL0DVmd
95tA2thS2Foj4rKPJu08Jhe9//EA9I661yoX/LPb0zY0aRH6OeaBdpFXY01AvGeJrP/4HfFHOTB+
Wt3qMgYB9u9vGNzc5c7aFStOcCyYIw6uMNfl63L946c60MxJOB3X6RR7OUFgpgwlYVgU8hI/Xk2h
9syZRIwuCcamknfdtirMoWjJrVy+pV07oz0rwLsHZ8B2ICkQSo2WmZp3uRPWyfHEZBdQRD17ZvYa
7mO6rnbImtvnuIbg5g+FCc5ENzTgFJh6o8/oP9iBVGfCNQ3hPTmrDj5MQxdUZC+l//0AoJBE+GHt
+2HyW5Y5CYRb/0zdiROH4XuUUb9/eeeer2lnRnuGsdoRUNwCF08CLYp1HTxpA2v2fzyIpg+QiWV5
mGx7lmRCkEeJrSq+WRmAQUMoleQteW0TnH9RHW/WMjIw1RUXPh7KOFeJFm0t2Cp9P+RaAh/aV8fD
5xjuBuWkR1tB5EQ6SabIZay7a9t6cJTlPUgFRR4PG1OM+Tcgb5cpKuzZbRENobq7+kXVf9fYqd8d
9bXzF6cC4FCoPJUcRVOn57NhH3cZ/6wAD+9yBN3BMbIigAofR+uISJv9knfq3LkBHrBPaubmZiGQ
Ja3BL7SEdTbwm/yJQh8vhAW/TJzX1TjVrkYj/8IiPcfZJZKmhRZpqj5Qm2pCTLJ4ZFOqQUR88BiX
fIvRvRce7oDlaj/Ti/CFK5uqO42BQ4H1Y+UQohpltNis96fVjj3T0SFsfoIwM3KImtGqaTsc5w/s
XDneXL8dvL8vuOKGWQi6p40qexrcDB1r5rnQaOidRAbpVv3jqM8RpofkkbB/Bhn4BE/vI2Yilby/
Xe+0Bderfy1V41MsipvtkzfjqhJvfnqX3I5fFIAP+xl9E2jLRUqgL7aD+6rrYYqsP8ASIyc5U4sd
B5mpet5La2xnG40fRtyLxz5pzOK4HfwgO0oiAFt9ZccdRnpLicIZgf6APNjQ2nmiNxS8DHmM+wxj
kkKvhxAHUB5FWOhaiPMtghOgi/vhaQWEjVmy9n+FLghFsnPgLcLdkrH9a5GMrLfW7lXiRg84qwz8
nHP6Q1AU3EYzfEpEkuRbDRL2lYctlO3TM8NruUh/dsHg2pXNQX9OULAD0MAFLRO0yKSAdLv5LvD8
STwDaUaTeXg1PaouuLvjPHSwUdK6EgoMXCd381+a6KkAQqc/s8Bj6aZuDXK+SiqbW0tW+W08CMEG
zgK7QlXbBHD7d56nNHAU4OaArpuliFLAYwcMpuqnB63/bvIaGvITf2NLcDk7P37ooznkV/8T+HJD
I6z/n973gxsMeuGotn587k65wHqyjyTX0GsQyvm0XBIhb54kqPwcNwRkJLJ7RquoZObTDG/io0yb
1uMal2QgrwXKnHF61UT9w6L061wPWJQRsN/g/tPYqvRXpTwyBQdRSP58OF0ClhNQXN4NfApbal3d
uxUva9Ry+tRnw5HxV7o0NvnsjjVsrQrkHjMcyQlIAHf4IgeoM1mtovNGzBiZmVIEkoHfXDdkq9MI
rTJJugzzOAQWqG3aZpxzX1+pxOpFSz6zXZ/yAsoY/saHb9urCJqJ6fHjC/4xN4YG6Cr2agW46ks5
LG4DbRV9Sx7HSHLXObLNZNOd17uJG8vn76apgCMoaiLWsFk4Z8bZduzGRuUZ/njs41PUJTRIOluU
bOg2qdIJROdWRO/pca588BbJvLa3BJ6UMSZRw4jTgjxY8+7wS/u3pZq6g/2zdnqw0Hox7lVrf4HZ
PWqIYrrxROR1hk3EfKOulyXOS/gtgs6uqQiwgbpQO7O/N+O6aGL2BsGw6PIjDk8GzB5Yu9WRU31f
6honi2ZxR28+wRIEdKNPku3IiLdjZiEtU5432IlvWF4voRLD0TzrtOLzvZ5FLb3Ryb0lTXGxfX3G
rBmc1GPNPXPvc15qyA4Uw+Pfcr9uTIBUGn88148ITrS0ewBRTmfG60KEzE6NKQsYBktr/fFAWr4+
ELgaqqJauym300/emtDoV/F1cd4++QbD+4s8Cv3Tpc3fiq1e/1JkO6i0Gjv4/7PidcbtS16r1VL3
izyEGjI1zioGkvw48zpwSKFAHnmX85ruFyig2HxNFY5Hg3FXXInFXTCFDuceJSpyTNUqz8UIEMUz
mKfi49joFTPH/3BqeWTwlQJZ1RYSNgthb+mVSdHXZaNjK8dh4NeOTFfGk3ZFgumfFBcxV77UYpal
+J0qOgnCEaG+kSlPSZgCv38TUNFVeqNrsuH4BPu1UQel5gAjUzQCgoyXcb8d3AyO2JICu03TlCwe
xAn4wYicZyocABlLlxLP0p17OZL7KaEe2K457FKSdKAAvyA7OnmvVafQsw2Omq5AzDUP16VMR979
tCEgRIgb2crXLJ0DaDC+NVD7VHErzXE0oqOoXyymBdCLRsLr+GrUKxIqicaPrJ+zf2VvQTOle7yS
GP6ePE3MBsU2Tuw5rO5EiDOdSRgr1XUd84kZ73Cn85afQvonHAqfW49fD34Lm5mfy6GVlhVz5Snu
Xshf4x/GyOjXJSID9IJeF0B9iOqu6RlnXpixQzl7VWE+wjGBHXYb8MOorVwm4VOYFC1EZgBwFfNv
yBJHniPr0QmnbnzSG70eVsAsm7iB4CgCqWtU6L5OLTtdtNt8M3YQhaBzTJFFVSiRYDTLJmYMTDxC
RSgNRaF/OJWlNU1+dHzINCqKmXGNsZgvlt1HpvT0m+cZVVUuIXT8OiU7+G/ObOBMu8NcvK/Povny
3zhKNvMaQ82dPmzxpCu10Y6JxXIT8fbs17XZL3iq8N3fjp6l+Eak4m+gzGjNTHdtOcQQaqGD3jrP
UrkS72GujjoTAyGp306tWU4CInivFrVlg1lh4F0x7hQGbvY2pHD/sY1iINQPbcZ3RZgerERfOrMr
V3YH8AWotqma3y54kgfzhgDcQKjqwvzrw5Jp3WON1FW9039ohytlzT35iae7EADSOSEhEzXVW6+W
MxWELm8X70cWLmBsqjg0gsDYjAeBZwjoVx8D0GS2TvasO4pnOFojHpDnAr53CVKdjls3oL0QV0MG
UyzC82A6TooDznHV6UBUP57/GMO99XtJD8Y+7hEr8xcaEvKKltv/hyBJUv1H3BjSHiakr5fKzpew
6b9Ow/Esix1BRmnxuj1W+Q2fHV5biUJLL3JzGIBAr6svd4FW6/uZMsMpXn9gCf7usXhiDh883EYN
lw8njVQwdTxtkK3l0GOyUzplirsMHMrwcGxTWDKQqBCyODVDh68NBNMqwcl9RbX+MP+0e1WzYhhh
ju6S51NGnonWGJblzAp8FHEY1nfa5jLiMyarYtD7qySAzGd9FIgUzj2T1WFLMnIoUgZX9GyLYEVE
YfUH2bSE/xiiyb5Je3wYo60/ToZ+antVYDrB+g11bYN0Utzcgc5+bbOpZDnVwkLMeKLbRnkKl+iZ
ZerPaxzb2jldfefxa/F4JZ83foBbDGLO5w2SFcGO4KV48ltWQUDE83f/3+yCLBILGVBBxXa3X7b8
bB58wyh3W+NM9Tj3VylpMD8R9z6aXxXGy1ol8DVI4pi3wDXAc4NeGtedcXb+4OTv7YFdFcdp+VHb
jq8cImJ7EcBSavUGwg+63xzc/X/TblupqOH6JcoNEcS9fozCRcEpIXU6bMiBxpERf1ru4IrmdUA5
WAUnP5y6Mia0f9roap2m+d62pY1gA7P6llIDxSwjWm2Iz3NBuFOsz/n9fCM+q9tRt9burkyIF77E
B8xaBViKRlo01X3A1O0WQUuyJ/jBNVoajLuYASSabOSltap9TQuiY6k5opXmRWbNJ29q9TiYvQ8f
AJBifXd8FbcGGnAUFJhHsEI1XZI2CbujfYPcu0aYJhfRJ7yNwLoz0lcGt79x4EIo0xAQpwg8Xq05
ZsQ8QXJaW/hyMZZZMrdZl2ks7vnIoR3J61ACilGvXS+dxPxaWLZFAqsgJ1V8DKoBoMsSx1CwgTyC
gKVwj0HVJqtoGjY+jWcSUsqP5sZbexG5oPPeWfC8i3x4f9dNSjMI6amOFGP4d+leLfUWRpgNDP4g
+QpcVR5fYwK79seRfDItI4S3WG7qSSBDIaGyMRGIMRIjEpnMggX71pNzjWlCqQ7eNoiv71Q3lgUB
r3WUY2qQ7d80M6Pp9HiEoUSwafnuqQV35zshn24AsxKyiD9395CnUe0EHrLzWotnGzT/VShy65QO
y2JmBneCPAHyo1x/yq5/Jd3oVzxOlerBH3Ru0mIjHjqsppWSRsEACCyLDO3HOphOnjC7nDvCE314
psexkvMs2IOV1Uf5A+xm7nSCIUJ2P6/fdvVudHsapDaY58iVcRM7TahNgn6h+VtX4cVp5EWtaMkT
D/R1cM0m3uuN8T3V4u2AWNEs+HgtIf1W+YBKYtFHCQDNAHij6gZ5S5xWHu8v+6WnpN+NL2ENsf4z
njrA1PKDEgMRG3LlRFu+b0tsfzv+H/ogDaLcmdqd9NScUKmxbP4w0my7a2ptBIrpOEDU/VOas4Qh
wbCUcrNrDPvBFWwl8Iy9qrW1HCokWji14yZTMuoasQNOIFj4FR1z6qDLh0JwEGMygNA1xP/Ja1eg
/wdHsZTcKTmCLjPX3FXqgYnAtwq2YQLV9gYKq7BwqGxlKjC5tZJV921bJQ1WJGyi4XV8e7MZdbFs
0bx66dB21xkoWxVYuFNlXfZEwLxAthbW3yWM4Sq1O8u9mT4yKdzz90xHsCRZLDa8CF4OZ1gF9y/2
75l/9W7jq0OtgYrYbt/pYTnjl2kNxEkmw9Mp591dMDv301WXGfpQriW60dPJWRyNDVPCXln7nT58
2wJm8HS5VcvvPj+KOmHp3wo7d+xynCwauC/7UAq3vj9gNTV402Tfyaj1KKI4QyCM+l7dQ24LK/py
4ARegNvOyr17xc2QdoQerUIVcClMW8CRcRaYdWCtNdkWv/Gwedxs3YSyRl1Wy6oHnr4SJvStQOm9
tQvfMJtov5P9KrTfMOrVT2tmtT1j2Fk/9158mwzwxssnw4G9872Xad5JPDfoXHlEpTn1E7jnvLEi
6H5Xcz/2x7+RRiprRMeeXkeJFFuKRR6hejGn6Lp8x6Oov1NASykMiTPloUGph+JQVxcKrP3prbgF
KtIyFCy9I/ErTHo4AMEjQhGBrB6ZpsT/be9SP/Nb+/3Vmuj8Oa20/ebdWIs61G72rqQAzIK4i5Lf
3zdVL+TXuwzbuiYTHVBfn5bJgeEpDxvdtQoR64OPX4C3Blhm96snPDaZCB3C6jEd6iiJZb3G0Zl7
SpYeUjE/ooCHZ/yU/9MkdLLLBoWzKkGtpeLuCVcQ7Y++eiGz0U5pYbulRTyyV9FrhO6hsNcoi0Nh
s34+LOCyPIm2kLlMxNi0X7O8pnEnjRkQlevIRGiluUkChC0bU6hEMC2qRtK1F8YDgECWuC1OB6Ng
b8hlgnpHGozdYYPIy1BS3gXTA2H7iIGZuEizYF4xWu43c0bu5sJjbJ85QhHdZzvWNmDoYdQc/LER
E4HLnrKmk2oil1uN1EDsjLxnBhaZ+Q2MF6revrhG21LtD+qHhD0BIP84jHL+EjpEnrG8ly3jEXQd
0mDUFtKPTmYq74OHtmV8Yd3n9F1bqv8/NtDLFkfo5au/lXU0HBMaKEyMbrjF8fvnCXUyBeZsce7a
lnOoLGotHYu0T/lqrgWymW8izMZ7kXrbFoOitrlvFK4ZdYA8zEnLL0Gfsig4M9IiKRC8QQ2b6TXe
LRDq4tNOnVDvDTmm0KM+f/6vOzYOBF//lf293J8epAL7tjr43XOSu7hpQeJKcg9B0RgJjYz3kpNJ
sxIP9CIPNYc+qnhod05e9sHWz91lqSSC4xmKjzhSVDyREtR8Xui+eULG75hGBhd5i4vYDJIJ1XxY
6Nqzs0xCNOz0oLIwhlIPCY/ewEuEBigzLzQSflXnewbuFy4XU6jU8iPrs/XJv3ZRRjzEt3gkxSjh
wHKimR7qfoXVuEpamuacOsb5dtbKLRXdi2DJ0pRn49qkPAYvGzVCIVDUKYJOWbYDofVwsSrHxltN
jFEhDHaWsHNevxpena/W51VxOQ22VvbWjvah4YkPV9QSagU/Dv7tu4bZiMIMWCW0GX+BE4hk6WbH
qqdYIVQgmX8vligl5WBglItTEOqp3WkH4Vf5A3ix8FQ+IHY40CuGACv+MybiU1v0DMpY1MLbPsNO
+WXFvdJmHi7otjy4Q1QLoHRHHG9DfrSZDUaJQkVAmyDg55+4LkHxeVJOzeCc5MBBULCnxwnKUhYO
Tcwr6OC1Xp/vKk4jpoC4FUIph+xsO76jSFpRi++fa0phcUcSnVDUq6CFVevV+/ui3k5JRQkEiZzJ
m3B3pfPhBS6emlD5wAxJ2QzVCWRuyWdJAW0XtWJ1lEXFSfJEhTpygApXvq01O2Ld6lu9QCVoFe5Q
rHJP1bFiUC+RvEQ8wnzLRLJDOSaDEDQVgMyob+lALTOFBTvchOH/3y/DML2f5wijzkhR6fC/kG9o
QgGBRV2V1U0eOk9OefwP1amrkXueuar4wSwJpExCdsBCSLHnqMeKDVhxehKBSH9UOrQGJbupc4AV
lexphr1veuFAND0CV8fz8BQlCwAA9kIyjRfVmnq0DoL/JACL4I0KJr8LKGJd6sNLBf9KkwthtCxI
5Ed/wI5NgRIDQZqlMySyIIJZcx1vhYRpNO7akziOZJYIODh6Df2F0ESmYIGypkfI/n59Xeohq1mv
aizyfHQX9VHUszGZI/LT71DEKdWkIcFrlIK/d+zNZ7j0Re0ODX4BeSUquPWZBHHR8V05Qao/7DrZ
pvV2GiMLRtKzSwMxR4TkdmNMWKWVSRx6tXAhccN8DbDCN3HkMO7SlrjJcyj17RBgqVgnPTNN1PJq
j62xO6OnBwk0/iSA+js5K4TKXoSaT2OXP2IkoGLZsG5Lh0qzJ6mXUKEZoQdQUyLQHJD+VpPFz4fp
HvcR/znx/haKzmM7aSUHwsFx7IZjlVJZmxGd7mbQvwdTO5fIRclbSlNxWnAj4vTfZKCFEVlCoRse
iDI3Nrmz2l9q8jUWrPLdq0pPOZ4zqLMH6BRtxYigeVGK5zDzZniGrrMew3BZ0+5NUIwpjYDmY6QW
TRdyRunw5IUXSIc7Jq7oYvcYwipg5bkE2M1TyONyaP8EtWEfGD2q22L5cd+o3P614Frbw1lNbPb0
KdI1r8zbjOuh6oWgmTwT0sS+0ltDLvHCDSu8mG2TQU+yeaALeGVDuaX/bPLMUwSg5N3wa57Ckk+d
vmmYsiZOY4lgnPauShnG+maCkkFrhhD2Iu2uw13qTWXTAIOBeoWtPigjfyGXi7K+T2HwEE9xUZfU
iKZ26y4HjS/11gpH7GI4Ct5sxnUgy6zkAyBerfHVHKGkOMftQEIRyNlAMQ4OdnVeUTSNjhCD5Wl/
gg8SzVy0MvWyGOWZwG2uBxDzzNeOCTugND7sTuIdH4kVaOh00PyCbOb5/nYspAoBMvSPJf/ZUXgN
wrEbas8wCX1XvrSn0crEiyWjcLFmf1eEoFF6ahO+NKiTIZy1ET2W7IbvzmOW/sOuO88gdQ6Qt/Pr
n1PnMSSwTkb3BMNoO1FMUvXyrQQNY0HvbhaL2omq1O/shyJwId7F8Amr67mBRwUSf0hZtzkL/mMz
jiumk7ThMRiIwTGSwY5wAEex8JoAU4f/h2YtwtHyYyDlPNZ58AfkI2saAkT5dS6e6+VEEB9Garji
R+zTOryI96ZzGALPPzPpq1+MS4sAONTWsUSG0dSTrtlgR/1Xp/5Cr3OC/tzGiUKBp7dSSGAuwFau
8CFirzQvbh07ywckHGLG/tWrXNxUhjjUro6cIv3UpdoZpd+mGS1WBn0zdzHP4Cj2gjSqT9IOEPST
7gsBMgntjeZqEyMkA89KM4KwkTuYCVFgt8oZcS1Y+stwZ4/3ekE+GvpaWB+E9tLrfF9hYI/hdvbb
7NIj23gU4jRcLveOqHx8P6gMUYiax5d4tbqaxJBK1cpJMGM3tWzLec0bc212piDaz2rj3GdweczD
3z6z+f2kb3ykS2v16hrE7mBYGnm7QnieNgT6fmeOsGeZNvcviZyuKFfxa0dkgnIA5LKzte3pVKXw
kDFWMHvhjO8H/OZhB6QrAVTVbCyw88M9O1U7Z2qpGANVZbBw94utd5YUKYRxUsXQSYvAKLJYKcj6
BC3smzmv8rLfyvZY/oOjFtWXWkTVzkNEIVQLKVyuDAMmNAfn7WopCNiNgEtwoNbDbaToXbvd7IIG
MAOculWiBOp+OlfzFKOCp/GF+9He5V+PNGR861SKPq2LLhTfSYRKF2dXhERtk49aXF1+QUCkI/hN
Z2L/M8xt3LqbWbhY3gWP4ylzHiDe1pgXngB0OCqcQ436t11x4PY/aoKJoCIAt4ME723lwy+l9OWS
OpBTCwA4eTbmwjkelDgF6Hnp70vZ+RmcE3BkcD3X4Mb2tMAtmwKdnSm2X03vBfo6/HsLgEuwgf1b
N9hfyW+OdeXheYTwLXbZ+J3FEpilhCdU4Ffr918AiL/+67cSbFIgSWmqQmghjMJNafx4wh7HD03W
NkfjV0eBPOSUWF8gbCYNIaW+mIX3okgCIxgwalG4P4zgrSUBeq0UqhPl4K73NivrwwPEFaibpMB+
bn8SqTLvTlUOt/EqXRBkqbjE2RhxNOEu/V0JOOHkXaeiJPDVhvDJC3EZ7AhnGsCMsAmDnbHaEh0f
EN/CKWvmw314QY4lwEXBw7k/jIqB3Jsh22z7n5bR4aAJeP5/3e9bUZ6jcgo4kdYz74yB4XTGV0Ay
VJX8hVixohfLg4GYywO/kpB8QVmbeW/pM+TEh427Et/fQe1KdHoecKAZ/dVUaHEuQD4fNMdWFbXs
4Rchf6UmRQYam8bp6ij23n/N4EJ1s0mrwURGWdiz2I1AMLjgzS+POki/iUr9lrW+KMPD9xCeLxRb
KYFZ3AVQZmrPYpLXDY6W6+hi7/fFYskklfwGaamFGT6O+INCriXQvVYRmuYMFWUkDyGSQn2d67hf
as3AENqjM+0ViN8nKoFYn9a4YV7Ii2JwEbhetMwAgqiC0FS6PBWpnhceiuDxC1gWAfJz7NoVkiiN
CYU4eMrYqiauSS6w0ozgcjUU81yHLwsup13hVupbYNxHdEe1VaQ8hwBquc6pAzZ1HKAD9mLnYm7S
QmlgJogZoynaOPKpQfcm9PcMkHfsG/5xwv7c3rF0FscNINh8HiKVGhARxq4KyuL5wn53LgM1CKKo
HgVuOTQZxSv/h52kVD9qZ8r9Sl6ik2Qwdosto2+O9KC270Rj4Q9dIWXNL1N5mKplhrfjlr+kjyEA
PvQ+b9x8Dg/th/GaigQIo5XnJuEAMmxUsgq5AGozvSa4WDSrFrz8bU60h018G05pb3s1JXBLkx8X
B4YtdSWMtsp6dr9yhzuEeHrJL5059pBIw7n2QFE2xF8dXf1SaSei4GhivPXYVBfAviXJG8I2VlPB
+YzahYOfmml857E3r4a5lLBXkTKLmYAE278ywnkLEZiDc7nAZif8AfPq9sW4pQIY3mMj+QmS92gT
3E9OKiUo2OnJKuFcFfYT3SrMXKjbkMIn+hIN6u0mNZVojoKKozdVgFmtFlWWyicXWayt8eaqmX3t
3KGURFjyeVn6JoDBGQfCYGCKShgPIDR3+yovCtnpwmHVPWjqP6BYv6FEl7pV/LyqAL4xIztnl55x
gMxogOgTWM1CeI4tmOxg/aZuLAhtR1ramIE2sHo0KmvxhKcp7Fy6yv+8hQQwbrq03LBstIHNRfxy
IevU1ndhFqlYVhLeU7izKQ2YKJD5FyEH3s70jY0IhhWMNbZxoML/AnT0jCC2nWZW7Hk5TJHp09ya
2JJWF9EiFhpe4heteRSxwuFQQtQyhPgvlXmrCylSSiqG7B3RKkhuR98U1F0XQ+LtNpmPYss4nJNT
CiPwL57jcfFUT590l3lUfGrh7fgvWR9BE/9xjgzWVaYRMGwi6RPR91XtJAhGCmq0wWU7LwKYW5zk
L/3RnTGtaaw+xXt6iX3OrtEvI+IyxAoaZyU/No0R989MYXaYFopEe8LyVmeyvxsCEbufwZeGXCvk
MG58ZygGCojD2W6j9nvQjXBgaX4xep9UzqLJSw5y6GR6W3XV1zC8K5Ce7227jNiagFF9oFLCUMmc
z6xceewc4o0dZC7rNosuE3Kx+qPHRtQu83993dxaD8pE2fLSynxdHYI39ItQrdMTfklfxyk3lxjP
tA+k01TcvYZJHzJcrljKG3DIWttpKZOzsBc8FqJ1UaxDXffzP94SvNvQbxeVWMZ4JmuCtZ5SdqmU
FeBGlfIN8Uad6uf2Oi6ugR+obK7rMV5VCePsqdnUBevFBeJclkfV/6gJBoLWb7CIOmufGmYwKYc1
cG8kxxTg9DZR4Tdh0nrusLcw20srQ2g5Z63Kc4QjMIao5SiOf6mH0v9bYrA3m/0QIFcgPn4INg+b
4MtU2ypPI7nBFtZ05yjN8gFYenL9xyt5u2zaBtVSgCQyIOV2enkOjQ9JfwjRQSYZYhvFO4xKlsE6
C4CFjmzNi4wPblBsG3n19FzEO1sTTj6s7jo3S8VGt7W2/xUnJky5fzxA2sZr509VAMx3FljSt3P+
dqpgNKhRA4/TJ8NQZOnVXuQKnVTCTyE8yi11MWJZKWDp4e2SqnsiOsKxE4ZdYD5rtisg+2cMz462
5Uhesen7SMmU2XYQ2l15rd2YJTuYe0F6/fLB89k9+7Po+brKRmI7s+1BxIqjWb7P3rzOqylAik5A
kBnexFmCudj6+pOEiyyFIX+30Vv4kRRkarbKxwFfJkNP2FgCTrGHDjBcw/Hb2mvKfX7jfGvfTsze
VPlFLn5Ihxoe/ZIsJwpyochJm9b6pdE4kkkjGFFUq2tomidFB4quNw7xk93yC+RNAABiD1ogYv51
l9OefgFm765Cmo7BhqFOKhqvog6s3M34kopiFsxdWGwqGDws97NXP/ljy+Bei6KTPRxkZHa5c1Es
+wBxR7gu+Zajn/DVczTB5bRnUJXe442U03bPTfhTPJpud2o6o8WztANOEKNsNQdI1ICQIhuJSoPn
O+UeyuqtG87Qut2GQhS/f91gEG8saSY+oCkZ8d6+DMU65ckDu2LlH7CGHfwAQyvzglsFzF7l6l1t
pL2MJ8CcIG6txTWTuUdGbxoIW1FnEwZTg8qZXC0kiN2rfldmyFsYNfuPC2YRVu/S4QwTF/cbgT0+
+a2sIBAyakk96azZArlN0LjJTFz0fFB3F6ZEvW1yM86ssX9vU+kTOert4JWpuUWT6Wr68PaF5k6T
/Mt/TzAplcaTpgdsbGg8OPcIF3GV1u0n/vXAcTs95yveSS8ZAexzZ6cTRpSvw3Ls0uGcaeuoEX42
eL3dXB91qAlu3Jkj/gFJ95jRmzWy3O81PpEILNuxF3Vy1hjAWy+Grw7mWFvILu7CkVSOMsSO0ckP
OlxfRFcSdL+3hsBAPdZpaN0+7a+y/yM9ZiPWP5YLpzgT66hfkY4Iw5JXcmF7fXcdwWNVAXOHSsjM
StoYFH9Dv2NEK78wpDKV5fobmf7S2LnF1lCo0ar6Y29nYoxEcTt/cq1bv9Oqzhc9sGURGqxC8hR4
8LnGuIuAKXdBqTakljb8kBijQCe65tXnXhQHa77gl2iKw8xAndEuw+mitopPbz6ASTdaDBxHszM5
98yrt6kW11Hr7SIHJai8j88I9tPBPjYLNM8DIwqkVlCZwcWWzi77S+0hbKzu8dFtRhyu5S+15zfD
cT5KBI5AOopNhc4b4/xCjzfkAe2pnjklOqsyjWPHesIk+4JfXEPynL9CpdHbxgXTklRlZ5w3OOLq
Dr+GwYX50Ot5vOQGnScti42ndG4MWOU5ifFHI8cDprz9OoeKIhz1i11Nhadj9fjfuAtaDLW/1G/Q
MMc2Cg0aliAUa/NtXsfep2JsjXYnCy85nEi8rksACyTTEcObeuXfFp9hDrUvNbad1wrmVKE8jYz3
T5MWjdn0TMY+0ZZYjV9sopwSJwU1erBIPFmQ3/lACtKHzFcRDztwns88IksGAGSoV3WgsJrBOSl+
7/ov5wCiPRNl3+Fw2TkM5D5tlGYZ9q+waWlxH1xPv0KAsdgfTYrvON3PDDKa655qa7QMbzqfM999
5XwEgrO+BY6V7xjDWNJrwq6jChDQMkqG6LQoGTaU5/cc/0CAp+yXuqmpitMvMXXlqpVhHypxyX39
VqK/jznytInsFuN5duTSziq2KkMwbWFGhl7FertRffYvECY2SALIUL6huEHGHxByyYzCe7Z9R+6p
ndrIq8I4xbO5p0iS6/clzJLEz6vFQ1n5Fkn+gd/AGY549XL4tqGLWVONyOSw1BEt4e37TGUxWxFw
0hGaBTUVdsohTnzxhlhF7vCdZDTTgUtKMIXOLxdPtYJ8jmepLjKJBphzRWIlOCku0/yAHmJZ/PAB
vuri4sQapcWfGtRJ/mj19HYN2nHZCM1gv/oYr+VM/BBeWb4IOWLZF530GafEDin1b3UxaTCGR3xW
kk70GZ8mxFkbVFXp3vXdP14xXXlpp+IR06INmHEZ/WQT2YF0nH8o3NU2ELiW7bexDS18ZSJn0tV7
fwoibYGIJuP3U5msS8tcS1RXnrl1AVg6FHBqQ+SDvB26V7XE7JmOaL4odh0ikY6rAe08ECz328fr
XARaauhkZ3mP/U/Sf1IoE11kEGyqo3bSnSmQYXq6wxlZLfgwJProbaMoIjxtaVhONWr7sKYiP+7a
g48yuyIMATdcT/SBX88ZUzVFPvKgdxA5IbRCs59iLtn0SRS9sSLKB6M4PE+XstEiiQXbvSyKDi4j
AWvYzlIo7x44jWBMk46XR54n6NI9siVyog0R8imE0ATRJfqD2vmstKfKhJHELesW2IlXxFr19xx6
jPvlzp72uxDgDJOXNIBOPXwqnVLfisNWGO2YK8wjjXcwFx8ac8dDalJcOAk4owBqgKdj8S1cUDEt
2pr1hnYNhQJmN1Ti4fBQv4wiMyj9kdxYLjRXoACEisSb34ebo9Nd2bbKCqchFaPGTjm0DPFzbJqC
iieBKrRA5hleY+ndxr9FngY6kJb6RqlEPnVRUNj9s5tfiAFD0ayUHrNv5lLfGDmhw1biZkr7Qps+
8+rOZRjOzIcrgd2WVy8ptKlpZMEhtxeXpjiAMm4FOs88nS7CjaJL2htCo5186fy6ztknRB+3q8VX
QMjV8kMRf3JsSJVuSDpom9NRUtktzLlSV1//qDa54JVsWRMmob3urJSgMad+WNGeZtttTBhqXDR2
KLa77XLi5jQOPp+XAI+aS0MWM2fYx/sFTwJy4BH82OUhemo8MWm/AMc986gzH76SC0pvyGOhZ0K7
jXOCCBx1MYrSTQtm2jjagkh77SQMXAISg89cn6vjjU9oeumNHlYq7i84usuErnO1nHNNDw5sorr1
V+5S7K9XAjdDVkj97/IRAnNrwstL31i3DDqxmyIPXGd/qr/r37vjk8g3Rhc4Kc5LH+aElz03CVER
bnS0gyg9jYHmW2YRCoY1XFxT8tVWmyO6aXVPx+1ZPSUC+Ik9LRyahUx6bc8yZAwt/wfAqN9C9bK0
1HrlrFgrXysD9nmzn6jAqJPvBDFQafz3HNpMzlhOFrHdeGEEsJXm5v4SgbFoV2ifwYCba+UPWbQc
9STgI0+PbS8mvNdGppIqNaK5CE8JH77fVtLMmMcpSHb2iDhzuYZN11a4jUS4u1S1voqtUpzv5cs4
p+GBM3zcPq8G2aPo8iqM/VgaxoF3Urrnj7/iL7Obe//E0LDTUHrA3NTuN1KlMOMTmRBK9nRlLj+9
EA+g0cuN5QH6+ficjnikKEVZymh8GVL6Q/5IpTyWdmAFx0ay7csbnEFW8Wp/TlaaiqJqwE8k94qz
IDFvZ8eXp3S9xAkFWOCM+uZfeDj423LzH1OWejI2ybQGjt/vYqXxqRZiwOrwUh2M0hTO42Dx/Sl6
4VIvIxfjEb2FHwOnu+h8jaImbP8jfq/n1/NJsSLeLwmkTIIE6yF9phiVH3L9OOXlp0h844cLg6NU
tOE7Z+glyp5SsdnKWS4exK3fGQPNqAFy7PP5EG0YrCraqqoe1zk9EhBz7v2DPC27YzgwW6Qw5i6x
LtlgrL/fj7lz1P9y+qsbMj9UvtBIpQf+Ce93r4GEzW3+9d+d1V5ShpVNqODJWmEW5OIr7itmF3Ke
OEIcpFeY4STppgrdKbV8jD+s/oKn0stBt8CjOELzGptnTy81jSni1Y69TlrFAYkIwgVQM3xiwdOZ
lOK9dU6yDFY5+QEHETDD6662CmbLYsln8XmwoI3hU42tP0h8N5FFdPMkwv+N65MUaX4N8wPPW5TC
FXDvpFRJ4HdOTPcE7ZLEOtgSGq+3ddplPEjQWDWsqU3OgQxwr/hjUFyQtFrNdMuXrbyLeD4LTWoV
cFcgco/XEjnBbzqhFuYgRNS53vlrwpVeaZPntDqutxSN/xw0jsFAXn827uxutwLbT9ZOwA/bJB7I
6/0THUN9vhrKVy/wQH/4gX67dgsK24Ka+P45pg+MHIbAAwc0nE6/Hxdj1CyBYnSIw85LM7b5pXkX
VD0GFhtOT3r40ydCHRvixyglBsfcXHd+i6kq5nJ9zHfIJFAjpSvDXM/qGc2mNGNFz/Qfp8K2GknQ
1gJOEAgaUQIUntwNz3xugTKExS2plHVxenkwWm539tZQkT545/NJl5DpxcuhhjOXLZSi3/v8N6gX
Hb+I5SoGcS3phNq+nRF789RZzZ6m6YzCdpap9MKH/HkMxY2JVO3LKuDyVhgMyCaTAWOBy74MHDP8
5qhunrf+SIMXSeCTQkMjtkysxlTVCorG6wXVs3YvE20LEfNTBWPa7wedzflZLt1Db9G3IEVYRQp0
lq2Lia4CThZLZxWXt6KjX5oXqAV6C7Eo15vW4OJVgnoUb1FCytYn5wKDPuyUUVhGTofWYbCo4nqr
AgHjUSlFIKhQelJwXkud12h9s8YT/gDqy/znu5/qRR7Q+gNY6ewyh9GlZBhxAvsKJBHxnNakmO3y
8Z6PerxH0XCK71TX48ZMI7vOWE0ka/rRayBCmy3Ov/RLzdPQMvDp4RhyTfD9CZjmG5zbUiYhz64O
zQXwgU37S4AjgifU/S7b5/v95GeCQBVVV7i7pUlhbBynlWsVzBxM6Ur9HlyzpHKEthorUIMthUZV
Y0OSTNn1ahv44j97MOi3W7+2RILqwtyf8qZfx71MZjO7PBFXcrBAkpYsl8Z6iibMZ7Jz8sI7ubey
yuwmKr34qjLCWW0iBvm+mbZUi6K8njYnR5C4Xx39zykJAK5T8B4TdJ/+B1yDcmXi4cbdUD0j9MJQ
imsNMTLiNuCaoedxOD6ylhyI43NZu3rza9OnPLT4U+98XpVuTIq08NX8ObS6TK0FtWkJ6yYxu+oF
RYKWoFqsmXk43UB/+R+xwWrqBKb8G7d+hdHX71klbON2bMYWTV+QAtOpm6iKpQ6Aau9aiZk6QncG
HhNQRzR4X8ac/VW5NNbydCcbjUh+5eyBYnmzFMMy6Nt3BFNUnd6Re6ODRdkaOFV7DONJdWoBL3v2
7oXYH2bbTYdWdfNFgNrXe8ySpY/uqsfjGF+86H9NCbqnWVwQ3DxSG/hy68EwuMZqYBJoMwUNtVjo
8AnSEnHNDMtJXNchJchH/oA29iHMMfqqH7+jpGpgUDLcxMtMZ4w4wfmcHTEFaef6iAUafzEFyH3m
rA2+ygEkQJ7e/uT8+/h5q7St00bkUw18ngN7xhCGP1vd9fjCPkm724XMu58i0FbrIHywMI1dtnCC
WTWqfM8KjltocOMApZempLlesqI7nWR4Pva6BmJy7F7okAw1CkM2Ak3z4c2fRUDHuLrQvUtP5U8+
o93Kvx7EPvW2viSEhBMwfw/LnJivXcJu7PKFzwKoDGhn6hQVM0O1xQ/p611E3aCxDSjrvvUU0Drj
PnmRHfuYh3Pvh6/yDgwn4AtZt5OW9gYTwUvMS0FbvV2/ayDEZYq6m5+ti49jJ84M4Re8GgPwBRZZ
mfddkIV1JO4SJczzWTVPTZCFkH/VxovnkcWB0tluxIUAlvfMS9VUdWCJy5n8XRHXFKO8U0JGKLi+
bIuwAvRwnDysHLurm+WfGmvCM8bhJaQHjFSBiNE7xRq8qIh+iSZUfID9gb+llvxZQPrf7iclogFC
2BGFv47BlY4nMXquOuesRjZ/giMBXIf92E8kx/xmfVajcSfwIP2TMG38+aCmbax/TT76CMNlqBOt
HRDwxT7tQ8RMFRtPiuBbedg0qwSRjESAygCN0BFnoSzY4OgE5wESyM4OzUTfdsOci42FAq7uEzbv
EzSheB3FtcIZfv/3uAW+dDLOT8SPTcVlm6E4aZlipIaGNaIpjGlfWh30hgUhD9PENEzsImp596Xa
It5deFijhorzwdhuPy+a+dQlcTkeXvnagEJziVjxwBam3ZMlCYyJxFMopHmO984TqhWTzb8JGsIv
hCFahEKxl/Rb2s2buerL6mYK3a9ZvPxLNYN99KzKhkDv5EIrVUP5d2fFSqPEQxR7wcjICF/hcsD1
WSS4fgc99CeUKAeGnZBnbHTHeLAYt9WO7Flfjl9Jw7An1xVhL95+YNsUcov831KuG2Ic2AA9NgK9
oxOl5opGom7WIHZZ8cnZbbu5jZVEE3uRel9YUTSUx4wAtcy9bysxM2FTO96BqrhSAH31ZPuCJCTb
YD89UXvtcr+iGMs8a+/t+FY5E0lsnvb2R7R6wFZJQkdVH78CGuD/PmFBYxWBhmaXyXSjmm/mhRad
rNxPzqqe8FILrw+qe+ltUJTOcDqo7aDFC6Dn+ha3tpWSGrR/Xsak9VXHVvx0Lp5HGFk0vJ5s1gou
DYeKq/DBoITG+buUj/f2GbCQrAzlplprB66YbuHx6lSwy58EpViFhm98ddOReYlAn6s3m7FB+BIO
r+P3uFnoCm95Yn//D0cHQ/CshVa79ooewNSuEgDE/F5a+5fAaV0CzjZw2yqWdm1fjgmGWNAAYLGM
kHBld84vDvtXybSIZCcK9sgF4ghXllmb20itRdWZv2FXSuGQdlN4BORX8c1Q3KqH8kZgkfKgo0pj
SpWIqdVOBkKlLxxT3LIqavJS2Z9ROpA5G2039Z+xpym/McPfloewcuy39KTIgQ/FXsMeShdrk2Z9
6SHx4XgCPrjaXPNaFU/YgQiXwkbrmV87M36rw9i0wGWbv3lNjHrfGkzzHsP1gkbjWaajpEciu6V/
mhA2dm/lNM8MaCWkBL1h7TrhVqEdlOQFWXoREL1yQ24ES9RfYvu1yRVRnV/A3ysYYzrvpqHzGw9X
lHf3g1bO/mNmn0aFh2zka5GQ6Rx4CrP6TmZf7Y5zCqYoz3BVIko9X3Lf18iw58w75SM8JYAD6OKO
1CYdo2abbENpUPL77HHgHuSfyv+fVt8t5kN/K3ZcA0cHGGmyTVMb9fX0+ZqQsZnflyGG51gjR9OU
8SOyQfTV0GhHwRkRD2B1tGH0ouuGA633nXgA9ULoUJWqHMcSQieXfAFLQbnjsnDysVensxsfm+V7
f1qu3B3wz0GFIE29iAvc71sIMLAR3vCGmbKjCcVc+4nLnnQVymftNeQ8iaFUDdt1Ed2x6ePNS7Ve
BoZUI1KtJrW+d0ipUSJDEUX+ije8wqtImi5vbOpuAYrHg6S3ZX8h/BtewEg0AQWSTYsU+g1oU1AE
qzc5xyr1E0btkIkYSSmZARg9jwgvKpXOJriHvuWf2UC/TQjTg7nYoLl1ufm5jilaMIX2SlDXtdl0
UtJaiL3pJg/nnvHJjJdAWC7YbBUroNb+Lgd5Q84r1sKXqCpO0StZI1m2gORSrxtnfngvgyPFHWEN
qB+BFQ8sqy/OsTbQF9OKax9aMNCI7OGedd4K9W2WZ5yrvL5V/Zx91REdO9fe6Ahq6bK5MDpoBVfv
NlwcFkbsov+gkbNzL0OnIATdxfxU7fpBcICbW2ZN9TIlU/6ub6gaAsZleCth/tatRI6oQMmOPcUR
E8fA3/+hv1mAaVXNa+VOdIbaU0tMPEL4Gb4lVreFsdGL0JL2pd43lsy/bK6PmINlcCiTc9Lse2GR
gPTCgej38QyKB5jsth9rcx8lazY8nDief218znYjKCDAVc42jE/sia5FWK9rD3/nkyAWjdcA+EAY
OOoJKm6LbQYiX7L8HsJTeQ4AhhM506/yON8yUqeFV3yDnL37NXam1S7Zy48TnFpssB9dcJIYo/tS
snWJYs+IxPaDLn1GrkSjuVn36X0IKLsCqj12nzGalGpg9R3P9OrGLKr7AFyW+wVgN0YZsc2AxNqd
OonYCDDcLB/DYLsxBhabAWg/jhfs9fw+ClGqQhuy4BiLIUPDIDpkH996bIyiSS+KTkFfou+WQHx1
HP5OmlSNd4hUcWXCI5/Hv/kHYyDjG4nF7+SsFuZZWAn0IIGjv4I3LvCkeId1AagWKg85ERP8zsr/
dwEh+4gLxgnuTQ2dvF38sk5I5/1QUo9Z8/+ceipcwghKybVXYhYDPLjALVt+r+QOU/77kX7NFtOm
w290jUxXjISIn8b1mtW9GJfrIK2XY1FT/y0sAHwP9s3rhdY4TSY4eMe29R7EqxcmstPSfZ5U1nFx
6Y1pEQnDZJQsNQSlSvIR0X4+K1QXkt0fDV7iybbukfe/X+dXhaWQL56rrPBGoCPT/Ay2bx0zCMA4
PRGgTXqA3GW9WOTUoUhx0rWLM6Y4K9DRuGyscV/X6w2kpVnJ6KSrzuXSiKLHgcIdCTy/yxnEHm33
MGpyWjdUYXAdaFMYMltPBTaMXM0pfQ/xMA7f5BnqSQVBI/TueDWruEFyavCJBKEdtMAxvZEMmTkN
hj7CX6HvrpILz2ODZOOi5Y8xhHlLx4q3Gzv/rgiuY1WT7ypH3BIAv1DMpEAadtMz/NZts6PPbafH
SMPiJwIbcYB4Rr64fYffm5PznMMUkBrJGNFIrziigiwBMZqjxw6MKzMPMCS4Dqte4VTkY4078FwT
cyqWEc3ECwNP23H8Pg7lmQBZd1R3vtQFLxBFUaZh+l0Ux6B2zScyEsLefOTSNN1luVEyyAEW+5un
qT5SLTRkQjwZfw6g5pfqDclGebENpVzr7xuxXlxc5hKCPFomgQeOXYOKcJJ8SZjr9zgE5gGMlYjZ
8jvhylaL5Kz0Swr0015yYLmB8UFc6c32BLrUrg6/FCRE3EMdK6E7xf4v5IYy0J2E09eXm2vnRiOP
88UpXZTDfMrq2vLSYaOYokY4a/ote1NCHPLFLG7oHUO1FaEvAea5KAuph5R1IuGj8scziTJHcGAU
qwDyffzSZP/sH/VADTmh01xEI4lv4kiDpIPZhSDY4/7cJ4FSr0yks7JRVU01pyMmniWx3zXMOekL
YNpdbasSVXM3i+LKUX5BIbXdeRuJfxbTN/1yOhfFuUuBqAa1y16rtnRmSsohQANvB3o2w/grfM1+
GmD2oz2p4OUOWXNjHiEpZ+CWE8E/slF4nJUFmRbP/Rqymk6qxEBHti1L0pZ4vwu0ZS2COh1l9whw
ZzM/u/Sj4as9/UwYC6GeasYaxn+jn1mhHWhzxiYs2s07QxL60SZmlhFv7DpmmPVd6AuNWMC2ZULF
EQggcdN9Ol7bGR/srccENWR5HYWUTXBHM8Tn5YddYETJYH3xz4frOgSBAk1q2ka1flcqGcvQ2gOK
pbGggRXnm1XgeemynksxyJqRz2VmWIOM/EYPq09XiiJp7x0xN75XzQqTAua/56Vi1+5rXOx52VCF
DJJuTmZGAOo+RbXgdPFmfa6j4ulDfXnMu/oybWRM8zO1nyQA/2N4SlSVWcq+3pFpoULZQmJBAAv7
cxaeJGklPskGhyKphgW/B8P3eeSUisFvzi8z5KiVjLSqJQ4g8dhUMFnaazOjJ8n6px9d6WqT/ed4
7p3vFldoGIvPO5blZNhsScKQTD6XevQ5xjSWIA4QftnUmf2mgni78RoMmUlzeztSXvTV5IFA/Aob
Q47kImX34EEu3wVZj1qcm4ubT0ByxxGLu6sFzlEW49xHEkKUqadfyDynRveq3UORra448dSnCD7X
zj6s4gsdtb6l8Il6lmJiXPD/mIt5cDG7aK7nvpxvYe4M/0oLFp+t52xgbQnJoVceLC2TYFVMDENf
xesc6lRRYyM0JZ/CqqM8n9tYspR2aR0KLbTmTSMaXbDn+DKMEwsqdeXv48ljNH8zvk8g2VyZ3Pq3
Kpw5gZyCqxgxP1OXRgZ6J3irUYfUjwLmLjyougPehgiRohS0ZBPLlkMItg4TXscAmECYrH546nIY
T+EbTUoKXhkv9reYHK36H8FiClSB+xQ7TidsgbiIuOCQBgoFeWy3fxDgtzizETASewQdELUux8V6
ibL3VR42vrhXvIuyheEnbBhpYTdypPou1EClcLte9wBu0aW1GUPB2SJMGYgEPVkWP4DCGFLDiJw9
D4zEHq/PLTkGTtshwNnTiTfJzi6j8TfLPpKVWksrr+fMRvxkbYgbmB2ybRkM/rp11E6GqLAT0YSw
SggrDlMwiOfB/T3tb6IbhvTXCfNWWzN0IbP+e48O+OKwxxdp+jmkmSMbMbukBg6PWlHn0Ohy02R3
sGb2PQNWOukpxwofghw9CGDIWAv5E0QNxjs0CURd0wa9/0ym51hqa9N/5P+YIppfhqQTqMGJKccl
cMlw79YXg2GW0ExNSHmRtMyIYOWpZkYRHNiKLcf0r99C6AXfMCSfVr4OkYStyJGQhHhC8w8b9pFf
FuRsJL9Cr1NZhZmstoppUosejc263Mc44gh5/YEiapf8HYNr5SvWEO9WPrma3/Ktkk904b/z0in4
mvDghGvzfs4SrYWzsWplo4WLe2QJ4Wl65I/gNrmhc8D+eMolF+ZsUlaTVPhDtXDrwXJJXRdraVdJ
BPE13GkWKMjbOFi4/qce6m1sJyOCFnijKJ4B+Nlf4Du5lFhQpbtrFWN06POKo9jrQ6/UxmYqMjS9
R+ApK1T6BA6xLuMCDijmTnwubLg5/SQf9kqXXdK13BQ7Jtmo1RGHAkvR8fjE+LzkA9ZfxU3LNAgq
HkX84PcJxQW9Vu7WpLd/pYKQzPBXMpR/XQlXXmt9XJD2envB0HIB0CQkZwRmoldXZBOD1mc3mvlh
VFoi0jV3C0YatmvuKVrk7ZNNfMUcjDZPrLoMfO1/1y20G255NnPjj8S+f1qMfAdGw5SvTJ35f8kO
eBXdmCRHVDC4P3tNUCeuyQ2GyMrJ5mtFtU2BsaSvj495RHCox2OxNui+nnZvUU/DUj0sAOAz2Vnz
GWk1m/ESqhQ8cgNHE2ww9YRVH0Nvil5Rer/wnxijp4xScpOihKbyeyGgrzEMyyMPlmy3+4B0yGzf
0p+Q5XYLE9DHj+mpX78uBCf/R0SKy8DUEghKi9SgpJx09rGZ9T97hLCal7v6LPyil42gmTJtC+OL
srIXS1CM8vsGKAtyuqlnFizKXblRumM6wJtxST8ldYRoM6HL1MGw7RCXAj8mE1jN0VWonJ8nzkcA
zvj2uHML/XvMckS5pIXvxI+rH8LythV4tOKNeWzW2x+GADbOTOU4VGQJmrinqNeh/wMQZ5sXjU1r
ChuGTyU23QhR2HPmLp14XVLQw//7mRgPcZ42vtdPOM/XmOxGbJrdFoRRG2OMB6u82Q6jDJ+C5b8f
EhqtVRn7HIpepPVUuYbcbK0OSsPIgWPgU4kOFLQao78kdsfUWsO0Mu+TRAa38gMqhjexNAu6EVPo
oqhX4ltlG8whTLAXcQ55D5FOmJg1CACNBwgnrUl5BYjBC0fXAymt2t7pyW7K5/c7Ixvi2271hK6q
IU+EEhJL+CWIeOy7mBXRe2PsDZ7L4e1VjXJUWBYp+paYMDJ6tRq3zBb5CT7mXzN6bwQWD2h9BmAI
lJzYjpwttvlMJZ6faxGPTZH0ac2gyCdfuCyuKncHVfYbgOoxRZn1GMoBPR2TVa3P7IHPNVqrihSN
UaW4nn7freCzYkgGSm2UtMCgdNJzqIf22Hke7mAF2EIhwx2PkkwWl3ePPXwqAM7nBlaf5ViCJRgb
lSAlnYpTBFtVKAVd+VrxxHtfsPngmyVUkGnOT1SNiDcGhmRHyuegiwmEBJ2CTAIhLhqMKHBho9O6
cz/3LLXkpjpA1VxqbtObvw3wSFluvWBQoxtLne8tdklBQjFyYLqmZIAxyBwHzqWOkeLyEkA1cMDw
izgCDPlwsjFiiHCcq/H6J0gCun3HV8jzVXeNxbeopmIlKHM/OvGcawfyWtu0lRBsu0QrgR0tWb/y
Y7D116lvprhyMwyYC6cbGLwPTOAIEl/J17BeJUiSwYqyr2Io5QUcTlRrwQisGr0fJjWoNygJmi7d
dXx1QbDLcZZt1g7uW9fiCCQpOgJJ5Roqusgvdlz+d+xsr0sQvp5BFi0rDZXn0YE7GSkaTSK1VLQ3
GpzeewGRwRpAh3t9xvuR+8uE9/Cu+xvmH32t/9aKbpSz3s4/oYAsclQmIOSwPLLrT1x3EiBjDRPq
SzvcePMlRLhXO59D9JyxOjZ9rq1iJncvEjUCujaWjR/OvFi/LqeQMymusM8jYf6Tk6Z9oos+MGuL
ztrwQpyAcaVdPlLLb5HIv07QGFcNdCaxnQnUFwJOyzj9CxJe9ouwBsORowwfmN6QjdBT57t7V7pl
mTUgm5gjxKzXq08/HBnR3lrDzx28f0HDfkwIYkU2oWFGCS9bnZpYs/LtOlsAp86c1Jzk3o/Z+p5o
I+QG9BIwWuw/cedWCCK7ZuG6+VTj8ewoxRzSmZJg4llEPoMPIHQi4XCG+URPoYWACs8cvgrEUTez
vtZ/PNmhpsaSUUhyrs7V4K6ZBOSodqjrDXep4vTnffHAVK/vD0GWQD6DlrDIYm7CuiTc95VG0Gk+
t6lBuX0wWrkCAEWT2LtrZQiy3+gZZ2LnA6Pl5hIxfmW6HVu4qdOnZ61+wWciNwICuObp91R0Vatu
Xz71rfLRq2L1tBqEu8MROjDE28XTCV70EqBiD5JBhjqCUfg++pSVmSsI7aB7ksTtIF3a8wNrAQH1
iOy+ZyIGBIRx9AXPfANYYz1T26ZW11TsVUqIa94WwhO17GrzCzzBdg4WWq3zdaVk7muFM8S3GOhO
/aloeMxXblhRkZVS19lgCSEBGT6RibY5sUzmkSrcw51feii33CBMV0SMSPzXW5DPF5MTGAMreQ1w
eawdwybxv9GhYvxH49AZChULUa/ldlOGvUiEGgB2Otuu/RRiYx8Mvi79N9+/31mUbNQsrwxOUKLO
5XahjYxSvXYEtk1TAHk3dTgK5hjRh0VO3utv453RcWdKFXdjeeY52BLp3Ripos+HZ5VDVvzBU25w
c8mkK98N8Fycvqi/Ncc8llMbbJt8LyQ98geJFy9QchlMqwfRQuaV7rHFAujkfLEaCPF41h3j+rh9
QKQsU8Wt3ZgPNNMobjTifPXKs42uvWewLg4Z/gZfsZjI7DKDq0hka70Md4iEaf0de4VX6+bzX91k
ZNYl9pcS2g5xjk8zcJmbVhfqDkuoTxn9B9PmT9vYxbxgSx4sLb/aBcpaz3SU1fd7OSJ2NOsvNAye
wojzOFgW5bQgEJ03xejloIRGFX+qZFKOn/jW7zBbMgjihGcCeOeo8Zraj0LFn2lz4NYWBhlPGpNM
ywRTNJeBDGdJ0yp3HxYF1Zdg78XwpfLCcf37VEGJi55QLGSYfE4jHrMvAxbuDnvOEYOPNxU2BjuP
oKRNa6lYVee0i/fjm3C61NN3x9UNQRZ/SNGP8bZEuvTHcGxFVp7pgAl3uD0i44mr4jgg20WH7krj
1Y3KOF+jLvnsFIv/2L8CSluFBjfc12sX4MxfSwCAqvx2iPNwnV02XIuLNkhn+ZtI1yU8sRYk7jZr
4dqRodWnxghYnL9KH7Nd6YPrr5/ISAfMWXxYNUnbM1HQ/AYpcQr6NXK1nO4btg/Fk80AYFFiQrlq
sWXhZpWe7u7QAEf5P1aONtX4Cv/PdBEFPTxnaLXHgSbE2cetJG0C/4ooIEXqgqhWCgQwb6CfEGgv
fmhEi1Eo1qVO1t7/g86M4ftGsP5123UBUprdvwEk2L390PGgUJiMq/HjBpaobbaMTc+DNMeR1MXh
hLByxcV7spQ+A0N+kFChwq/HQCeSQZ9m9gNmDLcopyPmoRZEW8YdqpUMjNUTAB5UIb7/F5X6M2Ar
1HsYKoDgo4gXpIzuNfpHQaW5nKw77ACYXjj2Ozxda7cZWd3JhOZelMcS7NL7ArvxEO4DrzIC0o19
icH0OEfhy2t8rFlM8By2evVcocwLVS9NUt0JBKfSqLHE/HV4IgbtM/g78TQHRfU/kkqa82Y9ZiI7
fwMFOLHy096WU72Keeha8Y6k3THGCJbx5K3eLXfpwpyjpIhPm4UHxLLr5rwpJqt9ORIB6530h+Me
CeyI0TLXKyB5KyUW3aMyo83pXugYSIstFDEt8Xg1Nk5YEzec61A4sa91niMZl8iKiUxT51JWKUXW
qlFOWclnUyVQFf0S9MJ0bwCWbfhJog2zYzag8TBCmjUGuusggGy79GSraFMLzHs7aAKLtvvR4iJX
4PZp6WH6L7z6/y6hLcLDAE2qHnEcCqHI2M1fR/3yL1HQ2m7fZpBpodSWyzwuzSU79RDu6NZ+UNuP
/6AMQTeiRUUnKgfnYPkZ4GlaSBKZmRANuO/Gm29h7v0709NxO3XctJ+RcQLhn9Ts9YzYjE4Tq6dz
C+ovgRYyBmSXQyXqtfxq6l0kaza4YGZV008JsSOfjnvxLC1Wq8/AlTDYBNPotCRN/jv0PH/io7Cs
qr26pmv5lEWMCGwtBVQuPiQJugzl0HKhKHiWi0dCOkLc3wnSQ0YhhnPEN+tscxJXBOe6VfjFlKjp
RlREaTtxOycVk9N312uPmjJWnNoKnmVCnVsBWNwMLgtcvuYfmNjLJfx/LrzfZa3frasop3cKQ9AV
XyBrbigrfTp3ZhmpSIM+2SOMf6CdrZifUx4aMP2vlVTUlwVo5fGjz+RCfLeGNuF90XC0eYu6t/mO
SxPi78fJUgR7LCtE74hDECpsUcutEPXxz89WKW8LT5iWqoEWlcZXEjSNwFXgOaBfVvozITEcqCn7
185JHvYEjl+8Lybb3t6tsR184952ZO/1A05DjNCsb9Sh2PzP9N+eH0slcF520f7O47XccxqqRiLi
O6lc5qSKJdtTeGd5vcgdGZP423HZP2BB17F5sTEWsOan5mhhO8Y2nnTvzWdqoHqridSNGm8P6QIK
HVnzl6DO0rXotxi6t08JHD1nOpNR9DO8cnghO1FiQYAhJYCADpLeFPj/VzYhkIOZlkLo0s5qLTx/
4H9reOLtpW2pPbMZ6xj9jmlJohjjKUcwGFeY1dUN2qz+HoXhvFINvkOohaka/wiBk17h/SQAI6ee
Eiqw0mQNLYY7ZGkejfy1xj2mSaZEOZkLwM5h0JO9Uw7Etq2dEt8gJT3u4XSQoX7NC6BKggU9q2nZ
aVE/beUFHDvs65vPNtgrGNBRMn+8RuF7qtYVmz5zRqpEi10bLD4dZvc4j2KLMqHzHOSjSizdo/X/
KHtUiAwtR5SrOzdKJmGLvgWZb4d79emc1pIAp3WCS1/hnCtV9CSWehMTcoI4gh1aYetaenWpt6/I
KaR1Mr2c7V92fbU9hAr7PzCEEar4DB0eiO4ck6QluHjzS59kjV2yTGkIQN/Nk7y6LzdMD5irGGvZ
wZ23ZHUDbtfDtT3dYm1sOGjGMF8D7NKyqvtUF5ODBpvZFyWLFachNzX3DW5OaSWMNkReOo1agrQI
UmfMR3TfJTA3Zh+52VqceKCX5VrJSh1X3AxeYUvBQ+l8BtMwgAKpFgSBBMiMIEXWxnyMg1x1Gj6O
2J3qm9Ej8z5HJb+WMo3T7cDL2it08zTqWZrirVqTKkzfiOY7iVPi7GqVjmxfryPo6Ddy8xLZhLiZ
9HhQNc+gKqLOMvLswWUb9MhJOG9hd+Y6Nj3KvvyuyQaFYXBSZOsTjOwPdyd1zTWVdHc5eq7WLJBh
bHAEI21givtqITdQu9ylQDMmSefMIPcakRqGtcawUgKu4tutr0Np7FtwLqgFz5gs+x8xNQ6UF5oR
+F/0XqetJaSkzf4PddNEi+BBN69hf99UzxZMI+Tn6rA8j9EKGKet/m9th1OmWYNYQg/1pmS01ypd
1h4dOxrK45QNohc0HLNNTTINkrwGYVXZsf7y1S1y+mvjr0msdiXQjyfGvDrOXT5ENQQSMkyPxk1m
WiajPfppxBHGhG9q0VHkw3dtSpT05Jiwfkpa204//uFJf5HZARcaylo/8Ud02j+GJLJ9zhL2GEAY
pIlko3peyoI91WB2odpRkMbxTlDJkbTw5H3rvs/1wgyy+hGI/byIYBGNOL3DO1V5FcBTKXxuMsFk
Q/mAPYTxFvbJMQKPReZuYvIE2aSxA0qG/PHf9ZwRJ70zZtltDzx/5Mer9vdJAdayu59Pm0dCvMR5
UGb2PMxW7gWlMBBOD4qTIhz1YEY1Jhd4fBdV5TdleWAciHv46MYYw0juTf7oxzFqXqmF0gwRZ0M9
mIrBVJdxpdxvZmisPBjRnGN3xqfxQIfCbbleWdplCfP/Usks5TY5mEEHMsVPYzALAFQ807KAD+hq
xyCsW6NRqrjfiMNCvzKVZvbFqimMMOONSELHp5OcE3WEJg93e/jj3IACXOKCkjGJ3gRdGHKD7kmk
BAB/3VQwjIm0soTBChDBHiR/xhNvqu6LYTp5GQ6rnZqdksGkqaCWu0nF/l+C75uRQSFt0GAVEeHJ
SnksJhcaDIrvdACRR7uQ3654uBYHY/7LKqTznLt3OgJWHH8E5F72nOL94V9tnwkSbSo0xp3OmNpx
CWJpKl82gldYLWmgPQ92g8hvq0axvP3oyyyqKJY50R+GEp+hrrIT39ag+bW592P7JIZFT3MsS+bK
bqy6da6tf6cqnWAwtImbRiG6mYK14yJ+/h+hB/mxPPFzKusIz4yJRN4wP/IwGJXKFz75RkERyBly
UbQAPqKislUAX5p89fxlqbQ/U3C8FMdzHMMEAJ+Pb/FSwVnB05NSTPERP+62rbHZcFeHOa7bdnIw
liu2kwJsKeODiAkCYTiOHHJMzASyq7+WbJxEQEKmInHH/BvSIjw06WI+yOy5hepgNU2MGF1sbCAm
gdLXFsw+Br2LjeQ7p27qwkzf0ecrX0q91woHaiOXQJP/V5Kk9v+41nvPbVnGY3irMIhv8aC0Hxv0
adJRM02rM/tddEL6gGn8w49db723XZOJlbO/H5e++n3P/FOukTcBERFIJi66Sasu/MyBqK1zMv7+
3TNajqZcmlhagBwIPJQUV4q/WeoU+7w4tcrwpVPG5G//kT0szfZ/HqRcpr3Xqa3NIs0Uxk39dar9
xswOkCSH3wXKolnUwe8yf2dWWf00tnQY5R53jsfe67WlrPV2b9y4cnLQBCoLw1R5v277VAvW8NFL
ShLmudw1bt82ejBIEhbeu1Rq9AZNaRsH8X81XRGXXI1D55qs3ANCA5Op9mVFKQPOV5oWFNt8i9RS
2wq80G2LSrz2qn3dk/qgfnxkvWiO+VJRdSNdBP7myw16kVgCqHZ7AV/kjCiLO68UnzFizo20eZN6
GDD37BjOiGHuN82bdvtwop4rGrqqgU4oAcqf7It3xd02LsXC2MqtdfRv6hwM8g7LGJIrtxaXMKC8
p4bbsdpzZ+3aAJrZxa/tBSbxMC6arzaNIEbRjQjByfJM/HWmDFB9NSrhwpl7fmxAt8pCcNwgnvRA
1aLbs5uxxNUKqFk/0CAMeOUt+gvXy+OHPSdv+Sc7ocqRJyafph9eU2Zfu5RYfzH+jSNo+kK5jS6o
wzvVAU46GyKSKfpTiZ8wdxQkjZijqmAe9ThOLX8qQeIiK3yxqIjFDKjOENpGd147v9ZD/955M8Lk
3vfq2ZOgIINEdOTAe0I9pXaDMGHqmk9HL2FcDiZaOnUiRyhc3oZ6ToixZEw0sN9qWGpAfIgVoxTh
EUZTOBqKcnajiYSoIyYCpVbNhCnBVZFiBfumLSn2uYUqSyPCmq4RadvucRStjrV4EnAyY4GxMBDd
fWucLmxsOJQsY4R7QX/Fpy0KdjRxJA1sOuVNjENjbenxENzX4MowifH0JMSUwpx7NM/jQnKoTtbJ
X54LK176W9rzf8iSmLm7pltekaN0L8p3yQER4WpjrweB52AgHptVm+p6UdHGhS/vgWqtXhKtMQgV
RTuxymSh06S9VyFmpdN/OFiIaNw61ZUS/BIFCd68lPSKwzqa0ciTlgn3unrUmAeqjeRxKkqBw1PF
jhirYqSI1RIBjyQt+09gKho6d05iDxj8YDu4hrMGkKsSiHcIp2AMfhNR2olRRmVuCeG1Y2M6AR+7
EJ7+eyVVYHRxM2t87UIGCxJKy/ydoXjh3Ru+wnFd/w6rqljygKSBxZoY3BQW3YHsW0B5zhmylu6Q
NcfxY8QeF8CA1gpVXx8J6roo4yGu1/Q7oZ4fuU0xw+OwjMd1Lcg0e40VMRSfM+7XkFrBDb+bv+hR
qExhe+yU7KaMhIQroRTthauFzvsNSPSPe14csNSLQqVNN9GaeNDSbZ3KvJWP8iqgppDWBk2/RKv+
/g/FN8YRGp75xaYH7Wui1mo9/x19y3mIpS+stKfr6Pd92r1CUYRamZf8JY/aQwGL7NRn2CmRyPsj
1AEiXmls6ChMzSod3fbs7JXyomx5NenGw1FUdt0b6kmtX0Z3R4msRiJY1AxdMmiN3X65QUFOitmI
mheDVwt3Hp1qaSvGOkht5BGaBlc7JUupbBFcL8BN5MwKVeU4T9tEs0Man3OAMcewVfLwrrVk524R
zfXy9lH6k++DjnnNFZNcYf8qKe106QhDOoMGZDEgx/q7+5Eb3sm0u63kCP0RL9haFzvuL4He+zYb
6T1y/n+YUTipq0IKBpd0ulCgyDiBLTJTLs498X9H8HJg8xB61bWcLcW3Csz51I8HvDi+L8gF5V3Q
YPClWuXv4YvfBdwLtT4Wa3crYh/gU94b6QEX3DFp7nbwGTP2CtROaBkuqpvI71vVCgQe3l+MWLqB
HeYL7p1+9cAdqveQN4AJKS6bkEEbNtgG+/4gHreBEimOIAqBlxuKm7arYFdihLGOxY2etuKY8Tt3
tTB1MiJBwa2cgWPcaAsjvK5dDGQ8d2Ls/zxvBzTqZlAQ4xlu5i21H4PC7T/NzhyPu6VoQNYbnJdA
QQTVll915nVTonc/uaoIiiwK7OvClw8hAKlCimCJB1imNk6v8rzOeXfdZ6OmDCm6RkqJ7aY4IZgO
GVUWWCgxbtMX5oM0iUdIp0L1ilN1+6r8O9o7uPcSkICGya+aDxUaI8xuakMLgUXSGXrbZtSYKCcI
K0eoABVPXp+TmkL4c7Bt3iQr6dLIlFS8YmVuzbHmKMp4nBBURiMf2s0TjUfnGBPfno5DaAx+nC+K
1euUSsIJjMUEEMeFjjQ3BqccQ8KYuFpD+1c3Ek4wdt77+CiGKT1u+kGbu8f7aggi4qz4xfIZEf8p
5sxjFcbokhzcZA19enyYi3Xim8W88TUHy0vjVQCrEX+I599zdMeyfRPJaQheTOlQ7z6u5jqsRN/a
rUMVDLUTllZTFw+NIQztsaFqYzaYhZQCkJA5ylYbV9ckwrOOqJKCtrqksd65T2hvV1nYwH/UoneV
n0cDNV97u93iUOuTEe/olc64eedJu2tF+gM0iM1hvjGB3yTzCujEE/Y8rjNONg70dGlAfTxi33Mv
AECS1a9u68W5CI7pmgEX0+VKE6ujojWu4zM5ugBXZmTLERyEdzHRq7OS9HbzFngXUVPfVQfZqFlO
LP+SumnioFuuUmmNJfgirutqe1aQ8C2IIpF1mmPmywJB4yVFEM9o3mVUgD0+ZQUqnTDxQkTwMQqH
02w8HyCFB3Ae/lr6nU1nSa/DK2OIkSc1t1aWoYxJICjpU6bV4eOkEvgW4cjlWSBMZoA/zu4i5w3N
/j9hdP48h3IPkaPADqYDeQ2RZdyMOEw0wlQ+tj1g87vvXrDowapKf+pws+LU2uJC3dl+GjAIKleC
Jpro+/o2wJCVBYGRQar/Pmf63wXLNdi4VP1HZrV/HX32DWg0wEQevwPAEsLLLGdsSWAMd9pWmMp0
NkbDo0BDV0ndSkgzoTrpR6HkpGg+CSbxOf+Bk5ulyQDXZlU6Hkzub0H7s6yhlWMi2xkmLfTMuSMJ
O5O33dQDOT2CXA4AHKZS1KZKOxiKUhXxwFLct/OQaWVxZMRVMkjynF+HfWjyHW86jk2vJ2qZfj+D
c5DLNv79mCYEhDeaq0X+K5FIi0GtbAdIIQRRi5wi+NdD+xDccQSROMFaNZX+jpOg/6BCO5jAHqQq
hw8sRbWYB2gdbmpmzS7cySlYTLIOid/gzKoTw2JzglckmspFSpwoFnAZcMOUPdvjRLK5RbdDT4SI
+dGchZgS0XtEHllpTUCCi3Vgq9L5NjiLkzy7cCGBKiVBVyLCx69ZRVmpOasK5ls/GldeDLC4IObY
/8dTn5ZcZAZgPpC+KhULJfrZmo0k+/fLzHq9/8jwPscu4KVTNs0bqxqbcAJbI8KwgquP/T9IdGe2
KJVb7/k4AmqjhpcnAVcxW+hYnWcaXZqWDLc0aqAbxVciJLowC12eEagJ6gBUNrV2KBX4zHjZ0nb7
bxkWMZuAOTwpMMg+67eSM73FNFLUZ/Wnk38V1/m/00ujPyoyydbA2WICoHM03y2axrKswfNo7YcP
DNHDWlRKwopZk5ybxZTXmUVDb0A7mICOyBdq6eXVFwrgH7YnKr54Qik/noa3pD1RYLv5k/8Ynolx
qJRdgaCN2adfsllqytxDunfsL9Ushbjdn4wOueSvDhUJQ64KF3vl0Zct5ws9dOlM18s430G4vkgW
3QRR5DdK6MFvbTgIkkGRoUqTpvJOsyeA8EIKMkKpODUBLds/vwtguJxQ99U9I5qeMMA1STnV8hGJ
vfXoIf/vL0AAtpUKKG8EDeXobci9X7Ade97lDR5Y6iBVT0lClKmimfefGrXD7QVeQWAWmj9vKqNl
cz4IfAdFfN8sUmb2HDl6aMDKFiifx2eHhvg38BiDlM38UW4D/wA5Qq/cbL4gouvM4mF3VKyXf5MW
t2WIZCf+83ojXqImx7vWblgQkmhknyqhBa38ek6k87Zq4Ob0+/h+4pWTGVnWk15n3yRnPIfhGpKV
xbGWfqfIVq59PgheKjctcq2TsDfoCbxOP1eoFwafBvnax6ru7mUsLaGHj5yxQuxc+khUSWJy8U9K
gTJgOzdhYp0P+lLRvfs7AQ4rFfHqt44gCtgz8i8pzAYL3CNfFGTaInKBGV5OFtggCZJVBDbeB161
dF0GtISy0lasUDpx/LeNG70Uj3XjvW4liMzN5/yjZ8XBBgCMuuaqKakMRuAIx4R45IAwvq8V9UBg
wORQI8+jWqWFR9KdP/+pCbEw8d7iTCvYKv2Rm4gzKX2W0j7TmClKVZ2IxfBxvw1l458AYeIZN2E3
KEHn67cWwHc+aOLq3GsrIiI5XLAkbLn3w15HJAxRPJUbvdXayQf5Nn2n+LTOB5wpzVCWtb83Lzoc
p3uLRPx6RMDEaDo1lRAvZxgGxN4rxeps/XT9DtreC080k6ms47SPIVbUEhMcDZ/p6bjBPVflQcux
xRqYrsUMA3jbzl+lo8oLFfMmhsK5r6y0tDJxzkXrBEwZgCzURBTF5i/fiDI5NYagWBBEzURcRk0Y
izRepX6KW/OIn6JVHAEA8QqJUwXXiximrJ7bSx8PNkS2lkjEhjdX7pkaJiUQ/ScbagOG+m85EcFa
ItleuyLqnAQD0nu1wmvGHUCkGiZthIvYurWvYil+GvOXHV++yHJaLHS6E7znPUJSRNpXvsl8zeDx
9mVRkVP6csnnB61bqwffB3yfkLjFGW22Gc4xrexv7wyaEJPR1cheFl6ACSsQ6aUAf96xL8bBUusr
PPVO/oLAK3j0+qHZNDNp8T9olGCWJ7jHP637y5BvCwB2eBUBSdl20GENUsUtARxA2SKVkBomGYcm
GSocVJW5gt/Hz4IfiYH71CHt9rph/oCyp1V8z/IVP5jyPxHdUn6aDcQ5+xiLG9RGpktGDTB7ePSX
aZllCOyicDyYJEFFBzGRhwheSfJuBGIOCQewK7IhWdjiV9ayDrNuC3jNWnWFxy8NcmwikAXz6zww
+NBBEpYycd2MJ0fZs2RbJ2AYV+ZZOaJsKMK5pSRILmARQLConhS9OsmpSd5pMOdz77GoL0PmQoeZ
owG54K3xEidOMzfptRKjuR4mbgq90EGG/3uRiOpudoblHc/1i9ML4GLQ/cSphClR0c6xbPagMYsO
KAlDrHcIPAsg3B6Mg0maHZ6YyGJl5jpgRR+/AOP67ZtoY2uzk6Fpum14esfu4B0DGV57PeDeMMwT
F7SOLSU1d+6saYX/CqLGzWrkLqKZqO6KwT1s2a4U6wCsIaM+/cA9i4FZLJCFqf7sQVVoFa48Sjjo
pvEwMvZUed8+M/sfzqxk1GFLC3tAt85fnjmCcBGSCjP5VLWbwaEU8cXEeBD8FMV5AMled1mU/yKh
MV4soVrye6mP/QyyY2UdAK+5NuCa0Lzzh6Q+sktRmrOYGuThN7W+cs/NBkmQJZeQ+9TfFIld2hf6
0ggPXpO2tKustIOxq/s/NJ9Jf784Y5jcRW8H3PddSAd/crNaaXm0rhV9cZjZImyix+aUXBp6nBYA
jlENGuJ0L6nvvcmGP36W1X4tit+tzlNxahfeT6Eq4eA3AuslP2bC3js5E+PVXHhh2OPOb60uRdKc
J+070gfesetHNF6ZZa1l63tRx+XfhY/2n2QZseYQ+VDOkdo4rtJKBwObpm69ijlFOGcRNBtw0UBF
8oMayn0nItZzcIGRzYfLEvQiXwNKlYf9ejmMzPLw/vdlvC2LxlubLvH6mrZ6x2YRRtUgLh657WPY
eazJG2qj+Ixnit/O3qCoxzXwz9cFFfWJPb/4N/JI+fcLegN0QhS2OLWwU5tJ6sixHNdLSIKS8Z/t
szH0wXlcnDGtLYJsAU1/cgwuDoYcAxAdiOiUReI0Ok4gC9r59nt0FhHAMbOjjXy/BwlA75IGafmr
FQS/+jBAC+XiLo2cmhuRcvoWYyzv7SYQEAzYXyDoCouIDlONlJAd5ajJBjMvcqFMfmAw+y1FZPn8
ta9aVWKIgHtSq/llKJsaPZt9I2WWR9u1tSqSorVxyIh2sOWrqiBa/9mKkeRc/LJK4qDRvCJKRsZw
/Yr1Nm+STfENZyovsyiSfMCmX4v7ekCxEnRCQMdvSlESFGQB695OvpFwZHZ0+UGmojtDDE9hTNZT
qyVGgcNQr+qr7pzLVtv6Q6V3QJCMGDISr8ofELTRxhSiRW9SmJA7njii2wRkh+OfTzPdy1yduqCk
ZgLh7qSdMvkE1qy50HFSP1ai5ZPaC8uddazZtF1P7Rr9hOyLINmsNnOsX+Dqj6rUJIPiggqm7GCn
IHHGIgXWuxny2E2G4qN3eJvZmn3C1ZAwQuXdrVS0lra+OUEcpqoe6OdpYSp3Q1nnML0J+sDNWSFo
oEf9I38wLMVJ7ve5NAeIDfHA29GBV/UCcA0JJt+EIt+rmsoXyWk6JsXOn8nahFNvjGC4vDKetQO2
7nC9ZcsoQZ+Bn/z9ScxchR2zcEUp28xG8Mrh3aguVmnS5F43c0gc80h1KwlQjfxsKtqgfmIENQlc
uD66J3NuRSLBf13cRmUfuH6rGumlN0fDqhWiNFN3z6bZreZcjG0HE204+mAgM72IlGJPALPC74xQ
lhOUFALWAymeNEL5FlxlEby05H1Bb7GKZrDicnkxqmSTc0uXxt9hNeOvhTEYgeTbuAU7b5BtXC/O
HsvwQ8aBXEjVAHqo42evw1yx6ZOpSAN6a1UINjSYRRe0rVR7NPxqbPVuxyuAjDtqY2iVYhZtHBrb
B8GL8UiEAnzJZSmzb8vEiANravt/T/XqooylhmzGvCbQbRkvr6oOBctvzJxoEMQqC778/oP0kaaa
JE2ju4srUT7qy8bs5LCDj8wiU7C/4fs3wiiaLr5lh1tTq2IgxiiSHpKf7T9bk2NM5YvTrV/OKqNb
mJK78s1H/udwLrRXM8tCeOwTp4fB5ZeAEC7F4aLCccm2EjVe2WKPO0P2eOQsgq4zv6f3wg1BOC3j
eLts2F8p81dA+yyoH9Eiabg+Qwbjib+tTiJej/vVsc18k9C9tudCuxJ7FTLcdODal+MT4UE7WGHB
Bj+DQau6gS1WvclFHP4CvWgMLoGjiHpwMsYyYCB8ZdXPEzmCF75mC6X0np8ZwtjZBmC6a72DZS88
ET0Am+KUEgLiTMxgc7Yi72qbzvMmurohAOepheMZ5p1VZWQqSYcIdnn7p8nvksDEAVYG3jXOo+Oo
tih1teoYEncEVans2t6QfC/OLCNR51C677hoe4MMWrEOrB3/wUPzJEo+YtmHoY/CHo94SolWwOtK
/rmeMQWTMuhDrk5dhGdCDvQZb6uvrHYRzp1f43CyUGi179PDuP4du+bLi4kA0zc4Y7dsGPuZ827E
BMYlGtiZvjYeoLodPAMBE7oSoVswC36EFbN3SAIJkOB1NBvE8mzV+72Re4zrVZcTBEREg/cBwKm0
ORkT/YvtvVmofPqnr6RLZJcEfcGa+H6V/CUvKo5B7O2ho2RnFMWotjtYFJ62uOYLyJb7EA8Afred
gx//i2kF0nJiF7RlJrvPFZsspccAoO+t0WPKB5VFBFOjHGCSYxSY6IOe7Ip3MJ3sNCs1zD4dv9dg
MVUz6qmxS985gC6cKWJJ58pNR1xL9WWq9rhBvK92OTTekJd/d9Vev/1JHXfXnXEpIjZiTWdBzP8w
cNK00T4K13sn4suulgwAuKbT1+LYZM+uLW2mMnJAhFS84tMLb7vPPrvd67CRrnLqi8vXLfx6L3bq
tvw0HZzNDzVw+z/pgj1rj1UX+Itjz4/S1CWd4JHzNyZsjWSLDaBZzieg9pucjh6F2kVYyxJMG/W2
1YJfnCqT+3m+XuLpMkNvvv5RWW10Xl3s8K7Lk2WuetlXJKtUYTGoBoEKw4k3hvUl6kyYq3A4DC2P
pSN80E49tJV2Wd/zTBeTvCsWSa16qhULQKFREeTp50S6QijqW2W5k/FtVfr3e5Q05zAhVeWR0a4q
Xh7qIz02HcGAC8h0uveFGl5djws3K2tKlU1YkMTvG0VIpfPttDPqz47L62Kkh5gfGdxWgs2rx+P5
gm0VNX2DMEop1cBWeEw6BdlluN2kxta08jg9MVRYcfxc93ePA/dEENDa5Fwp3DYz3CRT9ymZc1gg
t9lWF0EGTDjVoxxdI9NpYV11JN3REv0FGQ0UTrxd04FVptSA9jU15Quf1MDG3c23wihymL1iARZv
UBwaFU6U4zzSYrDYs07UE1WW4lkumE61khEcvSYowyvePbC+WXdUzCByFYOltcxIgXWkFU5KSuIm
oM3b4OIo2+wWQ3eW956jK1tkjj0IN6uSig9Ottydc6wjEOQqWP5aeSgjo0JjMkzMuPAw2J+evpD9
eTwEMs/ruOay3hOWR3TyDMPO1mSW44xWmnJEeeH7SQCMJIzHqla1t9TdolpgMAksHT8iQGcO9O4Q
noVkkY+DiXtuELQPdDdKiLHrV4tIe9B5hgjBwfVm4G8SkL4b8ltVjOE10EiFcKfE/oc4Bn4bzvqa
JRI8Oy2Lof+MfFbsvGpVvw8Lk0zPq9+lwHlQUZe3m6M+56os3WICKG85x814vypcBGjOdgg7VoO+
gSOQJtxgpp1tS9c9yp6CEr5nzFCBVw+egrj+BT5/z519XhCdwtYJnaYdamyDi5GKdk5pSyIPsu3v
0C9L4vuFwkBA5oNmM1lc5Sk3sCM/6dDJ6JziiNEtNlUakCjqT2KmaJiFfE6cHzl9CraCz7GsOUn5
AtzjnGKfPIHpoX5kBdqWcb+TiKjzC8GiufywH/y19AmuyFM7gJldipn3x41BXL7pBJ31UuLbROLm
9ONtwPcxLPZbmA3q1iO7YdXDIqq1DIQORBSbo8xztjzT8Sk2vVJyn0kilf3ey7bDgwhAeFqIkbj4
oNC5iwow+U/fTWC5/2kFT6dAIXygvBNgpnJdl/h8shxEzvB8vumBLTPpmFKPs6yUY/foIwM3/hdK
hO80N1QjMBm7xGu8md/J4rFWxYBJO9hph+1MOK7qiyUKGFIuAWRzC1ZcQwxw19bjbF+/+DyJazfE
Eek51U8gmwdhncHq8BIY22A7ceQWsfvBYYUG88R/jNXDpHk3ZhpBV6cIEyx4+w4nh5MnNoso31Tv
NLbKtD4tVQxpoWGfXOFegPxu91R+O8IsGeDaP3iSm+AmFn5krKykPtmnirEB2/F9jwIRWxBmONZD
SSaz2WLEINZ30Qib4bGFPaFozJWjjsHn4W7hc03Ng4Pi1Ckm9SoWMz6CkSFtyUD69VKZ0m3HLMHY
ZeCGfWG47tcv8wAFsF4OTvqmTVas2KQR3ZJ0XME5ZPZKvz/myeFV5DJGLPwX+4nQSKFtkD0xi9uK
YXSN+/rWvnNrpmF/kpZnl/tg02AClkom9xv5jCXAtwRTm4hjMXFEI68wlARvjgK0U42u5wLQt0jy
Ld/yFY7DOQ2eNxVyqogbyE2uWl4Xn9lh3biKKkJ3ACnxau1DvKujEhFogsea2kR/lppxgRyeCnGk
16vz/NefLT/dmY1v7dauAGzsaO5r0HxcF6Z0G+Qopwg9gOnmsC/M9SPyRoWQCLSEBCy1/ujAYyke
ZbeLbvrPHOxdrVa4jpCI78JqI11GLG0KlVEPh2a1PJXv+JSCM2ewvVnwCRt43H2BJXT1TYGqyUHB
yGJ0XhBUh0s5EaEKiqeyhcOc/qGEK+7YtHBO0TlcA7/OINCynJ5lljtLL5fZ+9E2dcQlPPrSXX+u
VF3gKpnLLtJ5Hhf2r1F93kGIIMkw6uNQ4MHDg45K3sFBSwkh3j/KOxc9/ZZNN/BU9qJSWoN4OBNw
gCHZUtTUrvVAb9rTEvjkrhPE81/Gw1woY+kamafnLdG+GA9Lnd4AT5p3ef11HUzbgMo9gY+8iy45
L+Yu9aWYBe1LQMhQlUYoJ5Y7+s50cfpwFhHUhs41h4X09BiGqKscEllb6xhBGsyWI3Ge3j2hl9na
d79225U0URfDkR3q82HCupI1WvO0k2PqBYS7IxXKRMU3LPiYsm2PMUvY2nf/fkNoDVplejNIiHbB
iaD23bgOEmsn8fiOqlSfYfgXIBdCsKvo2K5Txi9V1kI62po+j6joVA7EjCBOe0IPqjFG0PRRbP+s
rTrEdJ7PlUkU9M18TQqBrQTJggnmR5Hz9wJZOhT3qvqUjwjaQcGrU1ZQ0tLhq29Pv3A3Xm3r91T1
3i3dNq8pNAInjmUho+GrEub/b5mhqheVOCDhFonqr1hflYRGqWLxqOyhoPtOf/SPy3DBiWUtyM3R
QzudYzAkCT2OlKXPfmEwhakSU5Ux367NUd05aRtPOiotcaO8DNgRIj36ScVg6oSybmza+PpJb/1Z
K6bx5E2PpnMYmLScwXT9/60PEcuaR/IgvtryqIw3cUBJCQaAGlnQBwDkv8lZtzfwjR0lgchH7OE+
RfVYUk3gUehwmu3WKDIRn6evCvh+zBUioxJwq4rO+G/NlhTWNCBE/jYf759Rb20EeW/B1M3lllql
VqR6gOC6cPmDh/jIhFyBoIi6IOcttQGyFCy7Rm+aZ+sVXDnlFHemmoixosYuvn3nIRyxZLOrmNjy
8gSZeM+GRbyTKbMmt4/ylqnA/CPzyuGcAipsf9JgtaBSkZMwUw2MZLt/AIaPF+6CpETNDvTogKcm
4x7Tnja/KnAcJJ8j07wojQ1jz14XdQ7CmqDUZbw8iGew/eu0RHFh47ET86TVtTLLQWLMKoW+YtV+
z3RlPXJ2xWyRbrDfWmjyBoAMmwpDFcloLe1RazFlvmds10dRskQZvyaM4obqVJSNGzMifz/LWQ3Q
9VQ2Dw++jNjb7zSBoCAxN3FEVI23KprJc2Z1b9ZjKM5WknC6iAGoQ5REQ/HpohbkwuemFsnf4sN0
lGeiz/HlTj5NzJG2rINw6GJQHtboUaxSoaFbwF1xma9QsgQKN2K6z8jiKhqoaSaUsWig7752WGh8
wQdgB2jpM7Ss6UYo1ZtEBBRf5CK3JumuLWibVfvuzA2VVbTRetetMqBzswqsXJ+KriaBtV7OUges
9shoXoSI+Pik94L1/Xpm9S7/Q7MhU7JIO4kb/SG+BF3KccLeUxy7t25nWPAIDK49gDmUDxl/T6yu
le3CWU0PYfaBwURtidxBBB14P8lUKfE0lPggqUynL0r/IRXHAIcAtGAAnBnJ7Yljp+GK8BhGTDlV
O6sbETmRYXorOLzvtwzpdhf96VcAWdWhqon2CkcWM5qG5eSYDtO9/O4om8rcLNirjBnSwcANUs+V
lBdPRdvHXo/Ghrm+LDNeJGShLMiaGeTb7GYLlUgDdRvW2yFIFCilGgVkC4mF7MjFWs10LL9+136a
O6l8BzmEjbyrhkQxl4/IKPRY8z5pDdfyAKFyvRknGqvuZVNpjDLnxZ/07/ny1TMXM4rgts2uZCHO
ioeHfHlkKFcoz5h7yXODElQr9wD/FeiIPKbYFqaKYaKZ7yJz8or913AG7SfPTBWP1l4Pc+KlNEZr
kuBrQpBpGn3eNXSwBuSQcXD47qJwbyqCW6RoaXkRO0ELKDbwdLOT2c1Gthdp/HpX7LhsMdtvJ4gq
/ZxqWYcHQac2QVrOHUCkbhVr4Hjmjc2Dj4hILweEONSk+YA8K2tOfmnLDP3IWi3UB/e1E4nFQSMU
4lonZhRU0JTExRkqQJcHCRnLTH7T6DYCn0LYqCO4fBbuMI/DY6ep3SW8I+ynARf+15FqeJaYF4h3
OED4meFGSGqclPb4D11mC4wgNzF+VLOH7UvWsW+4xp8MtzQbg739EnC56sQkGzkUei2vM1xzumZD
N+QGOAsKIsSNMztZdwj6vS6T3jBImK7uHusO4CZkJxx+7GFx0U7I2olK9G0porIH82uWF9k5tWAQ
/D6H56MhZ41D47y/bVxS5MAi3uJOkSA9ysiZZvQ2Rz3xOJPXG5xNKiziel9OxgIHnXRqfxc/rSJh
fXXeH/9Q8HfTaLxGvl9ookiw3Zmwh9Ou5JbJeqfFOU558nf2XLvI3aQ83e0NQj7zmwHWZWMRjpev
C8lnaEtJzJqfbHTj4dNKFh8RPDab0nYMLWVDQRalLbpeTpo4d+9Cp+mud4c1FMOpZ5AyEDT2tZ4+
ZGLBF6K1uN8FKiCEiWpEqlEL8fiLVGf4VAGwnUG0se2qvCAXQdczsXHDqgADbKGlNezyQphg4yk1
bhz2SQs3qa2b34VcMBmftQZdm6nBqA7/4GTxXxrCePZZ1ttPKpmeZARUmpSTJFT757f3t3yaXiE2
YL/N5hC8O3bqIr9IWMEkHUZx8uBa5SobneVR31fqqKqwXsXeTe3T85Dd84CNGtX2rVMgfM6Fqzvn
tQYvC46B+O2Rj3W+XWCJUKyeQTGt31EtFGf4hRmjVqTfQcYYuKYyGxO02t5bIC0K/V7kg3R09Gbg
n/5FuY2jzYI48M1qRONcrjCOuN8Vwjws43DtcLmgYnoSWVxNBd1HnsdIfSQ+y9iYiYscZo6qrFSB
oZ1+E5HFtDoKMnLUyZDS2jE2tj9aNwhZr67oVQ9uuwJR8EM7WqEyQPDoFI4keToAZV/4iii+iglp
xJVDVEz67mTnyjSlcEq8H0Dn5ciMxV0JUVkZh7qRzTLA8zBrPQuVbiQDKq22t7z767hsnMJUPYt6
BqH1ctgA5VJx+ogJNGqyA30jZ121SaCEV9P3DsBOArRRhL/iW+Pxq4NJpx1Z0jmaW8RON+NbW/Ru
MWac+X4vfLGz4PtwVqfKUBkuO9Yc/UNPfHPpC+5y/UldNxZ0I6Z11MyJ18qdy9a90YiG5aWW+A6l
gp3ezSX1bsyRzsy6lS9tcotd9ceTQLuOTfTSIVyLn90hd7kkY6FdpweTEgvK9hyjGTdM4872Fvjc
6JjYfhKXDMpFYxyIFFd+tgUO+gVEVv4+Nx7y4BtU1hHXPZgEAYStv7EDqyRaPslqtkxLGVnuuxE2
dYycCyI/AA//qyqo4qsbj4/rpnT6CXeiX4Ua1dAuopcN31aze+IhaLCPxn1bjYpJAW8ZSVxppWsz
j3Rg40KMO3F2+sz5/hSh1lMex6tUG3zt24O6htSpbHGVeOyZJ/97gCVm72Ixp02qiakhv1xJvz0J
VnfIWxwrCZt3aKewTm0BlWuS2iTkswWTBxLX+CxZgmFtMe0NfrLSv5uBWuDzhA11v/oWUvsJ+E4O
Bbf/E0Do8wL9KoHHZtP+Nl2Gd3Thb9Cg2LR09FZl4mHnVkiaKLl1Z5s7RCSMQ2ftKOJMwuavIMtG
K/6lyIGoZu9QTq8OzdVlmI50+CMsWLd9wR6IwbrP+2XjR5OYYXoPGC6URvOOWwE8gclwCi/pxSPD
/NWEiEmh2IqPjekk0kkA8HzENeJQevFItGmOpIT8FNWgtrBmZzBm+GYTRO4bCAxogODRDnqV0N+Z
cCYSN4zqGJ214ngHsiQp9nJ3l2T4pCW0gEG8hnErLwS7N+sWF+fPK1Ap9lsUQkR58dkUmL3AclB2
/jOTbT9p5365hIf1CwM63BVRZ2dqGK0vmRPwvYfFeHfSeCnwcdMSh5jfSwVImEoGha++quqq+vzl
UoMIkceda7mNoCOMFc5xHWJZOEXksI7DFz/kWdncJJZllz9DySPu4KvqzFfTF6z/SSGTnD7WL6Ju
EnUjeYmIwOnvq0rgZbBl3bxX3iqMV1xKpyn8BiTHvEydLXJkvO2vk5IRz3Bn/BWW8w7Y6DPrUYie
W+Zt9cR+Ft9BHtXLJ+i/n6fBVRfbzYJX6KTcOzuEoIJ8JObRxJII8sC8arxBVqu3PAq1gF9bMo+A
J/e60jstGBJpZdfmDLW+nVNtAT3HWNyZkIIiXslGiELfGROpXSluIjSqulkhvYDozxgtmeqMLBdb
Q6JxGrWvx/FyO6qJgiqbSpBCvngx9Fa7LfQngYglyMbPDGSQXpJaCY62fm2JKTegQ2vvAxu2zqjG
FKisLxpdXNgR8NMfppqgWqCarIm8FiXIMKpTITO/Iq5XOXOMQGGEtuxvki9NFjvVNCgMCFnaQjUv
Ri5B0mSKxbTPI6dO25HAXWAetNEjgTlmRauzUCsMyF7xa3fOLjuLvW0CQzZkoGJOUr1BZZbkOkM9
0OmhUAGX5CjSDj2iyb98PHtqnedu/ZMRS1+m5Tov4rNcWY1W2Mb6KbFp7Y3CEz1vq4cxvNbqbjaa
TwDntZsIajkkuKuqr/8qTgP6bKOCilXvO4pR1VG/q4rDkFUzpdDcrXcuLveYpuDOVfFonxM9+3ib
Bic4gGPvOxffqLgySmVETHCv1g8fx8Z29v3z2rH6aAF/CLk3UERJ9eP9vFQvOdjzR2YwJG3vsvOe
W/0Mcd/aQ+N/1U/24K3ghypslEdrhhHvmyoJ/kO1UEUmwxG3XNdKy5gZzFFL9bF2HJywwubflOXc
N/+wU6e54GbqFJvZdr84ZOpMBgBsPtTIGhsezrBXo5hhugfUf7QpKsYovGHYORm57+Vlt19melRG
0nch3MSDpeSq3XixxKTcBWZY3t3qKHbkkwr5xtz9FNlT9powzgpv457LMc3Q8cB1qzNDkfyXPNdO
/bt0AzHnNp81HMOAE7GJ3zUyTNwEQt4A3NuIq4+h5EfWRbqDqciDVYBkP/T/q6I/Bzg0EniSd6Wd
ZVUwiqi93vfso+c4wmEukh4jsFdKHHpZZuCok7jotQS6Svqy4fxGtqI5SnzL4RrTHgkgEqBgp2ZR
bipGRDTAQBup4cf/Y26SdSNfSWAa0P87WUEv5A2V8auN3i8Q6jQCfc3Bro0729r+dxIDFb9MhmEl
iHDaPOV+JUGmuP2jeoij219+xeJP92QhHSH4HRZirJwRFF7td5z6z64w7M/F8Xs+H584F1TuvFiq
u9SlPTu96AJ1G+mFhBv2xIps6O/zcun/InfRDQL3C4aqWJgUEcLyXsICXJY45UYFUVWzDsIA97r0
uWuiEtubVK0oG3dOQBwtbZs3IIAsvmd79uGKQDwCUFFt6cg4+ksGCfK37HKxmkZRQaQKY6cOuGTD
26nhsIUyfJV0ThCdINm4Az9fS1gzdMyPQRur5GPPuVbligEMCsK7ypOBe+VfwMNTsGjtd9WVnoxp
SXedwWxHr8gTTDFVaN46Tt2jixb6APjLP7OEM+pm77/wlWdFb6dA/qghbNXNsx2Kchngbv0/ZhrJ
v/VL44upmBfGccCMxBdsguGYkzRMNJUXL85bhwaUGzBWNXDrySR+kPf/KpVEMrFXbuSI+/Tm4DiQ
clv0nppwYOjjENRZJPx6cGIZnRVY6MubJC0wWwKhT+hVt3wdHDFkShNJ7+tU/OsYZcBdL6bP6e8V
hqSmXNxLh7J02isKRqgtuMcUBopM1wbls1DRLmVekeBm6HKauKkLjM1O/B3TvDl3DyK12W2qYa0o
8SaZQIjgVFNyTY9/icdYiqlkLtUEVKQhPMK4wmui4Unh0xtaJBT/AVn3+54F9bhsyL6oo2J2mx6u
zEfRoOnfxiI7iQ3WxyXu+bNhdhk5zQxlwq0c+M5bntOOvX96oQoesjORILtLRW8oG21jb+isNXYm
uRPx59ufO9G4FKmJC5rM1+xP7CDsdmVv0f80rzF6KR99amohwUyQry/KQaXSDr0DR+L13u6YBopu
dXgTG1bW3Xn5HWoNrQ3MJ/oeEzwnX4qYyTbE1ZL2oUjOFh1tGbQW7jJCVd30I16+9MGOsqc5m1A/
nCbtc6jyg9mloKMr+e9HolgLB3sb+9ZjNm+zNdSk0hrM0iHdsDBhb6/k4uWb/S475lPlahJV4JG+
Rl+VQDUJj+rghqHOvTKOIF4hzJj3xnofjKK1siHIyDFR0E1o+LAiG4MKSv/p2UbaI87ZcRJYjq+7
WuGhsaY4D5nTZNBzmeDXblqDQEISys31DqE5LrZRWI2ML0yfJrNTZG6G+4PjYePOlfzMvmvc/leC
E+2sVgvrUJMSJYM7DmDSbCdE0nRrB1N2QaPnTupoi4qtMJ59KXz7DfL1+avXKjC0kfNU8V0iV2Bs
OAakl1pwB/7Ha0fXewm71AWJSV/uK1Pa1ix0ILRrcxsfA62L3qV/mV7hJOrJc6YYO3SEXCyfRxXj
6xRLwcVpJdu9JmA2fpFPxEYtBHGTDmMLveqoOMpj5syL6X/SwCBQLeoFVg+72xdwb0eLWZPMdzWj
8H5zb6Ettyd9XtcBLZ3EoKe5okGCe/WfTszRpOs2HclBg7MR3httNKoU3bo5Vo0vvhzoZKTmgon6
IXh8QnbjLdAZ0aY/NUlD+Kz0+G1hfHSD/4hzx5El5UflH3eVKQdmk0LBU97W+spUNNw9Y1xdT+EQ
Xm5uxFp2RE0bPnKR59NuLLd3b+5az+fAwEYQmP9opxfk0iD6uMAq4xN8lrorh8snxhtBf73Flpd/
2jzhXQKzLsaTsJTYeCABY49Hl11g2jtL9SQm60Vz49saS+ukW0iwXgNh7RAmlepfwD1QpkMN70GT
Q1m3G11f/OmZCQuxzHhQtBEFvHuFdBiS494wHyZmHwsR/AsnZqKTyeTo2aVmNmoqhHue8RVnB0HA
jqZ8Oe9fkup1nFX0sOxQbWdst+kVd7JGyMpHSeiJOo2hVuZhH5CMXoaA909QxkQKPfFLk+I7kqiz
PUPmrHzGw1NCalPTifMI0dWp1VukMraAsC+RgH+25nqcFWmwspqR3Cx6LDMhPvKs6X9Glqt0b8tX
/CDr9Mxc/aM0u92FDGM583HZWCiy2pYuf1BNE5l2O/P+m1V3vnoW+dHe2RKdy1CWc/FIcAkc1yEH
Lo1WFYsc/6gxiRDIubIMvSRKqFGPtlo66GXLhJIXHt8Sb6rzSn9uszlnsAy+DJnxoRhnih0NNuDu
U6A4qgAfTrbYkpd3smnPKl41ZCKjDSJt0VbyuIilDwuFqIpU4QS93Q/LqDnUrvXyxzJpK5uOWRqg
+4RI4+uWZFOXLlU0HKp4qJbbaKd0OB5+ZhtRFgf5GB38I4sIJ04sjLD9Y1cd9bg2REOG1IGMVJzy
ndUqjNhzVkWrUJmWIuxGJlhTQPbRwwERB1lBqgS2zxLA9Aj67htIPVJQGmZLc4lMApac2SKiDy0S
RZFmktayrx5bioob+E3EdsU2HUHL0BBuaRT1cSDpFYjsQgTfhESoCin1YXHr7Z3rtosmQ4SyCHK8
R+IV0KQrKu6/RuoXhfxjmAxAk0fLeDd/q8DSlkBAh8YcPvIgWuFBSOiaY5YSCP3s4msAdinRFKq5
EwA8tTJO+3GQLaPh9EQIOCI9c2IWMnHozY96vC/H44Q50BGHH78KUe9S7Ff/eReR9yaAbZqYxjGJ
Y7LzIou8i8dOEh7TT50EyqX+94qR3IR6AM2tE3ECH6nck0gfQC6k7TvRZGK2KB6VzIxQWPixzwz1
DkB/heECJjemckapmDzII8fNtmU+y/g5FAYZ8UCQtY3GhO83ID5ITdX67inC2LcKD9z0PngG+OI9
dKqlZKNpB1a6TFZbi1DnF5zi+pPMLB7E2p9DC+c6zlWwz2brphOkr9BlGhKcOIT6f5fMxyqRanFN
nDyAilxsV0nHVgPzaT6hYVFemBHfndAkMdQwBVQRWnxevsImV5uafeYV+rIWFwEBmtnvgrqhhU+3
V/rpjdMmUZkGnUGbAXgRTkf6L+COl43pBUQ1yI8E6183Wa50uaea/qXK9v5CLEGb/6UTOpz3KfNP
RS9Zc18ocX6CQ+VeTbJJGUoFUfQQ6Tn07o4EC1O4BHHdhsugOQEy0EomAyGlurvbYxTZ/QpIm8Oi
KmkcMgYB5SFO2jGkNnT+b02J9gOrYJItvSE+H/8Zz+uBdJgQGTR5uIf4aa42XUBa3d6ZrTFrvyBp
VRc9vX97uCQtUDiUmoiaSqLhwqvwyrC1wWbwm0SaFEAUqB/EHceuwaqdPXvRDsIi46iS/BcD63Ke
TiVOkQPpmQ7e/YgXsD+kjfta1MS/yhj1tAjDigE9jzqXchHn6aUrEC/sX4yEtUHNJUfzXw1g6I5S
pXBNnyzs2Y+m0cOHzNdLu+rpXTHI+EOLMf2Yp+NxXRC7FsZVcjUUSTDx9sT+AYeld2+Hn9tPAcnT
jrexON+nIpATb6CJMICVWqraKwKOCoR5jlcye4IRKrOfdijjEcs8uTgaB88Bzl5lLGNKkcY9qvOW
ASWmRyutJo9o5/X5/1POeCIeQJpZRWqUcvCXSWcubPWpJAE34nGQ9SWN4v4efiyp8Y67FmBuSCty
HGvLAYlci8cL5PH7wNfnYR4ABZvm4I2+ZcmICsPtKoTDnvpsTBF9q3Svm2dxChF8bxabVWXaQLj5
M0FPtPXISOV1oy+gZBIWgHr4bY1UKuKxQNgL7Dk4KKBVnWJesqdqN/tZ/zTu0hSNy0L2PsZzq5ac
0ObZHNxc0KOZE7tajZ0Z/BwvPfqwqtzCc/p3eQ7qw2AS29yqfTiLW9DZ93fkXS0e6pd6IY0R2w5F
L/0+5o93QJnpiPq6DjfxUYp2MmBh28ngXfRu5+FSgjf8vqjO7qVni0di81WgrW7MoQapef2x3DIY
qYw54NeCcKEB2A2QwvohK+6YnptpIrZjHCGqZVTvP1wa0VGqNNeR0Bur4IKKrOrbI4zUXixYZO+P
hRwtxBsNogjQ5zn50LFZI5GtkO8pDPpzfpY6tv1/s6cYFkbMvXUxgXPFHMOXAk/ZUpUC191Ad1YG
W/zOSFpjp2qpkIjsr6OirTyoAbIWtq1icyWPW89hUk6MsQGIgm0ncgFbuns/q2cndOfcO6S7EIIj
2ALi9SEROR8lTJdgyWes1Mdu9TYC3SJ45p4UbXf3mTIPwjQsizrT9C0GmwDjCD1UmjeiykXyKlKj
hw/dQP1sNHSR6p4DWr5ciFdXsndaWmhKb5N6qPyuVCD6OKqB+sLdoGoWufwKb6+S963cPk5ZAH+U
Kj8rinDLM1GJmOOqr86MhagUinuth5N4h3XX0gk5TCGA+W2pYEdRqyKQzoNaSr1XENvNVVbtm8Nk
kVB8ilLw/J/DkY6V6nF49YwIs3Rkv/TRkmgVjeDuJhtydtgRiZRPwBXaoYqsyFwTx+YEkfIONlbm
TDNUZ98aaAZHXkJ88h6uRO1XegI27QmPNbQn6IXzSjn6eeDCOFU1+ggicrd/xyb0+360HAeMhpA7
zi2ez83WebWWZYGOR6XgjjgadsrGuu198EsBiGGNMcwmUObGBBd0LPPz73zkT7SNxvs8GGhAhkw1
2TxUWnKANkT2Xi6P90vtHBWBpI1PczaLVm9RgeVIyWQ8HvA0oPJ5NhkfdKSTyKo4eb1heFIZwOC3
vSJWI0OJDMFvi8XEwGUe7r5erGdt7EYu+xZs+j4X1CvDVSBr/bTnXhplkaVDKxNQuysTaczYSwHy
T/P4xPybhDWio3yNvxQQbhl+OrqE4erXRpQIj2ppLPqPHCUIVaHQzEjLq1pXD/4w7hW9pVaRCI+r
viL6p4AiENCKIPfY07KjtdJMdTW+tRaAAI8jx4AWcYg3noD2jEEY6iKtmMuclOsYEbhgA25btOHN
uyhch98SUtfrUWTJRW2ZH6WS3G14IvgUfs61Zm1sac7xTqe9K2gI7fwsSBg6s7eQT+90rvVRnsDJ
7TunaE1Ph4HaOzLf9mPq4Bi6lqZMz0u/N0nG9arG7pyWOyCrJYUBTati2rJe24KiC8HUsIPum7dY
LOeeDutTZhuLAiDaonSPkezFgVe7biELGbcLBB3e3xAigGbGtoC8035RTg1L/+EmxjlIxJV7XNje
QpYuieBGW29Dk8Vz1Fi7XJXoBqAcSVzqwlcFQpukssSj3jlIHMnT5XX3Jc9M/HA8W27AYqIwfXXb
36w8z+n/bwRPI4Q40L4Jr/UaHTJGjdNVIF5nSfvuDGEiPt+deZogW7i3Yvzv4Y3zM7m92NQlpCOS
BDT6B+ql4g7tXQzSQnxE/Z2aRgz1B/hEnfWXDRJ9LmRIW5Gpz0Ui6/2CLOr/DJsrC7x6n4wHPJTH
mdgfz8IxmkEsMfnHbCN4vUerUF8msrxXF+J72jcyiN+h6as219jgEBOPhPajW+bc8Plr/GPcAL4V
Crx2IA/A6KgxSydwAwQPV1zadRJGEoPRcVsg4XUgni88UySzCUOy7iPBSctxI+uSAvTen0HyI08h
70qhkuYUdwEG18Oy9QLv3zFXl7cu2w0zal+bb2o5IlOqY/M6KoYWJfR2qp0WCvrgvz5AgSyz/p0E
k9ZrRWMj4Mp7OFmmTjObjVX7WDppt152sP7ospKc/IHVeoOYFDzyrsu5gKtTDl/rctE46DkiwcWl
KHE5gqlb+BWsFwi7A0RzyReBHtkpF1DF+MEWW2r2GjVEJywXmvReW/Re96uHtoV6lzoEwZEn+Qkg
/HdbPMO4K+aYMBjwIuEoy6VJPmNH71fRfkMrxKsOSUCaV+FN7cMgYziPaJbJ4KkjIdQD7gFRPzNg
dfJfgQ/DyHXETunVAY/8nfqHCg0EWiQAGrNvJckxM7+lNhtjoBBCYWWzlpKo6h6Y/9TJCBqVku1a
a9Y28LKPHbLuI5EeFqnMRF7M0PmGJbXVnB5+RIksWzNXS+T9CWs3w+Rtm8Al4fug6brU1ksvFSeK
zXjTcLu42stt6iuCn7mbqfXYNF8mhTZgs6PFgdnCx28BQ1SghE/1CsRicq1uz2D/Bkqzjz1ca7Q9
WFq0R750ebJiVgIEEtEQaDijIhI/8Dh0mD/tiqiBgjRfPXCKHAN9yQW6TN/bI93g6OX3ge7HsIB3
dErACcCyZ4IbUENl8T/W37y2osPqDkY2vU2d/HQ1yfbYNdHhXm7r+dmpZQ1JwSjWudOvsSykiIlU
NkeWo6efIeX2h69wFbRxOHFzzZ7JIdcvRq6zy9LRhAX0aCjbdt1vyFI2YWXrVI+uOH/vzEmW4/Aq
8qeCWtv3/yUttMbaEvf+wOCADGzPvn2PExox5HtjTwzUVLPO3SIb5clLY2mMmj9RbLbTNp6HIdC1
Rks0cDqGKNaxt51NhywniFk0us85Ov9R6QyVkKl8sERLV+2Uqb6nQUKujYNQP4xMvVseCaj6Gg56
gunOAfS7L0i5LVARpCU3ZtkSz5ikZFw6HOBlKllmUEL0O9zvE0uBPNj8f3XFKUxWxinDm6W6m2OS
3nAhuPLjr7vDHBJY/sxCAziiCwxAH6f0rwOcNhYV1feECSqgxV8v4wtIW6QkSODsj/SCZBCvwnvU
VoX9P1KgvPmUAey1Lx42Fxr1wzrw0g3F0fSVM4XmyGkT48ANDOy6EViX2h4Y+r0Ke+X86qIwBbn0
YWIqaVag5bZVWdVgxaI3QwxsECwMEt0jl7HGYsdafEg8R3gle7yxy92moq6kg6yTUpL5eS6Imfe1
oGs5hs6x2QJ80OWnGYGbg0to9V652xcNNfBIyH2ApA/WBFha0r3v6tUz895n4dfH26J3fCi6Oqsj
xqS0g/AtS32SfLw3D1aXrXvd+ehgNqWiUy/jfALQ3Yjyv6t9lTa+ekSm4L4pB1cB5fKBG2XqCQYp
GALRbGUr60m1a6e+cN1mSEvQAH6yH9Rw0i18oPrrgzt2Ips4LmH6Vxj0ZmKNjdMGc6wvp2Tx6zcg
p5z+STKk/rMvXlPABRgHqpKYnwl1O26/YLNbZ6FbNF9HqXW33h4H+UR1ANwg9QsgQCDBIowedXwE
M3UNwJajVce/kHRNyoZMA33fL6ZeG6uEWsdxrqZw7S6QBkDv1VnZpN2dJqaMOXEnPyZZchlbzB9i
l1x+BnbhyScOf8nQccgs//uSHGzvt+ScIBFAfIUdMfgyKOoTRParMC0wgX0YAZR3GBSmT2YoHLo9
oULazRnNWLFzuq5GjnpseMC2ZcTtaZmZkgalTF6GYOYLji5QnNXyXDkl2aGfVXCgByQUroI/fobG
In3/nqC0LQhXbowsJsL3xUVrRGVWgVijgW0MhkR2FfHo5jnEpuy0a4EgyAy3aDOPv+5vmhpukfV8
l7HWdkjjneTJKHXKqM3aOJqwaG6INj7bLVgM8Sb0K4UMSCPxiqRYXd3Qe28k9aa0TUAmW5dnTjLn
ZrBuXf3X1VZzYkhKYl3u5fjR4uIp4wG6Ws5uxTF1gywDlpoFI4AbY0KtnWJr5N8RQhNEDWrXB7qW
LyLGHdvZfXNIVeTZpxQS0h57rGZZR+5btTCctcoIe3sJpeILsvtxnK7xV6URkAD7466DVicDpsrI
RhNChBYPO8N0JCvAygGonFXnoRmREKvQPkiSdIFx1RU81mPXow+AOGqMWWpJ1QNpqbv2mvSAD+ut
aGzd5Xdi5DsCHrtl7OZ0ycGV9n1/FkpD8wmKVM3JzCWbsFxBPPxI8sNtw5TfHN22+l6OZwqT4//+
5oOlKQQkDt9BT2eHqMNzTUO0O3kc+TplbsZz1xbf/L+LSUsT0JCTJwwe3HuxMdwqEzZdz85Repux
630cVPwVafumXvioydBICc32d0+X4FjiS2Yte7KCJccORHOIm2ZXYpI6MwIlRKmzTDrN9i58WKbc
VIe7qQ1pfCn5yuQe9FDYQbkYWRxHikqhmEghLan0ZcGrim/TTdeOLf7VkFe5jPky6GPPHYEzrUJB
l+tdLOHy78RtIftpFvr0J0AyigAzOrPlgLS4qGx2vxyjDA1uDMeYJ31IAJhX2TvHdbjbl+8QTXde
pvPhb9yAveR1URGfwhshlb6FQRxVapSKYaMtQcMUoELqxOCtTkTBU8Gc+sCvLBVd+MbkANcgj7ms
KINImukhXMKt3bVcZS3np7a6AQVxRsulP+uwnd0jDhDBj8TippG6V16auFsFhm7NEcL6a/lQo7tT
cgJwEhmH3z4ZytZQXCMVdfbr83X7qCOvHEG8RO5tIlzSW4e/wYbTonzuDgkFO79j3NRmejoRfhq0
1PgTJKZ8R5FOby9uuKftQjfjmPp5Hd2MXtG3E/fYuwI4INRD+JKi18jaPjH8Uxq7sIJKwNcRczy4
ptnACawVtQFl3Wz/BrtRRmpK+V18LwWvFjFsrglkjVvX3m6mf9qmvCgwdbMvOq5n55HVzqFgUWDb
CDu62CpoxQKLCtTbr0AHzp/AzIAWordQNprYi7PPvSQ6Fg1MroxKt3s9wSuOIeZaOhIIQkXVvV1p
ggqiMobUzStyF7foG0tfhWCspDs0qkoXefDwEBgGWnEvSbmrxZkbto0kecJkzsSR7WaD8SaECYkW
k9nIngG+L+aad6rClpXMj3dfElzl+O8toOjC2L3KV6OjW023E1Eyg0ix4BlSV5SxoBrqRej6drtL
YUwAdCGILhDzUJyAODZFcu/hr6mLnnroAmcUS1s2Gxg61xfoi+SLWmVHTdtFnUrJODZG4knf57cz
HQSPM4QeKz6/T2B4i8PTg6i1nArDcV2SoaLZS3ar8jxxAGdrqoJd/Yu8C2+1eZVXQsD1M/fqEZqk
QUrPu/WXA33Jae6S/YK60KOhX9wS2fPnXEQ2HR7ecMFdrPFdSeeFIRGn/4g21CuwJjCak8p70o8T
jtBeNPUcU7v73fcNlx/NN009Y9D7Vg2JN0JWnqkrFdGRc+GVjhoLEVD8GXAG1n0/AnSd8bAn8urI
rns9Z5PAqwU5f3eGSNJXfSB006x5Ix8H4Ul1LZXEln47w8UvxphMTXcN6q4VDqTB60WbWH/ERF0+
Q/rombyGQ3BNA2ReMd/BLJi7gkS4Tf4tuLJTkvEo3adqaSozxtQPyHfpNVNt+Gj/hRu9xxw+she3
ZCZ7WBaRcyX3VbUZ/hYtFMKg8ra1KfGE1WaLosGwuMdpb9JtUk96od1PkeSUmlK/WuZFtU54ilHi
tkie9sHJ4UtQlQmojdEo8m+dfHxcS78YeehBpsImTdBTAmT1jkPN/sSy5xnx3Qb/PxQaieBWLiG9
D2wDrUOW3j4V19+J2hZUy6SzrAHBans1JyR2QoZsujhINgIiA0F3g58u5QLId9nTJU9WgYFn2r1/
vybRS9q8iypZdAn5QZKoW+wqQv/CaHs7wf/l/RZqMXBP9NdKfyuLk/xd/TrFwbm7BpWQyN88UUd4
C9LxKNORfL/AbOrQdl3kqq0zoUKQcJpXKcHtgZA2ASrIv1QrR54vFpd6kaua29Y4hPnnKYZEE0G+
pHY/VzPjdM9dMYFXUYYQK9xVxlzv6GoQqFcuKIz96kK+pfF9HUQTVMagfCX8W3Qak5tfuiy19WRU
w0ftDITKa6+RNQh64SEJqtAQaYFQB3CZICX9GA+J0DfTnEeBIx1jZ42N2/X07xq1+NzoUXTM/jG/
RqFPrDCIZNWVTdd8S9Id8r6YRMbMR7xnGoCqMX9mMNwpB40gyUlzd8MvxD7ANqOJsbbmom9QiYeb
PkutgU5LpWJTv6aQ0eh1Xk050S6hsbiqGpWmOmkmJl0Z8o6Hgs83do7xChYdic1EMeXLLRY2/M4/
k1QNqfTXwuu3dX5vnmuw7LqYvKRHDSMPDLQAnZiLr7aP8yekU5keRzz2MaGP+ViwobgBydbzUFAv
jzxphMEPDkxFpqgsgvP1acEAjjfrcM+5mQE8knYxtnVwdMsRQPF1SyadPw0FKJe8OJdUPAIAVQUA
t8uAVRlkR0qIRe+/sjQDwAP4Q9kv+BPPMKVh7vEmf/twRpVJCUwWrApy20nXqvLeKMUJWZWnUXBO
MBnMiiLl+g5EJqzM/xt/cET1hXt33LMtU6UCudqDP6tH2xjp/kgPQFy6aMn24Z7CrmqvrT+BNZfd
LaNfN5hroSqKyX64mkQvWhUNhZ/VQF6vwMIBE5Ld1d18K0WWiTEuAVvB8IPaxPhpLlhOwrIcmlhk
k/Kfe5won2GRwLRF8GawlxMKzXW5rAvxT0V09dxJbs78J7YHZV+UiWqHWwzA6VA7Idl7pIELU+u9
Qk8ZDsPYTBFkLMV0E62XoJI17gZCuLMxf76PmjAJHNAvIKS9506kIzY1SPpb3ixsNDzFdcKDz/kt
T0PuQqUV7kmgDAvy3AntG0aJ88qq2bF8EM1TbMG0wl8sxYBV1wzOmwgb5lJLMj6J4MZXLnqqgmVa
iM7b5rhLpje7fVyumBIDZsgRNWeeaQif/QiIJ8eyGsSrjWP4TP3NIbXtuOQRE2A9AtMqCVNqk01M
6kA/Gk3Fa7uNWlrJ3t+MUBUnXeIpcy0C3KIQCZkORBzHGTJTNKNgS8MUcuQ7MYcpuib95l96GLgS
jX+kdy9ybAWYVcJZ+FwqyJOhV2GS8SysyJIrC6XESE3AafbjFPHAMYDL7MWQ8kLFa1QBmRns/2cO
OvOepuZTIDfcM6wiVTSHKY1iwwFwyj1RJHzE+fjAaWdEEKAm4BqLtqcPaE9gsMH8YLKcn4V0reQy
IQWrhaTOpdVqUhzTwXV1OrBuc2emd53CH0jL+Mn8hr3YQyxAfSNapL5O0wv/YNazHROMt8HNf1XY
Lybt90juho45oSS7TbLPEvXVSEPp6V7rRJi8bsSWHaNSEHC45a9KqvPkYMtobJeUYNPPed7f99Ec
6OK9I0Yv47VUqeSb5Ko6wkfk9gEFOvjvUgXZP301zM1c/1R7qri61Yr+xG0FCzsEUPAmsa0Ba/mE
TGkLps3bdLFzg0gNrznX7YMwc4bqrhCzh8ZCWKFT0/l8ghQpk3bO2yvdg6wwI86hFPhFnYxBVcPv
CLtHJD3hrNJ9FgfHrLEUgLC96oJ8M4xbg0sJDcTKFULp7qQHFH4AXnISXIIRtGqNii6tPpCgv4U8
84LCVXQfKA7stUm62ksdctCHo8ZYry3ippKJTifhMuYr2N9Fqrgj7Q/qt6/8O9butTfOTzgwlY8i
VdVW10ztK3u2x0c6zxnRV6YEccvrwW90blSPI1Xr0sqXcOf9zxwRN6+MI+1NnZG5avjQXvCZ4JsF
XRqZONUwhFiplIJXdyJ8txo6nXTmdL0xlYdTBE0BcRd9IrS31g1Foia7/6M1q/kj82jH3pf4nuc7
EwTOS5QCaGSoSpcDzx7YRbqMtnoclVbBMDP786z0COsd7i9Xjf4S5AF7fkm5JDjMNSJmw4IBa/Ei
RIt7UugvDlTLzZhVs9k6hh86xH7gWFUwII8YvZprW+bbb0rgkMjekpRCoPG5cMT1w8IS4SA8UtLd
tn8pcjtPQk4DVi6VAFAKS1ieB/TusPSSYJIBjgsjtkb4cY9HS95rm3qvw0gKF+1sbOJ871ArEILO
EF5LPbPuxT2ieiP0LMALquoRaQYnZP3Va9vqdpAOSapWGjxB1XzHDc/gWvrtrFJ3c/yPm8DiCX4/
pYtZvO/XnJ1D1AVwwghkcupR90N4rrbaF717VJmozzRbG7GSvGx2f9WqKAUwCcj6CzFmtCA1xlsv
Zpmay2aAiE5DCyeOFaUuiMSIcfZ2il+hyxfcMxDSr0DQ0BT9ziraqbGuH9lhIDUshxo73XxlB15P
3vCDUDVKhSdluxW9NN1Mja8wIdli1z7CrmkrEfZyhffgMtvB9eFCQH15ji7M0k43QI6MKFfWExbm
KrDIq8rCrPg0hZIHVSfvHZSSwFq/yr2xCUeJMwBmYaSMxRdd4omzSwVbsSGDe66WzxR7BbXFoEVu
yRmJXWaxpWOzXYj6R6WHnFL4PdLsfSc6LrKNOuA0NGooceEqc5pHQz8dejQBTQ3kG3vRtA8CTPWK
FkWdhlpOKpyW1Vq6MziJnMvOZA3vhX+AUg0qmlGaVFqbadZ0BCOtNuC5Kl35cDPOAWASGBPaCDCW
nzw29XWCCpaDDa4eRnU4xJHk5F6o4CObfYMrfD5n+70X4tmEYJkxeJgi5m3emCoK8imdKy0wFmrm
oHctkpScNkAT2D7HhF9CBzv9bARzojqSV9uIK7CjK+bXw+F0fAbc19BM99ZQ2AWnzzl5HLVRkLNv
ofH5a7w56C6n/NRFx7/wDlaYz5M8x6vognURFlrU2Rw1zlJj0G2E4Tcn84OKo0aI9A9B4RBktkHB
bhDNnO7McAPK0qnqupGN5Xx+atCaob2sj6SQIom3mlqIlkKRG/3Xgscci9zqhdIb/xyOpSIPZaE5
Q32pcyCexS4S2aSdTAGmBSCN1UNmuVRJDl2qcSycv+ZmEzF4QeUc4hHmhY5WBs1ECNUFJ4g5M+MZ
2LWYwUF5BaTN/QauJ4RQclBxY3ZArgAi403mohfu2IHV9+DmIHPNZ+BSXkeW0A/F1Qt1BV34BDD3
gOIU3dTI8Q3JdmZkAi5IIByNmuvZ3KB7+zp4bwUnrR0E/2A6nKLaB/qdGIgn3Y5+loh4zgt89SiM
cnYkaX0WTQugv6GWQJQ01WPJAe7pfydmLc3OZsupKb3FlT4nWDbBMugqBZOv8mC1N6iHOZQpP9E0
Whmq/HYzg9PeaMCuXgUMvWazFvjH1M9bFG/MSRAs5mGY2LU5LcR4Zce6d5YScjgUUniQ5IhSuEew
3lc9rWktS5SX9GM4cPe9IqGAttm0OfIos01w2mRbCoMw3Y2qsfu9ssbZ4jxIVKWoF8opIhZWfvUA
mJFudp91kpJ/2tXzWJtv+deFI8w+FEBkS1TTqmYdXRIcMpGveVW/juOYYHXykp/nIKTvo60FlZjN
QusqOHDW9lAHkXO8qyZuMZLGYpLF5ac9DzLGDHr2CjTuOvuo76p6nzxj+VuHFgS82sAJn/yQWxMs
WDDlMXb+9Hs3ha3VqlOr5VsCJCVVh454GV35a65wLNlP9IOpyZXPbhdNQIGXe82SYAY5f+/4tcNm
wMjTWdWMQtmHD1UazwsmkKDZo+KGJuTKSv2zmdwcABA+tdNSD4Ub8G14p8JUAS6eo9DJoIfNLW4U
D68i4Tsj4bXzsLVIPIb6nGmjVeE3nAE98mH3qwl9T2h50ZzgkUmU+4+iMCLxDZbvTYWUoZQxNGyc
qRmyfyLvL6OtmQVyD6y52rqUOdBGmhF8lYXKUFVXb6Qaq7hEBBgdgTC3vnm7T9vrj1JL6MKIewbD
iucovdAk9uiQwieTyCU0mcUJFAN0PlyRTU8c+DIlxbLOexPChrPgtiOAyzNV5cQxd9vpLFvg3lwt
4PSZLiPgL2DRZxeR7GiDQ7ar7tt0bj6CIk6bRFH8nsn2iP+0XUlGgbgv5KwDUCtrWVEe2UwcDKMv
JvUB+1zvidX77BhmYqhVvhERV6kXFHlH1ZocVz35Yug1vvqcGiN8IZ2nUbq4kKfgTGv0U3cpHwe3
+NUD47A/+vUK6wWvOBxwe/t7Yufv3Sy1xOT/1jTag4p+kuV43di6wAT1/Lj6kG6co+OlMVhYmhX2
LHX/grnFziG745P64/mjvgSdqWato8htGupgHIlwD6URpMkk5t/AO1RcUbadCgj7kNBjYomqNNaf
V9oll1oHIX/S6TxT8ZyS+kHvfQgqIKGNWGf208D1Ebf4RaHo8/g5NdPHh15d77Z/0o3x2qcNJ398
xTR+NqjiThFYKhd8GYNKq5pYxQQ4RlKRxL76yaos+gQW4XGaO/jlrq8krGgkW1mbZVYByxPp5uzH
nlWXZUNn+XoIDD8g2ssSpHGTZOYWLD4rbv0COykri/L+0pKop6ujrW7L3fQH0foBXhO0qNq3zsZj
204TY+tFxqdE4NuprL2xEiDKLgCma8XjUq8/C8u9c5Lg3MO9+PSObq3sU4/CjPIEVF4YQj9GjRAW
NgbrwNf2R/5ZF7mtwaeHgPhtDv+vdWOJ+YW7QVz+SDZm5P4OOCLzRaTyarhixh5QqVHOL7D4Zuv0
aYu7uKQaPiGzKa1VoLaNphP7458StYmwFk4hloK8bjTDycv+mQCsAmXLvLgphdBX1s5LXIc/nBbM
c4v53TpBZUCjyCf9lH94aH/W66yy4V5QunGdm+K15zGyXHCBDgFQ6Ap10OGDkSYp8lGPwJ7EscQl
bKxpT8xg0MMFSxkBZ1SheXIyKZl2v178SkA4D2988ir/Kv45BMfSkz5SmT5xAzPz37KFFNramQ/N
Vwtb+Wyxlk4GLdKTMiHqQXN3K4OsDwtlvqEdPpwos1l6RN2MWdl92MdhaXlQnR54Dayx9HaZZc4g
ci+2x1EDm0jKRX2XoJ8udd9/M/opXK2Pqtw3yqYHb0E7znhSkKJnIE7j4VWWhQPdoHSbvP3NopxY
jf0eqMbGoSjdyf8izEjiHAg13qp24vaOBpm9+59VR0OWAHAqmKVemLtGgRuj8D+Igbqcf08aDGLE
imYHy7kZI8rI53RO4ZJkIuee+VazFPP7abTf0RcRmhGuHCp9Qr7V8xhU/UjbhKi4pCM6dYD0wxmj
ndogk2Vz3Duf2/NQN00ND/7uR4NCWqfmBjMGpb39muAsgRJznpge3xxPkWKE2gr4IePz3DIJXt84
zRO10dlQuK4cUWriWWIAG0FL2teMIXH8zaIfnSVrjYUcYfv2xv95nM0TqiAZDR2Q0xIFcDZRr77T
sXQnNBQ8fMz9Zt0myQR4SqnWYKL1eXsMzRnB+VRuIHTCThbxdzefS5hHQsBg1qfYmzhHV+Poeh7v
P0+zkRzevH4+E/2vHBJSlsxP+ywkecyT2aD5b1i20VhnRyPQsLHEsZCdu40Z+9NDYUwoTx94h6jZ
vZ3yzmVYeY7NLdSjHg8UDEhIC3N91ZgAp67seXs3xDn9XLDXyCYNJbNtZ/nSoououvelLwubfmjW
sJH5Nbc4/V0OdrnGKrXyrjHgJSH4I/OordzR6/groL2y4JioFYugwGeoyyZkPwPNcM5Zp84Ha6iN
l4rSKes8FyYoOQZ+QzC8kn2q8v0e4BBMnfHJIhpoSZHqeQc6X75TSSqHdq//dYL7dhAL9feNLHGZ
quKiQ17kB8Mkw1yKZVnVRDAyTbuXT6axLel+B8rj/Qsu1fKKpjgGjMstJEKgl7visKJxdsA1NAYx
oZpGZwuSfiKEqRsoi4dqtcNxZbtobmfi0ixRAoM8h0b/zOAFKJIfgbaJJh73pq9C/HOxRKEuTBx7
BwanV7ipUnlB3aksrP6BjcGqMGqJygCwzBUjPDCUEGjQwH80tkPzHHIVjgocQERUkGmfkb4TFex2
1dHTCUURKMeghN6QfXD96rR0C3e9/Wov5gGw/Ae47keadRKZwpdQ+Uctm2k1EIsQZ//Sfwj3l3wy
zP0FxX0p5t9DBemkgnRk9wKx1/oa3wx73Z9ZnpiCA1M0cpZQrB45OpOj5GcRHBt/qeiG7/GLlmgq
Yp0iTjqRJDOGpjfTuWvjqC/iUsaAkHI2q7qVTe4Bl5v7iWTLJuRQyNUrKjmHUfsnYCKbO3qwKrF6
5/b7OL7M6xD92MYy+inUU3smk6uG0+/soxLqmWcgrWs6SjG3ifkzPDKmoFw4XP/niuWbRJAVYCOr
nSP9FQhcZuNU+8d9w59+n2xEybjfMIgPhY0F19Jb25jWVA46uXLPckmUuToaf7/7Y2E5uUDAXvyk
FlG3EWiRUPJxiK3YgUSVq7upMs0x5b3wuJjRCKclzsrVMUy3zDMz0VKGZkqWdXmkhSbqi8F7Z8IH
IqqvxT839z3RejWxQbVR3upp5N4Wt3iPeo6VOlrMwwCwZXcPuSK//dDTSgCG6DWedRoSQTUQywVv
/6iEfiIUrEoB2FQ1h7hdEvyZzJ7M59wo66KqMfUF36uJ3uiK0aii6brZwoNXpSh/2r4upClcj9I5
dT8hNQ1gETQYiHAytlOqJ37fOQabZ1yv93r75oqydmZ7ObdjLc04EO0lqy8UAc2GL9dyMuyirJOj
xOnEJG46bp15hsiEb09j40PixuLrSOyr1wM0JDFdK155BiHWadNL1zLc3h4spVQLAWYHqFRXeaoi
dPcEnei803pDu7/CYcDLvxu61iKfgg+mnhv2qA4omc//FmjwTC5KMU5cSTpFjJVP+syRU+1mXWaq
LTi05cDF1US+mhhHZ5o2PKhJl6wbi2tTNa8oK+Wd+sJkUqXtkVDg96tmjiulmbO3BDAqqMGUdxpE
tCEHPRVpW0OF3lJrbuUMybGgb+v8jaWfmWk4xEw7Qj8peEAJKzk3ovBu5ZXODdoflHM3R1eE7n9p
VXt1/rATvXHamj41yH6DdWwyCwUosq3fs5fttxgmVaIyTG8/cVETGRNPCdd67pRvRPpQO7k0YMUS
vlwUxGIIT4uy8NgFihBkZl2yV5U0o0R+uBPUcdnOtgZDDjm7SzMrE3simv2Ik5MlRKnZoeGsJw5B
n8HxBBSEaIv2o43T1dQAnWjDW7JksSTBKxHg1OmG3b1VH2zBCyxbMqbeuz9ZQE2DP/XDxH74RHdF
4VUqt/fx+Q869o9DprdM03kQuqd3dvLR7nR024vEa40qi4HoG5OUDf4tD3xg/JCpnNn+HjqBZOR/
5KRvtqzoolwfQVLwmwQUxP5R47Fz7bs+zZ0N4OZokeS6j2aguPJV7mtUeBVWlpqwRA9Ea+pkQniy
nZvhck3uQ0gSKZdDYUuZaD83CcpZ2L5ILCL4z9JMeMc4CyQ9u+eNoQeH3tTYxznAhq2yK0+75W71
ikfCOpHSnFSVEACDO+RVwNpRBXglQ6H47jriFpjIJe59WGij0YdEdZ0Y6+j5yJxghH4MoA0e8wrK
F/VIq2PbqsoldtvwA/zP+uLNPDu367NUuk14wTMSlY6OEPPnyx2f2kqYSZwnUCEZGAMCUE7grHPh
2Tz4nQvCnr7RCHapReVjRGQYAU8LHUHv9amatK6G4BCWH88U4Txpog2k5iasHknz7RnhyiFVYZQy
UwuDaON5FV0O4Ul+Eh+Kje2iSww6BwOTDiX7XTCa77By0e3VzXHNt5OvLMUzVRMTgvl0YCfKcvyE
45YKFPN01uhaWCpf7x1rppAfYbIDq13+S+mIy1FQnKJACXg4zTj0klPyq6yU4iFgnxOTXtZymJyp
ZkUIilDJraws7WV1Ow1+8Mk9WtNOhkccLkvRMgumbmAzE2w/aWCnEFbXUluxIGr6qr7RV8uqGOb6
KKurOSnZNI2zAWc4FNhPI1hIopaYzMS+k5jdkJaEvB9aKYzYZKv+sFfIuZ8oEy8UjajG4TQo+1RX
1/9fAzo7o3BYAS1T/GL7Oy9kCWUDKOdAgj1YwuFh40mJH0OJSG1frx9h17A4giMedfZSwS9axeDf
zPF/nbPqVEVV4GqASMObP4mkJFwA/DmUGQn5Abbvj5dI6x0touNDMtMwMjI3Bt0frrRMYIM6rhPK
UN+yhvMYtrHcImn3ztQ+1sDT+2y6rY1AN6RKgJ02sdaUNPZmtukM5XQrlWExVhNo3QNF7kINgONx
aIgglwgGl17fd12JoGDjGjS4ALsJX4oWQWbr1Vx1cLc9uAf11m/ChcGiOSjbE2QeGDdgbr+yvMjm
IY3CVM65GlxNWUhN0rjDiw/66Kttb2V/OpvHW/SAxT5vBY3oz1ZIgEk84d1zEa8NUSpkwYO2gwhv
kDFU9OMD4IQ0Dzxk+Rk7NQoRNZZdGSilSC2GM9NWFbkn6LolpCkfOxa+r1v9decFQUA+9beDNIuo
FzjOWSOZl3cZQB8fyRU5KSzsRiOdYWzNk+5xIKu97syEpES+a62EQrSlD/axILBTaO5a4yqrGKbj
UtLwyaVL9PeHhHTvhfbVZ8vTGlhTQnsRltjtm5pD8GCLROfu67q+li7elccwBxh64ruiSWbHRoGC
3cteUYS3j10grP6rP+I8SRzubWU/9de8tlLqDmokIh4v4oICJ4TXuQiHtNE8ODP/9q9Haokc5JdG
1iJoTxROeXzkpXJ56yYcMIismLHXDllsSYKY5HmwuTSCIslro+pUn2aIBXMTNIqscWbJ5Yjc7K5Q
wWXWxA0WHWEKd6BuAOZI3pe3Bs+ltvD6mjAScRbaWXOmX6whUmj0PYduXNoh5i0EiDH1f33txB/D
oflU7cLdIZ/PeEQCy2pulMr7zmbbdpE3PnabCFytNTPl3RJFSfR0hMXv7yEsNiFZXRPjOEMLNzja
H7Fqy8Ixz3g7qorEH69ikB/uKHe3X+YV2MqphudVVX0imgD/rfvQQ3J76ztIEu9GpJ62/ysC2/7D
Jr6mRc5nbYB8gwrsEyQwVRaajWrFLNiDzD/cf7rFHds60JhzBNsqwMa0qu94n2paqMa2pu3AFxtS
a8GkwT4d2P2WhevsY5JwihwkyvV9Sui16ew/M/8nqKZAap4Ck/PtOtY77IwmdUVX/uhuK1RRhZon
2sTWvdwAK1lAQHWdw/whFtkhNnGa1qYfS7MQKmtp4JLffAq/fLT4ltTHKk82jbbd2VLpG1T2x1QC
L92p39WawuX2tK/mamnd4VpKwLNEpHvx3nrFkYcKQw4sYh1HEK57kOGopHLFMqf08e63DCRZKrzY
xSffIEhh8S+Mu6D0CmTY6QG0NtO9/jdMbJBboHTw8VX1f+PSHKqcgg/f0XuH03aVcNYvyo5yY5CX
Vo7Dsy978aZqA86cP1cNLAKMUsQz9IgeTQJMNuy3Bmmuo3Ymh2zisc9/w4+KL32RRxF7e+12opBc
ZaUTK7QgXPhrDNFfhOwuKq/aNrt/fA36/G1g2DSlajJR6bIwI97NdtfXBZA/SDoFpTCIAU9uJVJT
5nalTLTUPqRzEzvo360k2Rs8DBfJMfGwpMo0VRCuH4+Bw0jFVuDtsPPVyjjZiw92nNpESBZ3tyNN
3mhbU2ptV5gA5V3RY27X5Sv6GIHJyklgSYfEPKJ6Tz8XPtsXPu8BrFLgdgiq7TS3b0e+abc6CPbR
x4mFuDrhUq1/pOlslxAVy4qgaabX6zMvqzGrBjlYJUT1LFdCteUMkNV2qFA198L9rQKUzz1ysvC1
jOWulG8E+KfrWLhpDfS4zDb6udzqvbNZsHg9uJAQyQMoV8Y+9+I8A7jyFwWfTduCG6qi506sY8BR
Vxjms80b5Wl5t3FjFWJ0C0EIBh5lo/56hedY9ZTeXC3mMjeJ4YSNqafaw8h0ATc8Wrz3NFd6ZVh7
xBeWqzUCKIq8NRre1bszUemi33440TQXj7YtzTnedCuxV/lpLp/FtY7pG5RNC8L1Hw9/YVPs3aJm
0cHw78BZtfusIDSraeiBy9pLoLMZXLRNxxcar+X0iR/oKyqakEIUWFQ4fSirMyJOsipZgb4LQDml
SIp2mjpydpmnfSXqEWUJiqDufdIm7chdTDjECPbSbwfQ+QiNUuV7UXSWaNK59Bbjab4Rj4gdkac4
n5nTwT8D0D7qy9qzN+WHAGDDEEK+t8NwkyE7RUobqe6DqV5aR7oRUwKhn3SFLNHAa4I7G4JbddA7
KIJAT6rrwz8bcE5tzvXTprBB0wOHn/fo/L/VRfijOcVfP3jxmJDabKwSIuWpUE93wWT8N5U9FDTv
/rnaBHLD66U4Db783vo8z3+tdGcN49SnHPGe6byNGVBX3BKvp0RCLr3gdpDFpaMdlB4aZ4y1zJXj
D7gmq79flnPUD4xWQWIDH2XT7OpwVMiKFmQO9sysjECnUsoc8XYuDF7NfFyH+AM3/tMbCRdwaDHw
HMMbOcBBVYrh3etm8YEI02zoUmNl2oLxHwpMXzmGmoLZrAJyOB9GrtoVCSKhghRP6d6AcTNvBgP+
PiucD0DAX7j1zry1GpGhqcprVXsMOq+WrxTkYyK9lrsslXdJQNnee33pjb+fI+wVe/yVAHVH5nto
R7Mc3SyTFePmPhyR1DgZO0MyeZlBzJtU/46u0F/EGlxb8b0zjZjyPFNeleJaMlZO846CfI7BLnKG
EH+n5ISxxDIN6VBH++ciSO6WvVHTI7sgR41fBXYT0Es9vMxsjjyKHnqBfy3rIQ8W0hczIe91CEsS
CfDXPNkEU9DzWn6Isb7K0fBrslMMpldPAo1RH8WM6D/HujaBL98u6umgxo6/jjy2clvMTUJBF7p0
pv45F7+KbqGN5/GyWWKLrl6OgipsMEWdJuc9eR6di7FLqLNEk8ce5+BEQUKfKJE9Do0G57yMc6dc
XdS3VaP8WZJIwmJsiKW36yKZ4EySBu5MzSNWu4dMcC+RSTAC56yUZ+QggiCS09jwGuodTJGAVIrd
oYDmvv4kdB+LLs2XjiPzENGcRjEQtP8eVBsCwA8OFBBvK9VpVETANqfQy6ZPtbVtWPzFC8F6wl5L
RBSLgsN4yT1z1qYs0E0Awt+zEW5f13lSEul+sgSzQnh7Q/XfICXWNDqIl6GCyRv5U/uNfQRjMG6n
gBfmRyW6CvpDXkuYDUWO6NMr7QlcAhBzpabmdLbWipHZtJ89O4nnRXsNGuGU5VQp658QSQ3n+By6
ORfbUQWxR1p+xsr/Ykxcrq2h54XJUxBO73AazjVpmfWpyEM3Xh57BLmzoUcQsvkTINjnIwKXIVA1
8gQm/Mkwcau6xUn0p0c98pjK5w/R54Edom6UkraDDxgExjg0sKlF7dWXviYRnp3gdtCtYAK9wEuA
6LB3ynR4VP3YkgN5jzrb5bTPWMU0o+HrBdxSfp01Fww/fYYhdflzn5KVG6DLu6r40QF1w5bE9kHu
IsnvGCyfspww4bNUm5mnqINcoRPLJwzBPrpQ2ReXt6KgB4sFS09M0gqJr5XN6yru9ybxM/WLLfxG
h7sI0prRlmgpaJIASX1k7oyBbKhbEtFdt3Vo1aECnQ+zUQH9wi9ndmcD+kFtOZ7lVXGMnKkxREEM
581WpIewxln4evmJo9VUnhA/WBinJmZUBbeaSugU59d6oWbBPVe5Njmpty2eyFDKrh1nbAoSyEsw
kjTpkrNo2C3mVvj7Ga5pxKCJx3xMfFyaXuJAGSKvyMCImQSvYWY/mPqlH8Xiax/VlEElMQxxeRp7
rLb++lmTRn0yKostsGBQqL82d545ldgaYz4q53GeXJgvFe89pbpzgeL34TLWDIXOMLz2Tlec52nu
ZRGsyj6Hi7yDlrENcOf1fquxMMcKWD3/Aj/xHzp61rJXlRV45QaQMDCInTk2ksHTnHEt0dynF9ks
D0R2Li6fToHX8VHUKxFMkIhnFePPINbusfwumjidWVnRhshZ1ZqXrcgqhVvMo+OVgmM4TT+le7Sv
H2ah3nBHx+GYxpXqoE0amlLe9a1jAehBWuP4dI/zpCZ7+QQwQNdY1iSqC2X4fL8HjLS9H+xIdG3Q
u+qPfh+myM0uFPfI9dswnSZ2viJeqsPrs8lSG47AD+udU4S+XVa1xKfAeZ+Bfk89XcyCFKmg5Bn2
HfoG8tvBuem1lJcmwqMQ4oiRw8u7iXMz6nSpXYb2skxhpBvSgjIFeu9wUMuthaY/OWeok9v4+GA5
J7+4jpIOxTRPJh2qPg38a//Oi/N2aGeer/l5KeK6x+7FgKvqGv6PBhiPLqjgmVwkCKQFkymzkeao
wagcSdhf8/kUT0ZZMr7y14lKVK0WzKIz1sqdkSXXK9Tt4vXUObv2wMC+lXziFFsyU0GIJTx8ada9
WIKMaHU3nxLcBH5OD7LMctS5ztsMe9anTxJ040JYUOw0Kor80BPBw+tGajTCMUw9Xa8ekt0fB/Ok
zK0kxPvHVO44e1wBkMm21nESX/v2hrFCeWwmaKY4/s4tTrSfXnf5zyr1cpfJ3I4JlXYwnN98vPLi
XUtFjmwElgM8MtRK07WVnTIRSWyGPCzeq3r/0uh33jM6MqMIj5VNO8xNsal/rsczZ3MaeiO1I+nq
cfTuZcxdjLYCdXGdaPzBWhQeKCxp7FO0UbeZUL26FiziH3vjpn0cif7kCqxvb0d8oZN17Fph5uUV
mYCnxkLwKihbx/j+3ffBWorp7ikEOVsRtGbggia8M5A8eK+yu+IYCMvEO/2Gyrrz/xzi/VKpCd6Y
tsRMv2zkEeCnNCcuss/LR1rdJfqWMKWfh5/lYTS/SiwZVH8gdZsxGDWElnymau0dduaB5zaIuvuB
f+oGQBv2Gqd3MZD1jB+NufOTvG6YKUf7V1Z9Na29v5lq05VxatGSodPWLW+Y3/T8DBgLCuTbNcsL
vxFmaev5nNBn8P+KgbGTIRVx5eoDvY3X5XwK3X3JjO+clHZhQLba1/8wivdcKTLmp7HaBUu7n/2v
FGWoDPwlMw+t8p07e8PSiikLIbskAO14ZZCG2h5FHUjjsGMMalG3tFX8KWfVes39Rsa4wMsp2WWR
3gRmPEWbgUfzboq3qRHSsaNR0vfZIwbksk+P0Elu5xNIZOY1gvU/jwUjB9A1gRZfRyQbAJNJ+Wnp
D587IjvF4BqHaSL9fRDVtiKiaWWASwqpUuSjBExvRaEQ+9fuMcbJOFdqYp/BlYzBgJyPcVnwPvY6
e5W5qUaipZxP1yYP8XdQrbQHtFYHgVZHmpxSAg82/nig7R/s911SQf1TqBVeWEa3cT7ChnqUVpb7
Yrl0HSe4ZgCpDYyvY4rd42q5b3nrYOvD71c9t9ccwcbGkfqMcSw63FYxIxYsp9iaqYeGL1mp/ifV
f1wZJ+2eZXgqLyk0Ixc0YHKev/DOofSLTsX/XnUy3wcyIenE5LE/cYAhAHTUVZRkssZPeLpSJCP2
Uvr1im6ncDO5osYzbsUk/k83EcHmhhl8JQ590Efa1zTgMW/BXuz0zA3xeAs6LUCp1GJI17FLCa3b
o0gftmlizMJDqWy2xeaNJRjvWFzPvDMdg0IwUuvJ9vfgHXLHXShZ0Jl6hOv5CCT5kkMGyD2cGHmX
NiI2H8avY53t/BI/B/YEzAfEiP6Gd3AMndaOp2cKy3MOYLBQdsAf31FNtKEzgZ1zc5AU09nepZOC
VBt6Std+WKYmEtfatjmFVDWIfUeQli12OEizvjeYwQXqIzU+5zD/7Gy0pm2WNIPavaO/yvsOW10S
rYtK8xH3+70eWjQkYGk1jC2RWKVX/0XnQ1oJ8ks8I5PQRZpjbhTE2uzSeh4Q51RtcndnDGpCQZXa
9O+aJ6RrKimARqwzx+HTHIhMuBRk52nISmgIEweYOqnJscVYnRAfipBMoOadOAEvMlDTIhXA2n/t
hN4KBs9UN8utLLt3vi4C5dub1zCN8w86ivdnQLvyzZEePG93edTHAI5GK0/7/l65uqWMzMOyuQOK
JHCOS8OmBRUE+WFcruvbFxVomLOROtgp7p/DWZBVg0d5I3ljBAciK9x+XypAgtKyF3a+QqyLx0qy
ugWPrPC7Z/MMAmLk3ZOHkYk/qCRwAC+EMWH7ZK4vZlHcghCPrUDzAGRXOj8V828gCZm5SJkmIqsK
C7k3oC+9sDb0Z0sCjDctwknuQW62WfgjBvUtCRGwbzAN8opqW4TzEO8f7eLa6DTZ5QvWtz46NDid
ERtgDxEFpklOw6MV97XrXT2gj+8WpjrQkfRhvnz5d3a1aHbkg9/FoNe6g1biNHYsQaylh7lTJXK7
Pl+IbPKAA0UxOg9boHzmcAby7P/1RUj0O/VoTAYksQNENcYURiO8YaxM46VmEwQL/E39wUCmpJwp
2zoaLP/eDthI6m6Ypzt5gHEJwQljvO3v/Qjb8x9Gi7C2VBA4WDa+5sk+U+dLrd789cbJktFTgDyb
OdcQw5yDfZtYHUVAUuYYz9GcXvhfhIzfLgGZXra3EkF/3Qy42mTbalbgDJgRr6gWyNoX436Dr0CR
Imw1ZcMB/t4OswmQcxzvMIxfMvWCXLbL/jGG5TscI++3FQMS+fp+tnmRgSz2fgetmq73XkCPajHh
5ii3doMH5OlyTAHAT+uz/Iq+yPwHdsHvA2aXfhZC/VT4/oNICod4YfruuJ9HhmrhWzhyRgnsHKLH
e/bKechE4QEoxrDdVbjcEaW69/yS7VEG/G+KhzrdEz4ema0VGMe65bAtwm/QfhTDZQwa9zOh8w5M
STfO+PdysnjI6W+Fcs5TBMDOe7kIciGuRtiYr99Wl+46Waf0AjZh45zn/cflzVd4vEbzioUL5Uag
P8K1Bby8Fmdk5uG3aRfl90Bv3MditWwVaZpJTmVELgjRzruH8WUYpzKA5dVT8RLjAeLaGvsvKYwi
Yjzq3y57yYCd9J37x2sTaBAI5dCR1RPtQcrfKiHa6caNvFalxiQBwVD1pWJGurRjZlzhHMkVacow
cvsYw5Uo72GCUEx6lRNi7jwrsLq8Zm4cOl8tcpgLk3vx4GNvn7kbz3bPwxFkGTw+5hB6T2Tg1j88
lDsrvgJ8pjsd9a0AFJS4w7UXyR9Dz0BwwOBSb13MNukzUPcYueXllOmIFhvabHtPD32V1ml09n2Z
ObKry2YFMZwmSAQ/XHk29A780QXw80IsQxdjjG3rtxzaiAJgqesZiLELP4VDh+ZlnyxeqOmmzEhY
9s8dqWZ5w24KVughy6gi7FNN/hKqM9m+3tT/bEGuUWgn9lEO92IQ/gfQB+tcY5VDrq7h1JCvWWKJ
U3L+N09KpikfXgmWoEh7/vjR4oHwV+CqIMr1obJN7uuF9RP+sz6K8kg95i8HE+faWmUjbHLEQFvh
GWlXJargk4+zV31vMP46BBePZ2bP4GHWFTsJ4bxDTLEo21z7I1ArptPrUnd+D2CXy9DXMUZrqv1Y
nNjnaGt476tL70XYUguOq5wO2WUjDjB4gk1YGhbwQB2NHyGBeFYDO//wNrUYLRcqD71st9BAGjuF
Dz1bvP2QmPhfEsks6i/XixDjaKQ5ck1ZBdGj6F0gbUON07jFe5Yv2Xn5ZyojGPG7pb3GcHPTnJWq
wB0craAzZCEBtvgrqjgHgEL8EkF1nWY/cBYRzsiFEYKZBuNoHG6wZ10Ia/OSy3U0b+8iVw+DAckP
y/1Xr3rIpCZSg39sPij0NmMDhbqm7rEnWjX9/7hu8hhdvh2jw+V3fXgHZczlwy3V137Tli479cpy
P7wJANYzJK+L7SJjqIq+rkVdDflUccWJuTBjnm2ina39oOpACKSKVerUWSyTCcBKyvb/eR2kxcMu
MePLoTi9rvBhbl0atbiQs98KR682XS7Edm5SBCRuiw+Nx/82zbDvQGK2nntVxq5g/Z6f/p2ZHIrO
5WRbEZjvq6pXTCqUU3kEDkVml3/9qBQABzcs2/w89wHhLLHvuRx23CqeLM1eMtHR3v6Z6KR+2iTA
CTKCtpB79TAhmpemYtZQ6GzlDQFUuSVGTI0mIIindH8GQZxUxUEemlK57Wm+6LI9ysBzq6KMBORJ
YBeQCa1ktab+qaUffYJzzghVVWHCHUdprhvDVN5k2D1UCM+lR3Otk5lXIGnb52bRv7RBwnaU+oNC
wZ4hN5wpQ6jnwD9Pa94Te2CFI/QIs8OPMZ89AlwvNpWxnm1/ph+05K2q3KB732Dp7Wwb3QB0OiZK
wbGLy8ZWK6U+sk9h+282mgqOyt274D6F98tWQpihMHVUGeNIsGjUqLQzgGKPS9doWGIlGcIGtXHZ
Z0EtLQ5ie7C1U1rSGtjowEqrpEqDa/vXXCctjxQN9EJCbMGllCBzZ0sTTSVzVPnN3QBvVHSXqBlA
KOzgOGy1ilscBT1BA4FimdpM4+AQs0F6uCNE2lf/esKzizh4u/dQn4zHPzvdHrpCGhCL8R8b1BFT
huxyXSSxbqRM/xGC1Q6in2xmM9ks9Z/KDI8ZsdwmMIgVVn0sGh2tsdBBJJWEmV76IZDYz5cWIl/l
VWkuMlCp/Trg86XZDVY5WZeRWoaAVMuzsKZv7G9CnppKhzg6P07BkhsOyda82VLIK0A56XnSLDDy
wBVTSIqnpWatVkwrKldKsYbbmtZ/jAdN+7uAlUNIm3sbjGJQtiyqtSoWu2UUxVktKC0Sy5N7plp4
S04gxzzxPLyUaRcwIYfoPQCOLl6KNE9hQa1hQgAB1SVhNtwSxTMxgqCP3qfK/PtCpoh2aYkwIqJt
7meThpaShlicw7vIAcMWgUgjSNLwV4D4XAHCICfKuTuQrdsVtoJ4a83YZd7fW5/9WaEYAZNdNPH6
4t/wM5Ye8CpNQGXA7l2bI1Ki4Yj87cdD2IN9NjGbCgYiZjcvahVO2k/M2GNQYfkEfcQUThcISvmE
BxevE7JlZZVUi+vw8/T2tz07PdNJ31hw3muT0fPY7oXqVnXRKBZGK2A6wf21WjurcI0pfR0yxhEX
Qcw/ToMVFIk5K6HXxNz1gon5gVpRLZI89ITLFzWx/sw/CKpJPoY5DGzNwETOAl6kRt7us30T++SA
2ytzYaF9BoZfM4zku+8sPPvayNrIFyAICjckR3gOjXcN1Tbjlv7EeL1Czh1BwvAI1rv5bMTSY9Z+
wIwAXwbUyF98ps9X6tL3flFhp9lpgm+y0oh0WV1fXOP3kjIIz2APpm2gzs5Sa30myBhl2VpOQX4F
bd9Fh8+FHtMGCM530ok8WoxFGRulUxplilPcYEH7vh4MI6TZYqQhtgK2Rj5oC6TcgbeKGvBgi4Ni
zzvJ/4uWLd44psup1+Gfi1c+88SHQItBWcGdvXcSOvajRDsuSwm9DsHgUpl9L5fGxyy0ShXnVK8w
lyuluc6pDTkN2mjYfur5X27mLiDM4qjk7l9C91VaRHnH73xi5lf6J/p7uxdjxRmulzqvFr4jbTv1
RIKGAuWrOrLKeC4sG8zg0Rl83YSSMI9QIBQCCqxMg9XcrBbIfpISzTrBu3drvL9xK/8lsdypf3Pp
Fksxdio50T8KBRfPGIfK+1WvHYmVCvl/D3n7+Uxc6k+wHKqhNLDoDyD7iJGcKFEIoHRdNMeMfWuC
/GrK5SWWvdYjEXoQ7t3htMFai1g4RhC4oqKNF+/Xd3I5kMF4J7IizoLiHEFhI54ti+YdXmN56ZO+
/5B42nihIUntYbdqDXmVmNsxmBxeWZDEUsaJM0LQBamQIFEQ4eFq+VtOM7hsD31YPABUsQLdn8lO
kGA3bL/AmM1McnkvlR5oBcQrROTcBTfXRZcQqbQGh73CVWVPANoF7pv32dJi/XFU97Q6T/phMp6x
rWWzdurpTOoh126h3VzmDqDBOX0QhajMdha83NkkdiHB+A+gYghWGLc3ueYQVCbBd+AjNPi70CcR
6VcahaTCN/qNVmPeE+FZkiLqeP7802wGlfReZ7Lk9yIRawzOBol4vXpxmUlBHPFmS/NjQ+SRaYRL
QYaCNIsDxlIGaByyWh8UQW+otwAlcz8ffeKlJRE3UqBxxL16lUHjK9hatpRpkyxDxf2d63veiWjO
/TMoZFnedAsnswvDxpmRJ0ruUbYftn4ulxFcZMmqoAhNyJS38fP/qkT8dkktFM2wcr0DWBesa//x
zHHGTIiBZr5lAbFqTtIU7+oJtlMvu+BvWI185HEHG6epS1Z8+GWjV6jtQheuad3TQxpb2IDwrdqI
dQT8WbaOjPMQLFAVir0n5lgPKYqkMpeRMI3ld/vMY2M1LqZRTsDFBc2AugAlrTs3z+OMSfa7vQ6I
yZ86ub4wmnAuQRwrrFiAbfDtWEjzK99mH7mIenEuTW5K/fFh8LmtACZ3F16kIvxpC8BLEO26sJfa
bBRXytNRXtIJHwbAQRVqUmiZpQm7BVpwYBanOas9MyyKqUu1jHGJkwLVjnNTUN+gvnlIAVQIUjQP
YJ2mgHRnFYR3HrnpOzTjqJF1BtyQTZXmCBcD9mVlanZbXRiBB9z824SGjQ9OukLG3dU2081qzsin
TMRLBDVocHVOsEz6L3hDtbVzUAKIMznx/8lZo/f5dL3ZQocxzHarIQD9OKINRlV3WYrKxZm+N3kx
FQiulHdMbOY3es7BecaiJ15BTjzDwuvk5g/8u7k8R56OEUX0ttG273eqjoAMODs9Ghp4/OZUwsQ8
odhFJFrngsZ/xFgm3ftqQbq1Bmt5H26bfuk2dSu+ryD8eeY+3V5eRHKnaRCZvSkmxcHuEj8y+bVV
dxBmp6VCqFgcLk5C3uloz/f8teck3hEyteS5LGABm1+B+fHyU1Znq72kT7mAGE89Xh2T00QZRwAw
axNE+GSdg4WtfBG56RT1ef7GbcTGXkC2FBFKzRuxbyNgZJZg5/ZgsNJtTHXZTVBOg6W7YFb+fhEG
if04UOXtoP3TyFIV0kuQ/WEX0TyvDCubTbXRk5FDIt3/VvmJodRp/6ZcRxFpIaQRiGREuPzJvvwJ
Y1VviBS9Mf/Za/TtJAdklPKYqH/Pbf2EUAP7Lvaju9X/2J1mNj/rL+wrdPwllbrxd4FqrVwgaSdR
Aj4V56sTclKqUePN6cIvd9GLiZ5laAhpI9Sw3qaH5tIY7+02ChTwb+mGRTxVXaofpe+GJd1xqk4X
2KPgVjW1hiGK77O+rk06JU7HPBaF0XcwqFoAi10F0233dUcrD95jWYDdyJidB0O+4O6D0nM3uZ1Z
PzOQyccmuzLJHhiUuyB7cc8lJ4Z3iyT9DIoB7+oQm0PyP1j7HMg0mzQx9ypjfPwoQ7CzlEuAPVRk
yvYQUz6tWIsWrKTvCSZSCHjBCh1vsXJcSiVvfyNMyyKgfeMN5BBmbvoz4QdFxtkWDgHJtmEagpjL
X/E7FuZSkph5dtUBgw78+8QS+97JCHeFkpZIPzi1m43ehRD1rNVTU3lxEE6ER0oI2ubwUe17kUfW
A92FKFvXHmLouwSmOGogY+YHZ/J91/IHs9xTKfkhaIyJF2fqR9WAe7YYXp2U8YbwOIhlllaDCahI
YWN9S8ASYJgAukxdKd4qVFtSIEBewREAEmcMm0FDnooaGr4sKUv0aNK6yMoXDELi1DvgTvKfUGyb
dZ+zWhhwoG6OC+k84F3plFwpUsRCermT8dAo4mm2H7BS5oAk4F11HNUKByayu7S3ESdH8NVEoGLH
9aSX5JWlOSGaVg6rRA5TXiVrxqvLmos4PaaNH5e1LvOSpNT5UC2g7RB9W+GtKgHKmSreq731WNR/
b07GMLIWu22gVPtgA4RQeQdj6s7V1Mf1zmnleChyIH8FUmHOge8BeuTqzRh0gfzm3ziYbALEXCo3
c6Pjiz88cgrAq3NDn9oXI5q/vpfLNVJ+Kh0G+6Aawr5Ew/IdDe2fKpphl5NSS01SYumPJ1CTinaR
4K+H5ubFc6KITXvyTTntJUyX92144kTh+LDGeGEcS+3wGjk3jsOxRPD/pxOUQ80NUc5qrXKGByNJ
zlmBnSREkvmUnicCBI/0M1Az52wA38U+uB4sJIqpYG/bN0ki6aunsWOOnsGwCpdkUpok5EzVyaLo
r/xW+dmod/1YW24zY2kQuI/NJjAEMSSHHS6tmWT0FzEUs8ttzrMPMVixcf+jqAhL6NTEh3QrP+qB
2K27QkgtWs4Cqsps5l6GcPPFDQbuD9whhhrk323HxMohEeZ/unXnQLF2NZtQE9UDr4K1Mhyr8rRQ
2kPK/oltUXeBhT2OSGxlclXmosJLktOTVrBjvhIjeYndXkRNzIa7a/F+RBYGnlP1eUOpFJQtAdd4
on+uSvfBMN3bP2xa9PziQXlrxeuzh8HrNOXCQR8xlB966N+D9M8Rm5Jt2/yiJngqnj9KLp8viERa
jiH2FCgNvg1xlJZjv65KQcT5iUenOZyOagxXVngXtPCHFLJ9KEgjsU7wQNaV29yqXf48y/3hggaY
fuc36FaX75Xem/l+kkvMzZLbnekWcf360dW2qDsa59KWUeH9QkMVzTm/VG5FwUfRBvQTR4ShYXd3
Q55bzKz2oaROMZD37kMtKor0hX2rMm8wV7vgY7ijK8FKFfCeKw+CZX4ZJNn7imkgx0/vRApq15RJ
CK/V7waYMSdKa6KmxqWfGHicomvaEp5vZSlqBPIWNTggi6kQt1hwJERIzNV2BXpJcMTGZpH7Zuut
Fao1shC9EHogtK/RKF8CcER3jfU+wkt1sHBWg5lelh3n27iuoXUF4eWqT677tzRI/ZpdextvlvBf
iRa9B246pG3XVqlvhUlO2v4TUOPaUxKqznDnJqypx3ZCFpMgYdwYybAbiv1Rd4woOxyMIJJKBdSL
xYT5s9aB/BGsfFvhgitJj0uos26VkzHAy/S4wlscKqsNR257lULReObxvZh6ang+daSiS7CFJDtX
fRtT8slhKFeqJ5u2QjJhwKxrFyXljsUVhYm7Mjk23q06oKmXiyTmu+2bMI6UdVKgo8XxMuyemPfO
Z4vgtk6xjTMyft70yJ87CH8QwCOe4q1TJvGCzud/A74u7j7mY6AcH5cGbBvraYXgc1P0/y95JE21
U9yqNUy1xVyStnhOFjsCH7bw+HJEnPupmhdLhRliTpKFEqGkm/Yuiewa+zmAhVvUrxq5C3QTcbcx
AdoC38y6NNl2aqm+ShH37s8/2Vza8d3dDRrYZNBc5oHg8BHZtmBH2T7cV/U4VETbsvS+dBCB/tiI
T4L7LNGVNiebPCB5/MRYAo460Dhz8dhdLNbHPFYXsRlRNlqaTZspq8j0/XGqJoYtqWTn1uh2kMZD
/ky7uLF9+71Z95ZgTSAWn//sd0v6f4DKfubrz5HLIhHPGn7rRFcVOi+GEWswroZ7/AaRD78IfYzK
tr7Ncs09KarFL0Nbzs9f/8XMfttpRNryvjbuqbWd/uKj3BBQhQAtE05YeHYAQvxyiCMUVPOpc6M7
irNSZzrvgbQ4hZFeHcB86WuqNwwUD1wuHBgBjCq/YHkFhjfG9YozpCQyT92OD+txBh3VwO9Ia2bv
oEfoS9Vb16yOm9ElVBpUy3Ngzoh8KtoC5njqxwm/MshBUtCnurxgeQo0+nvWSHs/7VuEDwwJ+vtB
WQEN+IR8eKNH1j2stVomSbzdtGlQ0WxpnAAoSEVL2D/dFd/lFnYjyjCBs7C2+QRqTZ3/nUf7pLds
ESIyntrOkDbq3GYoJwfC74cftWtOYQ2JAZJG8KMNOSh6Epn0FNscwhlz4m299Pb5XM9Ir0ilfICS
MNuY0CtkdsdYJR3seI+km35GrtIjQRu+JFcbK9AkI73qnRbggqFUMgQqcITpwEivKYlETE/uyBtQ
un/YYeOrffIfZtVfOgL1fizhPtFJPBsjcCNdiChVghes8QSFrtQZiXbHm4GU2pzVli9NqUP0iYCG
g39wVnWR6vK0la6mfGwZ4BNdHxqPtPJ+D1a+nWptimMMUxbBAdIkgcC2zSuzxJRH/0SuOFIYD+xg
0rXiCBkEsayvprNElJwfehe38gEgmGG+uLl49m90ZTl20yAb9Bq48YNgvAhZUWndXfquVI4uV9yR
y24+ofy9NY62VAeJZUefk4g/UrQZChESdntVdLcM25GeEKH908QbLC16ccBjOgH0vE50HJ6v7t0K
oYC//hJFpP9F4kUM3g92VTQtc0lY4i4j2qlysay88duIJ3BjadvF0PyUTSZQsUHILJs7czrBdLLr
6qT2qcmhTfldH7EKfdpaHgFupyxYQPrXjti0BRo0UBAbANpkCdWRVZkDQTikmKZ8Ue80D1Ov7YZT
ltE0pW4kKThklGM+Zii8O3rgMiZ4NMCGdS9o+vd3HG68X5gDu0BF6RqC0UgleKGJtBXD5ldRsh0+
NqWnHIkwybsOC2OfU0cgoLK4vp7NGQeJQycnM0ss5ffwqR3GZwT/v/qRbKvf0NGea2+tbFslCats
viY+srJCz5EUMBKVcXczEWYtreQ2x5ZkjAqGTA+/tICJr2vjojWHJllLixYA6Xj97xvc6ZZk15g0
3iE9/JelFV7rPsvDUoxtYx+u7fIX8DeWwmYRAHI8BwcaQMASf30zDQxJkYUxuytD+yMDvMEd+l8v
geni9vdhhMAcXdu4FXRxLlw5ijiLG7VDQvK16Ke2Am+B2JXL9mzyrP4NbT6k9euxGZcEx1DMvJeP
tvZPfjvnGJqpIOTPwqt7+xi4cH0+z4a8gRSjSgrfI7K+p32ZcROqmCbZoGwn4LutgXDnbMx7yETD
iQocabFx0wKbk8q0YB1uSNrf8rTY7cIPxtEhpXu4wdO+/JOaGu1cqHELsI5E+zuR2Zo4SaH3eHzn
YRezsa0vDfBXLOFGIMcJoCTX8Dxka6nJ0EHPUW4l348ZzKywPF+ZBQJnlX9OEn+pIN4vi24tj4MF
ie8F8pQbMH5FO16pzIjDmydd8yyOFuXfpNJ2IEhvHtS/viEpMSwu7wXLn6gpoYOqmYq2Cif2JpYH
wBnU3kKJnKKSKGQxoI0bVNfQ0j8Qai/aQQ5cSdpaj5e7EUQvTSAVOYfOUUaNSiRIxu5MS8M3GCE5
pEhnOUhiJ2WbmAoQUsRGklQlNb/0JND+BlTK/6YKhTxSkMQzYsazzLiSYnPoz4muwETnub9UYN37
TTMBKkrGCezKsIBsAoRSRWjiJsYxJzJTZ6b9UmIv/OjvcYnhVzPK9jXSTtYWdipLYR/Tn78ZL599
n9/Y5YQuY6esZVAXh8Ht3gyZ8ikebl9smBSe62tU1wIoqk3CndLXT9E9flhTsRcymY8f/XFOkZWY
k6IYABNorPoHXQX7nEcReFsi7fritQUpu3gljbwnWcCoKyMbCWwxeFErRdNziDbUHY91RswThNRD
crmW2o2ioh1vpoq2PrF641N39NztaDGdvqLDSY7YIDUR0LSl0WCswGi5GOu6bc6LnaVVNKVKVG9I
CWimM6asFpQiwCX+JlYvHtLSVZx6mIwhPlc9+fLb3FuL9W1dEG4XJh0uxKJQsqIAz8/gDHcajkPF
rMd/2TjnSO2NIWPGGy0QYOKXBrKxm5OY/MR/s13DtPKJ4hNfsp9Sr13DW2NLpjVCwISOArDFgIl/
4r7nEaCbsAZ7VCjXLikdzGqkz4GbljLGatEh00sP9MNR9C88LdV2nGW+hWA/94PItlBuc6Y/TNro
Y4yrUdkJopk+q7WEbpALvGOvN2Vd10y9qCFj2t/0GUMXfShgQChcgcODovuge/jE+xjRT+4TN8rV
ar48FgQf9aRM0Tk6B+6N/gnpxAxkELVoWxczwlKVV1JQIHJa31pxLd/y2HYfaatzkRNc0HVeTMMf
RIMfen90NInPP50BviXlG+XRBt3iU59jw6kpuijwyo/58mjm+/W1fgMDo5kHXpwOUx37iysxzBhr
Wvw+oifb/KRI14zsgwnuDoVpSGj4YnFApAyHmgsXEDi3IAvUp5aECCJk8H+1dfEI4ExfAJwEkEtz
SNEvLDqPXv2yppGbEQC7N9HCy3VKbky0onAYeEelv1qJqvRuM5zP+jkRQ91ka6tc+tvIZvG9voD1
PuZ3Ud0Z95r1x86lpWAZ5ia6naDBWDxSzdOrg/xFYVOyPP8QJf1pehtMnUL+635Z6f16o2VYS3Vl
M4Fv4DlQMrWEM6R1AwMJO7irMaUIaxJsRKw3CQ+0PHVwgRiqqDIdefeh4QBC84xv6S2K3HciLeCp
bdpi7RmNboSHXL3kVWz//1vsJLT1jbx36kvWc9NwIc9DBqE7w5UiLOtBoDrnyDLjd7EMRI/KwoU0
8zhMx9VRxGdXM76RFAIrVFypHyaULAAmqw7TTILMM/Q5nzch/dKhj5wwkueoMiOfojRoTJ3PpTpy
JivE+x5FSddBL5Av+0teVN6J4/IdPkDRO7H9H5LdJojFvKkxdwqe2G4VgfFXb31x8Jny+pbOxYJq
5+SDJobry2IlB+hOYoTQIw6PHcfc+zKOOr/JVfhoU00puhv7PQw6bNaWBQsvxp0NzOrEpPiy4gOy
14ucF5tYN4J52zMfWBYOimda6g47Gx0jzQbK2efXeIEiBkEeirTXX6I25PlnIkHZatYYTxLm5hlW
nsOm8O9+9kNBPHrhKM+e4p6JfjaH2EC+qRbq8oxTOumxK9IF3GDvTvz9Ulhr33LLOKdVn4kPvLpx
aKTTuxtPdpzLqyXpFzZ0VktVtOzBpwwSXX3lr/mtr4Q+axeYUn7b3DHBfeBhGGLdJo45LhTpGwwx
Kt4hK6q5LVw5cDPhdM//QV4LeTchUm6/VmO/BeTqMbSOuccUlxEaREIgR19HK9nAcv5nlC8zDdfl
1KSYg7baxG21VddiBYh0rfwWDLke322KmNGqCcQZkmwU/fq1gQwV4eixyL96/6K5bp2wcaiYUap0
RquDBpS3zcUOpLYgYVNkENn9pDT9m1PFWjVpqjxAaoCArSllj+L5WyEuiqK6v15SXKmwFGbIkmqr
FjLBhFAYM3YTzwp5cjuMQHD+Pp8jKp03lm14077spAYjRV4BoVMOZH0gO201tV9Mha8/dPesusHT
oU76C/6m2SJ6a8kajf99CJihm47CDWscNYTScOa9+qUvln9l6Jz7InbVxhLvAwOj423gtkQ2SX2R
Ac8BmWgHhGR91eYq4OjmdvwG8iSuIeG6b/6baSj0UxipPXP8cXNdGV9vFYB52APjc4M2bZ2o5Z6X
89/YwY6GGh9xlJw1CatmypMkj0Wn450uulJ0u+6QCMqGyKoUIlvuB6+NJeON9iarUqcdb/+1NzS0
3+7H/bhlp4IfRJLuODE5lvbA/B9HFzh26NOoI3iGp6UenF1gW5G93pU6TzJ2E6iFaabhnXJ8epDJ
f9vLioPl9rmIo+uS9luXmrDwvI/CL3Uk814yFdJ7tRAhvR/5LQKivYtxltdnsprkhRhBFrNAvJQj
Dd4mRbEwkiYLzjpQ+a7HbKgMKEg3BrfiXpPDRPw2gjVWpqr62fnOLFPVmjrgiNRuv2ZAjZipEbzh
ftZ4tTGx4f1/UsY/VP8sdAti9R2YXX7+HvZGVf3j546SJ6aqB35/SfbVj57EJ+yKFXrJNHoiBTZV
Fg+xFf7NcKM6V4M7aG8mcUkx7j0Pv6G6E+yWJiXli7rmXraymGl5hFoQtikmW6CvgqkCDLpqdIrC
qXVvhr9wDNk4kD+9nq9t/gaUxsTQ0JZVgoutwUnGzld7IaZ2cRX8/Jg0LhtAmWaxHcrZUp1UFrZq
Gjiek99gktTBCGRm+Z4zQdMfT4mJFtbr2RpCb/k3j73WIg67qjfByb/XKwABRKPDcGDTAN75/sxC
7IjkItimGpCx9M7cw+ZcpRQD2/NBOWLe3HmubUsFaBGqbPog46KoavJcGERieP419ySKjBsTp1/W
leonPPwWa/I3kpYyBtUDx6QjQhZ3lc21otTilTTaZxI+YIroR52rZ8xZsYyAhll/CG2nXUw6WHiT
TlcS4b4SBIUJb1GLdKaPvUBgPrWylT3PX3srIpWwA8EhVUfui4NuvTTfws/SR2JZ4YBCP3xa1Dzd
Ol+R8FXiI0aL09AZzQk2PAbisuFmv59LHr/5gofIuN5A4r+KEd506auvCvVTjBwYKBM6IbhBaNO8
KmJZHNB2pParQMVVCrA+0AdYlTF6yOMuaAfm7uCDH52ErBjHlBlVJvIdIZJER42rZUpLv9JgPx9u
Qc4LHqjktwcpw9byI5a23LgANwg/O3utJfmDzaY8aIYgyxE17K04j1Uwe7bQxq3Io09EmbhXO593
RQ2u8eHOIozUOfzeyx6RtqGFTmamAfmV+JQaJADV+mBspR5sV4kG4USkNaWqzyoaGn+9ddn8Usvl
RDyfiru0xI9DRgvMaZ31AyoVhF1KUsD+5Vqf1MS0g5Q3Qg4Uk+A+COCvnrZooGMqLxo5WdLynhUA
/rNt95HEzivukhbnqOmxJTFdRjj2NB9eCjepuB5PSZC/Bhzoq5BcFW0BL1thtvr1FJ2At77BR0vm
kyDwNNM4Qp0+q2J9RCUorDE4Q9RBYaSanpWvq8zuHCF/8m5aPUFyD31E0LyCLh+B9FT9WGIaWyv4
SJ3CqKB6PvxBiRC3eBEDnY/EKDAh6GW+gXILXCiuP3eeEVBSu6v5WZDAdMvnSg+1IpxWnSKrID47
4yFTCknWO/qrMmOnkN4Mc1DxNnV0V98fdb46NRu0DWqkAuBMKP3JowhjvX7/D598cc0ZuTuTy3yS
i4hrZ63bq8RxfwNjHTw2iAGFhyF6zhxDcOLxxCEuCgo3yBrIghAkBJS4hrdOgQPbZ23Yzf43QXtY
1LP34KKjt4ZGPRpK/Whbw0eiMgGlhAI4JTqgCGGVc5G0qOMOLW10EL16zePLhPF5IhrCpvn6qORt
sL+ctov9Ayl1cvcbHChDV8vnfrfvS4dsaJXeqAE0yxvugPVJVGoJ0qaXkylODD32vvL4QVsUrcbL
kd5m+sqvO145UUITENkijPwfDDCkBuX3bxcs5xvt74l2cAkPw40H7XW2Ks1bZL2yp2EDu8yD1+0O
18kj19EBhqreQ19y3DIWYGcl3j76DeoJrWXsMIGyVidnmwa/d+iMj8aBxAm3gdE+V1CT39/vJOKo
RVNzzVdkBh+CcIv+QlT6XMxAsXK93wWeern3py/t2xxrHTMy8GioKHouK5jacXCBAclS5SgAjTkd
iha7rjqZOKEwficmea3JojA4bloHifTKCuBoa0YwsKLB1zHL3nOQ1kbNZuK/hOmPJNYcusY8WLE6
UfeULqj0K8GiUvfjQDloihbbJlFe/eBo+c7UWqgs2dJYYLVJvEiKR+oLCQijqR5HDGkFtmyfH5z7
fNafyQFmM2u7lF0ixOKI8HWl64wfJoUn3QKRouuYBmm8eA+n/hNNYuKrdPcJxMNrGWnslX6DS9a+
243ELS5XNc9cTX7oXREMjnhku/2Rgk+KDOPxUWCp8Fl4d6KVhU3jatMcC2ziviLryH+rG3yk6Z3k
wmlHeoWM8E+EzIEeUg4ER5YxwtI/2Urs/Y9QaGfjKoH1ynTKYspLuITkdiOYgRQeAvf7ruGSrg63
W6UxTDsztUxn2B9PV05A/vIjpKqNtDAjiE5YzU+IKS6RaLDJWB1kVkYUFUlYvkfASYIh+nykmBg4
axQHM8yKjqL/1/zNTvY+uhSUw+5+PkUbcrHzNtFk5ewJaL5Sn9aAMxdZZZCAmIcyVv4zL+bWhqNI
RX02qAepMHL4/WL6ndADltKW9FadCv7FwjbyOqUgjKlk3eKzhH1Y/Vj63v/OtXmOuKmZN+WjXwn+
p0lKdjDVhgvcGgMnogD6PAVeaRTwIfwdDUh69MJA7vonjdLMGsSHAJbT/DL2ioZUSuPBvJkWROhF
gEfMS2uWfGu0dgc5+qyboMpBwCMV62zRGtPKsk2hjUFPHPX07+cY8Z9xVUOf5G0MdgN+Ei3R3YDB
1GkqC8XqP1hq1nB3K57WzWWqTLvbV3UcFchLC4V07AAZDxWnQUnlWmiib/KsyD1wlW5GbjpoPzij
t0jKmmVYOmCI1Ri2yP0xpNmnvY0d2Sf1AfihXji+/BufRthyPaDEbyHVQlPmgpzFOu2PMRcmZFG4
ecROcS5tqfiFppuFScx3eW88sxmnyZS+hGBA3se6o84XxCPXjFMMZOaJ5HYh+NhJOBjpgMe3VhWA
OrxOHmMg2QLkSmaBSKMstXBP2QhR9LmgIsi9ElNCfatk4d3PlvA8asXsObEPt+NVFE97vnaH76gi
i9W2QOFson6zvcCdu+E8xAoLZGWD8bdF4Nj9US0MT44ABHZwgrRSILcYZWbDNeiEyVr5VbpBzZye
07NcXcC5jlMyjEXJYqL6BP/xRnrElzw+jK3albWSoZS8ftPfJDEY5VIBWKFbAJW0T5zcFvraXLQk
aKpI9UUHsAPgorRFYq9vczxlqVmbcUOFdspsonA3gArAcweqAl2UtXbjPxPsYVCuWOxqXn90tpd0
RIUoN0pjygFBpzIkve4X//aR+IUjJgSoGvJHPcENApIxp11KiSkGqTRZx/rGGo2C0mqbJ5ALl6aI
u7JV7wcueGvrxg6gNWJBZqnd9bcgT7yWL/0VrE84ppL+4TMm4NTc2DEb+V203Cv0WNIcsJ+qfMo9
8xto0tq1bWaX54Oa+ZhzunR6foeaMrKQ5t+paWTODbm2Eo7Thj+Clzf9cOmG5Wb1f+1V1iAt27nj
OXf3ylvASxiCRCaN4wYNzE5zvDToQmwOD8xr/JleHkIotUy+f/ziexxSAtVLvcQxG3rYwzRMbTCg
ArDs3LniP9tx9FuloUAKUh5nE6XdUwHLcaoHumgO+Xwt7+HKKkpXz+aJA+Hrt9XitbhP3z1kKmqf
hPgj7Kh9kJ3JzBkPcM7LOuKBYNaBSCon8UzxAMnKoWeQB6cZfKsTddbRMIYNnvYMby6/XHFbKH5y
d1vK8WFIoCD9/x9RhwdHVK8NJFGcLHoZeVfS7dCQANPTv9lBeDuUHxSKjfwp4ABuBqBS2Q4XmRru
LpZSuQY3xABGKB+Yv0E1wG1n2t9t1rndKGL0UiQ12jaKU/WEvXrah9AJpaUyWgrn9iA0GDdsjVtA
F2JhcatOyKCTctiCNjdie8z+c11DI70tUkZ+NhkvgW2npONT7FEmz6VqTPTpo6jADfqkqgBBay/Q
RDUJG992uG3aA5hZHhEo7SZVDm6RQo1l+V+ptTtUm7twtv2XlmGGKR9AcAhf5v8JqZYaSLE74Nrg
Hhy3Q7pFrR2oH32NyYGTdGZYbBqAhPS25wLotdRDYsxxnl6y7+S9ZJ/4BfL60jukH3JIWQ2DqPwN
/Wgl4WU5cEzxE3dmAOZ3kaQvuDIqSDZyFNjHPjkyzstQKNv5x5m9WdaTVjspBfTdLqy0912B3kVF
/FSxyY4B92HPw8ZeVBdwkXxmviiVM7OQIYiYgtEFEipGlChy9HI5g4XzdvjQK+nbw1Z2qagE0fA3
AT2gsg9UKnJxKz4fDk1IRW0uc7kWup4UjjR4nsidBBozYasF49gOcM9yCjuQPRq+uRi9fZqcCavW
UA8mxUDiveD9jx9SgTrA+NFtnVepWNPynhWUdwpEBVbe8+3rm90QRVxezuQ+gsyp2FaM/42Et4FH
pS0D8w+OhfDQ3qPmj93odB4nAacvgtXGvWPcmWgN8c0sljKWeyJFlOKO9M4hw3+5J36FaRqCbLeI
R6qDdbo/U6ioWskwBOgBPvF/tqVp6dcKqP4dfVxyF3XHr+YLCrG2Rq82fvLDzSrdmKoGICY7Omu2
aaJbDOZbc8lkWHdT440Igl8YQpVitc0UE5hzgyTRoOOx+CE/9VvjVwui4lhATLDDh78CfumV2z2S
aOei79gPj2ihryAVCfqOkQCz/p5MY3GwJuhHhjiGeM/bCc0IaD+aWQseoDoZvHCv5jUQ/cymnQQJ
jfXTysxZxxw/s+ckPl6LmqB3Fd53rOQs3rZQAPWlKI3FzNUdx5tQBLZX6x8CrFsEl3buysSmOshD
i7c9D+E/x9xI6Bs8lajbLIhphC4n0RNifz8Lm9OoiA3lE5J/OL+Xs+dPiV3Ag9OEMqc3kG3d6kls
nfBOO6nKY7SxOLzKF6HuS+Run7vJnsCpYVlZWL6SFym+ztZcTwMMKz7qwi/SRNz6BVwbq65+n0RR
9bD2K2iowNElSWw57DeY0ykJ+gUkJgvEEz+hB2AkHqQhc2JHfRglXyBkhGDUJdx7+d3PKjiNWcex
saJyqIVx18RdD4bBhLBhd/CqWNMvLm7dPP8pSCFc2Z0WLtTrLz+kLz/2h3xkPZytpwMf6d5AD4Zu
VH+vImykAFpo+Brcau+sS+bt9GKnyAjxl6yc7A192rUB+8fPZ+3SyjiOP2UIK+PMnn0W/jADg4Et
CybGm8Cmn6mws/L2mRE1SNX0p5lONA/5THO8a9DTGQu9TWXpwDbHq+S0qwGsDqUrytEYQ5aZpDjc
orOUiqf+WTXPCbtjT+L3puevjOfDmWvNdxjfsZAerD9XC2SBPae2NX8jMYldXuGNYa7U7BRY8AzN
huv+v1MabW/FV9KzUjzdUKKg5u5RZHum+5JQ7GWcjXSyF+m7hdt0VN+nMrlJd/JlRbRgch7tMLgd
J1334z7R+GWW8RKoeUp1idUCCnqABCAnmXhknwuMVyBGGFxUz6CMia4w2Gxh1jCLIBw//7VyZup6
Zb/ubNHXSdCJgrzKBJbeZnrS0u8vhIIa4d8RgVV86gnkJ9qB12Bhw4MUWLsfsuxBOEePFbFR31Oh
7ORVI+rDwPDuPiDaDi5Tzc/Xc+LLPZvaxpfHUYZMoEPl4g9JM6TFOLRkTWFonm5XI3XJpoJi0AsN
SYQcObjK86eBsoLZ2BdsXtIK45vfjrdkIBS1lSyCVKiOBWgVzptvgockFP1yAT0YvTQeVwtxKgmG
d4tJ2pClQBGrxS/JdKFSeDPq0kxkFI7wdNouaSH/kE/tfl8C5UuwxBJ8jMcZCEe6LeoyNE65FPDM
bBOINyP6FWlPgpyYpMHGzAfl0v2bdS9SqElL9vgG+cErJIWKZbWN08Al1vVoQnBem1yL5JjdZ29J
YxL+e0BUHHLl9hofCmkCexPogmvrlIri9wfVc7N94HMa5ZbcjWQ4NXobtZSKqjf4tenBx9+4sILY
M5SA19P0nzs/JQeXlowA6WTJebkL1EgWz4GNIAXGifdg5cZqJFf3PEX44EVcEU8pl7HvfoBTBeAw
/WqFe3JowubHIhjYZunJJ7l2vPj0RlZ7A6rGdvPuHEHPyd1cgvjUaprjdCByKJuC5yaKSbMeXeGJ
Lbx6k6CgSX+RpRFwpMLaSMiQl392iS9iLNDgURqNgHwoR+RWNdEQVne2aNWWK/BBItRQvZbgOw39
NpBRRUBihJZd2Z/1QVTETtaBWK967375v2JrQc+/9ax+VSNvKXZThMk9mkDER6mYvrBZB/yOtzuI
W9fWWHXQVIcxCSMmhv19bjxjUe0Ll/szwJN/m80zDpzN04bxez1wAOJEF/3b8zm3z0Y1y8udimgm
Hor8XJuewLV2S4zkqZ5WHKx8DnMJtIZ5wi8rgHPKU11jIUNI3Cv2gqq0Mj9PMG4PoEqrHoyB6T5e
tAc10FwK6Oe70sy0Vq15/KtA3MzlYbGajJZQBna4Us+4skzY7NFUm4qr/2/xnru6uoI0jxZpexQC
HGWjVG1RmFWthezSWcZEL3XfK1ZE0DmJpzW7TMIXHoUP8+3bm0Hmsl06F/M5WT6HY2mGB4JPEGaN
c5wjO076iz0rKdejLWxeYJLYpbgefxt2s9rArkLwjasPDzrxfOxETiq1hihHX1FxnEZAkxvk2Hcr
1/nz3IWiEkoGUweUa7i9DrwwtpPNzveoRc9tSbabbiF/Z3PILQ+dr0Eqs0SiZegIdqXw1/kaav6Z
elunDrxkBCjyTS0LxZUc0X6SwMKzwJftWgMTg7YRmwo7SpSzjIN9bQszl0HcdBIl9TDTJfkAxd8L
UCLs4RU2hno2L9BruD+q9F+/hwrtJ1H792oqKQHd4JZ9QU/qSZpVH3P9dJX1iyXOqweHmkYlSHCR
koFAl20hpgTGrooV1q9VAqz2WiuanKJXXpeWrSbPsCIIb2LWZsxf9QZIsYesv/AzPMxHhv14WXh7
td/0AgUeeMP3FttVIUfJC+aSSbtAu+CGbLntwBXMQ/yXLRaRayH8HDl1wU1kdt/3fbNmOHhk2Ih7
HwYNLKGksfeoZp/QuCSuR4kRdpQmkEPcMojjER3hchhGVHRuuOIZruygLRFkLhrrUGF6yIh9G4KN
T3HUUla3oCKDc9AcnrmHUATwfki5vnerytNiFFgdt1hcT2gvXi/OjZfANjMpxOsIQMIGF/0UiGQ/
6up/3XW1Cs5sEHHpHEiFK5BVV1NZtVHx+T0xK4thl+n8CxBZDvKXEdtIxiBAuy1yb8jFJEpVhvx4
cfTreDMtBPmHrDN69BUvBUzdoam6NJfMELcP1lM+Td5BTWwzxHSenAmoaq3p3w6zxKHD0B6imMMQ
8F4gCuYBmUcbI9jP6JFU5w6/wjfQhBuqFIRAKtbH1G/8dPfVJNqT1cyBkqdMItwESiSj8iQBfmOu
Q6M9uWLznGhjXXLEfPj0zvysnibEGLpUcfSABvGqFr0MGwg+SElavB05nJtJ0GdU2oTh+P54mkEx
DVu4x74DR/X7ChmVi9ekeX2p4HltFtotVD5QqMwF33f0L/iKQLpFuOmu81gE0m+PGPsVbPgNAn20
mCRG+h+iolvEVtoovJaEloUTH6Vghnz8VYhA4AHRYXP9NxVneIueq3G+u5NdqquXKxcR31VpW/Me
M7pz4VzZzeRzMBcXUBdH1XFsJ+6qNz1xfODS9I3SoFPRqaVISQz7ttaPbQXEbTQKR9CNbxyUeLYs
5DiCo+PfOBLSRM5o9w3eIRxCexqfl6ok0Z+KMnRPb6dSbmBjWLLk6ajC7Tssk850dvHBbOdQK7Jr
HJKW6C0A7/Tn4NTMh6bSO+wuV5/uGaJCAnUquZ5o4g7l4khEbj5bER/7zvvf6HqaNDj87JVbC0P0
wRlUtatLntknxiBUCxrJ1NqmBdGrxakolSXFV6iWJE8UeoHot/7r0STg8JWoheTB5xzPB9MHLPam
xSGQNlVRoSm8auUSbCO2hooEtMwog5CudPQV0xzkNWa8p3L0Lg/KFO13yl8bQ8/uhlFmQeSzQAb/
njenxceq6inJy4iz5GbLY7HAbXbpsR07DpzYXtfSq25izYN7v9I2n78nGmi5pUDPB8OzZAGip9XA
KxzT1AAwmRqjjPzLz9bp1mel5wf/ypJHwiv8Gms2JdIddXZds4SuoDO1fg2VeZVWD4sImMsoGDJ0
9YNdMuCk4qKmu+PB1mCRLfCX3vkw6UU/pml68SFrD0lQr/0z8KVvL1PCCjJSuRUKVVLP4Zploo66
UjMbCdvzdqIOPPGpY9EGXM6BHYfAqOxRIYeFcpMlPFlmuMmYK21zt494PKAtI+6oB9WI9wk6lTT9
ILKcb4oG/0bE8pRwXz2JRgjxiTlixnjZcmbkgzY1c9PV1NtLEQyfkmaiVGWEUeXC0fCat+cPRnbT
c2mkgkIjlizLMFoRA6NW1Tpf/70AgYyjJVU2mowEP4JnjMu4Up912S6QRWBRoaZ6MoLDd1ERro85
p9Jyl0g3QdQFBzCYFt2rvQ6bbV/nOORbHhnKGpqUSbiH6gs57L8nhdw4xUHjxesenrCDbuqcdG52
HW0YXTLk9EzKFAyevOrSAGFCL4QKfUUJGEJ8RzoEMcb8j6378vAnNtMM6dnosHP42oWCLZN9jbyd
yKXSIp+ieoKwPM7NxGrXENaWdcbDpYpUQ/m4YExbkPP9N+L6dpevylZMPzQ8Wg8M8GA0Q+0QZul/
liu793MQjuZ8/Q06U5Clp9b0IV17LCNf2BqvF5uAnmjPahcsXQJjOoqRcbMEzvrYd0x9jZhAQ0BN
eqJHUNSbpJ2oRcV4yFGCks2drbel2swBZok575JXr91OqYZjNkU/9Gob5bLOcHgLsc6dCdHQoEr5
X0leWzXXaeTOchoFCmGAD73eK3ayxn0XMLMjv7W9WOVDyFn2BP7sYiHzcxvQikMCXq10ZhQ1p592
6H9/exYVWPGz1f8rXEE8YhywLtZDJYylh9GJIGSkks5rVsWiMbBqPP5buXuB9+yUEZunkUjTldSB
AUVxOo3v25IR89T2HqWRqo8Fd1Y7DTl07FCelFVj0pB7PfdY2gvNP06J9dSkf1YiqK/LhIU5YXo6
kej7CdRbOwrPgOxKmkwndYgzqgwV68j2ZSfT9d41CyfY/K8EFvnKOjcxNqrenpyonUsdQIOV8PMp
3bYD2k5Z1uiQhOH82Qy2U4rWsfCK+fsVJ6qOy2svc6GTdTqyldfGh9gUcxDGA4ujnfCDZiX+0zHg
winMzzeOqMpMvetfsKVIw7zsKzUaTCHz9jMgXVOvXvP2vtO0JDGJyO4q2ZFVBW5zCDGYZTjkS20o
rsfakDLF/rMS0XWrebhUg9pOhcehGh8YhQRYChqkrRXfzIpFzNGHsy3hQYpMoX8zB4BZWhsINpo8
xvIsMR0V1hsMTl6JaKNv8gUrIwqfvTGQrlUCsLwteaDyRaHYmE9WeSHE1MiIz0elQ7sGNYwoWGD/
b9KJaiUc6LEczbKUFEPonzQfFvBp+JtGmtu2SlzzYs/9OVL8oTAzfywbkBIRYZ20QxqGPyi/od4h
h8ZTv1sGiN+Tu3sWOKSNWb3umB/wqBT0s8yXUFIHnKF8DEZznW7Zk9EibGYop0Wec8roSTuQa5G/
8VllyokLGy9rVcdbaJfX8vQ6GrPRbV883s7ooVR6mJE2sqJiDiEIQTt+2tbBYRjHSeTB7iX1NMc+
Eok7yXZ1e2EWZHnS2Sl9C4q8vIuJV5qLJukNyr3/vwPyKNMD++mACkdOhB4MbqMquFM4F2ozf2AE
Y0X1YAMckhQFrgm/fHR2B4m7gpvOe/8wi7dxQE4Y+AqcW4AyAZbnkE2mEoySi6aULCGXbiIx3Opu
/bivn/cSlPnNV1lEbxvWh8i8AZRwvQe0o/n2jkNFVvNJG5dQ1PInB7+Khp6CGwEaf2TRZqbULC8E
6DL2eLG1uVIN/sX23cimr+v4cE7BIYQe2Csxm1KZ9yfyN1uq7t6OuRYEYrq9jOmnTxjIG03Hr04s
FaNGyrYKj9w6epG/5Je0062zHEkAG7cja2VZ2QsMoL0yBGXY3gvUZRsBuIwbxdwtcFLoPbBF07g7
Lp+oqgFbNqLnpgvL0XwB1Kxcv3QiFg5EAKpgKrzamFkf0JgrZuFUfhMyJqPwtaisQZP+aIJKc/dg
6b+h0jNifMKWtojelHaTW7E3dej/SB9F1q93uTqHOjCeCdZpP8vQRDNtT5oGRnJ46CAekrltXASW
ed+z5EHlkRmCajzCktpU2QKoLPUCsCs4UoN8ofXDrMtZH5ahUBdP1qyo4M7opz1JErG4bdZPLfpP
aooqJF07yKV6dSJPpru6M1kE6hTL0mFpLaPJmF+ynNxJuclD8SnM614Kcisg36UzemehLyBe7Hs7
xp1oXp1Dh8BQrUuh8DjuS4eif71espHupygnfNwN7f0jvH3DcMQiHx5HVBHsqieZ0yyBHaysFBwv
OaK3Zrcu7flW6S4TuHmXBW6yB2zDkOuTGqjEo8DO5hj7q1Bi13kHYlV69ILcr1KuIzuRB41qqa80
mwX8KuKkq8BjNFw/p2UTCnjiM5YW86ypXtJ86IomHXvvzamiMwGmIMvcaj/hbeNJUtyoQ8synKJJ
1V6SA0QDQrFrrXnySqqGvKwd0z6Wjt9ESCfVRz1O3BekDRu8f71A8k8AlsgG3vU3mhOxcnj1nIeR
+0XafjdV9dMGy1wALUYZj4IRJfGNHUS/teE8u7AMPH48O5WBaeT6AQRCfluiZDE6TPxydi//aePy
tUMTjhWn0mEujdbsfpyVVVZpm7qCPcuIr7D0x6lCXqahsG8rMeJ+yIDs9AH/fJGTNr6/iA2Locv9
kWxvRGYdCBJD0a7G397KDBkr/HSKmNaKYZD4n9B7p6HttCHXncqbEeVPpYwEkmRK/FDnohmEs1uL
/8rLU1EeQQN3MmzTs8POskgZrUlZDL9DQnIamHX56YpWj0lVBDoKjsiih3M+LLkuowZOi09mG4yr
q/2sidFb3dS9N8/XLnNfHyKdhmm0M/xPawpeRUxWMRiuikbYZLbLAqOll6th8lP2W79f+J3ObyXV
XJjyLG/5++nwOyuLQrvQfDrxc223n+uF7hirgh7He9vvGVkhVzsuGy73eM5vTy2i0sr+/8xPl/kX
IFC8qLyq42zlwGYyYlECqkxPfHzutwM1NCwL67ruTwpVF83rS/+bxRECmXKMBoIKdy0a+e357q7n
CUu6tVtIQcjzd4YGdiZmP1S9WiKZejbgXSKVdLS5FehRxwNA6YI+8g2ok91J+XSxg4nPgqj2k4lP
Mh0zxaWkQilK1Xj0qS/rcntZRU6sUEkzT7EQC24+L/hPmSDrIZBtD+aaOitMWF+E6v8KJf517uFC
AYhjwgxIXCzlS0BKsfO4VFgyu0XFImdl2lT2J53wSHQLAEoT2h9tLNOWgt29CdDsbPdvKw9AD22O
qpDU2QGH1JQCjNDv54ysK2LBazWCYc1RUe/nKTuJujUKaSlgFXEPke03xNXEAOGXKOUKnwBDSFfT
ZozfNAJ51I2mN7gtsHIzcBMSVrRauAwLKSHO7lNIj8clVniHX0jMh2ONMa1WhaBFF0Ptm/dZHPBf
gEDA2bOgi4kcig8MNUc24wIVXpgTvrCihCMzuUb/0I+4uL3N1Qs6rWVqFeeygjjk4N3YLrKUjoup
ltQ12KUIIKz46lEsLE1pBYS2hrOQ56uD6UPcitnuGOpbJzan76ufHW5kGaOVqcaRpiGxg3lTkP6o
I2mqEaIhwl6QdUq7Tg6t85BXOSLusiiT1pqgvvtRChgbMzwle5d8uCLXlO5Tt1bIYJr0wUifsKF0
o/9pncgURWD4mnmGd7Kvws2bRHRZzCJNptWg78nUAoZ53xIWRLxANa9LtIBTt6ep/UgZa8Wv/nZJ
JTUNnA8VxWfa8xmK8qhGChTawVa2XzWxuOD/pK/IfXcWZgXP9C9dLKo4blJkZ337rAg4ARwX4RhL
/ggoMYOEs9ykJYMOfrZ1N0rJ5UhLrAt0+BMFQ95dUuQmbDn+k2bCQU6nEBnCoinOa2ftEcP2FJQy
A55YCI3qSMClQiS/NfIOFG0ivuzGmh1RSNiHd3NccoQ8bWq+m3TS2FMWQSJZQhfswxVe19WqFvTa
45Tx5GK6U1q5wI3TrRbKikMdN0s/pxQYjh4kODsMfZl3lh/5WML3zbxgraE6lYQvjunPqH7VqIr6
r1l6kWlEFuvXfMMWrdsvrozkNhlxF7BZB+OusGXMXbm2D0kC+l7YL4Wq4tsBAbZV07H/d5g5DWLJ
mJNH6+3+TWtIbmJJviSTVa0xvxPKdnV64eNJddNHM6JAxyoOjRFIPxo0Ca9vIGRuEnNTBOWK+UNS
QOrhIoJ7tfU+JABw1AsKVM93lCZxc+A/LOjA2RFfqBmjFA4rFBVnWNUArE2KZif/jKtLhRy3tZKJ
wzCpn17U/E1mMWRrn6ZBBEjZ2V6utjJOfhc/R4l6gs/LFPYGmKX7V1AKReMDUTzpoagJPowWTzck
QnRoq1uC1fDv9Wayz5AJRvebfJu4U6qzo9yjlQT36Q7VTFjYOUx8CIsh3gQMbZA/folspolUlyV+
uQm1wkoFNk4ekUoAk43hA4GjBaHb9tdSznvna+Od/ZuDFUEnoGtXYFgIH2V4jbmDHSRv9hVvINGE
+IgaoslJmqC/kB5Mfmod0ae1RS4TUC5l2j38y8hTkmN1/akdXISZVy2yHU+Iq4VpKZTvuGWXWRf0
w2M0GsdnrDqANi0GViIEPsCAzsqKsP7W49z4zFu45QCBujRhQGRecqiV+W93Qc1Re/ZN8C3gGmN8
3CgTk+nZTBmQl+lD3/ZUTCjrTUUmpZOsfZdMHk2Mq8P1vhSpMlFppxCPxnVDSLcMx+L13IhEOvlx
6VzzX7ElnVKPthd4OMjkQTkyBCNpjnYQIiuES2TWpAAjuTcmuRjUMTTjkvYtwmjTX2uh/nPe7wIx
xHHLYZQFbrKgCphuyytoB2fs4uXJmOLO+CGeN3j8UuvpnFd102T6ZnB+66A8Lwym77de2/tLFnt6
Ayf8tUB7pX0S+dhITNb5mH7sqEEvUEmW04hBdjRC4arGn1DP43QP/Y4xiz6+LOVrYL4196Y5qczF
6m2JXiBcTUmWVy+5SRs/7FMI9M1MxKON6Mc2MTfnuoLwnKHCUqtP2MF+ta9j56QiW1zu3JumWW0w
8hx9ZPClQmIrBkyVGVDnMFqCu42KF1B8DG7f3LxSESXenNFEZ8LdxXgksBw2Cdf7x8uBh3x1i2dc
vF+cnqFGL/JwH17f/cwv7aSPk9MUVeblM1etvRBJ7CVZEzloGxbMaeILUbmKK5qc8C+eRdEyb87t
u2GdNEt/YIKSB/SgGebZqIfIRXnHL6eV8OK+VhNde4TxY4NNohaWxLfkZ1kMU1qHVvnMgCfuzgc6
qb5JOEXb7qmg+f2K+yKx5UbGiJKnUUBLMvEV2yhy7C6iy5+1ndweacYV/qnftBP37vo59l8Juxkj
unHTj9Qo6SmZv6P1V7aubeFcmPRdZ3t+C+zwIwgy0Xm5mfFZ+m2OusXcpS4dY3+goV+TU6EfmdHP
RdvUkKA5NyQnj+hyVegyfixFK5Ng3TJ0lgb+jXbywvfQPUwj5x/i0El97swcZ/7nJh6/UC8+EH9K
AaXQvVTj6ca3zgFZWpFB1YrgcHS6PFjN7SDrrILMxMkfiqnEh5R3mOqFRJFolkgArjNOtZfF66WR
gOscvLYK7IEvN9Tx07d41CDseaSMQYIBogfAHn67jf96tT17yQzcnbcupqw2hD7pF7qBS0fwQVrC
9vbE5wd2fLLR5+/w6HzjR+sNR6OPoH7Ic3+K0xqj7jalh+dKlFOdveF4kYIegKX04zb0PyqtzsxW
iMawEoummy6+tV3/zkBYWacJOZ+rr2Jk0UKftGalp7HZUDXlAx9zANBpBXRAYDFF3J861qpcF9G6
Ykc6xNb0v46n+dFHEwj8syZQfiMN3F69JodvWf4Sx1cbh/ZtQ9NwidIUjJd5TlP5S91mbDhDvzcF
OABYlFm3bkVdvvJK9GL7D6/rhPigTn0Qj1qLip7OjO6m9ioyVvhfTM0fWqu5jBToOO2BRiVGVrnn
qCI0gcyI5HLtJK4ppZE6KHkAb0KaXjBVZDxZqJNrG6aRzH1OjntF8AnnEq6UvNTMR0iaPJfbBhMU
hW0piQN+nUxwCbsRNUkreXdUtO6Eob5EIZ9RO2yFLuZ0pPfN/87WltjpdkAeKnjVO0FGKdaIHDr0
hGKSdP3rwPeuEOC5UX3dPVFWKv7OwSUwGXvmKdBIYa5VDyRahs1iiq2fM9NbNwGJtZ5vyz6Su8w9
EE+jmsN5u34YThR9X1Ndg8U2sOG1yGxmmfZ9qQl7dfj7meSp4mTF+oDvBOkMSdo4mEhCyM1qwI9+
BKGPQlrVOf/xmUZnmSZvDksXU5GpoeXsjMI2U54hy+wvChcNd8xbQpVFYZjbjItkjUPkkDqCS0nD
e/6CEDKjg5mZoNN0QNK9ZxFszIQEhOvUNUed11QJK6BJZq4Tho4kR+Q/VCjU+RNP4sq7RlZwue8Z
fghfxo/wgbNPvB0XZkRQIZri8/hCTjv+h4P8bWDM3GWZcnYE2YGxhHoL16xinZcpGQTDlzaT+K3p
win7/ZhMM0tGXmnP/pSBIj8grwJKXfucCSBMuAEit0fw2lWItpQXDWEKQCtwmljfN7TyPQ5RbnQf
+uyElzca4MP82G32kYm8ibxkXuRCaq9W8y31yAhT8N0Ch7gEfCPEeszdbqF8viQehUcXuX36d4Wo
Sj3tARwW1woaozdC4FYQ3aVxOeWlCI3Fh8JMbT0JSRyPU3Pg/qu3Il0PHFOzPzlBxONfbetHP1hz
TcMxQ3MmLo0IW0ncfySM+jH2BM7wDaKPRDg2B257k4RjY7wKPBcAJ9MKNvzqzMHibdGYhDFZ+CYv
mqdA6vnsc3EfRdw1iEHA2lvkXNJOPZ2s0MhoBMG3CDN1jEJ4QF1ICtfNVnDzT6PgyHxlEnsQrz2c
oq9oAqTez4KQ6HmtG9z0Zggz8AVSU4YuCFDRgOSvFjaNRjMIEew3SfOujrMviryYrfzYczcvLosg
2Org92OpEdVoVseWkcP23nWKx+0xeZrG7E7pA9rWN2hX+QocnLMQFGf4sg3uf5grZ8nwnnJKnoWG
5bTIJ+bXmO1idgZIUgTNII50Lto6XUeP2j9GJRRyCRVQls/gsIbyf0sDvbHf4zKgJ1SdRCbjuKt6
Djznyej3G7JKOA2sV1HHVMe95iJA0i0mvJ4gnfw4WTj6zPL00f4aqe2FcxRyiMPlRqOWEjeHS7AI
0fQ5hdSb7BLxBbusWj5ixSo7+DAX4vPe9B6T8GyBbCSYg1XExG/O1WTH56kMjtzfX3s5DOELE9YH
NYXMgHBC6vBnR2gSPuAoHdlmVVuEjbr0GVhTHIptmFEgs1BudMFTaHKZvF1z4M7hgUFOAdJhVULw
8h4g3P/KE+l1vMIrVBraa/HI8NsIN3e+NDgII09/5Wk50Ia6BW6XZbsRp2XpP2OqJ3dbrvQx73OX
GX/8eKxX9YuFS8asD5WqE4bhTizQLwtPYyYpcfgKLA47I4+u7ji2XJd5pA4TqOUh+C6DydZHvmIe
3XWPs2STO5oVOKRvkRd2SbR2Bsjg6+DniIznCYt5McT81ph27g+BNqSR1me6RD1hmKd5oaJ9Se5w
G+cErPgp6DaA4XHtBPXw+v1SCy2O7bfUiTLKIVbyVRiDv6IKSUNP+hJlX2WfmDk1thHv8MCzhpF0
+V/P3Yax96u2QYHmAav70UKYUkcAboNQTtfDj2gVkz4fRymwMoe+swpO0GbPJTELo8EdvXiR4Prt
amUEjtveEdW8tDqGW+dwJYMCEgjyGIPXJY8Dn1yfH6X0E6Q6SOOHlkF+EVZshvkxzvXdIVqxapL8
pbRlKyFll0N3qMlLZh8owlI1uF6W/ioQSELQS/VuNUZJa7u/EaFLJJagVVmUeZICx4UEqLhXhcAS
/9/Mt7hRfbTQqpP7jQc/3UtEma9GB+0aO1qS9b1hyWMERMuc5usVfEo7x0CLY4qItLTaTVfYrFUj
GfoiVhMnzhXTm01GSCJcNihgrQ4V6h0EJIW3n8engmnmmFTkFH7ugV+oWbSzEQelWLeYX2zsgxMD
Mf+jeGBYPqUZvT70xSGzPWmYzgfkUJMsMsgOdGcVXOdOUSWMDJY56i/owYCLzPK2BilP9GP2nORa
XKji+u7SSbKrs7GET1LhLpJf7suZWgE+HKXwtwT7rzKq9sHgBXyUSIctLI3+vTofaPQ3LwwqGgjo
INglLmtAGecP2n7YsUMr4vWvX7yBpzcSdnsivyfn1pq+QlweemUgaTctlcSBNK8pPnxc6xZVUDdo
5q+F2VtWIwTcnEKEQwZdhGqQhhwhv8Pix7SF3mC+v9W6DaeQYMVV/LRLNOoCVO/zjUiLQcNSAojP
fxyuUL2bG3OBbHfcPl+XsNZ67lILaCH5bM/8aqyFbQ6UMPt7Cewrm0sRkwYU7n8XvIL/tv4xCrGz
ugOZS49uHPNqKYVNWLyWyTPSFk7h8jmtw4ya29oqwPgAOStcIsFVMdkWkp+Yt+I5mFfZuTz5UOfp
Kqli/8kccc+oJkCzsWCY/8KntGV6N5fcVmfQElUVoeHGjAPcfKLofuTCyDH8yBFRyukNc/5tEbOQ
ZC20I+vpOmpahjFdplnCgIn5IbahK+Dx+lS/oHTA6Lf456kZal7LZcukUFMI/Vj9jOcazRbF4tt3
JstxV9uGPrzB0b+1YMS0bUfSzAEPMdKQs3W8S3tMABlF6Gsnq+EPrSN/WvSqpY1OKk1+qMNqOtIK
BRH0S4pE7bCiPeiB71R1Lmq/E3bOsXZI3XxePIdh8vAJWAqmbA/6X4keb0mxJ4MmIG2Wrmaak3S0
MI2E5uLn6mpPup4D255jLN5v3dVFMD99CrEhIeHDoj8TEK7+jRRR398HOJCUM9NDPvxrYO3VNqvD
cy0g8M/yfPt5u4s0ukLrZZMG8XvSg4Et8OyKRRA70zwz6ucA69jjVcn/MW0aLfh5FmwWwau2i53J
/CroO03G8AVMM9p+3TRq5fqXttodJZzR7ZSqRuL1ifpKMojmAaTS0jsA27pwrl3Y2zO59VJ8Z22d
RNNZg0B/lxnLXAT/sUE/a3M3QvHcT0f4KTLnCjZPhxV5TohfmVXXDGNyEP9EZkrpwBiLEBb4KPN7
z22ypB8B7n6PvWVI7RjioBxBLDBfUO0b+6omnPLaxhm3UJzt6Ni/cR4pSUqpw7Hxmjbo6OFXm5af
jHrCmxa2QF6V7Om1+qn2NdWfniJeWydgIvpkrvVM6hZWiJylTaj/cTFKpcC1gd5j/Ei2vgSA1obo
g7+bRUqqEnngN0S/vW8dAX0c2dYw3w7d//qOyanrOhvz0JFg0zau8/owEO1SiVytNk1j9fL7Tujt
M30sqRrg/2apESMpWqAg61iTSCW6TUcBI0BDsZ4HgIjQ11Hmf7iZeSOpth5lUhv2mjDGDIJNlpim
X8wK1iIkTfMr5uX9lii3WinAUgMJEVkI2a6WeTbWPxCNrG91pAnhiXtbxvJw3neWJbrd/Ri8Tk5q
e2tgTptgFRayNCmNCW73+3J5Yry/J7Rq25ywWVntODzTlZYL9FPepIRCpFC2kkGnlxMsMR18P3mR
urAbskHAiYSdSg4H4oA1x7/0fN3JND0J0rcqQkJyIiEgCNaeh3tPuU5SPmpxaTYf+ilvwsc9tp+o
7p9pjWSsZXzktFs9VEt6gT8a4GDyhJ5rq0tAL+Mhs/SkEbX9I9Dgflh4E7iTvip3t2pwjGUjiep7
vlRZ13FQZFT4Gir0Mzd5mososJrpEe+ZSqdS48xe/2VecQJ2IKB+KZgc4+GRm0z2NyP0XTfrIODo
laNRmqjWdQkVwkQQoEc2sgNDeTremUYqbqD4BYdMPOmNmK8NQc+lojRcvSqJz+xKLhgD+bqVVP64
gSFB5kzUykcA1zu5U4+ln9EnlVfU/7p0R/xTFDIe9gEUZj9KJrPNXEcPJ1A+IY4Y0/tQW6Ckc4X6
YTy5xHdW6kxQHbsfyCWSnNugTBrshSt47ycQfkbDKGoOQyJVTmzIggUbBvN3dWJgLtU7Jerg0gd6
uVNnKkiSUEAAz07us2uA/D5hZsz4L+FiyztwB82h1sZ3eZ4ZSc4CU+MYTShyDAOy/zZ0lqYwLEJc
8Oop9rE76zjT8VLUVv7Wl/KBI78gFTksjGLqrEhZOulQLRl0xwSnA0xqSJbE6l1cE+1eHYfsL5id
ZPRmoz5ijAwgU33fu/7Q1JtxCBIbHvnIfI+qhpQ+qHYzvNTOeWDnvKEbgbJoBYz6QtZLxuEqLqzg
dhFHPc0qzHo7JeZlt5z0diQ6P2HAiM6iPscBXjCw3M3ahbbud6lcNll+bTE4lXBIByDlYk/HieFt
PGrHZIK307EGjgtnEIh8ltCW5SDK/XsLx02cDZSrpyFtVUD0PVtoPn+PCYGy9w3SQldct+/gjdof
1QzsnuepVRe5WTLwE6QhZi6s2qmdHDWxjE+S+V7Z2cGHK2K/NG3OK5wBICxzupi0//zPnL/YUrUj
Q34J5R5LTTX+KR59TMu1w247HCKuwSOd3Ng/+X+5QYvDXZvgEQa9R9yPO1cbsimx72rF4NAY8Wai
9U/E8BwnUbQ5dvAQHBSm5dPxYDsq6Qab4DbX+EwuqKJm+AK5YaD+T48tqbpNzGvZ29CRm8XGyBle
8aAjupiwKm+Bk5uDVjuOD1Q6P36gxj672Kk7RcgrelmiQ7mQZ+j7868y6hGZCo1ZOwaRGYPdREYE
fiY2PSYMXRc7M5GoxEK9l5X2FG6xCvGeSr2Y7VUMXo0zTdUT05lnRP3pmqWmPqv68gqilKuT9RMA
GB8kWN+4zuDx+BE9XJZTZiFZFajdkkfdG/NmVkxdJYCXFCI/w0DUkrTUH1N7GybsMTcjDTHXsqPf
lvLsdBXrlbGJuxonmuj4OgW8puq83gO7XyvHlWzMjK17mX4Kol1CHumEzYA7BZc9pLseL6QI3gDF
PmOKo0Rcpmy3RYgW6/TuhSF72QfeQnPa37esBbiv5FJgEZERsR307wIinrLhkRu1/y4fPTQ4kJ8E
NubaRuc/ebmyYM7ayVLcFy4Z1pHUtOfvgWQanWz/hHHw2E/a5j7Nzm1P8BTkieObJqROAjpI4DWS
xlMy3nCFOk9LRpU9FUyloIKP2LV3mtz0gMvvtba7lAnK5il8RmcZtX0iaR5t4MpVqtwOwiwY5isA
vB8k+fbHUHwt+7SLtuLOWs/OQKK4LspYpgTirt/LsGuaT3mdjmI6dzMiOgwHzxNdEgOBV4/iE+Iv
aSa/CrkJ2jsLoeZ/ntWsAVGALCtD22WAEUOqA2ex3X3sBcbg5IdScGrH98QaxfztkZXUWND+UEgO
C3YueHf/i8YelG2H8DWZ0ViVZ3Lw89kHHUvNr3LDu0pY2chQMlJpj/LBE51N6YGwIuRdSWIiD+yq
9f4ifJE6hWU9QdyPg4tTIOs6XTHYZRa4eqto2gQ0jzCw6xAzZQYp2uRUg3TBz1bmeiC7t86mNzug
qDwgG4G/XCl60SZV8sDfXaLJf1DkqZR3Tvuzrp1tYlvm+LzdtvRjA1kkrZPKcR/kyufZmNAk9CGp
Vm/05D6AfHAkGTnw9EYnflbo4mmggUu7udhXdZeX1FdDk8GFDHbEQ4JVboHxpAeDPJab8Jhj9BQM
I13rmpTJadrH4RXyKg1GU6+RQYED+T2cpz3DvpXPzi4FKp2Tgddxm+HAteNZXuPztYVK9PZPKlnE
6XKUySQR97+ZfJ/xbqQxg7iNwn5gsiGG7Wi8IcyfyWJUIjwcA3u8sK5EcVcn/ce58nyYo2nEpL8M
KJ9XYvOX1YDq62n6DRlp5mkhkQLYSBL3/nUPe9klX77XYPtPy1D3dQtlXphZlJFDEGicUFdoALwk
Is3UFZHBhgGkQycuDpS6C/bKMaaCZCiUhFxjZxI/DggrTK/GF3aGUHP8bgiGJA6lML7vT0LOgK1W
pyAMgUWtH0nDLfjXUF5PtMDRwJyiV5bxRhteY3X4nCxcrZwMvfgjUrhGWLK9HM4Lpxi4zHSdZdac
DNhhUSG10rDDzM12+aPyqsynpTK+R+WGabw1V5/wGUbkTKRQaHa0/P/0RuyDlB6swRL1cbOW9BiE
pMv7gmRk2IhFAC7+JrzuHtVA+kSApaxz+hVGmna8hQhefTSLjk9Gac2Eg8yeJXD71YyCl79WjYnH
vjXMu3FnmIvFjNHXI7vB30Tsj3woJbc1Qf3HYoH/tRAQOSvvMfw+w2PrZxyL4yO50vBKsC8GsrOV
N6oj2BQNItUwebV39qC6cj2RmnsuE5ITIrHXYRDvCfxD5kDVkNdm+cALMnf/mRYoqv0nV/QPQCo1
haSKvtDqTT40dnyCsHHcaBv+FmyZybolUm7+oH81L7tvUSlf4Hq40FYLX81qesVURw9tT/gfh9xy
w4lWVzgbQxfqFi+EpJJrImDCvabBEA2cLACcf5fbQYW3P86YIy2hnWPriCYVS3oQx5TMz5nSWCId
dlKsOco1Rd6dc/ZxJETj3FmEOnM8kChWQG5/g+aAnXs9oposTsjU5b5DGT6kvl0J7JnPoHzINEoL
guwVW2c8r7YRSplbX52YahHbVkrRt2BogAbE7EtE3DtxPdF6yWJwJquxHyZ/+cPGbK9G35EqLWP8
HxGlQNYytmN0pyeYo4ROAzJB6tmx3F22XeVh4/X6SCI3QoYR+VehFOf6aYpR/BAaFWpEe4ayuCEt
VlLS0cAcCjr0NnAfP5pS9DQm8QgQ3H42nd2U8JNt6Z4a4sXb9snLyp4gk+9HMk1V6HgClQBjLnsW
mfheJTydiHNvUH9+01yzg3lkqsWSr8/kaDp8yw4d5R1FTvNvoaJdgl9UYV70w1Qqp011lrs8nZnv
a7KUcFD3qFrLKpQH4eV5VcTZoxHC/i4ajzKNnxu9AfY96Vig8ZXzAHJJ5dYIqYGyH5wziL8dV2ae
pmO0YCSH71CQAMB6SJSXguSBCDDUIP5bdF6V7q+/0jsUDCcSAb+4COJ56j2rLTJEB3/d+EJGKFto
O3F9oQdtQOc2IMDo0UzTyAeOj9xdkj0kVbDJAOIYUn/Fw8rsThE/zeaS0vh+m3I1ZO9Y2zwpTxMK
aKymAuvmRp07DmZvXWSto5flcUN83cEgowMcvmCZscwo55htimkg9A84RSBvBn3v04jV9spx4osl
NX8+Qjs+7D4rDG9/HirYRQ7F9JAuZgawdUjJ3eEiNfjuUxMKGaZrqTy6YW8S3jbYneXkHPS8Ce49
f2WIiODOSdwuQTl38W5q5b6G10WIrQqXLQ03kDWgKW5dr8aDg44jipaIs4o2GDHb5HcmBpm4E3rK
j+/UbHwVEuD8btCmibM3fp64Ii6d3ztwym2LIpRBDFojswXnsHH2oF7iZOqXYJxA/9AoHnJekjZ3
v5mFvxSwZt0n7Z7l5YJ0ISsXOtFzJdM1GVun1I9btfoRUki5TbUdoGb0XyD9SddxirwI7M7X5kQr
AR93xanaXCZVWUz2Z8wZZzEc+JBj2oYLmQKyKmPKVdfGdtYKceNhwFVo0gmOyhqMFMCqRT/zBu+6
a2pJLzHKqaZQIv4HhE80klVdJgXDQEXktHGxVY3JB4qPuhs8IlzbcKi/dxMOR1kPRsUEWrMflswQ
JgOnof/iFsG7s4FUu/4bGKADCRfx5BP0+uuVl5XkLlmsP9XMxIcSbLCSHMHooGQp8zkCYwR54TRY
zSilpCVfc52+AwSnzksvtIq/wIw8i4zJl7UjvHB67NBjZHmkaK3mo5Y0w/yYIad0liUyyy27CJtj
XZZJ/Y4YHF420b1fS5cI7P+A8xdfKfIvScrFMi2VsoVMrjdIAY89HBFRQhFLpH9AvHrH2fd5w6gH
1EyIN/zWczqoP2ZI5Y51KCUPaN48rWa6k4oSBCAmFZlP1wTMinxZtFzgeeC8WnbL0ILhpOxq4nj7
qkA9fiOYYkHOl2ASOZ9ftkjHaUYOX1SFrMGHlc7QaVmf7YRN5Rbxaeba51u/HQR9YidrAC8ywbw2
50ChSb1qe6C46v/UGeF2vLUanslCMlvSCwcPLZ+YbFueXMFATQ9Mp1Y3etkYdQ/nUQ8P1piGMYad
28Jf6RpbrLpq5ASNwHkjFmsVSBpPnd5k+OmWc1YEmyqMXQAOaP8m1KaW5CBj4jQR+0Pa1UU/ZDwt
w7b7Fchs1D8JLgvBJc0fZFC5aPhmmr1FYcalKSSVLJWcbQwkU4Z0PsKjoJnnQ/BP9wIdZXo8D3IO
uGuLbcFXOOcOic3iHmoQK61Jk7jcr7vmznly4A7Oo9vfRUqcICRa0LiIkzvlUHOxj9Ed9SE5+bq9
jB0UnPxvrHe3/JlGKeFxq/4LtZNNBf1TzWKckR2roWzIy3ueQo1PEft9PsVzGy5utqgY7E9JZQB4
ZxixmmwSAl0niwHfXNaUoDQDxzkZyBklJiut3CSVDPHaYn2uGjOIH3Jp8XE8jPmS0XrLEZglVGNY
wXf0c6/wmdRW6wcFEDLT6/Rx9taLT53OvDbVX6nHnhd2YSEISofW3aCvdBmp17q7DaOlvWIpf1dz
7sOWfF1+EcVRe5UTe9alQ0YWfxptvs5sYG9OUJTaKxRDeMX35TiGYK+BGGj/DEuTW4yOuEk7l+Xr
LiqR0KieQG2JLah6UziWEEEhMwUYW8WHZTRChPj9QPajMoNK4pb4OsK7IrmgHvHvh3QD0asvBT63
BpxRgzaqH8/ag0jbhM2dlB//0ryM3A/Qvf3omPsqweCJtSE8yDnDH5dDcdKQzSXZIE9iGACNHMc9
7tgNNACz9zVuaGj1/14M5J1snV7UKL/N8spq9kJA6sj0EHz/1aSxZbEGibvSrC0asifVcFxywwDu
XdqWSvseVOibUu4YlKCK9IiIY3EQgxvigrYO64Ey2lXjwRopTdAOAcpMsKWmNP9I+tGsrtfL0iE2
bAkkS71rh6Qx3SjnxAgX4lEgJplYIAh7yxX5jFZ2RW5WRBLS3GFWXvHiZ6FCSoSM6bc/UmBy7rXe
f3GyurMgmW6QTXlSYSFpjS8NscJu6qfr0skiHEK/6Lj30WbHjWz37nGeeKzSegNmTGmMVBy/dV79
yP+3h/l8CMC0eC8h9jF0IOy4W13PkS1jDfansknpbISdb4JeGo9j2dO3Gji72vfdhOj3g2ymDrcp
MgkW99sDEPiqUvpXjCKlhNiEDUCKjzf0PZ+e7ROhFIMLw58QomSuN9Vu5BZuRWGaoznryvp/owx7
VY/uLqP+/yhnqr817gNaayvp/CV4+ncEPUXxJ+OJBkHcqLxtsoyzpIv5y8P3k01l/EqvBew9Njt7
eYzxaiVNnj0Khjrhf2qbf/qalrs4R6X7ActPmnz50Xg1K8/Hp7UwnT4GYsgC4HZEwQS58pzW8KzJ
/9xHLxOoFRIEhoYInY1VMPYZdfTcNfeGuVO2do1vuIqT0gdnNp/pHmT9QxgbSqdSoQwZUZ4HnLgf
dYKAzVPDVtCjDIRVZ5zDOu0CS4CNXb/yd5jsV2lR8AHMELX0feUkLlhfvWSDSSfE8XnQrIPUJBQ9
P80sYXV9QPKu1NdA7wisIibd5SiZKeNj11BkxBvq8R+HvBp3qRpxK3iQ0URvJujnWQVg5dIquk19
dHJLLUQ3i+TsKUmLz62NZFbH0iHbAQ+av47f+pdNPG7QAuD6n5xAHmHKJ/IhWGSSDBQpJ+upGic/
HUisl7t1De12YLYamQsRE4UrfqcEzxH9cQG0U2bH6+3rBBWKz8bFa5yJ2cqwq5/A5aoTSgu9Bjwd
bDO94GtmFEEue80cPDp2hsDDt3vJep0xtat8XjJg2dnDny8FVa2ZF4dkYDStxeE455APZ+6UG80W
SBA1B2MBvOE6MG0rKAAx7uFPSebn4/vYetj2o6xAs1CX5D/Xnn625Prvd0OuM0PJpBXw9MUEsa6w
tEXGsuYYptYXKNBXzP1zuSv43fkKcR6n7WK1WlDTaMifyR406MDQCil6jCjZM05BO0pDCKlztodD
EiNa4IYoRbyJQD6bKQGXFPbNvXTXCKLzXz0R/EEPNXu8A0rqTHdBxUTq5Wz9wMLvBN5rGSziWx1m
SMUJrE2+JJaxhmlunrtvXZH7jias6H3nE95zZqCSFQBvEKFNMWAM4VTSfUrBGYMEmjzo2hEEsoJs
KuLgARzsvU5MHvbL6nmoERNybTnuAOEIq/NZMBvKj+6J6jUhP4v66Czd+unT7dUaf+gyTmjDjrTM
AFNDg88HtSbLnHS5pUYHiSkYb1YOAjx7iENvO2krIh8YI0V55PundWTw7Yhm9ecd8w7pTTN9PIW/
RZ6M1mShmp19MjINHq1kFbn42adwTTDb1Q/UpAmOM5Wf9NV1oHL7kuzHaH8czsWVAH35JJhO6XC+
15DdiXHUO/XvfN3EtrQp/bItJy+Te7DLAr2B2LXTMBXZ/uB8SBS7RNaQm7hSM93Yw5ZMB5pl+QED
dIkbh8utOduVdcW3Er6MjZCbeKRTxWUsYKH/f7Cm6j9cR/vUfZeBKA3dcBfu6VbtIo9PtLN1bt6W
I+t81EeCzWsSNA1UBkMwOeMsl/M5Q1692v00IA3g2W2QlEPPK8c3bXiX47ZXOAupi7OnG2DT57HO
m1CqieTcUYDSfaUyciDu7AmnAPKJApoFKmfv/bfjulMU4OxzK08W4UgyPE6nJUV9dUZI/udOLL9L
JXvNDJ2yv+lq9AEGQhFETQRkgymB9yD50bYGJAQcmrO/ZmCuTu+aCrVSAxi2IiI2sdiKBADymSy/
8zbxgQJHWO7XcQUIlZ9t0O6vyu6ts8Kcwh9/0uwul/WzVfwpJQwp1YCSYUn8uY+2MRel5ElzjwNr
UYLvYmQwJvgs6yZeWsolxy4uUH4pOIfuXmmVAk+abMywyZQY+zo+xT8JEzQ7ilX4xJw0xjxjqdcD
ilUji4sMAFii0TtJKjHJug+vcIHOfKe85kN7AhgzXy5PHj/ROcJI34Xc2kjFSw60S2lowzkp25tB
34vlYlF8Sm8PsOC7K1ZbQYB8BwfYL73ueL5XL/mPCBDE96ZjSPZpmINYEIhB4vE+Pr15mUOM6+at
SUWntl7aCunDSreE+hBa5L+W/70xQCqjnDCve2ySH7f36sc8dbDhlp3yRa9sAQcP4FyKm44zGzN9
Feb6ogglVOWJaM62O5K2aXY8/aD1SszSXzgqP6iPX1Ur6W1e64SU9OLym11MMYym4wo9QyomI5PV
shkeq13HFucbf2BdPcifFk1rjS5PenK5w96lv/+Omuf6o57qyRCJ7xc7UKQ/AY/nKBlwCEBQhfMA
brRfQv58ahedcS4Z0mfm23zvw5YgDBcXTrDMfvjYaVeYBvKQmTS8NwOAOv54FxUN/HOpRlmZA+U9
DRMNcQ61mY6eZYtOPkqgSw/XvVBPO162ojFdKj3ME5yezhaws0ShjESNjmKe5uhdn1tUGXdwEDRz
3MqLXrFxzeN9jt1LlbQ9d+dd5VEYxxiNjMgCNM7PUxC1eqsxGuJU7mAHdJ2CcoAR0nDasORn2vi5
8h6AQzfDPBpvk508CDT9VeY+i8Jr76cWCjR0IXcN02IuLlGF8MqJ212hI9doVWmaoZwCmyErSo4O
/HZeUM7Jlo6sEzjb5al1EFDWZCGJyT/I+ha6h1b1t1WNDr1nLeSp29GlsQgOJpZl3OBBMFXMSLus
v660deURudCkkZrx3HajUXzSgamGxk8XVH0Jkj2BwMPrUXd4juHr0smDyxOPtqEBSsLf66IZfYQV
cvPU3TgD4uGsuoplgKBTuC2o57uqnaCqE/tLWPzef1W4gfpkX49gpd2ih0udeONrIL37qDtUkSLn
wUgC3Rsrp1ISsrtsjhVAg3/sdzVWzFlN+JRvXCQqHFOUzVgeMHQ9gM7DMAg07FtOp9KblqeHEGGu
MrbNN0I/QWlMM/1pXkbOEMI/hVK3xeeFcvJEMZFjtp0N0FwL0yHVlr2jBCElQgMsLKtTJy9XSCM/
jl9+W2sCKFfjA1reaIkDO7kCiMDOhDNUGb8sNBJITGF00tdIcqDLAh61cbRJfpWa/v49nf1zQXxv
rOPb8Au+gupcutSodL+D0S9q6G3nceW42b4BOO++eoPfWoFtkqsaqyxOZNj8VNsnql8PPAHbt0Sp
JNTcbX7jyKNjvMBxON3KBO0RveWgZOBcnXpQbB+xdE/zhTimOKZuqAcWF4YylWsdNaDrTHkbEGSD
eHMgdeu4QcXVqaBqGsjkSwWT9cIhLWemyyitu3D5TN97hEIYQ9Nhqyn4SNMdncuXk5WsbqwNGl0K
RizJGdwG+t41KJyrl86rzAlBXSf3r76PuFT8yKNbDpecWSh8ljZxvzpzjfsbrWqm+kJo8qiv1pjS
Eg+aa8ePFDPFV2y/D9bgX4E8QRe2yxIzZqIsBDPKVy32fgfKl586zW/9kFQgaEvh+69l+b5OyW73
FAKn4X4XxIoPdPLxFconqb2N+8C7xy8g9OFGaPMRbjKIAH1J4lQD87JKG8iQTL/CGUOHW30U8dfS
U515VZgiuT6DyIzqLgW9mGBkwIGxBqMRyaXqAz5A4X481WQF068mmzGwnGlrnfCMZRWVBU8cegLe
WzNX7zCGhBtOG8YZLy2UGXsyuxiQzov0o2UK705sl6SmgBvQDNq0GoQdyfuMiVfTAWgLfcdyPTZ7
Z4SvtQruwa8oNIynTNlnyO/hJ2hlfnN5t3C1f5Mev89C4MA9Cm9F1Buu7KpMXnBT5zxQOGKAcTTQ
jPhn20JAi+Nz+7aBgjd2u7Tz/3IGcrpWhPOPmOavMXJKUDSKQrR2if6VdBPaWXcgXJn1ZNJSFvG7
rMfZGlDWIIzfLgnbEQqAq2xN5/EfzfmJwC98WeePN8ngj8/lu77xBQMPfiJZI941fWbGlU8JKj7U
hbz1l85lcma84QWiOG5yHX1Ek1PPKJGVvWiWC5rSMj80QP2Sj1h3RgQSLMlIUi2ISpLRh2ZLvTCE
Jkv6vZ+HFLinO4mFoRcgE/NHEb1bf9zac4Ou4rVG1O3EXTjwE9Kr8NVhEfew57HNWlqIn10jOOue
4DszgyEou0e7Ih4HuAE+6ijTjH0ul0FW6AH1/5kMKyfi9midA00UvCraFDc9jZ64q9Qz2PBgvv0y
dY7N9ojQTPLuq76w3VB1ZMqta3FSbbFrqLPyeSZMYKv8xdUTsG/lWh+K2Dcn1Bm0JTAxikphrkH4
P8qs9j2M5f3XgWx4ljg+b/GP3Q8jKMLpWU621j2hrLW6gSPJ/TVMvQgaNfyVlvLffLlH1z7sz8T1
sG0F9kf5Q2JOkjnWRzgqha6DKW9aoWC2nkzR1mRM+JBb3G//yyZLQ2QlvHT1NKhK7Jc6LW7TOIMU
cMviFxTYp5s0SDi3aUzxKpvknJxNdtTg9vIGukPGkc0So8mSqNCa5ecuhArcJYvk2Hph9qi/kns9
zQ1u8LLq/1mOv/giFqh/2RiWhPDWsi+3e1mRJPIvyMm0O7/oC6coK9Gb/yNxP3PgRhR+5L2N3OP5
83u1RXW0aa4bh05WBxjo52I8CQwQkBTMSaimTc9OldQcpaGKLg06zRLlFQFO0uENZC5RjC8c8U88
1JmfRbtmLW9Oy7vi40euVoVUlzlFcnD38QwPlcOusl+zoaXbxSCszPOKL9YBQ5Mhsp2Z6ujgAUHT
rW4py2mH15DJcjd8xo+5DYh10nYMG+yC0cl2rNvWBHaZle1Xx88c+GcCuf3QeiaCWSy5M1QHyNS3
qkQDIAOCiVanUPxRo9U7MUTvGJjeomw1wZMnQvMPqEHa1L3g1dXpkZZTsbkkCXYjwymX19tdrb86
Owxy+ekHFtohOEd5cau0Ebywu642nKy6p8EEIFpsLVcCvXtuboAMGzix7xl4QftkImqtdzS/Ml9R
0Wc29Png+Qxbn2e4pfk8kjP3EmGB/Uk+pN/Baqnq04M5BLzCcR6rM9sQA3UfPPkYhJE2ptscsYNl
NUccCiLROFLX3Kp5Z8i88Y5UIlneVu0xMyxzp+QderuG1dP1Q+1LnFR5rFBz+Des3fYZig1b9nb3
yGAW4eVBhsUI0hkDBjJA5qsX6VrbefRDMLgMLej5x3lqn9ZCrbmAhspMWAjHFPoSTw3muQbqDeY+
4sQfhaRzZAvbhcj6bd0GBBgsnT3VI9H60/q72UX6078SvVS6A3rzSiGqQ7fyW/AIhjuTFbFXzuMl
RM04I/6nbodZAbF9y0R/yehWYZZ8pr5veHGOtUPemEl39vo+bHcvn96G+TW6lbc1nPCvmQ3DFeBm
iDgtgoZ6f6RRtbn7J43J0j6UUQ/9NvEOJj5YZPyQRgsNw6RZ5dDjCZ5JCT4hTRr4rI4IcsH6cVoc
bOq4kMHXkRzKcT3w+pe8fFAJPY4YlId28t3z8bmwVDjm7oSxgIfOldBm9AzYT2WpYF2VcZPOBUgw
WiqvzZqljMUcD1sgHCKFn7xNN142SPcdrTaAAtNuK6F8ub+RO6UhFkDLiRGazBAGYpxjubW9ibvo
ztBFZHgYIMpwtMl5J/m60ISPBzzd96SKdVCiQRmrlPAKyShq0J83JVLeot5++xhX293qqfem9pWO
Ek8a82hGMDT/a/x/SfgzUvWwas8py3Xy1Ej1BQtw1KPkoOSXuu1hAU5+EKNXO1JG74V/kjPxjVbM
vpkd/uYaOOEtfWGkYIehnO/MgYx72eRYLMO/gpz9fsRrUHavLxRtOjvHJWRozmbAZn49oK4p+LMf
JXGws4CmB4bHVcru+vXpTq3ISG9XyDyczqgHwvAMwNx7XfuRL6DpHhWQoiIrePdcuxTvATAyjWsA
QMYplJuzcMybSjcOFii0hfZwHev8likPmNyHDZdB2QuElZKLZU3BYgUu3YFiTRVyCIz9CVB0Rkga
5LRasWF4EpiymRWaQo93hU2mnt7hsqFKd//JaXnoBlty0WQCiEfiPrsTo0y9UDmJFcJLLZO4V1LR
1gcUHPl2ECL5rUaShVCTLf+FGkZSkQGBGxB0wzkpeW0a4CmvWmOi19CiXrH+eZCmDoXc5J/Gh/6T
9OfhQzeuu6GPn8LDHpdkSo8KjSROAV2KdVSrE/dLqrAMziyYsjKTlv55rf/r+zi+2pJTF0ZUMesr
oRjY0DiI+X03iOPrgWGuhvGxp4H5IdKvyyh13dkEWQP6PaJ1Vi6ulbt+DTmZQOTUsfTLptMmNfig
jMJxvz7VRF11O3eeMQJ37AecfKiYjEv+ELmV41dEd63gHz0AkVOJ4TvPxxV0Gj4RAx8TmT/Cknnj
bQ5fwZbePoxR4s9SeiplpQ/rKEAJAymqrvW3mxrlv5CG6+OupD/zRF8w3NaCQFUrX1xHNKSaHNH3
ct3dFVvWT1Kp9KXbAcTmV1yvt3aTk9PllOvyxBqizq9vdHYfxa+FJxAkswYkWnjf9BvoO5UwzDIp
yI82fnulEFppq8wlZATOK1hUkwwrIUDm2CCWVMDUf8iQIrIov7Urxcn4S27Z3CbGN3qhPNNbc7la
9O/6MA+xS8WXPUZc8YctsuwqcaFEIvvW/zzbJB3DTlfgSh4OPNtGovlGsVcdIZvb1EzDD110pr3A
uktup/QRpWbLromsHdjYXY8YBrk0qtpygP8jqd+6mURazUseQWhGbLplXp9HIpjxzUsMKY4f/j30
2M+GX5x9u8izksLKxFM+uTn36a4SEzxzWs2Aj8rcLnpcyl3JCFN/mGMWXQyy78J+5G8yPqweP7tF
zWkA4oq0ruQwkW2H5GfldvQs/ygu/XskHPuju46XgKOvN7WTwmX16Si6tn3/yLc7v+lGmR6pRy/G
qazA/5jiXMOoZ6NyXZReC3z8zNm7bdrxB0p2DNUX67vJIiKCd2dXjA1GaEH9WV5NKYcyKe0xZ6Wd
+i37IlulMm9hXUYyD9MuvAaWmQNtUNz+VJc7cGe0gzNV+O9WS1w35AiISSpzkYygqYR1qy4zuIyM
BqaCrctIjSRf2325l4xLZeoYNbpa4kZnYscr9kkuqMIRaC4oh/l63jmLBg49dUnUt2A52QEvu7gw
l164KB5y11nBcrxTnhviWZSNmAfzhu9naA6PyTBCERXlwb8Iaa/VEgZ4u7DSJfMxWLNW580dVF3s
P98yvW7nwWBZQSENg1zQIl7xtEQr93vY6X3n6boy0q9tjCfEPzo5yoQtVS/cdwEA+qyo/vrKT3IB
6NUrheFPE/7Hd/qO59xh6pPDRsOOhtTyNnDDs2dveWy34UT9TJj8IrgAfGme0tXvHUf0G0bis8MD
sTCsTrdRV/xGIO3VkNkRszdVtn8vJS39cyl3cYjVFWj88AQFKmb3Rlm1oxfy6rkIDB/vY+Z+8opA
gIAHkeJ2COLsgGQbsw943Kw6opF0aMH3CSpod1ZyGsdZ3mQhFUNv+hRblMGKZMZfi3rn9cauHiM4
TVgaeBOqp+m5ME/66kcGz9SvX9RAKQjkKNRb9DKbX960krKu0XHVzabGV7KyQ5z9s0j1agylRO7v
uaZYoat45vSbPEeBUVGQMmMs4J8kxNyANeHTU3lDyuKsk/7G7rjC7fb9eVZXB+tLdQGKl4YcuBdm
giCIOWTB63pRWeKMBStMXSjEyowIIYAhvv/BUgNVF4U5YfdkZwXpbolNI3c81ro4g4Lnd5SkwGAJ
+nIyPFg6CDpT7a8O7VpBtQbqW9cGu+GxmFeKsvx7cZ6iK76XZy7fenVraz2bs/RbwcHY9TO7x8M0
q2nIv2TnejMtQ1vsjQwEj3ydEAIcJ0jp6ZjklArJEPAxSgukKf/LgVrck42fY8y51OdbiYEUkl5n
698tyEILk3zO2tr3cSjsPJ6nuj0I2+R5TTE6J+FbwgHaMuh42Z6m4wrxLtUIbd32vP7sQqI2aGCD
fUyrDt5MmbffLz6b+l2bIk8C85jdy2ou1i1pZmJa7saeqMxZ4BcSjUayklOak7xM3wS4l9dR/Hvr
2eT0QYSgXyomjlCetHeCHRS8z62rJNHC53UCw9e05738IQmplq+Zp3qaBbhSpL7uyuuCS94q7oTJ
UHKxPOM38ZtYiW5GYV0W9iG7/PF2kPP/eVkzGBvCWmCiKuykHL1L4K4ofM4nZVhqj2a2+lBtxLPg
9fbYracklt/SF9ld51lqyMwVF4luiEQg6ahhChbDiDDRIXQXsu7S3CwfIUl0hSH8rAlTcUAul8fd
pFeWpmMRY+zSHwB168E9plhLx5k6Yjn+FapmS9RT0M9Q6lPcYcaNe5nff+HJGaGompKDtTraam71
fVuifivt2vrh5xwSAmPMraQwZ+Z5ERBcE0mkh4FzDGpEdf5np8qNRQozr+GiVNingnAc0QhISaRd
UsnpsgTNn4mguSfhMJDQT6zfvQNVarkYVVKayW4hUTognQReP5B/tT21GEDvsVhtgjEFJZ8auPyG
kxzelK2jZ5cbdfQwH+7f7WrJ028ct58SfRPp2vRRno/Jhgi2OBxhHSEf5hD4DTCaXg2UfWn6lBLh
mI0ucDXFUt2KLhObECNKpeVwUDcfy6z1Cj7ZwRtIPbMdEwt91l8QDUxWnhVCMS95NixwGgufTLg8
rpM7p4m85fx6BFr/z6iCBounuD9ELcawbOxX7bo3mj2QNYWR3EW9QRfsj9EXzjElKsGQY0RBBefK
QEFFTL2ryOmOjy1ZPkIhJlot3cFln4OaMeaZi34T8RJAk9E+UEXrrO8rlw9+BfY4eq+8jJs0cOHo
Nu0lu2YXC+3Bzkz9cU3Ob3SM7eMzMVdA7UgyVll9vsW+NtUbmPiHDG4+VJeeFkoKc+MxXvWU5Nnt
Pkuf/svkWVPmJabpYsPejC+hIhZ7QuRXtkWW2ELJgOkwbsFIkaMpWRNKOx8ba7KipPO3+eaPA0VI
GZ2PiBCjrzmD4R+A7ewGL8nv2cU6NvEBClZoHZ0i2q1sIELtmi3HbT6/SRB+cqC1UPAxQlM1PJlq
ora0Mju1bTBhrczSOQXh89sZf/fytLkjtxVvOizvdjxwqLIAaBWruh5/ZDNUpCFdLLT5A80pAbX1
4wZHld0ZuWy2ZWT2Q4qRk9kdW+1eWco0VeBEhHx2DlsaVvi42jpM0F6x6zcCEmM60tPi3HcUyf+G
Z6b/12wUt3E1pCabzTttD4HlZTDo6ihJ72TjMfrDQ/FSVWjMZiCaugsXYbdsg9Y62cUyiIVVppwL
TWxeNzF3peba1fZpjeSnWc6/Ax6hOEr+MAlr2gUqkxdx4qhWvhfD7+v5g6jjz9BlhKCNlSsPWUHb
ekQkKb8Bg+TjKsHg/SRdMlUkA4vmpYkMgsHmZKZpdXMTXcOga4CulUDWv6rDusf6KSBd025nDp4T
hIRR/qkqEc9jnMvJ63Pj4ihYAZdWa+vvcyjHNJXy4fZZUeWs8dRLw3bc0Igq7Eblozsk/L+MKqT8
IGZgagb/mn5+9qfOku2E9zzqoi1A9/8XV21s/+4BGEm4hx+7yC2z7TEJ8w+cYm4DuAyLh50qe+Fa
8jF1s/iAXol/5jM4nystJKiiI648/GUQTuMFW4XdyVdLaQhg7y0Uiq6rqUK+U/+9aA6HIMMBihIb
k9oSoctajUImaciGEreNv7oA2EZyy9g666n0mTzeYZppmSfuWRTXiYOjFH0ZYQjcofy7HNCaGN89
TQlZNp30Tsb0RdoB5rqD/TnGQ9Ahh9sW7eDHeRoMPTP41TYnTs/MMGvnCIMIoEFMfzMsm3/HLfTX
SksKer7PpA3xn2bVHavkWOZt9KTmp8faZEeD0LoRmNzPOGdCQVXTKVVpEZXsvplaeL1/dIgXz0Zy
DaK7Ag49G18sF6fIFCoZ4wsC7R2h5V3O0sOy9a63jjRbUFykJKf8FDF3FC1nfncPRhpBx46ibVGl
zR8vuJCCYczwgUtHppYQ5B088jB6tzsqhkmGarlfFdOhOEpPUN5Qe7DQmfwQirFF2KD4k5d9urkY
ah4z03e5ozfPPddumyvjC0D2ws/eQzATL3fmesakjMJ5FJT9tP+5PlSx+PkWBdBI0U7VFRzYQwTr
VTl0OwONWwja7nJw7F9gJnxICxKAScF+5dl2oELygfCekSXkQSCzJAebwl0bgPJvKpGtIQNoqKU7
LJYl7nXG6JBMKz5XwBlFsRJDJWr5FWe+5cw9JsEV3/WD4zEq4qcabc7pmOt5ZxHwBYIKMrc6RTDm
CCGY2OlQ76ivGcGBqNS1Gn3Bo+eO4VNZHWJ4N8pduvx8/P3K1xpddEujJilaF0ka4Jk0mwKOQOVB
yoqP9a1jzDp/c0r//XXDC2kYj9GEGzbRdA7xFb9mU6rpIjQUF4pkLo0Z9uu32RcnzZkrGwhds5Sh
G5c61oMjFIgJD6flxrKYnM6HpBBh3zYkJALgvtz7kJEvkOD96WU21TPkM4kyYFSX6tt+a0g8LB7n
FTp+12fTtSN6+Wr7BtL5U9X71afZCryJAvorAkm3U184/dwDnsEWXkQHGym9E0qmhvzR2McEFfVK
xzvA7Hb7giwC2/5R9TgOpj/RC2NAeIpf4NnHCdknjCNJFKYrZ88cpidMKdDhr9eb/Z2UnKZX9nYF
NmmP8nljEftMlJqquqABt8lT4b6nih2NvJVftr9wg7jYphE0Vxp8W3kH3edEv7XQk4MemEJYl1Px
5y2BnuL23uEssVjY9ev6Zt8d/4knOpZLADohLKzQAJ+eAIayjRCVAt2Ixqcr9bGUPmrOYlGJ9QBX
0SIQRAxEAu0rROTXbvq9XEu8p1+a7P5XaxXkjFGCKjKvLG5nezwWp3kKRHJhNs6QncKlak2FbRaQ
UioYMmJtc8v42YUh6cZwoWZcESLoFl1zAtXVwqpV6sDUaUE8+Ws4+FnUKGrrzJ9YlfqqXWkhsnDl
mmpE0AcxI5xRt28IL+3/wcJrrvSAI5J0NduFWG8fGfXCGdmRcIBOrvRUb01I9Rj6KWwwp36gQ+1j
44+JgDsvq+iS19af4kt8tFcIVTmYpX+f8MbCrsgG9gWM1Bemp7o+Dsyrzfej7HMTo1kSROUCw8C9
Q9wozi06UzTswYQHhbstzHCLasuJ8dtjNx07gJAa6yxRInzYjoxcltNeOB4mGnia4I5FanZ/vpgp
D5Rv9fkX1+ijqmrqe6wCFSzhDrdkpmeC/SPUh/zVI+5+tShKPfYjGW+gSdy5RF2eDM/0vgJpapdC
EToVg3D2bPDA+5WikpJqZZpvG1Vde8mPelwXHB2Fquli/b/Cuooqaqu3bLR8h/JKYuxfPBbj8YKE
V0y1j+mPGvwIAxSd3AG72dmTBl/Ca5pNJWv7mUxh1C4Jie6EJroOdRpIBIB5Vi1o6odlxw1a/rTG
2YSnWLRgSfXP1FMP9WdoB1qk+Xu9NVPJDoE85uUHTjqVfZX+3xJcUbur1yeSRASzNpak/HSLaYin
bdSfgWzvC3MncdfFcIFX0+OOrX5LSawzxl6pXdsiDWfvkzlFPb51tg2RExrG4RraUcCjFgtRfrgv
bHtpIarAZ66a+vYSByRnQkaixzAhb+Aw96enklAi6zCUYH5G0XmdZKUEgM7fPpH9uivAeUAo4ElC
irT/vLxhPJ6aawwttZYd6XchlD8JNUpASk1jLBBD5WjIvBnXqDqvmT2O2hdkHnr70iCwi1LxFUDf
BP78AgXXtVNEnzZzIhrhRhfkO1YIWOEITLul8tQEKWHPMbC7ErzIji2jMAKw5FdYXhADtu0mm2Vg
We1SUkokIElycaSBeqxdmrpVtQOeDKLnGm3fPUO8yyLij5Xfk7HEB02CoDL4ALLrD8tVP/8BlJHN
02qpIm3/WCMawJv/NPhStrvTe7Q0bBZ4GUgINuML1vu61iIsYPA/nIHg8xIF4RXCmLRjI7Atr7GH
pjxY0f4jKBvQ7OYNQDy2umNEZ+LdGX6xitD+wFpXcA+sG3NjlxLdLUxCAjJckzuMNz6PG12tyFMZ
Or8iLWE5r4BI3a1zfYE0iHgMdNafTfxmgfU/3DwhGCapMWIntnjf/3zFzur0ROXuc+4h6JRf+A9j
IBJkG/tokMWesl4YRaswuBlqMEaLRvrc/3VbKPPibmMcPscVCkorghCsQ7v4NOqkHTP4GDwBBpAC
6an8AHY5OqVXARyHjGP50QrZkzDX80366M67ZXdPaKz5xkj00CYHkukfmFEXHfr8CgYi2HpjQHPi
JjKVkk6tGvqUAzCB68a1xFY/9HhcXqAMf/V9U1EQmrI9gZJdDVuKqZz9Xx28Nj09lReKtB94Gqfl
6a8hI0eFzMb68rxr/DWx+4ie5+OlegoPD8SHqf1o5JX19CshA64RbiMHQFEInFllcm1HLBM6WrFH
OMI1xfyX3Zx/jCJnNsYfKb//8TEWX69GZWpqR7z0PsVvhmLVBj8J2rGtX+xQrXBUIP0ifvP9A71i
K2eLqRCMyqwOW+3p5y0lyJn3ow2zXNeWDBOtZfLbmaF1MpKZiLR6JSPLJEOydFFuzAxeWO4/3nAM
ode4xMSANfhVo/yng7SCQrV44Kfz4dMUo9jhi3H2mOBKlkmxNMq5KJ+73vr7uuOe/9wEOUWwwY5n
efLwfuAZ0IY3AwnNAbS3VhgY/43rKY/c/G/ynWBb6mh5ZWrz1qVP0AS4AQe1kZN4PTWRHB4ARPfd
ce5/o5JzFb7fm4FLKsBHNO+uxvbhsCwwHuM1JPaLXqpuc6lI1Ik2a7IDAICqz3yaDASDomNbyqxm
b8R/K9rqvS3IyWhAEaGJL+2rpPmQb1yOYveTrDJkUVe8gsMXS54NX5MyHSDQKd4ViYMaTrFIum5l
uzlVVgVBEAcbZA/9VVV70Kn20KQioG6qzbOvyOqevi174l1bPpXTw6JlKxofdqQCHcgOpjw4iOrL
Fl00pImz7tbDacqi/h9nIEP7NMsSkNmAkkJ5RGEkXgCgk5HZYljAfkSOmFlKdTCmFwH7pCVGpjka
d6JNGcLakn+5syQgCjIgLc3IJuXKY8LDRNTGDbNiAykt+Mz+C+uq0/XdT63fh04W5kroWgyhDbov
iTdDP2VedA/qp2KCeU9M/03ZlaQGLDKL6bPErcsvTnXSXGHsZ9IpWY5NQI85czCiKbLW/4zsKA9k
Eqt3Lu/UoJyWzuSek6P0OhB9MwIGOQ6jERQ08Wirs27JTUMwFe9vSNpiFrgcCcn6s96cNsd1N3nB
8UgManWc5AM4Sr8m2IMcaQ4bwIdA1XQ+BRkL+NSkzG/RT6YzP1XX/xXmkVBQzFUsemxW1UuzkwrU
dxxvkitaYbPCw0X84aUXJBTGD8N+TmimBxAe6/dcZRLrMsmlDjZ+5+F6UYossKffYNllAxzYd189
gbFCPbEWqZfoPxqlrqtvDKfuKuXHSp/FOHW0knUFlY7SZg7CmVF+N1pcAdH/YYOhV8Bo93HPQovm
EjLcLwS/6hj+MYjxJ6UofucTm+yyCyClR69ear77XV96bMoEv+REBbRndjZXmMJyg7UiOFzdI7yO
cU2pkofsA9bj8zdvGiV6Zxn71RFxLUucbuewOkmd5y9yPLHl+7R6aEoKy5Gcs6i0Pb8F38mi0NIl
LZC7duorPxtogJ9UKaky1iFAnBczYdBxFrlowAe/OX7ZbJ5O2ysy7r/UNxmQCqt6e/oVfpWnvxj/
3dVzDbyf5l4pQ7IAalHEojSkPA63ubzR63Qoige6N5jwi+lXYKXvYIqJgDVaG55C7uQ0RPRjICiP
0iTvxnZqfYgJuXVbxUJF/z0UBMVc7dsLpivu9lsD+hrXGsSf9PuPs/kEQVvK/XDHQMGHM4/I6Qx+
Mb0vv0d9FiIRrNNRmEGbo/z0kNzCMGLPEyKMvPjKkLhWHCAzSie/rgl2dAgWJCczAH7A1HFn6lq3
g8B9IG7U5e4FGmWxF+PN3jmCkUlhPOuFoNmuNWE2nwWKei7HdfslDCHWKJuh1w8apy6Ne/afAkvt
zincwKFWU7YlURKe8u46DG+NlPDck3yFy6IZqD3lNfvBfH1DqXr0xFKtn+hxu2NT3ZjDOLxCsZX0
cSg+kyg+9DQScmV5m/vXSp+q5xYXMCD0KXSYPMaeQGq+M4bqPGm0Mjzt/98GDZEncVO5kDYJnyfp
2X3IpXsej5rzU4sZ15dPcCCa3cI4OL+I16XrK3Ai8aWAD75Cz+H0XnC5sPyzBg3QfYAhennhTOml
zmmhLtBHHm17ssPzbH97MHSxkCxNMUA9NoovWDjn3km4E1T62uppbN6zG5p0z2BHB9T744Zu5RJf
QJ8FWmqo3kILmEda+MhEjTpt/XVaQ7Tv0QjPUHNWXWGNV7bpKbiRN0TUNNPdP7v34+jwcUaYPlfR
oeQsaEGCWM4XF0SrSZqVc8s/GME3fLFCs8aCiBWsoQVhZMRmhQTt6T2EZqltfcrELB9T4HEPIfev
VAquWD2Y4u6aYh/vCH5xlN1lSW+MAPXxavfH7bq/V+YXVYlH+pAOsuLE/7Dsjmzg3DQRDKaac70q
nK4umBaUQbIJGSvXN3k7GcxAvy1JaaFbMFO9eJfzwsOqIVkdf8EWdo99YMmeL5jMinvQt3TK1ArA
2yMkTnFhnUh1pO6DOqbhO6fLmpkYOe/lAnL9fdXNpkWi9GD5+T+TwGFxQVPlPNBjDgEh3H8eZr5+
eD2SGI4xvBjogZQOQCqB+5yRkO4ifTm6T9o1iN6xeK61XYDO/Ls3rF6vtCOfuqL0H1HTNM6zUlTi
4GEy2C0A2SHlhtAKbE2poeaQv97oEvp52ubB9zmLMJ/0LoR/zu7Ol2htMnHnCa3h9iheDY3AIpVe
VIWYVEHls7fJvRIQGBTs1zy9PKPbTI4aHBMYZ6HxtYaiMRuHDPog+o9nzEa9pWlgTyZnSfgfj08I
s6a4sugPY8d25dkYRf21HPi63RreQg0/+67b12m+Aa1UxkWltQ94RByw65MLWe76cQ3ism9hm5OD
API5EWijWsa4lgH8oqP6zxQEnDSgzaRkxCvtPzboXHWBPHcZQcDuCzdSDK8a1AMNk3eQV0gZkRSF
MrAkYWh6m0R78uv4yqQri8a7geUjarGMa1V+7QjyPI3vTz3CNdx73rZqVscS6EIOWQWuK4YosFvg
nQVT866al0B2xshNULDvX43TzSCkG8tL8F29qA41S12prlb1iXMI0jY2SLMDLBXB88CAEah8mMzf
H4Q2kBBgcHDKQAEJnvuPgYRU/B1xjXrB2Z75V1d3WVGACJoCKI4iftayTUpfTtprW/Olw0TQLnNc
2bAvJL4mHUa+QwGr2iq3aJT5x4gkgSYO1ZqoUOeGGI0+u0Dp1SaOKsVav5LFjDyGCiZzNp7dqyt3
gY45SmfHxtXwpSUNPsJr1L9vA21QHkc1snj1v6wNwSNIr4M1PmuXyWh/GNTCcoJClHtXFEmg7S/y
hQNjJ/6IMJSrI/MpOlCGgxJJmk48hUk/+dQvqoCT0KsQMlzlBqQ8LS9FmHPfN9qGa8ywJQeR9+1i
KwPNNWPemvd/kGpyy2xZ8B1jhGRL5TCxhFaIZrm6WXv6ek0RJnBTBjrw4ZfDqY4c6ZHK1MiDOTiX
4UK/o6Fi58/74Emmk2A4WCwlaqbV6pICsTIHbcNqmS7Tzv3dSSjjaM8oCTtFFFeWtsBiasKtlfAR
XpdHtGpD2KMFo+6p9Y466QECPLwi3URE2Nf0ezVJVpfjyZxdoVLLU8Y54H6An64j7sFEs5iHdZcj
p74CKaHUOEeHbXjbMQrdEgNLq8/DktINomU/fvxKcwc47KTjBLPcsdQea8Zh0Q47JRP/Y2gsocWp
OPRV8t7B1WHvLq9VhzLDOBAdW18hJrlxmNhx1VhLuQ/Dub0IX8Ils1JQ8LYfCtRx0qduCpRBLmKt
iA1/sSe2Yf3AYeR6uaAc1Q3Aq/8bGH/m0x/3YBDED1u7mZRS1ZSXOGIsgBnjeZMkYWmXNXMZMs2G
neN99EM0aILkS9O95rBqTnRDduvcYVoL91OjYdQqv7NK8/UGl4q8NURSM8nVdGp2t99RrukUnY5V
MNPBlaPiRJbK3F3s2+K+UlYge8VJFaFCRqe7Lk/+QKGlgIqeN4wEmaECOgiJNxX6ZsE3ikCrDFI+
cVgCrt3PjCUdZ8mz9yST3m1VO6usCxJX0vYmla3TNhWJFhmN/LojbXqMrI1IVhAmdIONil9ytv71
4dzHZtf1JVO8fvTrMN2ZlD9Pa7eRvfZEG6656snA46DaRnlcm41qq2H62vnz5KwkhKV72XKnlM56
RZmM/5rbQpba+P9pCAZQxv9sm1psb37nfQCNObk/8clzt3uRQGjxDuf4ay06Mnijn8FgBasXH+2O
RVhD2S1Ra8zjQ6LTcIAcgu3SMTURu4k0XqfJgwZdNaC8Vdb2mFZboKkO89lHFppqb0c3uurmLO6B
p2RNXu9oiJ2urdEmD+zwxLzVMUJepIoo8qtXfr7awCh9vkukuFo+0I4YjKBHO6S4qJkrhoB0ibbS
CyPa2sF6Z71RT7H9mT/Ah5DSTNceX/7LUHkfEb/UYSQsnyB+75TEls3bLTY82bSP8Th0TTWYnZYQ
/O9jILesuBgpMJR/d1wMksJoss2wLBF6jDuCdauFmNVLRjDdwQ8WQJMBjbIEoruq0YFUurqA2k+A
DQ65cTwDlvGaPdf1HjGUEKl7pWgJVpQlzdxob37ApbYJcALmZ6oEUIVKDw8RPGGM5UDvi81T7gFi
0AsW543DWWeuAIE9tf0MKIg98FN2NJMe3jCoMF42v/vQVeHWUopOX//YbDgLMQVfGXUEEKik9cOc
pd584LzBJVJYQTy8J97o7kIXqh+vH0GJmLZOrdgxYWaKe6xqlZfvpbCa7bLRcvg2CA7dkwmweA/H
UXGNxKaEPoxIx5XpIkxd/7oLyrqOlaOBQeU8QMV2IZc3NXdaFU/3NB+MRtmSgvCWD34rM68KD4nr
G7r6nNXsPaRUQWexFDnZ61JkQa07CxYZf4dT4jVBoBf9AEqjeBrc+QlgNHn5J++SnPuXq0qgFr0C
MW7YldaLAitinUmx1UOE3oYE6UXXhyTLZIgLNuyR7KqYq9clQMxsNyPlHuMGR+QV/jOOfnAanczp
AQxIYhjhDPSrL1Ym0+Yu8kyx+P0Kvv+42PdLiNOVGyCvUnygtNnSrjpECy/hDZ/CpOwSoNj9KjlA
6dO+nqUOYYNAnJYdHMSPzxFq6hx7n3yP5yrBPBCJAJQu5RP6dLLIgiWsL5Xw9wGoCeMSCN9Jeiwg
cojlJBPdxWKX3OGG2QpIECUTLumYgK9JqZS5mHaBeeINub+lW+64tFjtPZe6s+sTCAZJ5Xiy7wza
L5zX7mnlpwDdQdT5J0vm1oknhPjxNSZbzuyVPJQGx5Jh0zm9WoyN4KRKAke2mtFfBgu8sn+uWYJ6
2iL7IcMuLMnLQM4f6tvsBnK2ZvGBMfGDouWf16ZRUcggiE6lduInkTinQRvQKqVjO/rQql5P3uwd
oeBS4+JyOd3jAeANkMnl/AwVCOEHB4RTUF4GO5VT2A5G1qum5MmExgjOeN3d85OJegE0Ly47V+D7
j+CIUPHyZMxocEtHLn/GnI5IU9gYTX5B7a/rAMfMW77REkePNrAUFgfaOoVmdxVR66GIiLclRPqO
VOTV3gXdxaaJfLEuNEmsARJiiRxd2UMYX37z2W+AFxW9DEkPDZHSOw2NnAKBELJ7/49ObgaLIJTn
WkPJVtHR3NLJVD9pl/RwgXP/ZxFXTEuc0ZZGGNM1tWIcFb+T18bVmYF34wKEAWwbregt9gEPiXh9
CxCruVR6Uvuyd1YK+E9ECFuBFnJ85BCuf4Iws8Nx7fQyXSs8u8gonIEugmtm7dVuqOXOWWq8GZsR
fnc66uJVDvDTkVEsybCGSFLGxdaG0i9zWE80fbULyF6T9U+iRgAgGLw6Tv7Hj6ZK7ki6N8GgMEWt
kZUN+csQhT+ml2aBaIe24RoCSg7HDI5xy3os3iI6OZIJ87j+8AgzZ5DhxMyV69u/E5NnMtD7PpNx
94zcYk6yxpBNPgjOY/qwqI4xsCZBY4hEFmMtDjt7ezcnSGRZTrc/5UrkjZ5e6DNHN/HCifmawGBB
ibG1lJt/aRtkg11IDlyLlwQE1Eghp3wgVz4+kTR0VQBs5IRAIzP+rYNPjHK2TI6nHXMw7aEQrm8O
W32508AHAqprfmfSl3BMwJThgv9w2WXGr87RqkxPsR7OX6e+OlLXPrX95rIk5hguQOwc/GJGlDbN
1QxOTlkRSwMoIpmUurpQky9t6iIWvDEj71UhsHGXSaJcoAtyzquW1C1TItYL5A8jafert+FFhOm5
WuvVEP7kjbPDNEGcTQpqbHnAhJwXnxkuvck+u/Env9Z6igXSJIawFbXsuS+OuYBUGk9a4o+TMZho
tCHu6n4XevHtYbcdFCW75TTSaqyp+CwTZcRZshhU14ywfcpH/UL8fe5NT6xL6Lr0vR2DrJiKgLJV
gMyliPKfSTHhoDBUqNt04AN50jAyzuW4UNIn0xdQSZVGIewH0NQTucg4oaceOe3Kxgjf0YuqtQtP
9qupMXnhBTQPdeUbopWdPyB+WOGAbPiMAk/XzSbgpz6P3MESgRNtjL8hXmUBRQBsIZB8bmhRMQZ3
E0f7yGtMqHsYaqQZXCLe5GsA1l3/NdakiF00FOwqeVt6R6lvrBGIqKbElZTaFgXkqlat1OyJCKYP
23dDpq0fshDazVqcRoTJn1T9FuLeHEerXEE+pSeTVXzVNcow75Q0YP+5pIPeLFOxNzQiEJBlwXTo
t6KwQbGpOwM8ws94Zpmg9Gcx8WPO8oYXE6W9pLYLHtiMEPgX0vJr/3o+gGxIuX3I7o81kRVhXkCu
Mj/DuyxW+PjX68G2XBHfWzX1YWqxV3zCmWVdHoAjWq+8mHHX1FZ5bWB+VKM5xcUFH5uvk8+zkApg
Rn+wn5qOIbFBDHLPo0ZnAvyw4NuNrSqfNDZBRar6kbwiuNZ9CHCEHNUc60QNa1x1+Y1nMDMhg2gN
gBEbUURGFEuUrlzhp0fXekDzUzLowYFjl2eUQwrjvnpbkzGTuYG6ajCY1Ei8VHjaaV9SSknOOIkn
+0pjCU6xZ8ZSW/jM46qTus2GidFS0YMv9FH0BUm3O/MR/XDN5q6JdFuWM74NOXyk3DGxFHbqe6yh
peJECOhAWALUhv4PSpPiVjzzJu0d1py27eriRHxWrFPeG33de5/wXbjijL5xUfBUohXdctCi14QG
Q5MF24U9NiKjGPvks74/OabS4f97+IvuDTV0NKWtp8diOQF/DlN9NsExrPy0JVRN+KsyfkglE31O
0LIglxRdBK493q6CrlGSE4FpwzjuTSDqzPDdV2zaE8kFvAgVWDxACesjqdjcbtwtxmKoMzJQQbul
1KFXz8lhgR0TIHx5bNxvSQwwxfDYHkitVtSpU1nCILA64BryG5hN1M92GAthUIAHlaiZ/zQEEzAc
PvN2/vlU0Gmh1YjMKjfjXeIMRzrvB3RCErhEdezYBHdSW5zV4lOz8pJqoKrVepB0+CCZgSlQLDjr
fkceYV4+7A/ImlVsujV/v8Jhkrh+yvhISJcxtsvm/F4M2tM7bFNgDf3uLw0q8ZKAsIerLJUj9r1c
tniGWHa0ReHzpk7sboYw8vI2UxX2y3vBO7Y55om5IB8nG/IRCxRlbkTnVNmk1UWGOUP4osC+MVV5
sr4Vxbjfy7mIQMXt1JELsedjY9dh+LaOrd+odBMRc7JTm3RXzlNAvockDtHQSHgfypiU+zZ65twj
SZGJ4F2VTbkPIknsAUslrmobIyp5WKcBK4S4GYVqa0mOAjE4vaWdVIWb9AbmyWD1R5bcymtKy3Ob
ZGvSH/YS639STYa84IfAs9+8TS2qqs0f4Pm9BOIq8aFIQOMZZlslzMtMYBtjdRUgXD4pzIltatjM
DnuJl2RuGTeeCx2EsUMgjz5m86I2Vax4YL3HU1aoXi9NjFgjssELVSVNPQD5/+nCn+QM+Foqa3GB
jXKA2yepDEnLb4NUBvJiVKu1JksQ8domLC7NOz/ThcYpiRz/iDDvOeoJfwAPMgJDCcOsw9A4giBU
iieltYu6mmvVVdssSAOY6Xn0e4fV9DqQJYAND4KFtV1YxXRuy7s57Vgu8xK8HjI65GbQC1IPzyLG
0SmXh0e5r31x2UNgxXsD3W6L14vrlZCHwaGod/fApBSxXoLN5SK28bZKIDdva8VR1+1X0PVHHDSe
DupBlAObAe8bJjxKSuqXYAxh1AOfOK3pISP2JSifGJlwxQ0SNtZEHt3CQMN1yrDWr5BfPTHa0jdD
tl/qgZH+anshp72pqYdLteB6KbbyISo0EfxyUrzbEUaFcd3LEZd+9g0Wy5Zme9U9IXBnRoRhH3oJ
FQwVbUZhUXCWkW8Xb8F/SDK0RDueFBGKGSuLTnvCHr4kyrOujiF8GlXuObwTvwSiX1cZ7uEp9DGG
VKD8b+CtlZIYNf3HFrciaoNyCEYnL5MEJfukiEDlK3wYuSmVmqRtaJwSm1g1EUIrHQ436mUTWsUU
00U0hK+Yt8dDZ6BfmEgoN1hPCjnfgo4W2D3urY+cuhYFlD1zOks8Ko7/HBPyj6b11JHIzWOVxNmV
azfNV9j82YSI8WHG9ZONPok9fwjHoaexpc6bXB4Hpl89vDoWlDl7WzpPQIImh4bxAxT4cryRbEGZ
fF1TD2C7+hs29U72UrJkfoBGM4M03imI3nN8GxEb7hDrlQkAPVTFOeiWTe2U5l9irPmGD0NUeNoK
0dedHsl/i1vVjeffIbVWVpdmkPWVGetDu63FatnGPljxNJz7pUnFQuUqSdqSFe6WUEQwA7UACDdk
XJRtXmJVuJjyprPmxpWsoLOEFbCjO2oqluzfNPdUtSPnLo85DN1po9+BbAzX83TGM6C4yiTPvoxI
GwW9hBaQlx3u23ahf12B/YboL+fG/h0tqSQQ5Dx71QAPEipLQWKmu7heyujMJJKD34FMAe/LJrJ2
6F136i/ZqCmO8Mc64Iq7kq6sBVom6DOY29SLd2NVACJRcmSZyZYlwy/yazH03sTkE/LG0tFRYAh7
IN5m0zfUfvvoEPXjDIaLOTGMavUdEWQBFJVyCeK7UiMId5pRhxApusO5Ap4aLMpfCbuDDWxU/iye
kTOv46/wESUtA7kWwSmIofj7rsPEhuPOsQZlWGPD0y1H/YUj/OJ8qQEzs/DVw7Ij0meP6FroIrjw
KiX03Mv1gmM005dCisIFJLY/frdJU2JF7ZhCNSEkfCXgg/gAnY45jlS02MVt3iSBbryv2lBOxXyW
M9W8xJ2vxRGgZoRbnXztPUBtYdt5/1xjTXllm/2a8XQqYa6ChAoYewPvEyEpCSXjZbjV53aHW4QD
ca0i3TkKSxIBO31zAHU94xppssHbOWVgk55pUZiQP7XN2uWYA9pnABptlMblUifjDe+ykguHYRlI
2U/Ofq5wFpHAYGBnawoEuOWVdCCwR30652PpbW73QVRVWAW7+SgLBwcjNH9EmUTHTr6cg9K9SP3x
pzIHkDR6hIkf+G0MwTlPXEZYGGhLXobcP+cyXpOXU0MWk0C5LGTwDNrqCtOJ2ZsRtmSIxnqhZjzD
8fRdWXrhdx77ThBoRqlpgAoe3JK715W+lai3Ty8e0JrwobsWV72PFkqeUxz7rjBB6hDkCbNQMbar
GYwY8Zr2A5+tP4E3qg3X8Oc+zReiEx1/FQN5+JDR6acd+iXdW8DY3DlBvUWMzrb7oY0nd1Uu97lv
7AGLAmNPStdUTa8KQlD7QwvgMtMqpYOBjLd8SqkN26svonp9T7S2VzBpplSXaIjUDgQTtFmJxUVG
FJElOGBtfyJvN/fwKp1WDhQ537E2+pYPGf6sTdalUNOZriYk4bNcBYprmYr/as22TF4scdCCLL2t
aT7QMxychr2zTezE21OkclJ+90sWahd6vxrjD9/dkp+Rle4YkAf2nuppZNCV5hwNQHSA8F3K/tG9
8T8DC2fPc5d4mDRu2w2em5qeXbuJIK9ddkWO5v17DYgYvpbK1nFsdX8fQ7PPhRQMOahnMDVs0DZk
Cj7htPkv2xzxCJiG6c9xJ9Qdf/WoUbixU3YMdQuGD6tJIUPg7EjnQ8kiytrKRp2IJ8wTJ9izJu3O
BWSGbfNeL7edc7Z4aHCKFYCVxUQVvu24nKWnKYUbhx/4iixib5uSAy6WtNHdW3aVbNAWEhZAWEzk
TtWzyrjfeHb782awN/seYFyCsz3qfh0iZmrTqU+nKWUn4h58sdVKCNl/RHR5Nm+Q/zyVjWLEVvnj
HyJevNRw4ZSLr2LqcLCGaLiAmA7BXx6aDOWZOyoPHQRq9KvnIW4E5yAVs+RgkYdK58DF1SYTAZNP
sCyvSS1XVeMfJvHekuZZlMZdn+aP+REyUryeXcWfCVI0iKBu+CQptJQqU0e7PcY7U0qHWqXzLFl0
x+61x3JqNJw0IvE1b/erZ29+7XtmTDX4uXrsvCQE2fRQTJ/1UUYrXiV70Vzw0By+dhGALI1rHEiP
3hjjZRu0kXqlmh2jJjYZXFEbjX9owrMmKqASMl6Hhx4dASArRn+R2bPBc11Uk7AU9fNRrvblJDrg
l6m7Qi3+nQT43r9990c2PaXGB0gqJ9c/KOWquWmnbBDUDFtrDTkcyz18l1+nioKAGl+ryiNMsWSW
9a2XFb70tOeOXQ4swTip+txJVl90E8n9axRW4vm0MBD3BzeSEOP8wP67c/3L51IKB4u/RKuxg0Vd
zb1aDb0zED76nK/XOgMR4uik+cf3XBujKpSSDm4pJy5P0nIItACpre48rhzj+pM8NJ14q+BCcOsn
8Ijyfx/Lnk+DjV2CSJ908qfTzUcAhPsRiNLc3EMmIdwBCz0TbI2FecpHqjzi/kmsM8KO6cjBsgM4
P6GyDinj+q0aBDwuJeXSKaY90XPOq3jKHd6vCG1i0O4gwpFDXISdAYDq9+WbcMLE+BidnJ0gi8mZ
9ak/BveJxxOkRaC0BfY1j3EOlL4kLnNQ8yux4GFJzjmvvy3g+O8n3kaj4ldALyD/Gmnkhz+fzN5n
6GQJywWDFhx/TFPATIqqx5ugblokA5c7Fowx1VFXzHM46iJBN59DhrLd42szDdSiNB9tcPczrFx8
wDqvHvak9C2u3H/maY1li1NMCYT16rfPLLZzqNogRG5o9Wr/Jn3aFWb6HpubdkTwTsLQx44oecxy
PmUkFpD+dttnjFY0Y1Gqyxkih+uGKrF6vSnbFfOmu7Bc7kgOyKEyo9yx6PihnVGs+/GpcKGLjbWk
CazYMDcxHQtSBV1kXUjYaq4Jb2Nertg7YgFjEBavoIHM/J6FAH+u+iV2chK4QMttk8jkGJUVze5U
+tIjfJy3zBGwRMVA/dr1l+cHuYD84B1YMo/dHqs6FHcyNeQyCwuUcRWnQ60Zc/yGpwiQYfoxRPOP
1nhgCM0LftIjPIg5gxyalh6qO6m1okXQhfDl3JO73INRRUaAK1lm44N2hs6oB4qf+4h48zt3vA7x
2hvH+eOB5Nhddjgf8Dw80d1Hgu3kEWghYV6HGnCxtwGUCbCFSltUNONyCvVeKXKNw1eziVgECZMy
ZBgFeJnoIYveBm/XsUKEcRmlvkQ1h3Y0QfyyXA+ImrvslqmFWixQlU6XWfSzo99jdz6/h6V9GmPS
ZA+PmNXVEzmBQT+NKRLTlW3vpOjHiO4VmAG61K138N/+HJlq6+YxoHQfHlLXgXX18WxEf9RLnQSx
kADoexIhG0TZEUcnm+kRzEFuQhYa2okA88CG1EJaTlQA9mJ9AI0WQuD6WEWaJ3Qwps+ycLnr57p/
QpZNYSQh3wMB+CslUHcXaEsHcFXQjIV5DerGfH8C+Mj3oqoxLLRsbM8+jMMkk42iJK9d17zaq2x9
TFmvBkzrAZ4Y4zI03hfEv9i2BOXrD/vuf/kDZmt4YdiUU6nIL37cBHAWHy2nmSdHsGQsQ5vgkuu+
U+gr2mBaevHGJwEbziNs08q3Z0U52RPtSAP1lS/v++j3hHZ91rOnwrmB8CUImVBShRd7S8fJnv4S
b8SyvMerKdTVAmje7JwIc672aMjFkcDNS4XPdvEV0DJLGYuJZieCjUV0ER3vc3cIXHoUucP9Ls2K
5GLP+KFoNIp3+RQsAIJcID+Z/cmoJ10krkGqJSCKgb4Px2snG2UL9ne/61hRTvk0Lw7rr5qTREBe
BlvhQCTq3A1QhIMoKj+3xzxxDofURGfrczkNj7RDrdHs1T5SCVUuj6Yk1dHY4IMh3A4+HdWfhw7c
2pi4mAFYdLI/WWKuTeTfwImoKkbrg9L8sM2p22gCX5uSR+e/t52uuzFHqi6EUCY8pZXMNG9l/Mvk
FmsaJBQ463UoDpQaGtt/EBIvsBtk9pTeLxsAPvKkshQkkKVO2CcxG/4Y7UHdCFqWb6Bl8/Qmppq+
ec4QkLEGR3Kyr1NG9RWr1Y3B3uYG5aO99+8svC/DEFbmyJL2HDBRAjD3YPRrt2DjWLCsl1U05jst
o6oGVmuNdAafnnemqXf+9mPqlueExagtnsmrxIziHEpQSreQlPs/8LE1k3AQx5o2IBbKU2O5zhEF
Lnr7gjdej9sFGQbDyOwM6al2LQkWQHjKtEiPnsoPqDb5eT+rxkpXfD2RF22mB+SANu2D0FVkPyll
QwvmfqgU02MDztFtYnIq0TIwn/ItpCk8xPPj20DcV06rXFRmNXmI3V+K//2AiguD7By6cK9Xs8+g
xHnGcLx5TaZjbfd/9pk/yD+GaSXKAHFliVcUHWb5BU2qEv5H/yc6GOeV9yULD1bdYjvRHFeBlzha
0PUOwJgDpd+xDwIDyn4Vhr99E059/E5HrTCyV1CcsEiJsvRV/2RQqebtmjeBrxE3brUZFPM4j84L
I8Lag3UqlJXVIMHrDqonFD2/kmMI2nJe+xXhwoeKs5plMkrOzhSyyHy9U88HwWSpAlUnOs/T9pEO
ZY0NxciCNR5QmHZnUL6HtJOt/NB/uVTMgRsYaksXOgsSbl0e9QgKdR9bTIfQMEl7dl9p76yPhj/o
H/Qqx747VR5ySp1JBPfu5RGn0edA6ABFwaARbQ/9W2UWF6N+9EQjSykj0kVS+rWnnmrs0VdwH7CW
EmVd7ov56uRVSKtIQYfvFe8ONGYnpUdL5ZKx7Ofm78Q+Xbw9LNCPnBdZRkP+weHPLIdtdMS5NoPi
q2dS+3FkSQbV+RkJCU3mUxtmpY8sLA5Yf8MPvXM89ZswRtzX5xiSURsgiMNMkhR/qQZi4DdtxZMp
xWgxv6dhWtsbi6JNGdMzxgQCYYNMm1bbH9qVcoMLv5j3IGc9bJWGWHisX5TFv2UNs3klfSPueY6F
/3cPMt1vW+rCeiOJtwtY3ksSYgGqTWSnxx+krNYpUH7mCF00Ta6h0T8cBqhPkdBCNFoP4AKih47d
PiZWDmrUlexQ2oYUudURU54Wn86GF0uWlIclFTyoeGgfhYqe5jCDWYXgh7CDZ6wK7i4yDhQxpt7X
2vd+19cdKAxwanE/fabrGnDdFrMdlNd1PUSCMQNEXK3Ji88cGZp6Us/atgZN50ut3SwUzjSLhSTS
aoEr4lgNH/B+W+IvlWrT26dYVSQqYILBbaLp3JVcghzAMEWwEfMLrPVIw01XlFCCMwonn+/D61jt
CQDYsULHznds4fWZ/3XpwLFgcf2XXVk85IXTGo3IPHj0KLUyLtgELwABCR1X7mUFUFtFuuvglmUu
9tGzSXCojhZ6rbAGkf7G3dWb+MmR3Oa2BAvSFjRVfF8NK9tI0GDivTKZdcIExOLENCy2awZVtI3I
6fhm03oKgMhwbHkCoOYsOIt0stX1zVK3of8z5NdyFdvSEEFTWyl2abIFMNWWEeTGK6xEZHakgH5X
clTmEs7Ni3NSP7/KXgEZeZg80mvOmBOprYPOhSi2y2uGCzOZYJP8c0yNsogBI29m8YiS14ukvUnY
pbchzrZi2A5xEA9TnOLeWJmaBvB+6eVf0IC7Fi60ncf3IY3cUQxY6Nnnbb3iqRxnoZmenrDLpBbW
zeR+j2Qe1wJSmIAQkeeLDIT/nJ9zKeF2RPWCc8G7IzxSBdWsYDzIimfhr1/73gX8yG635LREsjKi
CoK1wAX5r7SxLOYInt/JljXIPF+nlc3f+5cG6PQnz8HEMnR/OVf8jsYKTEv19HL8b3Lzj/pmFLC+
lKJWD2Ui/bmheCDCIuwofpW5TCRDJ8oCzLRruW6rjuz7ATKOvzAOca3u4N5csDH7a3r49HBnjSwW
k6f7XDm3XoaXJaqSDnJXesBTcoO4/aG/Z7Z9W/6l6m1WEXVEsbPCqwxcYbAgQEMeZ5C/NzVT1Lrx
1/Vn/AhexARYP0bqvDrAotXUuqGPMocqDosxtaYr/G6sB9H3A7bf145bRkl6NNEVuJo65SU632jS
dTcYkpYZHug/ts7/rrW0xuM8Jlh+cHbDzWHM1RN2Adb8IEi5ftzjYpKwynreh2bwA4tC6LvBwnaf
Lun2YHqBpM/S7xopQfpDfwLt2Pcf4bywXi3I4n1g+dFByEAgAbyBLqpSPcFPkLpwud/P7waaxPDT
DYc8xhXeFGLFEpF59M2SGqw3VsyOZDi6W7RrmT/42jzDQ4kbsFAGR5BJKRfJNm3d06Epxfr8XAq+
tM1uApBTRqljCs1ULYD5k9gVzOOmjPOu0khxjhUBIS6G1qYnrW4UscYFy6bahwCI9kcBIuW6Clz2
nsSsW3gto1joWbcZZhZ3qh+k1QBpya1Tx/its3BS9SvkwjY7fcGL3XVkEWbNh2qXSb4BwmNHCi33
Fxwj1+U/Yg1FrwFndaSR8suGxQ89eyGWOjh55YbJD0Zege7BpGR7nnerY0naGazgK4EgSSa3NpSv
tGJIBEnUOaPHdUSEdQ7kELfqggd5trBGb3zGG5CYYrc5aV7UUYjq8/0eqJUOYxso5s+oZv4AgJPn
Kk4fjtmjcy2StvJqo8xa9O+zbsYWiUeBazgvvZp/C9nSFXfO7gHvzU2N5qGmgZJd5stcDZ4cVuCb
S+Fnmz9CDFNi5ahZg52MjFUTFSrzAVIUEHIRNFsfHlR+q8vkD8DF+Zs8nlvh9CfFolG+6QalcWRD
jLPGekfwSiXYwvuJ+XIt15gkR4RbCnPLy/UN1mvdHhEhBY2LIySG6G3LPLIBYIzt2BcgDLRFak7t
PL43ffAT5Msjggtr/KFChLv9Yu8Ht+oB+UXxe3dbVO+xlzaF3A2A0lYcxaqxaC/65+wV4PFtnJqy
CfB6OQsyVdPOXrw4eGglzFCMPnB6ZPlvhRmgxUZs5D/OpKd4m6VR+jdpb4xsGCaxMTnlk7N9NeBE
i91m6CLww98UG/SuYrnPJOwOHtele91lu1g3MfuVE9Zjx2/iSYPzAEZohXmnEuxsNPsgX50thVOj
5MnHGb4royuRkuRDlVWoldxreI2LpTioGt6+rRN4NIaX9oOCfrFVpErodxqRl9GR9D6TVvgHMMGf
EBj157hCustuN5NIWRKp74NubQYjo6mXZUkEOJZrxCUUAMW09GxieFZl6NRCCJbjGJGatn728r8z
GDPTOYwZb/br71yJx4AOYzyqYB1oNb6ZxVcqv5QHOPpiqxaUqOUoSDDPy9kBCZ8ufgIYgNmex0yg
0SIvuB3lWy5DtRad+jzrn7clrjPXBqWcV5psx67SZgDggoXhML5khW823a0SO5sY9kYnU+mAbKco
fIjrf5NgnFlMtJkOxp9OrfVsHCLWEJRuHgvtp8lO21w0VSAAE9O5IZqL5RQYvdHS/B6deYd7f2fa
MGwuGTJhmqE7/iW1iLMe/HTSKtab0OYNSsNZt2y2vU4JiBcsDE5r+RQnc+7Cu/ya0W2K/C7WKs7u
dPO6aYhNJ6JmC0Obm4Ev+j3oFXKlwzkwryhB4zOogCnneDSi/6rdy7zFiS/uCHwGOImLboIk7ImS
gStyB/4AT+6njg1GkQhyTEebjNi5KLa5Qkl9rY4FJEubIri3kChYiGeS6GfBjhBjWFba3+U0Z01j
Ymp5OZm2X6dzI0THcEmUhvYRNFywpQrX1JIfmQbQAdVPq7AutamzzSm/2AYL9uiUIxwIXsIf/OGI
iQmW3i3VB7GiBg8H2YhFVAlHZB9mvqyfvPCi9ujH/Xh3TGznTKeXrIKT0GG7Dta+zDAr5tcv1Gdn
R8Sc/xs+anpPYnqGMp6HYcB1JhS2g/e1Zbr99tbGxvyaIXsSyg7YVuqeY8+f2SrBJ5mBvF7Jotcb
M40g8KA1EiF27jLcRKMUKLGUqs60YCVqNnRdXHYz1Y67l9wZcqoJs0rHmXV+IGklSrwjneiKND9X
nHzxqGiQ782Sp96a4rROJSWdfDMF21Q71dItOKU6gY553AIRNvA8BfrYRwfnwq7UHi1aJaOPoBzT
YE5XhAHpIJHaXDdSRwoDjMTcQIfNWjnStXTlmq8ow0Lmb5ohluWCf6j6DILxDepdb9UabehN4PGu
z2LglDxvTG8SPrVM3fdu6Sdkxj8OXQ2B4eqjHKQyhKzt4czSVcXN036+kDK4qf89TJo5iKqtFIE/
n9KK8Guml5A/2jr/GkyFQe0X6+emdb0ZVgr4WTegAaFVyRAn5/iLtRGw7C5vrvl2CP0f76kk5+ZR
1+u7BL87yEKXbHo17clmSputbgMRP35w0E5EtM2mFuCrLhPelK6SMQZIZOOAtNHmcynnZQMCdTA0
vHlrbGq6iCRJNDt586gF8ZQ1NT1U+Tfb1cmKmgTPqU+ueZqcBUoqg8MC6VA3QW3u0e7WEvrPYmJZ
VxJME/Lt0zR7IIrfk9mDauz8ZW5C9OseiadAbNC+JW9pCZVDngRm+iTpl1oEeWtTP/79/Mo98JVp
Ck9fn16NMuVuzyDqL2B2xbPwXqXPfwRNrCPZJsvU92HB3yZRmlbhkSO8LbkWlrwr5E4N7dvleH6j
cH9hl01uW/Uru8S2dRilu6dsmg4gqC5EZfUQjf2HNyp74UFVBnDUIErK4CJ9mvPRnPwUc1CkogPB
3AwHsQfAvoDdqsA2dixV5OFGAttoNnYTAigSFmDs436kk0KBlnIYIoJGaIUIk4/02vF1HzeGiZxf
UFnqysk1jG8BTHeM4ySUeIR7KPdU/ge3W5IdzlwpGFaRGBCeDmP2JihKkHyIqaHW8gdGT7rvviVm
i8Pm9Q1maXMHLBFwtt/ptwaFwO870WxafpnHC8Z59evkWYX7DP7TBlnJRP2tcln/NNmP8EzANgXL
ZrcJLSzArhrpcBN8o0tCqRjWZseD8mKiHW2PGzgW6/mFXjNhLmOQ24kd+Pip5bl0t2gGaypc0IxU
Q4ML8jCVh3Pe4WfY9EPZHVd4pdRb73laJEX5K8uehno9HCZjyUailcrIy+t6i7VTGXO9nznmz5eP
myv3I8hXjHn6ZPmU7n6j7HxC31iLG+DAZXkXpNfB6PTMEL5vauqeL6C5f3tuUfPmncO4lN5nkqvn
VbmnuLEcg/XFF5bt6UjjyejHpO9bNUSLI1rm/NjkK8VooIpKj4bqk2DFk70F9O5THa2FHCP9ih9A
gQeTjPhrrfBCgs2blNtT/q/Qcna55ma3Rm1NYq1evfmT8yAPOEU53zVdcuZ2AyXFsXVdYJynKmy3
ahOuSyKCHQaeQckccvDLfEu0Ew4rN5Q/6pU3UnlrsHzf58uwA9yquK97mlpRlps4wwBy7xjWd4ER
TrEEpoDJhCzMCW/SdbjigbcjuS2NwFgoS2yObcaZGrhEEgMLmT/X45ayYczFh2jjkoifvzjleH/x
KXGhg7W1E6l75/TMswaFQJVK0gAhZxElrMEJ+BRNl1ybMPtgyPCm0RfctL/n772iIg5h2T6m68pW
iooHsGQP5JdxXsxGmZ5+0vX7Lokb575AEIRHCa+Tp1/BtZRlGQsfnO253BugyU3bRPzvSl/N4q5V
ylgYQBjIz6gEFGD8amch3VrLIG2fltJ46miby2FvJmO83k+2EhoSQ5jXJlKSfCrIsRzXVCztW0CG
GKubU8W+MK/Q1aNfuaQSYenfIZX9ox8P43jaxFrahtjsgwfgdMo+3Y3jpcRH18M9B2D115V476fR
uTtPLF7g1LhnsZK/LusUxHpqE7QbgX+LaMP+pS1wL3uzBM3Ne+szJadVR8knbMAFFM3/bCGVfzE/
1C98R068GC9ICC11jrPc9d4lIQrCrrfXEWBFCeq7Yt0TCKAghIcq8Bzz5iI38PpCHGSEUzNR/65Q
ahk59rvpWeSubeflvjXVYS7edURMH5E2p60b14QufLQYPvbTwtitK8xN+79JQ8vlCHtCFrp5AYNb
AVJLn4T6TTK+s6EEp7sBUR5OPnNXD+TePRdepj7ul9e3PsQWjDp0M5HLX6Sr+531waO1C5R8UXdV
EvsFPD2JRXYbo3fQLaMk1RYn48eqV6RErQXV7mIdlOxf2PE91oKdG/hUUrinRX0sg3KEtfHMupTo
kITBIKRG+1Fh9BGE6s6aq9m13ZG1U0Yz5zjLwSrXOu6iTqRXIPddFqN35Zd2rNPHXra0sAGcm9ZK
j7uR0mZ84sDh2DYMoB6WYobG7p3Llwp4ljNve22WMy/nnhausPRdN7Nrb05DIsk741SkQmDnKX0H
GFp4bsvFlM0Q9CMluiKj2l31s/wDpUIUshU7BIr6SACP9D3fbp3iC/KxAvhrne9mSrZMjt3AL3Nw
PFOp34nNMpvFyxaPm7lavLvCtiOW2vOyFITTX35HbTcIfaUnQvlr2bEQM88DUdBWES/wnixVMHc3
1utSN10L28/713qv5ZIiv0pwjvMFbip3WIP3PiOXEP5bAaQpbd1GO7sBQPy9Z2hKaAEesjEYbSQE
1x+31KfatynjwQL9QNNntKQEpCITBBF9S6djP2vEF0t2DQIROZ8AS68DVNg9UjMVuMU8gwvLt0Mh
OFtyoyPhD7T34c8a5meLALuUNH+ux9LRCguDbyYndRqe4g8vnRP/tNUCr5XLsssHA8oVSrRchNmr
aOO1YSNxn/ACtqgE48AunOsntygiFG1V7mxljYJJaYV0E5z5gjzQN9iH0Ueg0lZH/ncyk99d2sdx
YCUe7oQPqhYv7O5XkGJ/W/9V7Gs0nAFCQkUgfS+QI+qGodyZtj13s6juuP/FHrZMWditkYFjS2j3
lZ9btEBVOEJhirIXexFi8XxawKZ047hN2waxJm9oI1Abhohr1TeniHBqZ+r8Umqis53N9esXr/A4
izuEpiQ90VRajm2brsd5M+2nBSphOg5v5Bu/SJQxU/8YcM6d6jvyXgpVwKGxZ7XgR39AOMewtUlm
w8iq8eTvrrpKCeRTwrRbAGSpZb5535QXRAOZ5XB8QEt/SObm4nbMnAdw0lpvZWDLkvix+fc+n70r
P+kUqk1g3j4c6BVY4mhb5bUVIRNf+sovnEC2YOh1LWkAxtcm46s8RpiWZQbyMQAKb1lqusxdSaqb
GqMm1V+8jvhDIico4UcWHNj0bo/gcNEcNWxkRl4py5Rsqmf66Ik3RrMU4urOVd3dac4kLFa1NTNv
RhqsyqL5kjOXoHGicPz2Y4SNbDEXJQR0S+kgjXJYp9SiBcpYK7yD0HpTwfO9i+sfeXa4/HY4FNJI
9dycEnNjnw2OJH3eHr7M6uVfatAkp22hZF2YaZLPXsZF2RPjumL4FnnjTqbFg6ThdYeQRLMYsI72
mMT/QNyYPV/w4Rg8BM2DkuHpcsIuz1irAFwMEnQ0S6QlatciImXUFyBKldvHf05b77pTzV7gmUnF
hpXBxgiDWmBzkQgHj+4isD0MwBJSWnpVLC9qzDVysunVqiT3RZ7KOg7tjiq19yySFWhmRuQP+nOu
t/kUo8rhsVK2zBvV6Z6S8d7mp8FyCY8+7BKBQbhSTqzCoNaoGV+K+09+WGQ7k8neF2+qNbtzFTFe
eyDvHIZV261jTQ7fo8ZPZD583P5rzMovmAKUTSL2wO6GMF8VXEk7xsdOmI8CCeH4W43wOTTtbTb8
wHRHsH2zoTuEsHvAdvg1wcSHQUGsb3M95TkgsUTzXhk0vo8mgaqpl4uajM7XzuSR/SqNA39TeULT
sDhFYjgQDyIM+B0Qk7TvN+0J2BfOFW51P2F4NM70Iv8A53YpBBSKbJvkMtIfCVjSaTlO8jHmSmMg
21Tn9Ptp1wuJr9DuKQZvoV85trgRV2advYUaQ/gBENb5j1bHYsixMA/vkT41K6OLLJOmx9uioaxC
ppmg59goyfDO+sMxGi713Ksoruzm0C/MmtAh/c0jIob9ucbywkOwhLMp3mbLSZgeJkH4qH/Wajg3
1CQcYIOlGdcBQeZYRVpsew5sGOrqmqXHes5eumOgAARycmeqytCru2VSkNcd+Ke0DYLi1R+QIMpQ
GEICjJVYthC0jXmxmFfiMFJOtqns0OkaMCAsJ0wqPxBZ6n/QE5gzQfAxvR8zGDQowJ7qRccF1Ypr
98XIK1uKLZ9mdPmNSsk+J+ZlxCDBipZj7/mi9SfEHL9pxncW7/IGVfWWPykaAfawNc2d/6YBT8tz
euxTF8XiBIdkh/UGcFJUhU7lJMZ36XPdD803rWR7NC2dtpudD2h0s32Z2z6V/I2HePvXUgBYfc/H
CK1IKHbOPuF7dCD8+mdkwFOeZ4dq9EqKKCRHmE6JnbJPtFP9q48feUMu1/z+Zlfeyufs7mnWc5OA
Nm5/8NV8ctsviDrW57Htkwwg27xsRjjYf+wLh1xrAjzkaLNFV54JsLlVhsxk8Gp1I5r92SwEcq4n
gBhd4A2T13s+h1TewYILBLiusVhld5B//9GPtZidpVSybvYfP2sRozQdT/wPQm+XtBg8Yk1wady3
GXCs4XWkX29ll5d5W1owGYbst5ES3nhIOzCwDpVuOwFc532okoxlrtjUjXwzDKdAm1Ugvm1cxovB
gUi78MrcV04pj4M13EMQVXZBLin4JzYIReKTgh5OX3mFa5R8bxEP9ngc48MZ3KWzkus0URvFTTrt
xqOlhu8u79sHSgY/QZarc8bt9EvQlg9LKBDtH9maH2uJ9e5qf3tmLxloCrGMzKZFo+TlyB2Jzmko
tN5eHvQqt64yMRK8lxgTVUdihekfjoNybvwYvirQtwyf4um0y5M/RXsOHyCGTVx4j7Mh8E/ZCbiB
bTAScplEyAXg/leJeSjYNqlXqcQxaScZ7XBq3DrP0Zjmzn1DqNXYyYyuM9TJnWsgf7Z2ZFk5V+te
43E1LU/1GZSQ5ISxcq5FuB7WhgReR+pgJ+NX/JkRqjlWNGdtGohfahYTLCcQ3GOGcRyX9pgEaxbh
YIf4MPTnKGlvwU3xUKq4HV4oCYi+es5epJw1l6oHgTTuDtaQ5H0niAmDfZHcXJESixtlyZHOytW0
dGB/uepp4S6y8x0agEytqS1+nau4dCSLWekqF3aWqlsqUar12YZMznGkZwaxcgGz9ezA373k1rLB
dGytlJDVgI36Oe0RCEyGdyP0TOSfuY3CQZBzUPGYB747xeIFRLUCnEf/tbUHCO76YG3gOHj0lD5w
B3jEvhL5WmJlbc3d9Scztr4+5I2pilXAbxy37VVRuQMW/s/PC71Kgea2NCXRFrPhDXuRNLRhOGL5
btAfdMWc9BwZQ+U96GwzVA5NAOcXEe89C7ujTI9wt4f+Bl7xjtiHLUcbKJcUqljJdd+oNgQzSC5i
pV4RVPjZTzYzKdvawnfvRuFeRwUp9JfjcKzFTL2IFjSnf/8eceC/V0byZw5Hu2qRhxqQGMa/63db
ixRoqlZYS20vciuKvaBPc/lFXsOAuFmJuED7CDRpCRXfnDDKEzxWPgq2t9U//EUc1hu/R02sBtNx
vY9V1zbepbqvJD5t6tiZME8CxUtXSqhb1qnXdgwePLErGfYulF149SvsPfDS/8v5bBJnOsSwIf5k
SkIwkeCoskNTPyi96ezlghnKzwJg6iSKfjNl3tKmURHR5zmzDXq0Ojleoay04fGZ7eh5H54KnW3B
9dUvWvxD/0S1cQMEAppKC+Iv+3lOElrzkwetg/afB0Wfs4HAZdn4xinGRk+WPNs7cfirVhN4pMPn
hwPFqSJobr1KKFjC1f0M6jsaNK4IUJ7MtnhmPpjrnUEPnx+2QVJmBaOQFzaNEYv3YacnV1u750NQ
UZzQzF5/pRMgPI6IhT18VJavGiyqyQPbEwvZqInlvqjVH3ieG8ivD2hNBDG+x3S7vKEkY6dCAppF
brRHsnj35tJ7sOq5aLVKDdYa5eg5cZk+v0fulgCjClM0YUjLTI2VhcrtsNoote3aUb2OKe95Dio3
8v11WHjnTpPLeNEQQMtmEaiWHn8llzM5VEHNKQcMn/w0JoI5jpWBAP2EaoDv1ie+OwGSdiEAlZBc
zXvMgpPEeYkkiMtlg6qD+dAYc8eIsFVtpTRR9cODHX2E6gvRYqJbbZbXvBzlZ6ozv5zn+YvgzWbc
M5RBE6/soOr2CujgeBLh21FFEZfTCt7yTncHGHYNoILdnBp/+WiU/p1S8wi1ruFHSRYtrr3nhjaZ
/nosBcrXS+Zcnumtpr9XLvJ35IK/KFVVyt7RL6Z8Rb4rw8xT5nToEHe4/drZqw+Y/p7Lfm+Dewlt
mkzcApW1y3fpyNKLNCjNSNB72/TvyAeuNHg4tUDVsXVcuV/VUMYbDSEtv87cb3MX+uusO2av7OEn
v1KI5LwuZOu5lij7frV5fbA7DYTY0oKvkjY1/lO86SUA5+nIge+6RpsjCIUDt4ZZl07oJ0wU1BPb
OciU3tKMlasQLYkEgc14xHB/3DSqCFTPi4QZ+qQqG/6duJwjejFyBAssLvtJR1E4oJ/vAugvL7Om
5cyKke6vORVQ9eVKWhR1iXKrzGGWPQtaTuFH/VyDx9gJFrwtXja/kZDhTBmQvAjpNqQO0omnk78s
mw9LdNSq25K3okeEvuOhHjgQYpVBOga58VDIFq7Zpr0NwGHcdDjoxKxq19BtUcZ53bbndepu6v7q
5HNwa7WKUwvrwLK9HB3jyjX3Q9RWhuCwXsUfQswGQhMowJC4h2/A0HaIrTIQvDh/AkIPGAGP6/j3
Y+SyigM59dsbpYK4vxcgkIp2lPeyHac+XhWZyKz0gXXdPYQR2pcHis5eYWVaK93axYfWg1AL/kC3
eNoSkz61raG/J3Nc0c4AVOON0xClx3nmAyxRpQDfbUDW6ibwq1a9zDA+k7eTx5MVu0VcLaN1Utb2
TyBr1usQ4y66SNrDR6+j5Wtx7hosNLuqKKQCiUFUH6X7Iq3KM1ME9Pen0B5orQnVGuTP4RVd11fd
GNkc0299zQ0NOSwl6omuTR/uftLCbKdym7nHacqDPPgQgcr96eZf/RlDDQB1SxU21z9vxOhvsB1I
toinrcZKof6QNr20mpij57b1BqPlTpRLs5KHwar9SlRdTNL636Y5AdBg1PkwA0h/xrDlVLL/gW7O
Tde4zaHkoPQkG+UreQ6k/Avq8emN/eApu9+1dxVXVnNgAiXkK9pw0A+HwHktGetTgiQA2L9SIpw6
NCDkQhl6YYlx2CvhxDW5N8dsZ2A2IzUHmmQ2ws+LQUMIs45JVq+3XK6AjH1FTSMRXcpYBRTnP0ab
/4a2DpWuqxQB3cnQBKIYC5lsUzTuwxxZYhZpUrX4vUcIaJkIvNljsjBBQ2Ylo+zDdIF79R8rTe2z
JTDT4qBOOhsG6CbOUET7mkjFCl4a+bJ8TgN4jsjy7ebNUhkVzW6cGDrDC0DyHvLIjeElv4taVxAc
27vzDetPIppi4Y3mBuyOQ6Q64xomUveW9dBJRxqlrPzVYiIWRB510IYsSvPEUkfLs4njJ1agZm4f
R2VVgxYWxvO4ATSd60rsanDajc+PyRqr/C4TA5frmzeE5jTiSGzmnWvTj30uhgNTQut9Njf12ZKC
8FKG7FjBlw4/m5iCOdszmWI6I3A5MfD7nkW8pnWCzLyfRz494pyqSwFdwQuD2Pn7u1UPOOXGq+tl
N7lgY0Rd20NfbhT1pq6SNhwfUi9CT4FBrlqJ7qw+VMNGN52JDIfaHq3P01KoDqqwp2ABNNlgGVvE
Uj/HCpGDVV7lQX5IhBoNLfw5+Vxee47syH3SAt5QDJXnrUeT8plW03/NdUbxCFoWtZLr8zKrgUG6
svqLyeH0R90WBQLM3x/a9n9abJsppUdPueKtCWsplrrA/D4HfwJdeTdH+IScQgH+7NdyPApmLiyo
2v56MpnC/oFpAGl1rDLe24gv8k9eVsftZ234WOwQth6jklIdZDO4r8pX0Lojdqbq/fYubjO2/l40
3kPzpCKhaoZMp4y2Al/x9Ax8x3pwMThfT2Zha+ax9hD7pem15WyUxs7tEeDi41w0ihh8rngCgfwv
zOvy4xorZA/OxJSO/ziYcjXoojp89m/FoIsV5w70VKhM94+4BGWOt0zGwhmjXqOxD5nhZM9LxKP6
llbFxO+9cCfBsB7YOgbD1PXyqsKT24Hunv8yDsuy+88TydKyQqMALgawHfNVUmB5M/QCqGgyUixz
B4cPrnsElu8vXmS4UXQlkIZd8S47lsxJMdS59xaoyOfPHO0wXudiuEPoAN/j3ZDJB12l1WLR+oDe
SSejaY/b9PFmKE5i8x789qLlQiHsjvvf7+pPMJ3TPb7HuUBRWdLoroDQc24k5Q8KfCsTPAY4WbTl
FiwVLeMh/rZM+zkd1oefnOYKIKpuXBqYc9Z5JcBtX6R7jUvtfoEaNQ1ESZ2d7fuO4wcDCeQA5fET
lcPOBXHkM6LR+ZvUJW/ZE739iMb7fw59a2FW6ZTNaM9c97apNjDr7WjS6kyuR8gghdLc0s+fyqAN
JR42H5t+NtFa7P8ZAw2+ZD8Rg/+BuM/+nOQcOoi86meLWrVVO/8eMAGiGnWpM4Zu/MVerzujkQsM
AQKuKDe4T1OnLP8FGnILp2KXsZ62ZWydIs3UA21Cm/Mk9VwBPtCVBpgqMiAGxL7rsy2xJl1/7IF+
DBIx8IggLQqEvci3VXYpSAHU0bou09hLAzns7LgjySTC5iq4t5haFXjebT/o+qLtwxRLkg5nsg+n
REjbhfphPhX1haZWXWam8eO7St4EUMBSBB6b1mikoIYklgJFB9WBbowsbdwQH28zOa+427CS6arB
OOPIDxQHsi8jlu0MvCUvPDhuUynAKFa19dpBI2keRqOoNhZT7u1BUeQex4jtoHMf0Kd/tbWirvOz
oFEIOhGVMT8ohPB0veuPZA2xKjuyS601CxeePhMeSaX+q3s+kZAaY2Kv7t+i+xBdeCIeq26jK0xg
t32LzHXbRr0P3Ejso3r/sD3idU9q7WxdU5hZv3Y8CcYkk4/Ymgg0AVdGs3rz3JXApWURpk8yKz2j
F0ly8lQzandt+bu4DxZaMsl2jI4Tt8dIPL8rGKZ4RP3YQfoagQqTyuwDcfqomR7+50HHz2qXjE1i
ib5BFgsau86L3329IYvo+PMIj278s7dxyFolb/5+FRUtg9G04qL3CLuMTVCd+vULBWzmrBVk4JiT
ZB1U4ifmsAUgMdwUS90WZPKbdCxPFU50Oku9Flwn5wXB4F9G0ZmS7P8jeJNavG2CjnYZd3hsLXr8
NQuVzlsZh48ewv0bGpG2m57fQVNqrnI6qvDyhPUYGMSc1Zxh5z6uVp3JrrQpTdcsLhgHoyTgEvl8
hyk9VTa03/5cvVHDF/dafEvjXj5yXz7P/Hob8lNsIUwEnAe5PK2WPxDTK7V0rsdYF85njW+/WT4t
+nOBIyEMuPZwpxDvxJA/q9PTW12GKkhiYbRaTa+WndVgWnap9mzDZrr9nTwtIBs1amYDXfKLQaYg
66Jm/mfbog0I2AEw/3VtU/w4jsIQPm11yRKGGT8lfrB+N7v4GOIyyPmiGmSAHS3XRfzOmFI73B20
9P16P8b/Ihw1cfcSYexOQwk10b5yxz4DLxeacFpmkYVeviyZOObgTRP0f1cXclpAYCzXS3V3zFn2
NoI5V3FAAqIQR7Hw/Gt4a6K9wIEhaWD3617HPigbzdoCbxpalincl0OHvpNY/Xp5b56X5p3KkdvM
UAqK53RVp/yGHrQyFZEAurYA/mMwbQakboL8yYsFDybOc0w2jKyf9/cPwXrQg017nBZ6lRH/5cvk
UWGP/RnhVemzkfV3Na0TOrFzFZLxc3oHRZ573+K0xdi+rERg0QiAn7ktMAg9/TELQfGwVZBg1/PR
7OLUNqh+I/I2jK4Y0rU/uWTlVfWI4bW/bAeY0zwj7fw1H3blOIEArXFIHI73c8usF0N+DHSC6+wm
immJAKt1dMULVpCORWW3t+0nlgw4eORde+cgCd9MR4jrLgtoUiGBOTHanJQXSwiYdOddZmofQlAL
teG0Vf0gEgq4H0KMjVzoh2aXAfkxJtT1J0MBhV7jiU5vsKnPP5LAqCYuwtMaykPlsRiV84oHPJ0g
6V6l4C8L3fcge4+ORqisPRNfx/nq7e+vYcHbYQxXc2Z6U1d3Xksm88iF0bJ7s5Ae1pWtozxgviQa
qGqb7jrypDIUOEKvfpcEyr1y/2GTNiAEK8lhMIDP6v07lwJ2BR7t7rM1Rv/3+9jP63tKMO9FzM/0
jzgFpA+V9x0ZF72C/mB/BGcbPkXzjDyZRcIMUWRO3adVQ4ExpuefDlmhXI+nkhlM0O398JSj1qUP
SmU1UXGkFtgBEbmi4EiVD5VAMVabWCFdulM/SgWhgm8a8BJPWX0kRZJqlnOlQizyxP2p6cqY6JhP
bawnbBvTjAyadDk8zLmho8Wvn2L+SAbJLvLRaCtoAq2s354BsiP4W6LIQu2VSFX5R5k6N8P2CkH7
F70anZv1JWp2tVKK0NKHQvZ7dZX/SX8Q0NDzMvIydbfgPDwGP305LG9/8vCmP0gBgV7qHLwUiG8R
47MecPoyG2m6RB/uB0vkuO/c0g265KMTaVhURJlSdjxxGIjsgj33x5t5/G+k1SCy8N/S6bj24Xg4
NLzYMmkzG1e0q0NtagxilvQdpLUI+P3GlmcI6JnIRsfOlwiQhLZzjmqu9WeQltLcYu/fhLcgcQuS
XMJE0cunrCTC9mcPXu94saa7jzAaoBrWiSzqtaAPLh8iOS5ZqwHc8a53tK5NN/UQSznR2bDiS0Zg
YbEcDDF5OjN5w4zoPKL7zrgBLrbf+Yg9lSHYbuq72ffxRbKAqTK5++07tFA29w/RBRNg1o/P6nIU
q9kZMeLRklHnLDRoWD2RgKAXD20TGKpJRP2Dv+6n1TM+qYqpYlXaNBlNtKjAH4kq8jwo/CLzcN8O
MHwaqxz3Ta7rbqfoM96W1lWZF4Au7O4kx1GjcVfCZ/JhCCliFBXanoEkYADHcXRiNqHs251nQz6Y
vRll2dSAZW1WVn7hweS245EJhTH33BSQoDsmlJ6feI0YQ2dE5nK+RxLuW692gauysPEcodfp2sWN
/2rKMbEjkh+1QGFP3j/uyjTcP9ih+xYPb8ylpW90V9bJGDRp67QilZiSJHBvs55juR6jzMOc/DHf
yb53ano6181NOYgOHC9NsWlckDE80x7iqjBVdqwrDQMtDlKTu5M6lAzJ+3jp2vLadqAKexQ+4fhM
6zdIwBXC4lAwYN352OaSOx+bMGK5QX3qNjE3orbm3aGfRqLy2PS4npbJMVjxSdNSV/E3Gb2X8Hxg
DDBSNgGhDi+ka65nW+era8wLN60KYqHVAKM6fm1tmGewhdQ8qE8UV22URoThiQp4xc1znny7aGra
5v8hmv7pFY+hrFfFx0OU/lMGyV4vX4NAZO+2oYjlLkVvK9AiDw+2GUbd6tXuJlxe4AHHf0+tJlgT
N0LJRPE9oQd4vXez4c9n3191sZmNi2YNNM/tsRhIQJMHcsYaBS0jNigZI5tDsDYx0mjx3SfumiV0
y7GDjhP6v+odKJ3xzGG/IeGRDOaWANrr/TPQ3QcPnGx7h8dTaFVfZ9lPnMQXXBXNzGx3woJ2opc0
S3QEZDAefS8uoHc17yl267UQGbdlJAjn5UYvBvmtBpXM+4D61ms3ZejB3DiV/KHcuSApW2t3wPGc
Wcp4gepYYu1MZTjb66/YBIzjdfmpTUhF8YqcmDX36gd0jsR1SMyXEDdR+7DjeHiJoxv2cKTQbh2I
lhge/3EEpNZ4uWQHxSx7PQUC6HJscBpe/KVo8RClBwcAVqIb8+4XliXs4IT/tEVO/Qh96XhWsuzQ
rkmAPA5F14vJCjkFcp7XYgbC4n6BMVYFdtJvxsO3i1r4jVMbH6nJdUVgUhnFrQWqdVPtDxA0DLPo
ySuQObMU/Glhfwz61Jpvtc/bX/h/6thiew+rAu3xbO3kyhzaw8glZBte2tEXVWetdHxsxzoKrN43
c505mv5mINcqRuF6bMXqu2WE470eB6DqSm+dNwhMRBvi/6o5DLJVjFfJMBPCMg8AmP6Svxzwf2wV
p1wLxLjLPrnGUrOsKvUcdtu/PO8cgG29nUJ7sXcEJNXGwEIuI6ji9cGsfAns0/xRz51AloPi3y99
JeKoUop6L3CQ7Bc5QPd8s91cXGEYZAw5tPWFp1xwy9zZYCkJqhBD6zmxTA+l9Zqt4afjC+PEQYy8
UN1t4TrSLNx5tmDU2AQPrK4h2vO26WxXBzN0W8ySUcZTqSb6ChZnpbM8/hiolqc/v+x/QYtmUJ/k
g42jxzFUw9igJU5aQbmkZfB2KB/piZEvAkjp4Ma+I3oYdvCIi17QSb5CeQeGBMq0r7o0NXHV32Bv
YuRXzfNqbkelw3KkiIuLw1F63OPepLPJP6O6eQ++S5JGk+Y1hnsSbsAOIJ1SOEwiGzeQ/RAh0iUO
0gTSsgY5mPdZOdxeY/s4LFUoSl5JauSje6Nopnu+fckzBx3m5udKq3j0AY3tcsZAg31dn+BkSoQZ
8mFgmy+kGZMKxXWp+FUlR2vwCZxcdZEOp6swZ1RzgEv8EYWcCfGjPWL7aF3RmJsy/ZkPwXZEtM/P
cBEqgneI6LZux6Y7TukU+UwBsAMJwDYJpILHoaJGXKdxOr4ttEFMNZT5VJdMDX/IOCA82Avadpbo
N/viPPrVSkbBUy85skwQNeJSwNrrqkjcVv6zSCYwdlzOsXAcJNg07bDMtDBx6HCUyttF8P5PODR7
nn7dBBd5az8aGw2E6c0gHkbjWc8w1HQR8ynGeTCHRitSwkKiqJQQkAIcpWEfVUWBafHpq1HeXZPm
oB3GBbzM231ZdoAe/HxN9L1ZCTIzuiTPU9AA6agTGFpUhvoMKxM/nsBkRKvGiJ/dRfRgD+Y+uhw1
tWxBGa/jdud9ISjzpfedeUsmUkZZ5bNHYN50jNDLSQWaRgg8T3fvVl9o/Dlty63va1g4EMSFRtjM
JZWEFtBRe7r6dxdOun8ghRpuD7oJ1fILMj3j5NsCS9AKbpC23JD4HwMzSRpCKIw89R35FcXq0dBY
AtqgOUrGf5Wg2LYqg7M1rHfKbbI2CvpB/lg64NLqSANRLt6ZQvqfXUBvkYcomF4/i4bJhk6BlGco
Id8yF/Ip7eEVMqoCsA6a0px9aaoRxXRmMiV35sm1WdNRKA+jMMr6GadQlSiaUePIaot+9rcQg9bb
hP5Zwo6SBfVAxqbfqDF/vcZjTKOSC8JJSiivSkXzmw9TvnD9w9O8l1TxPoyc82kietEORawUCP9K
5oEpJba3g+kkeMQGWwxBWsRandO1Nus1FXblo0gbTr1m2SEEHRjdlPTqHU5+Do5401kQXcep+oI9
KQ1OsDrzJTzHGs2mQYa9GxBaMa02mmSmpAegA+Zljo9t5kuV2tEPD4j3GUOtjbaWaVYz3c2s8qV4
gg89yTvEhWacmj0WlC9V1fxNRxmMEU42+XZdttCRfemIIs7E+8wRTCFPYt9n9bymf2jo+s2Or3Bf
kefHLwaiGMgS2vTxveqadXDhAnI3PLhOZJl4wn0A0jJwfI5UfZGTacNSCpO/lT3IL2MUudZZr7os
NHKy7uY50FwiSMGrhXWZOTCL4PPXunU8i0j61HYu8r9VOO+76DjMCOHdyHwNBIhxRN7Rc8fUztb+
/uvCMW2EnjPaBzHKSkSajbxiQvZe4Tw7jHv/FHXXRXWOimsOYr7pbK9CBMWJgb3cp3LsuGMVsF7e
UWHZpsfr6/1MW5QYZJJ5szZjYWLc/NvQxIBcXAWLKgJG/KArJaMoNjebUzZ1bpzUzfwlJ9Pz4Cir
JGPiZqCppoiNxl66kubu/DS3MGRg2J19xUp5Uct3CXRCisU/2JYT49s2bQIjlwJePJ/3+8CXqK55
fnJqcmm7P/slfr0K9jvmygjv0RzoOVUuzFYzD5SW/lw6PouXSwyaEr0uPH2UDzUW2h2FOmBljtJt
jFenOCiWYVRD6jPKGCmfx5WEhmxEqoPIYKHnFZJ/+CuU0LO7/hmr7r11tGxSKyKeDodM/qH2g0HF
dEnnSRA0L4PkheFs/IU3ySpRhTSFHSzQ8yuRwP+OAN7vpE+wSCATFhwGvQS+4VFllFdt8/LYD6dK
Qilzn1tcTvg2cqddy6JZ7Dr7SySi70qjMP/oE6EEvReX3BAn/TH+kEDF8IMoRrru1W8+EHGYJT6/
wFH2xYF09pN5GH3AVeifDCDr9ejh0vpIB/CRS0Y+qcnWbWyELJOUwjxMX04Km6Xde2DH6m7+iZz9
yGg6E18i0oh08jS58x6Y1kBywZTIwsEQgLktNxi2i2DGOHypaqz3+tDvVB+Ja/dyQ40a+z1bxogV
dWbJd1QhGvdVPB1UTy1ODl8YicnAi2jhBD0zwzVIkp1TpK4IdOLy2T6AF58mpWElvkSkiYSQWKhe
ZkgCALESNRzp16Q2ibxglfBnpN7HpeJIrfTZWyNSz7NvN0+nr6MBdrwgg/NWdElHITNYBz8e7hk7
R7pcgASwIFImbBanjREZXcsXBiFNbZxG6DZDxr0UcKmu7xxEzldg4A2C0nWxJ2GrC+5Q38WqAPQN
50jmWVG7ehntfWcvcPuQlUVBW4xfejpzLYiIuahfTpafNpoQVAJ9WEceHJs/zHOkTpMdZAggKC46
ubuZUt6eadZCK3eYGcyGXaaYz5UYE5amtD2KB5vy/11hx1V7wN1U01+pkuDm0kIizG7TMchQdOWy
1E+qA4p4qYq1RkMTlKYPCtoqDU0FHhRjsUnoWwIVLSg2acS97hucsLYGnC/IlBcTsAqXKFREfNaQ
QfgyAwqLmD2ZDm72Hils5BaE3QL3c8iprlM8vJF/VnWKF7ZqJyS/XBT54raoflbrLFD9KURjUpcV
ZKOxW3BBRRfgyX/HH/wkMmmI/BwoLnQqVnF9fJOHRNkSX10OMR42h1svWwsnOOx9uEdAHmyStUJx
UXbYkI2GmGwkw1KNCO7jZxBXZ01YLcmonyT5hlyWHPZMYhE7K8lp77+GeixNUmI055qgSHhswYR/
Ikmi0cvUNKLKHbii2zidIPBzZhgYs7lMMc5wIoPVUAGW7Pk2Tuyi93tDakb1JDN9ycuV/3Su23Gp
sYFC49ZqBn/0m9kjS4Zbaisytz4K51EcS2i0brQGOwjdHCwdXOCryyCnARdoZIIFB1d1ZRd5C7ac
qB9WZIX1AreQzYRfYSg0IKe10hIIur2F2l7FAhfNgIwPnKEiY1SM82J/6NEtT/cyQvVgqcFxBVXw
/A+O73xMZ1DVktYgp5qEmKw41MJ12W2DiRSnrBytDLuKBjuOHJJTtxgIzsKXC0wBWlU5E5jWz4e8
t/qWBHxs3TLTgQp6ID2lKSt/nwPhwFvcZLuGKJkpvixcH3oxH/g+ZxLzxIbOC//SQ612mQwwrboe
Fkv3ADOTF1f7y7WEw+zBGEOaGr4DATsG+KkX2BY4tt0dE0B+TNR0PxxOKllFDdVJUR96JXwjSBcW
Pq/7br9jRk2iIDEQI8Pka3OowBppqwxk41JJ2CacWZiEFCtu8exqUg/mXO23GSsG30tGwlNEeo79
IyT9oVzUS8VAJn0yTKZncx9RuRL76yKuCl+YQjhYCjK1uw6drp4E8RghORHGj8kOY8qzJlp6OAX6
G7kRNAR07AqdX0oG5Z5rWbPlrcMikpVKxdFJW0XVyTEZUbLp02hWEMrsfCanmi44Jtv52Psji2kK
yVpEQYaIZfGw1y6ez2w0/mIoZSamI1YfSaLAPR1D7L+l8orzAIhvaTdlI+pH6F7NzmMec6yzoUuf
sgiaRSC7iLTha0+ZjihB0Qrba4a/NU1oDMVY2VWGFGBagQpsmWanocy5D1VlAiNZYlmwLhSPBV0j
Qi7vVDhC8iCx0XdIqVxo4fpE5De0sEroFbBG9q/J1QAOX/rQiI0jnTzy6re19isvefCZarYuT3Px
E/OJI61XRmhC5RG7SrJNB8xOGmEAjSzlaJ3T8OoHryQePIhO7g3vYXBsuJoBc1/rbBr8+fwAhPms
+oRSYJuFi89heBCrWOIyiEvT+zU3Ve1nduz7xD8Qu0R2dmx72t5k4Ob0GfqM3Jh/pfniMN0mpARg
FBmQGcaVMyE7OfzAjAI9cWlS8yXmYcU4HVI4H8cdDG9UMfYtitFdtPQiZYSJ2ktPDFrjB9XUybsU
aEdxhcIbGMb66nP1ZscpSKJEXBhocoFB0pQYZe44JOatG4iS3C9r4TNBFQAhZcGxdXpv9Sx7RcEV
4Us8YrVmJbiwO4BezDX+w5BMIEdhezkWjQc3i9R72mCHBccxIUnzb1ecg4k00WELIQzrt6rkkJ5D
XEIyo6KdS7pAOsHu+Ytppwkf7eWrT4NSU+y+ySwrEdNH04uIa1zy2hfVPhmNzqHzoQdzxiwxkiM2
8nKeQTSED1fmRlWLkapft4pfUCNYW4cIqv4QaRot1jCsOttK2efsCZLTzd62YwfKgAcjzBMTvf0d
CfYj8H/YpI1FYC0QWw5xpLN/iu72e+mpugq3Gxv5+K4JAlHabM/7+0rRtEOOg2FtoiU7SS1M2LY+
0KcA6FUo1/p07hf1iANS2u6NY2fdU5WQVYu0lL8SJr5DBQqnBHmGnY0EDxjPJULlis84bKiQHslt
62+1eSaVJn9Vsv1oB+ZrgrkeZf8GqY1ajurMXEaI7ncY3VyUXWzecG033SuofUjguUWI/+WVlel+
YINzz01sakpHdyyNZuD/Gvty8IwHITW6ILdLDyWIEDxO/BajVMn0L/VtCEogXyjPHPSKgeg2t5fS
zLHDM2kohbXeW4wD8G26KdDQSS4IPmhHyLEH+qm5CpykFled51jakM4ys6EYU5ZgYtVfbGafcPHk
vaPvT7IodzVZSI7KfNYZOP4PfNXkLXk1arRrGEwz2HN/UwCYJLi6CucE3OeOSorVseS0/ww4VlSQ
a2Sv93KJNj02gw3Xh7dPtX5jMpE5cnAG10rssMDR1CU1y0h0L7/TpopF15HEcnD29kIW5IQ3uzBT
J9UbQ0CJ4t7r2mwnUHzmGcO3UZz3xRKFNt24zd3AGKDKrrbpYLQ8QhTlKU74zZF4hvG9vIb5hcGv
unHyYYAPT853WsagoeCnGuyIvvdA64amKV81bj+3TWJNY/tCU7EcU1ptG9fiCwleeNb+m6waXjbl
Xyvqz+QFvXgxdvp8I2Dubbl0EhoBVBrVITkkJ47BTHK9vBafFVMqNdj7nLWLHTe3GLFufU29qiNr
5RVz2igf7zZcUTmmfyDoehQAjqkhC+CcXdnApDkQye0owOW3iU+YLgwzOFh3J9tOoOWtUQn+kQ9O
T5HKyT+3SsyhO2AoGD5valjErLJm8InDcseuFCYSpC8ZrKTzVc9KSeu/iRgMXAaCcPvh3B96cJKU
DQf0uB/R45ZUWLAziVc8ZfWMThRiDbIlll0W6fmr1PQT9SmEE0pQzoMQqyqiYawQlVE55dbx/zCA
0kufEs1K/bd4JNP29oRs92wKWuTB4CnOb+QSdh2edrL7BqAA6vYqI8p9JYyIUb3WFqZvnKikwYuz
CF332nu5yqfra7kQXObi6QIMP49Q+TxfVlf+SBD0UJc1HkXzD9DihZo9urqF4vvPUrAdzT6AmmsD
iyMeYiASz6JVi9UXAq6xwYZdUUIGkogaZdU9gWqRet5g/z7pB2ShyFnPptD8A0D9xEqy6YceBykD
rMn75aUBN9o0cedCW8ZVRGEStQ6fW+SmCruD2vq24hZg8Gr3DGXwRPtSdqes2lyqvHmFkTz08pup
dnb0pUj9IvuwEOkB3A7dU9+XCxh8gF1/Em7jR2WN3hGPBeaXZ/ZwTAad7IjR97BPzLL3yUOb/qMJ
PqHeWL/hPJoKLu9YFbLFsNqr85D1IUz9/7fk8nGjpN3e8zT26iVFg2SxOHoq927ztvN8oDmqFzz4
qF3XbHxXswoCKKkDFfJ4NBMqS6xGpsxV0GCn0kg01LRY/CZWN5DdrPQV6Jy9rUhB4P61RC6bmVeH
IGeb0NaU0ZRcnC72ZrYYdAb7QuHgdZq339v9a6L0sPGWBn4q9Q0MgWZKBe7AzTv2ir/0dPiYra90
Bc1r5dvA+Tn0n306/Ds6dKJEHIv9SViwUIMBckpHoLL23XzaJFMeocNSM95R4Yeuwyr5feXuI7Au
GEaOz22SZInHjN0Ca4ZSwN+7IClAo2yjyoh6kxLoPpJaFQiUjBt9V3Zt45sPjlxHtHWKCFuuhHMZ
s85V85jqsurlSzRgJjuk/tveQTTldewj6XVRRh9k1/iAKb+PSEiUiKDkGHMILKnvnQBFxVWZoal9
xdND8lcUw7Tbkr7l4MdYOKwqcLC45h+afktsAP94hzIsn9s3cW7L5B7Ax/ZuvZsOgW/8c6/Mo5LE
H7C5g+1u9R0mIQ/KQFtudXoDh54oI5z379S23GA86wMnZMy++Rhum2lxn348Px1NWcrGtEdXhR/I
eaQHDjClmC0/M5Nq0g4AKexKSoTMRi7LDmlDdBvmA8+bTGzAy0u6CjkoS5cOEIox0oFnpBVHPKAX
7VLbHldemN+CiehhpNZZOlJFIJLLUXCQzoOo47ao0miXV/BsGWvSPTml0Lgfyn2esQJyNlMpyFea
yoa8P9Ri+Ggqd5NiWHuzrieouCEBr+kZZG+olqr7/w9BlMZ/A9CjaucFealJewUhCpuEjSJAnrIL
K3ehGT6wrD3YfJPNb0uJwr7212YBD1EXWFxN2KYVa39sFlNxCy0f/mjapE5NENedWVJDPiOCaYhd
u2JzV/an/pdD/W6yzl8uMWTGP+VzfThRSWQwdwjTKtX/W+TxlKbLlLwYEzX5lTR/uNXtBbQ9AQJn
Z9A/I8Nb0wImyvx+IKI9pDl1wbG4wRYcnFWh3gbh7rrqRhFamhr2s/iYxiIenR8X9GYSf524AsMH
FPSNttkbRuhnCr1OWPooNEIkILUQH/IM3dntd1TO36DoFkCdlXCaIQ3VWFa29auOy0KfbRDPuR6T
XpBt5EeEEYgSviXRwhvTZCuVw5PRCMcr1/DfyorXiEZqCDE+4edMvMrOHCeQTkOj3TLgW4GF7QSF
X/N4NirqsBCoOgXxDB2OdlsWoP9TjrCJYZkIFgil/qtMVepYfe2TkUeAtvCRBckTcA3WCY+nkN2Q
X6SEwhfzTehuk5NJOfCpDZgrkxSxykdwidhkvSHpP9BC9dXDBr8ybKQzmqvF+BB33k/KDWZHGztG
MwmZ5qIZpx9w67xa/kHjMjKcnqPi2u2EJAepniGMCZZMqnMuTPiDKGqtdezFi84bYDCIaSkXKVWa
DSQjaA8h3eWz2sIiY+7yvcSLgxrrPzlrKLrvsOK8QSjFfkObyWvoS1JUIDDIB43oIc60eQvRb/UQ
deWswsUGTXDjFfVhE5wZdmu+F1SCbgl6tL7DRr4O+eFxBMZDjKhk7vBSbSqIta+eu1a/dwEESUAF
PjxVTxkvgNrSqAkngs6dzAh3hinnxy/LW4EnPl+Ts0DHhKNehqR4wP7TaGiAZWaO822BMRe6QtyO
0loPtAigkbu+h85Rl6gWkah/yHptfROveRDWuP3K5SZ72Puc7fOiGwPjrK+NdNebyV2H+MANA+k9
KgECqYeJ5UxUBXVQldj+gE8AXk2DiAqva4DkhwPwGthleq+TxoxkolUrZqy3ONQNkKq6t0YwNA6M
x9oeJ5sb9Un6WBNl7ydZlYLwnSwihz9cujDbBOvBu8+7jaUiiEo0feFNU988Bu+hXKWsWc+Z9r3N
CkxS+p6AX8zqvqPYlboWmGoIlUZpNoTKKeQ3K6f+cYIoRZlaiojHkEVtpZeZ3GSHEk6vgW3YgYXQ
//hOqfzZw+PbmDpNNA8q1QlPtlEDNmAKKV3BpagNQjN50sxHFmBz57+14m2X9FVwizzdlsn4jJ1l
eM3jU75KrrIt7tOSDmdpq8lAI/cDuSptaFFS1/2AroxxtWXznDeRu/NM6oWiTAqLiMK5rIO5OfGy
GraZckQLVvmzduViXNbaFFxDvwt9DxLPncl/cJa0sxvFWAUreAi845tmc0hUImd6UWYRWz5btboJ
GGtkAwXr2BsT/Z4RSuYxEwFre+qXuU8IuxGxXPv0oFjrLZ6LhIGkaL0vi/9cA67sBDdmL7PVetm8
WI0CQiM/P5XQC9bSsOoQR34PBjRUCYP/gC2D+eVav1kpdNo9XyymX7ySxvOSCplbhlMjXBEVS4Fm
1InQzr63ejXKVJF9wUspRCZ7NcHNtdGXrm3wLr+LhnwWna7pMM4cMpTyNzh/+kyoUvJtxEgU+zZn
IFXXrhkHq1h452bYEkfAKdj7OlBU/CAtXE/InOdyiq5qpQtaljNNRC35RICuuuochZBXTvKbuDhg
gVasHb30xtHiRXpD8A0YVhXsYU4bm7UEl6iv1USdrk4600hFokTkImYXVXEkgEosdSx9R57GojYc
s+ukKaT1Qf6lCiKKDmMv1Rn+8O9GOSN9Xm5HGl6bgcB2LkikMZQA/hleKrLAMRI7+aqjq6VK4zCJ
sgSwmMJO046jQgAtmysYYShOIfU67uKxYaYuNvzng8+9OnQvykm6uFCfoVoJtuirhKr/M+x4zG6I
wwRqyacITD7ClhlwJTpBKWwW90GurI1jDtOrB5rk8r8O1V3t/tdhNLwQ/AfR2R2hti63kXcrEXkZ
gDU7LoJK2AfDAGexZGks/3Rd2EQrJ6WQ8LB+oXyQHvsBc+nWqK/pQTKPVZ/CHmmM46mVOFfpeFbd
oDoiCxGrDgQ/UgEgXdo+UMluBP0k99SAKG0VxLc1cAIEJHuEpRfBV3ZfF0GbxMZHrCdbAxc4gGrN
kbeLQyosbF3RbSEdAZy4883SNDZCpy+7X4NXF4tIq3ZrbgY6qN6WQBNmJfDQZJE8fYYjD68Vq88S
FUfc0FJVVTicXrP39Cl59RMBSbnu9AHsfYcb9r3a9ar4SvnkBht6+xtoQhkHGFWeQBX2Lr84s7Ri
tCBqePzi5CjxAOwx/5h41BJJilLr2wO/kQXGjIYpkMf9cGSYzUznbUuPMKJn1JYmXwfYZXeUx0GD
Qa9GVkVzIAjdDBjTFIQj+Z0Rzsu4qM1LT/zuriaXwQtXGipZzx0ErOGVfqpO7Qzmbpt7UTrLzfTZ
pUi+tUKQH1nivQwwbZitCh5g2IQz2y+JsuXKcReSZXRIbSU5lgnVAckwQfznLmBOvw0OcGSLa70H
RELOxspQvicvXk4ZQy36glTMcKEKzuDxz9VmBajhBv3rvPpqmH61lzUhF6/Xjb2tRETcPi/bXrFX
oDFjjc79MtKPMw6ljh1i97rHKsBq3M1d5Kw6FaE6Bjisogfi6XUbTNfcrt188mHLfEkiNlyLihIt
KV9BC0VJNN8Xq4RSYoGoJ6wlCm+lcBqfUBq9ckz13BkDN7Eqq7BF4ci6aTqcjgo08tKuWIGV3NP6
EGKSWdTwDITML1BcAkptWTfHIZp8a9A83H6AftoE92w9E0uFQKERCk9iB8NjBnkgTnMDRAzDz8Wo
p7BylYav64WHc0HEjSh+B/btpeaFnjPo9Y7YpxY7Pw6AOXQeCzCjfvua41fb0N3sSPyGsWgpkAD0
l7CNThwE/GXS+zIW89QVkXMLMDqdMN/6gVSqhlG18KjDr2otwz6QH/gcY544yRs+XHBMrw3a9fW/
levqRre3ph8FahDHT0DTF+Iyb9svWuvICpcX2rw8cEfc55u6UDAoRSZGrEebpBQoVO3LHmdmat/9
uM7Pe0h4FCWjPJbkDMOdI8Wsv2BTKmS9BR3PDaFieibDKKLEOe0yJRh1qdyZJQ6mn+nWNwNChPnW
dwY06vLbkPaobIXgw62Kt0thXMif2t1q2ql4/7MbL8WKM3riQ3VaQ4j4zzW9LwAwdmw3qHTF8iF6
FtNUcFpJW2v36D0Yo9igjQl9GG/52VW0X4I76p1G/loqMJH/WX8CNnO2MoWueDzOxd9FBDCeidWn
VeLDr+IHJkp0OiQSETpQ/TP1bp4AgM4RZeSKN1mquP+5QumpKlsCkLpD1HttLksc8DrE7hNlZIP4
gyh6uqWDN+NSfwZJMm4aDpfgBMuAA1i1zDua1MQiT+7WOAFXtWPHK5JQArplBtIMnnrOzHQDxQum
XLsByFcNegZtpooUC6yhyPpiQmiP6MM9nClUSowNFFFxeixSc8Y6rW7V1Wdd79XcVhhg2Cw4cRbk
6Ims6h41JOOx5v1zJ4IyER9w+imAZh0u/L4mmVO4Ne/ZYt7xWMzKuxGh+SxihwlpX0T62ikHoh4r
stOF8j+2bH9vev6KGau3otIYxXDRb7SCVHCOLfVsSHoO7RIP0gOh5sReUe2es5e/8Epk4rnN0Gst
/IxfZEV024D1ueOJrd20pZsuhqJ58TYeGk7DJEzZ0kkhCqZ+ALsaeRqHvIc8HhC7y/3Ca8vQCUDk
jLndYgY+IPZqvnojj0JICwKfYV/YIFwpF4/NPZx4UT/gE5LUm5JFTK/ShWO1t6JH2atcpoQ8jPqD
vYtRTsLgofj6zJxVxJgUBS8Pa1N0PU2N4kqt7nS6KNbFkPler9PPYbTvQwSVDP4thC6y2z5M+s9I
QnOuPrKF1dlgHRVRu+jJoe+so5e36hz5U/D7rTSkOsJjqv44dBXSuOEYVSv8FFZ/vWVzRPFws8bS
gd1AZaEI1K2Xm9Xvj6vCf5ZzOQLBddAko9fz24qk+ntEcKYgwUxCs7+d7luZDe2jil5JqPBMUwNg
rWv+EsqForcFTTyeb+nsz8Na9irV5OaWJN3HyqxXSqAvuF33qwG1JUMnGEKr+Tr/T8bHqc+JxrEf
BKFS3+xlhL1rSPrsFWinaRX/2snQ0baqpX0dyr2V/9oph5emKpg7KBestYZhyMbcuoL9wVdlq4K6
NVdFKQN/m14Mb5FwLUHQBBn1/ljEKpCAXjldu90vzwp0OqpnikR7oucbQt5tjGJM1s+2mbJhBgCs
9FzmdvOUuu0TuTuqUlgOAbkfzObrfKVIZKAPSU2cSgtpXXbN0igCHMMrigDrBf++gjkSD/531QWM
GagQkpr9sQH7ApaAnFzKnkm8bIllQQmmSM04/T9fWnsgHpuzLHkPQTyQL3gh3OxsdPr752bbGvnt
NWTb5XXyGIlzVSZzyQcX858qJLS+ErKuKbrpq2lGXD/60x9NviMRUOo4EHQiLevauU2sVD25DfaM
mOHMuN99auLqU7wBc3YJcwch6+SosuMYOBOAwOTFV4W+GAMxl5Z2ODxjivNTj8Exbkb62XdvSHfQ
qzCitVMLQZcdJ7QCFJ0WDhrWU81TI/ficPBnVZchFPy8vEH1hFxOoTjHTD0SAQeMOV9fP1rI3FfR
a9vC0tjwnqQgMRKqymLfVFCAVK/wgktj6U7aA0of0kQbie5z3s3+pn4gy3ld1GYpXiASHVKRGvig
t1wS3OtxQaXQH33n/WJlLMkRTz+lZqNf6m6axbS5ZJtpoNZWsRLwRp+qTU5V9tfKnLlwGflOdnkO
Zoz5gUH2aNlFP4UW76jpk9QzWOJrQoyXANWHzyxaBkB1k2dRH+0OqpsbbkYplTi0TUVgzRj1Khe6
vZ+MnyoU/JgV7rzwmsjNOFcZed9FG5slhjs0yVLvXU0uu/y+lggCYjc5mJptdVyq4vIA4nfwT95i
X9Pl8uAwfRTjn1+mD4lyMYiwOGoD/Focqvs3JPRlydBDOPmproaejwZlNGQP6JI/Knz05mx94SJr
JXjzdmDRqo/bk2ogbNZcc8MBVFxbHaWu4+W6WxAMTL5i4iMW6Yf5OMbKpyarsdXaNfwyfxgtodFA
rnFGP+GOsbf0DMO3vBnWIR+IM2j2CY0bDj3hUOGnFewLyl7642Ug8J+0K2yVAFHQc03oMDBkDSbR
PSBAq/fsx6TKCKkoj5fR7c8UEkEXPUt6SaArdktWbpMt4LCjh1kAmnD10CfIdB3Wy76m0nmReNab
qdT4PEVNu6BdhG1SXsoSAgninnY9GZu1BqSEPjzix4AAfxgZD0vBQ5ZdDgnB5a7KDcYoVSRk680q
Nqhl58TAZPtq9xusuaQo/BlOh47hV7ZzpmPTKtml+RUv7/bLNyA437zciKPnvqYmyCmnMMBQDsdF
M5K+tGK180cXMH+XhTAy10+TfAJxZJvYdtEQ2sF6Wq9AJX3CzdDn0js15b4ul+6+j2uKkRjjyaHE
IRfgXVlKuHeG0BSCk5E4HQkI+LeNWlKBmUIelFEpe8USc7imox1fRWLFUCM8JUvb6tuil6UtFrts
7LP5jdMEhQQO6UWi7t5yJcunGV2bIYLS0ilnp0++/id9w7e3sG+R8Lj1FzpSSO+wV+tPyk+DNaAo
8RU98mKFuUCay5/G2KZWMpVT9RvYy+6wg6GJuap2gxfg+tgXGZ43fsmR+PL5bQq3uB59LVg3edoE
PCflYzys9RBHGBUOY1RlWx1X9pqnObAl7b+pgZCB2xb57cEDOgOGuKwzDgtO/xfqsmWUMfdH+9FM
ZZMu376hkeqlZuHtBacvJclDK6+FlREBirMYGvQWJVxs0mJy1qZcm7/+U98D6lhCUw3srFZn4xJg
PGuzXDaxto2BebO/1yuYyldQAdccirt1Frtyz7QCODuCngdYwO8eyOfPRkG9fVSbCJuFNW9tAP7a
dskSURRKrBBd7DK4VaJeJmOEubgCJ7ZyAzGph4QWK/hZRqM5Z5rKT5lQFtsSjBxkFr8OTNrtismu
ANXGpjqhpzGVegExE1tZoF9fHMUYhGZEMGDH03SMAs2S09LNsvusEtynlZD+XqkqQCuCFHKGUqMs
UqgNxtTegkTqxKzYtPRBzVgGKKTZEOMHeq26JvMy2X4nMq0/SfOphMKPhXkZVgiHnvlKC5qH4A+3
cArsRvsHXkF1LzOT8auzc/cqRy17X0WE5x8DiyBndiz+PdCEfYR3YpVhGcJZn5FN7OKUgOkNbMCk
WlpudAshIeSLNAd5n4udjzcmi19uHV8h4C01eWwHqCu+aZw9xy5gznuLCaDtj14Y83akeSjTFE0n
8xVaM1YPqAeD5UWCrlw9uXirXDYz0Flsvt/YYMn+HJJtSGR5X7WtO6UzeDLFtGwapn8ydtxPhL4/
UzFUnxmKr/bTFsrgtKSqXBsex+uaLbCCZeO5HvcYSIfjeeg3t1GbaQgkwyv44A8CZKDc0r8Ugku2
iCjTvRFRLgHEsSXHLcFiTa8xRqvYn9QQ0QMQ3zUyDkOfD5nPPRBG1Sj2dXl47Vo1+TNOJJFL6Ji8
u58vPClTIbAkvxIVicv6ThgSW5lpUhiMrw4oRKatPB9kM7ju3MeDDC0m+7x5aVzTfBDBkIKeDcKa
JgBPwXaW3zZWxbAciu8fejA6esFukmsCcZ8v3UgSEecua99C6+irCOoN6tIn1HNTXNpVlsMA5k9W
xD5o8wM4d+yJbbfIqPoGt6kzQso1FyJJcqOBIcvnZY14RvfHW0cQRalYMd+5FgXRg5pSxih2Q5Zo
iWom0qagUmOqe+yUdGG6TIj4cQW6znj5dgXAlUox4PrUpEcw1z1aNfHQjQyk5QGuoLpqbNBMLbVP
qSLkUj15SORrKdJjbPWuVbmO17amtkJq8qnFSCDRe2UQgPcf05Ro4ytgzc6KMgrMSJycZraMlaQF
ZkD0TfhKuUTxwAbDdvv1rmv06P9oNEox7+OHmold0iDSTezZaD1yWs9nRUmCm92PsfbMgwS8Tj6s
QTIN9kPd9JNsU9Zg5XQ+el+dZwUQV72N8xBiVfgkt5PcOf3NtJnCMUUyBvxalLFBPDXjewBLoQXt
1jRqKR1yXCHfON9Pr3Knqa9HuKnPpt3nTFioYChrXofzPf9dJqT2EmbXd7zBwNEK7q0znWM0zg5O
T/wWFp89VlVcCDY6FJMS60CE2lKUC/GGySA13cie2Er6SS7V2GyIjVUx4Rj3V3o0o3uTeVJCDhX0
431uHEYw9Nu8aDyA8AxiDdMYO0upzcrfryvDzQe0IoAhAqOiU2FUNXM8sNvp3XXnOqoxLmQBfn+9
0rxYxvhINx4RQe13FAwQEdSA3WrK+WbdiByaUepEeXXVgP5Pe8oEs9PYcTOviW50eOhjioCnVSbT
NWeSm5JCmuJlRh1ODqcKCQdrWMeghmz9laITfkZzpl1zihaCkNZ3L8RS37p2JAOkcXCytaxoORaE
dHwfAO8BFSWBAr9hSbPAk1YWo6Icwj/9BnQu0lbnn2cQWvkEZg3h+grRr+PsZUi2vBnHtydQlcYg
Ruc+DIYd6dxsROgXDJalewK4FupyXQB/RastMw/KNQo9+HNXfGDNfZtyE+7+BOo0RMkqpFit5JeM
XlzUz97DCH8C1455KvtvolgMKPo7DF5W9wngL+1rnIbTiVAKelCBkVkRkLQLP1HUsdFZShsAlgGw
o4moqN2uFQympfOUj32OeXwC674iV9fFJectUchqZs4lzZK4c64aeTu5gMUGoKQjVmjKksQqbzFq
ntvepoYv0mETLBpwrQYaQc6WgB/rlmOtu3xEDuHo5seerxe4MdQutTjOg4XGWiABI2LgGFk8GJxb
b0VtgELgX1wtVW/1x59/iKSaKdXXELHQ5akA2hpCmQkcZI/6QcSYLNNk6HTf2O52qPxNq8hIKxl8
KBD6gg+UqCpk4yxnfn8PHFIzFlu3vRLc6wumq0GEvpZ4qSuHdj80JFuFKGFRVckH9f64VxfSy8rt
EUeuz7DjGATywerwKBWKnDZoI/AnyIqq/AAeelXfGEeCo104+Pf2uydq8/osePyio5u4mAO2A7C3
iq6i+nMNFik/ovSgV0mnK1vKHzjWrt03iqXo2K10FRU5y3eKGiLqhnicJBsz7kSz0mqX/R/hByUO
fLylWWJO3AYLteCAoQWuGvl2ne1Efla+0MEuhw0YKp5ymt+YUAYjlibI6aZoOEg7vCBi39s8/yRY
gKCu36ZTT2YoKxZwj7UuMN/1UDAPva/gb6BqzWCBwwmirUFAsn7HMtFv/huA0OdDTVcJkqKfZx+z
cBknGoDiPZiqTOVEnUJWg9zG+Uwgh26tvzWEQ0EVdr/4pygF6tOK3SfBvWz4GEIlXxSc94zJcMLp
MK5TBQLKOW4qkUoS/qW0fy6aOgMZqTnFcDAaRFsh0nAIJHCI+EKqtXLWYaMPlQaMAFPoO/eZGZT1
jyp3zdacqY7b3wZbUNgriaJ9VffNu6mR+9NTO9bvKq4fX4SNDhqPPPY+g7DMxdQY2tRL3K2AjjPH
w/rDQCNe5xpMpxTv4wAsDJzoTxKCN67uqFLHtBHYvUgbUSk7n0rrE1h9XMl3m/NLVJm316CMZbgU
hjJkAFKUBNErcxiuMjICHSlBbi0nCdxI/QV6izHG6YH3TBBOd0zvCC63MOU90jKEwDFZVHl8G/Su
/10vhY7RJzrEncRDeT3ZDx8o2HZFiy+oM5nBpGRCCEkljAA03+G9/O3wkUe83VhBJCHDvijfIeqf
0PfjkHZmSepRWa2Hd+bMc9DGchxGgQCrNibz/Rhc9n3qLa1bK+E4ogh6FbfcNI9oFrJqzqI7UI0P
2JhhemjsVev7J6kXOFzJKsp47UNYEj9i+1KNIWcSQpkAhkMY7nxY/nepserbgreQLFV+GmyOF1Be
LiIBq0eAKrYUk96Cy1Woh+5R1rYRynEcyoLIlK+bG0WlSLl38h6g/IyrSrNoyMEEvEDmL1k2bIBk
1fv73AgMpW9H9IFrij+QV8fiT0qB0AMv0+AyQ756tSz2FOp4dOS8klp3njjxKhv1a36T4HJOMDHo
xIroHImn3R491T9nbbXjKYJsAk9dKxy0YvP/jDlsvwf6D96liVnjZ/GIBQxFl47wmdi8dUGNk+ED
xS/kphGCoSxZzxH9AvouoJ6dthS1E3fgKlA6E5ipUFVkR8/NlMXQlrc77KRhnPai/6dDDC0J2x+8
lDpTo/egV43EIA7AjKHXigAF5BI8poryChy2QKL+/C6BFa/Hwz6nruFWMvRyLGG+vBBsQvAqV3ei
CO7yq1JQfIfP9fyzf0BhWNYMnsgPkNUMdY2pP/zEwbMI6aQdqWMTz6dkaAVKjrgCQovMnwiifS9P
FYUgRemuDgjuVttFLRIiTz9g5SMSex+EL9F0JRg8oHZ8Z0L3nu/r/wUs/tL4XMqRF6bc+JZvTLQ7
+win226MzcIB6YyDjFO4OBQzfIXOuIA5xxmrc0YDh/TWviDHIAbk16U/tYBQZ1M0t4RvhLXKUzLD
fBXfLgq7IYbZEGuBPCCy0ZlB5gZ5RtoqzPdPKN10vX39qepiJSc2HhI840LrRj8gYvi+XqgnqVQQ
btTC0zPSzdlQ+/RvVhTenDdkCI08hij9t9gdMbY962BmRp7GfaPFgexatc7qqMUXNzcNsJSg4wQW
0xiQL/9G6Qp/J2MURe31KI8dNIRi8EPv9mI/8J3kMVuG8DHW7i3arpWEByfvHCgi7JWZ0p974GHI
pjHFp/GfE5IM78Kg+IRiFWjX1FZGzvYr1+N95gKQ05Y5ejwNXX0Uo082IpRsTovqnr0V8yVkdBNi
NxfnfyRPNqIwFFaG78kRTBVVGsFwwKq7j1S88TNuuO2CtVZuL8gU9cFRHxtwzR0eORa0d6i6wFD8
v4ve3hhaehXKxEGjbHNVljBuKjkxaC+VRclraZFr/G2fbeN7bitYmt/scXBJi/ypuTSiKgqNV23o
6cZMxEZIL1BYmIeYztTGX2OiVWV2SqrGtyq7R5XrL1NvSmTtcwiv4KUPQak76oacPZpHAyP6t9zq
VA13JTLylno4AZrFk+l6xf0jlmh//XS3EO6hTTgp+BoRpujryGrO7qEwIdsV8eebDUE96LAveXZq
gx+MUAJxF9jXiXQDC29MUH1M6anIe+pcfKvplvjvJF/q7uG+XDk62TAuJImvAQITk8rFcn9KJYn4
elbe8SRlDVAoaJdtYrS7HdMFYTAshSwCNimPLfFjg3UiW7mGijb3uhnQgAzx7VNg1CkdtBw7iUn7
7AgZ9bisuqLvFUQN9y+U712J0Ha+b73T2ufhwZ1B3M0cYDDrxWIWduMYgoBW8LH3Joo29t7+GkNF
2LIIp/sTIjf3ZbNHqkujNi4omckcK8dLor1+AJGRotTh733Ba70EkGr2G069/7oZZPhvpShI78QZ
iP/ULdxNWIGSpLTVv6jR3GNa/B+FxxBgFJxAc076pP46HW7aRRgyrp2j3RAUa/LNXwKtuZmNzX+G
BPdYEWlJVKQhdxDPw6SkHRCglmQpZfLTCwLpnALAsuvIogZOumWOy93ud1xI7bNfHT7oHLPYfSar
8FVj9+w+P+fmz5YuBOvQsbhAkj+kkmiWWS+BWJh+a2xfwvdaZ3uD+pyGEWysYE8CEY89XMN0e6GU
LTXngz8ciXtudzC9rdzQxAXN/ja4VkTlLxkC7gEkTDU3YpRjdh3ixjq0A9UCrANGZYAHoBeimF3M
pZiLVsJDCk/8MBJiOkDI9EPZ9veRin/G2Wj0sg6+T10H5KDm3lJMsFcR2hGtxrPncVXTzFtZyoeh
/dK0wTdg4VV3Q2uF9LlziDpKAm/FjkWrKxb5O9qymNAGd/tvxUsf89UW+Itbo86/jmAfO+qA5W/M
FnV6bDfGM73iP8VTtnAl+8AxYCMszaoVKhz3GIEvnBknIPf3Pcexb/+PWIEky+cAwBke3hsdt/0v
kQtmgE6x1oOFpc0XCvf2IABewxj/w2xoesJagJo28Z/IXmmpUSDykWVoNmZlnf36ELdntD4VSKAu
Xg76b1RLODmBp/c7k7ECa6oSSfEDdpXJZ88YZYT+8Es2G1QidXbXMjPCSWdPVEgTedf+xkZ5nZ0W
F16X7469jTpwMgKmTDVOcpmsPhyNrLgA0xCSpwnThiSRS+zjwl4SDHms1uy38xmcmkLL+ORk55mk
Jt2CvA35geRMovZ0BiuhVePHkSOEkDV5rfWd4aGSMMR6AgD4HDZ09wvRzVsEctnZQcahLl+aEA4N
aueTmPsTeVXiW6lUfM5E76M5TfekVmqso4UZbxrRYa2zK4FH7aMj9GtbevwY3+gAj2T36llZ+sv5
HHH6uucHo+bwRH7N0r0DukNcw1lwP8et1JWKJUUmniO20Q+ki4mbN+KUWJ4DgMmg02UOY6rCX1Ij
qmn5G7L7cBkAJhIcLuVYQ1ScW1cFuZlhXa/La7927rBmRfhNSm1WohwkPTiV/d+qVmhYl6g0EQ7Q
f51MzfWZd6BTePEV+r2TjcECyUw2+8LGKyclWFGgP1CnIt4R5PiBciKtvEfuMyz70i7j8YdRl2gh
o1X/mFw+u5nfGM35SVEflcAkRMsQTRHLKHmXtdfqHT3BvIeCHqWvFnvIrQ+//fETplG1asKnMrO6
ECWh5OfU7GxjUdWBY911I1i40DvURblU7X2Lam4ZRnsUCSEAiI+9DqVtyKB/i1trWElpVApH9qxL
eJyJwEW0g/hwMIa1EzG6WwISaiFOrUrfpt612IDK+mXQLvFZ/ain6Jxwo61jar6CyI97rr0z+hFu
yyMJtHjm1UYk8Pxk4+UcMJHiT6iNMP7BUM7zInHDEogzee7OYi0+LG6VWepH8r5v+geeLWel0czB
6lax+4NOjG2BRyeYRnGxvKLOrISZgA/zZv5fkv4DeJXLV6PcUfUy+IcSKHxwq9taAY1qEwcIYzQW
kG3gxVrsV+mtzk8HuJPWNqUAkIuGaAkAbVauZzg9cwwPhBDIXksYypRyTuL5jW5//pS+Pnx70Gkv
vtyTUsqdYW3G/KdOcD9YkokN4lEmkv7+5l1GuaN7Ev+2haYILWriAltQRF67XLR5QVbMchG+QWLF
gHJfhMMNPFp3e2+9biat4lFLDSjTdtpmIwtWjze1+YQ17R6aKtW4pkspsL4b+9LZeEl6RGyUlpaQ
2ndYkg9EZmTPL6kYMcX26SYAX3+qNFxoy/mUMRtG0Y5lSAp+6KEpykBES45nVcHivAZvG9aGrNz1
seCx8HRCCVIaQ3wlItIQq0kwvTjAASKeXLelozlwEqWlVzMEZ3yOqndjVPKjBMe/g9gRGsfHoWfI
wjmA/ZnitgWj1RhH5qyD+g6dZrVSdSuXAxjlDC7/xPLXO2ut7YuUjmlj6FY36cpXieYlJmpYRNj4
U1I1Qwij+j6TrRh5yOmWBpnL0ZugAIlrWKZ7NfpG3AkPqtfPY+a2i5lbkhUFWweAJ8iWzqHTz9mo
hAgboBzdVFBoe1DY97xloGV4NJJBvhKVQmkx/Lm5OXDxP7+CEqQGkPyTnDn3nMTuQ2ZSxcYnojAQ
z/1TeWlzd6RWHBN/d5M3UAb/kLXpSzAkSzDLCONMlEshgXFgJs9SC4sHSBQ7vQiWwBSnv2nDhMo1
ytcpmLyENPRUemCPXsBsouF9TEI/oV14xtAr+Lwo9AHE0jmbEA4iZiKQh4Juz1iikR3j7fiA8VTs
dKISR2oa4htKorpR5hXJSwS9QBgNgONaO5rYHVEP9iKjjZrsfHJhOlB+bafOn2isR7LSqtidwsYZ
btY0T1lO0/SRSgNaoWeTZmFVZkjmrL3IQBI/tFA9IXJeOE0MXYb9PbMHLP2EKkzHLW0EkY/V0Nf0
H04Xc+AIpxdjX40agsN3xBI9JLeyFwXTURMu1Tp58wNnMIfpFclG8bpj1jmoWzpgb7ZcAnFsyZUt
NxNR5sAgedUk/hfeJmAMImnz/h9QID4gBvXX8rprde4m2LJ1l1LVy3JQ6iNryr99Ox0opzWHJPpC
grD9yltPEoXDMhHtjbnjkXgbu8cEf/mt/u1d/xIZMmHomToRNHj2rXvSksDimWnXfGT18WrDjWho
cFw5SHHibLf0tIBMKEUdySiHyUD/833EXsNO5B/z4yDZUgFyt3Cv4qBf+8h2jYu4CBxBFeQo/tu4
eaBjmFKkdaJXFSzMHCU5vNdFzit5K9kQWPmp5T1Xef9NwSUNj1cEd/djGiyhfuT4Lj15ONIAizfA
3kfkoC3m9KzrankTnm6gKDia5xMsH+RsMTWdicROCDpDWh8kRG6akwv0IJA5Ee41nV9zBTRGH5x2
ceg22o5IHzhPahUcGyQVabDcvFbFor+oy55vBK5HOvI22333PMjt1Cu02SkAIm53C0DN98CuVdxM
q2j8xwcxF45BEFWgb448g7oA3J152uLY2u604bS0YYoRPaiC2B+BMyG1sbpIj+yJmej8ypZjrium
xV4ujG9DT3HSBjyf2svJzYczVrl4IT8ggtiEbsZZk1oJXRDwCEeztL16z4oa94GtrV/XwecUS1so
cEVXsEtS91zQymCmKEPdAj+fpBfAqNZCPmWxTfkIJfNKvIC5kI1IrlJ9i14AR5QR/0Q5IxXIoBhR
xCXxGbz73Z8oe1jddPDE1QiM67v+Qn3svCXGrtIx8cUzsoPXylkmoWVuC+nwIdMAFG5La0fVIUVy
Yr7dSsVeLSgzSGwIKcApASGimZEk8W5wKLerXgikztgYbJUaeslp6DiC0N7hZFkeLXTbFFINhNaB
RW67Nvq8EVJK1eAoK+062HN7UQ4Yg4sUEHRPSqmEGXPyW95pk42kcFoBYA/craxizv7M+X2TWFGH
OehzJv4ehlPIathLLEI2zGU2Q5+8LMRnQdSP9/OieBwwxYAzJaMUEbsIKKJB02/PSZ7tnYoiX+bP
OjKd4/oI3ZGxl9LoTCl9SH6JjK5iHcdQ/0+vAIF1m3N3yyfMSyevLiUDqRgSfMtBDbO1ZvFpkWjS
zin7D8uXs+0x1NVrLqIHAfbs03OvvKySuyDul2Zb1ms5WWv6ukFARq7ZRu6QlL/+c/5+oWI0HLJn
nnd3jM4ji5qqM7SdPfBKmofNzLFtjIx9RxIl33GH27VBe/IQJy2u7HvsKjVo2nwo55KjdfniglOm
UAMzVjPGkyxOBmApr1RxwiTiWlyrrLWr10MzLwr+J3CE6VKQ6v5ucsku+3UG+wRLYu0vF32LKqkS
+S8hbF2nstE9BU1O/Q33Hl/qY9gxm2SfHwPODLp/+SK+Pkk59f7vbM8Dv5ay1udJfkNuZ7fjQ/EI
/7HZAXgeCSUvneaQlJsjfxCVBJTcaFAJjCqxMv49PW+YvC7+NHIURdBa6mwxFLFqOPyw5zbV63Dg
HPJoF3IlC50c2lYytY/SgWdiWmAENM9Ya06W8qNzcNXP94zh1PyndtD5McMTFRzZzAjZ3hzaaBbd
phzEzuLbYalhMYWzGHlhjd7ZfBLVTpp0wYC5lea6LIew6yyxgKmHHqG+L0FUqH5Duoq3ZvzsNezz
1UcXWdk7nhMgEP3svcIWE69EoyF2ASVuKhT9pGVgxvrZZ8m0kyV+IjER0ZIT+T+ZJFztTMvlhz1Y
on/YOpZ5SL5bUhUcnFPnrG/2ZFizMdNTmbw8Mp/y19RwVpby65uyBxzhxiRuySqTgYjRBRtJ3icW
4lzIdX0esMtGXLzE/uG1dfzf9/Pr2cmVlLVk2233c30HLmK9E1GdNoVxRDqmmvJ2RtKJrfnMK/kA
E1baUviYlaCO2ahH0cTS2KF3RKNKcAL/z+ifuyrc4JqmFiv/wE3CcSaprngz5h2zRNo3mphOfXo0
55co0YhjOYSDefaIj+qxoRb85uB5hxTC8HnxZbPP01KwD2LMAwggF8qCNge/FFjos17zVhtoqBTe
mV0kCapzQ/YojKQ+snFv/f6MxLRjqY7Mzf4MBFsIQKghztRhPiKWyafk00cgOqIwgD1J1Z3BfsyW
/NU/1eX0Eu1UsrpZO4VpGdvYXx2fx1Mt1+XFTtINKCHs8qNkk48XVYH3mqAQspx1HCQIl2AZEAmu
gsUIU/p0O7ydeB4K0KzPAK1rY+lcbHpS+jmhGirah9vQjDNo1Vo9+TCWbznonAnqHQUF/AGKgh1y
ejIrFAlWwUiI7wpECQ39nwzwuGnsih7xwO0YY52FRb23mnawK+Qh5wygclP8n2T4l4X54FO/qGDS
wil951nuNwuc4nAAkmQ8keJZGLUXC3WVyubTO8XasWH9lam1T5Okh2WBZb2CZt2RJmJ2xkxzswAv
AuFsGFEEtS7NzGyZVJ9cMxpdmfzGkeF+BVm7i0juI5AR2YhSRscpEAPedV7y0lwmqXfZXmBqzw3o
kfKnXASp/mP036RTcbV0bT1sbMgPpOMRaOPMKHv+hMZaZF48L/JOGcOO99leTxoXPSVlKU07LZHD
V2apgI4qKGzOoqBqGtMzHfMMXvVNLep+pqHgpcj5XbDKvRnT3BnT6W1nSKK/rikXKGwdjFHpCEwQ
OmHI4Qq5Ku62j3YmYnWU0+pLDtQ7rZh0HX40GbrAJIrl4H0qo0Qyz/RcN5mWGPXRTEZzZGlZAcpq
RZey56mtNnYCnGUtEmNF6rC2CCBUb9F7rIpZKLHivksIzZk/dy20c53OYT9rZR+0UQ2TgL9+az3q
RgKNWAl/1MZrIohGqvERRoC8cP2r2fEonRmAQaTruNfnzi1NSxZhr9HYLla7sA3vzvt2gsNBS/73
v3kIXTjnn/MmgZUOqBb4H9BinhZhooJd0vl1dIL+BNfDVVa2ojnKTAO6yDmz4AH2/qMEFP/gAQzR
zvxQhpW9tqjVEfaMG3FbaUbFX5Arjd7/uiTDxqtWy+P5+BE8kEUDjWrsnKWDFai15PrqgO4JotL5
1HlAB/XsqHIk3RX3MeH22vv9LHi3SoXSlRN14NFYC0noZ1uB83XBzZ0bBAOJT1ZlYvYVl0ScLOcW
ebHx6EQWEJD0XVOmI4QYQHj2QFuQdWSA7+rv3UXJSsMHWJQGt+ZPHGl41ZCZ4vqSXPV/BXet1Vaw
aEtHEvO3awxKcIri9jiiC/Xu1IA1icNHL4IGTmidc6JjTomNfGhZT57arizIEeYpMFI5z8wS8Okd
c2dWNUmX6eGMHp/Kf6lGl5YESRvY/cFLT6WTYQXU+7mxH0u042/Dw74p/v+7m4NA27Wlvs6skKM/
PRw/vsdK4nx/Au0gP7ISpzYiPoOUlIIxmW/ZhlFigSzzCnHYINfvk6O0Y38my5q63SXJzxnef4Lp
9hU0r5Wt8s8xfTZH3naAdTbEwCOZqqBuM+imgcGECIl98kQODKJyr5pjo+xQFbifAVx7gJiicGZa
09pAqa6eE1cZYf0y+z5FF32zirBPlO9cAzSTtrT0hb40HzzF1N8UEpdr4mldzkxTU1r8QuQEh+Pf
tMbSI8InXf2OkqUEw7D4SMg4POrVtDyU+pFaqP+Ig19/nb2W6pFc1JcRqHlu62XdWphIT0SBroIo
sMWh5wiSe1L3xa7CyBnsW6WCTrtcvcVbcxjcWUYu2q+Do9DKSUykwVrFfATrpOq1+V5vzceubHpo
lSQl+XOvOaKJws/L+Pyp3XbKWAB75XbKbFdBYDpjdj7hMDQKgfu9c3sSBSQPVa92+L5bGYd5bai3
hjLO6Hee3w7GeB/CXMSFpdA2fuyN7XIU1/mVJzzSXsuxhZdbvK8BBg3nPkbPMOXWHffd4oO5CXVq
pYGM+G9/Ppi2sfBnCRN+qLi0oKFwWUacS1Y8h1pgkficyF2p5ekcSzJ15Yx2fghECWiP+r0P6ntK
luM6alpeRWiq2NnwphDU8XlhESTykEjO9HnuXbqtMxUrUBpKxKl/DeuCa+kR2TuoxtIH1efyCsm7
oo7yRtz7GI7obcHkxCw5gPuNSEnnPkBrrR+uM2pfFailIElCtUDeSTfDoc8/7FmIAwrFR3R2rExe
36p8c7ZuZkkUoEnh14u3YU877exzHlprp8jCrXoSQNA7bF/Tr/1slCEuIQqhI963hdwuMJPfWrxg
4i6oEzbC7EhaeKgZ+ROBG5N62vfL83Yrkd4StAE3wE+boXwHddlAHciH1RvVSFFT3dRA8bgn3lqt
LhppbISTmWi+B5/nLA63/FGkfasj4SbFzAJv9fZqtu7IvTf96f5yGSTBjnut+f1gJNaaa3TI1um1
stazPu0uWveKatyKXu3wh8NtoXf25+6Ob1yQSofK7NmU2LhO3GVrI6wJCVmd2EP5DSfSTgSQMwzf
XAR9xL6a39qXMiAf6WX+v+4VyWbWSf3MuiDwq9qBzYWLp1rK9PyzfZbd0uPje+hTeya1vd6mFtrl
fOSbW9a+3VSiSJF8Bcb4uk8bMUvp1Zhx3oTsL2c3ti3jrOzDIcvCj6JYDwN2Bmo783DxEIvQ0u8V
JkgwSUwt4ZveTyAhsVQZKtfWMrsGoynaFl5K691qB9YwQDBDKQOyl59MoMWe1AOHb/f2gDlVWLbK
u09PMTEtkRv1MJyL8SZ+wZfz3UG2Ws+F618AmiUz3eZIguDcNd1Jth6b791fllHL9E6nTdZVPhdh
lZXo9d9vBNEbBePW0gYhLmcpWBPxHbSjGKDIuBbBRUX0RNd5hjXKv9xqCqlHp5HdM2XavUHBDyM6
Nk/ayMYtbtecw+nrOAtrbLpfkxF0IHA39ZBJHl472PmNZQ5WG1qaK4mPOfj3ArqmgQb6b6zlGwj6
4/PmmTvBdaTXWxl00Kd5xmAZoJtMiZpKm4wQemma1C/t0kFL1hyXI9ICqBmHbxx4KbQh8M3x9UL9
EwbUBCJ838j7galaHJkeasWsxsuWu0qrNyUXZIurPjfBdLXsgIaqXy8yOf6ZYcXRaisct3QMbbjE
PFe2NO7UFOBebQ2Dm8jhzzQ6WRqcoHEbpgXfi+cov9y9NqpcVNbszqtS9oyyeYDucnxafyKTqoLQ
TRhYynGIo5AR7q4iffnc+W+l6BeB48ZbzzYCPmicjCfD7OfEHyvo09OII0pHGJO4jA9IRLDxdDnv
89zpLl63/YOzxUEp57PWKLwqJdvZe856s/DTSww4wYuqCmvmsVn9GrfczB3krHOk44a5FRZnQJ/l
LI/ARLoXVQKFoquol6G3r/7QBYJ3iS/AKneOht87sAi7EHomNqwmWZ+nTPf6Nbms34w5H+JCOtvz
hnmNSSSF9EI4WrkhqHnIvy7y5lL2MUlzP3qWQ2q/qsoHGOnMTNOm3zbJDKbCb9MCm3cTl7WFRucA
9U9aBCba/HrvALWbO/fl3WnQOLkZe7bRHJ91lri2Z3f+aa8d4m6vUA1FNwRe03/SMU9lzbVxKtpJ
juYptso2PrQ3X/z/bi4Pb8cmeZDIRbOeYEKbC+Ze24j5S0vAEx6WJ3vyfVy1hsqMZH4jdq+QWhaV
xlOkfi0fv7N2oBlP3pJNpOFbiWD9PLciiFtM4KJgKZ7MX+BnZm2Hqr7csL9zgcgcYd3ClxQ6ACAA
gEHwETzUtjccRnupp4192wcWd6c8XIsIi+pLeY6PfeEx+GnoZ/k84LqZkRJKiBAigSnMgirv+2vq
UHkOwVNAIaGQqbCeb4lolWi+j169R1u5PTRZ7xHlFTzCvErumujWHrHc5vJZai9cuANTg9ubwIwd
xvescopYQEGJ/3tgdwAY9Ulus1XddvVt196l9nw3uM+qxmvtvuCR7SbtBjBBF1tRdAJ/ZjlsS/5X
P7+/h69VvugFPu/KJJIe5LlXRBVaJ6pBIrWAIv3pH4HtsB1LUs2QX76bi0gzhgpUAH1yEHopOuHK
hg5xoZUbc95615u6LB21T9APkCWS6Qli5uFbrsaAlCmI5IXsNBsgAAPChCSwAp00bxVBAAj0ghGq
m6hcZzKEAdi0LOaDHBzy9GlDxKF3OvLkcTa4UQiCYpI0hbv+LLkDvwOCNHZkU7+UHEr6WKAj2aiU
pddmThFronOVsSspF8P/967tEg7w5E09S8fOedzAsk9P5Xspr9iWbfnF00fJtZZUQtOFfnj+jdgz
2fpTdLfEIoCJ8jBzbvJXQAa9BsdL6ARcrXVqGPXvmsopfsmIrTO2WTDiuysnxWleN4pg67TXoI0I
zQH89a32G0UQjfgxLRLcxCLRKagd7bukFSl+MQnJ+cuYlv8aj79LCIjmX1UOsgP/tT6W6ocm010k
aB9J1nC2Hpb6tPe/9KrHHGHFavxjtZA09HjzJB7+8/Bm2uUkv6B8JffHQIpPTUhYtbtnKQtHI9oJ
lwJW4tx5ya0vhI3k52YVS8+SKKfpoNZCgfZP95fyM0dNXp4E3RVlDibrLuWHn3Z3TkjGLrwQuSdt
Dtwk8hBxj5Y6lM/D4Wz7UhNwA0/Y6KS9qiFQfC0q5ScVFuVNtnqqhBWyFGLRGWd8aHrwdw3zH68V
J4WOICuANGtboAtR+r6D2jDnuthX5SvAHKX0BiWaeOS64Bh0B24aP+Tb72MhhP2bSJ7UhHaZSiD1
vGKvt3jS+Yu+Aw4kovdFCAPwOgGkL+NlIIdFIOY1iMrTrLRTBaRxhaCgbwaVEVGiO8Mmc4gbnv2D
UGux8fXmHK1APZWUD0I2qY6iRJ4mQlcox+nT2i1uJJ0TOzRrMadXkDfORE4238/66Rpj3qJ2Pzek
MwlxpWG5oaBlQgzqNQrnrFOArvsFCfaI7CURuytL1jn/73hY7CZbZB/R/7WCL4tNq6Vrb8VHxLFa
wV/jfrvyXU8sKWJgERfOqgYxGaNg6gpXlMdh23ZouewZIKd+9z9v4XrU8iPEUoB6K43BHEeIwQnu
Ccx5POkt9dE7BQ2A81Ofa1XwCpkYbDniKC73VGdH8W37kNZ0xNXsrcwDoBhF+T9V2zKPCEgNUz1t
Y7cUQkePmeFAKI4Sc7P6+qJYh6n7hZM6Tv2E/YtfaA98KQP8zCr1BPDhQztS/R7mf/HMVPMNz9PO
sO+1Adh52svgQFY/JVQ/YvTu8vNmcr58G+0Y+idVwljCmtMBL+qY2/a9RmQCS1fHK8Po4QBBsDCw
RAH+NKcyZlnPebGhszBA16GxlXIRnffcynPLSu9wgWGN/Ws1cHvxnXZaNAItIibQrdWhVjvTv9tf
kpm5ODPeQ7YwjjVeekNhn75SOqri1tPF6+wzxIa9OxcF1DSMOwNnxUmuLmGDk+wZrnqXkiSfNWPJ
sg+RR+PWaCIqNdHfBIB4VANdA1FOjBV+JRAn+zj8xXqHzp0EPjpxuM4GpsTU2u3gDjZHNYpB1CCh
R1P/KUkoWpfS96po05eNnHIhg6F9IvPZou7LEg9w5hMUGmDNcmcYXgjCEUgii0SR1HW2JiAtRKZq
cBXGOPQttyzJaz+bAvPPeDb1kXzR/kEdcrTxobL+BPYmlZaRv+61117z0v0oGCTm7Xgq8bQmXojQ
j3GasVNUvFi6O7o9/fGWG3DrmK8XfZuxrrPyseNki9MOmEUVjdHgnebBYO2AA/CZJV9q9SC1rJPV
3eh6vCKStZBmiZ5zkoD1kda20uaq+ihbYVCojp6QV/bL+NLY5C6fgsbBeNCPIWOE+HG84Z1YnRZ3
kLKyjgDr4eTjE3Z2pcYNPEQI+C5FwxuKyWXKqwNXQdYjwFvyOYeZ0jtrTtLwyNXQ00ZdHPZ3BpNa
tQo15ew0KvC6x5ZgZD/W+y0gRsVXDghbJqoohIYw+9cANpXdae/PD/NcCuTQNXfd10+/Rd0iNDo/
7LJ9wMujYalYRRS58y+dvLBBL0+fSc5ZsPFHhTCM3sPvSWSvUZq1TfGmWCM9TYQk1B1aZOVR233D
MfyosyWxW4RYNWDtcOFamrM2FGXMpb6MPZWbU6J16j+o+rFaW9fwGYbuWatKyKa7Kili3jN6vSaz
fZq71t8Y9voMr+wogkMaYgGWYfj9qVdbKZgt1UgJv7Rh5vZiuFJgE7T/jjr7ZXkBSMhxmDKvciRW
7j1w7hqxf36JITOv16UiYF07b+aYzkXw3ftbH+X2011QIlxs+rLN84UhU9ELKhlWA3voLaUKLmcZ
pf4QDANwYmsENASqeFPbtCp5rHiCQ4JDFaDmiYV8iHS9qGKr4NajzmSoNgHuX0+/+nbhmhNUW3F2
3caLlOEieg6ga9Bs1ZgWLSUUBT3JiBAcfSsNr04r6aw3qdF4/F54Nb9FwAj78VYTzJwj516jbE4V
6gSZ6tGqmug1Z5neBP0T3yOSQYyG5q1FAGZeAZh7sFmyZS6FoNYPhkCg/LxrjJXkoFv8a8sY/ROc
LjUpAeNP8dQWSf2VF/K30LFXNILjfWFOyik9wNQBt0+spSK7073sQd+WpQNgGDllg9qvHKViyjIf
JvyaDWMjXIhZieG3DDDEtxEe6rACgwQAcBxarEe7R+N3eUG/ukFQXCfw20MYclIOTiQeybHZheJu
X18aXXIg20MFSDhsq4CCuCBlRRSbWUzJ7L8qhBdeMNYP63p6GpeVNQMAg9WCvEFO9J9duAMCOGSg
dF7VA/DyO9qHY3jmyYetKsuyMCdwn+ZikTA3g5y7iOsEl2QCj6ZWurMzOyeNE27UwLlRP/vr+Z5g
M1fgvAid/pW7Dx12KW2kAArFrLlHy8d7y32HsjvVNBQLnn8SppPcGjWdQfgOXiulpjrKqizhX2JN
UJraLrPhuW5bBKIawxO+Jv7KGVjasowbrJxvvxgYBSbe2pmv5kBenX8oFFaimj2fwBlvKE9zILBM
VC71A+am+fHhdzkYy2jg+zmxt2VbvPPruGto4FFW0ZiWyfIUOEoA6q/+7OFcn9I4uq/ctXaUmLYP
kMSLHC4nRBVdMyz1YL1gTe16MTEDOO8MAS5tSqVMEHl3zfLW+MmxwoktaCIAtI4hA0jxU/9oJn87
xFNvLZil3hzTwhx8i8SeeT7kmF1ZiEan7PDrmt01xsUGDTGTsC86iDTAjuhLNnqYOpgW/50WOBDa
muAToFBtLRI8tAmL/7G6rMCUpOke5EUsio68YTS4mY66zbRQVYanQGREup3Ry05TNrrKW/GTfzlJ
gZMN8b6DE22kLAEY1+wfDTD7asCC4/VGOa0rThXQepciTnq9eAs7qb5uMu2kMdA6y0ht8T3GNAWV
5wT4kYiWblKBcacKY8nZ+t33adWXmvseijr74mlin5A6VVDxCyTMF2KIwkr8yGNdr4Yu7JOQfVR1
TVmORSZ1L8Hy9ieN9cycNCi9xg1U2M6OBJkF8PFWFvBtthTDKPbaEnd3W2ZU87uD4zqAVkEw7Mm2
Dxi1EUWDnvCd0G3I8hcDJNDTzvCu0M7aA7/e5RJwrPwi8WEq5gpTdSlvA7usCNnu/7dfA7MMjFmg
drchP4rWAzRIZguPHQ+toisZHMHGSPY6mm7tiuHgGKivwGFE323QQQVqW1RsC8eSXCnEv5Vy0oGR
U3lgGj3yLJ3SyWBZ/lxlIMxTWHaEqKYx08yFQJm9oranVAFq0aROLRvaauMb5eklOisFHwUgSeHs
9Tv15y9e7IQepSDwmr7f/iyXgR+Hw+B80dSBD6gzyZ9DPMIMy5ZqAKYuEvgQvyE4QZxdP3ve6Qr+
w9juCds+NxLNagf0U3cH+YeEB7odZA1m6xlDg4Kdd9IQVdXapazz6E+YfbttbvF+WnuCAV6UTHu5
w7h+79T+sEdZiH7KKITmNi6Z3nnbj7485SMnGPIfI+zFHN6RLViJKbNNWhxHQxAPLZWqC/XKZLHl
1+mgGTuLAAqOsaRPJc5OW2naQlgwgQ6plvRcr4P4SgFW6rifjv3HK2SQXcxVvPWRI7F3Cl6IgjQu
fwfsbkJddIFMwxySM1MV4PVsZMonaM9VZA1Bbv21xPhpC6zqpRr2NNz/mgUGtSZgr/k5Jg7uAVUJ
qjJI6uNP1KWq1+D2CaktYHNCpt41zHlBGMo9nG8N+zVdTNh2Bxf8gtLDlypTgXDg6EhvEGQl3t95
z/a+P4RIwmGSJDtsRfCJkuX2ONnemuCGMqbpNF0sRXq75KlLgX5QxthNKNB5PzvjWfW3tbWHsLFR
QH/hrEfy0bj6EaxhSSTn2pQRPL3GR19klAOvh3eoNallCpmluSRn9Qlgbh82+QaPETNgmoops35n
2B4xji+M8trE9FgbF54LR4V1fKLFzYzyqDGbFcyhPHXYoiUun3eMzU30BsGrSF0ZrduioAr2axBs
NVc3sGxj46mCgpyPg/dvbvaQhT0V/bQBTFn692IwoUsyDRpOTzKbl0M3it4+IvXTNkQWuaAH/goB
FAT0W3V3y1DDIiZd45j89bXCVlsCqVaIOjkvjJgyCOddJVin/C+sx/VAoK84l4qwZVyeLVSTOq9g
taPuIHVA2ys0DxIrJJrudFi7CqWcQDmOv5pTqM/R3SdNdZLXtv1Sfrr8ESTLTPTxZQG1xq0qAoe5
Br33VW0Tzb7V8NmPbyrBokE3FzefVRQHHcqZM7stD1Vc2AoiJKJfHpXq/TrGMI5re/0GXTN63Mjo
TCQX4yrbCjuL5wH5DvypRXdGuDpP6i0o7e2/hN+rRVi0wsoTxUku7MRlWgAXPNRaixxlD7WN8hvz
jacWE3spu+qjKtFLcZzBjOMOQJN8LJY/Wdj8mqx6qJA68MaLLzpIWAblP9pktpHGQQhD1zJ52bSk
x0e4LT96e+MIIq8oBbm4gRiSxN1FhysgkY1ciC2Wf4uWmVmMo3/YFX4wU1EFSLT2YkFGfCtMl8zR
/iM/e91HYBK8vF5q8ihy6vwRPE8JydirB4dfPkS7g09LqE90s011iNiPa0NdvbV5ocr5NmgUp8MV
PZl3fZmuJRTggzrTk1mfMPkAvf8rcSR9aJcDR2+9DjBHwejnkj3U2fpaNdsY5a0BBVBO4DtDpnCJ
huTZdx6Ib26YWSUydRPJ0x2NmPoSxdJjGiiqojRGmRFn69wg3toL3HJgoV74C1pD+kZJ96sg5OYz
jMGtvajEGSidwdBqlQBsW6r1ibt7PvywfTRE+DudgE/4RNu4v2wQb9oF1bqX3GIVmRDp35zc5fxz
7me5AQ/gEI84JlnpbIrLJdr0cV/oThG54a+j7tP3pvVtMPd+j9xq/boGw4ecAIkG9DU7ywFo3TFT
3ISBIaquvYTsMq8y+FiaAHyZpHmOqPDIoI0dscJg88BZYdGMjViAE6M0jD5KhARJPZHlvcqtvaU4
lsrXa8AvtquW7YeguC7ju53BjFR9INc+lgQbMnXwT6pJhIlZ3VNR60IFGbTHUa/eiQoCw02XHLYF
BSDVSCcB1edE6gklkkcH4bK7Pmgv9huPRObVfxg0T5kfOQfz6ge2SDmWtrG3wiSzqZkuKSEOr6WG
YKpqpg8no9ULjnAw7rMgKJtXckB/pZULKfVqXcGlMoYkqubD5qulcNPwzcq5npPlndxMLbEpIucv
8E9UDrXHtY8us6vv3QkP75pAqYEagu/RROD2lhokv9YQ6FkevUdNW6h8L2zbDsEvRKUEzX4Jya2R
kiVx9+KWODET1ApPrLNDv8igOe8fcJ386K0RH+6uH9IR5aYP30eQVKbVlFspjN6zwvipTBeDrScx
FSavA4HiusnMfdpjf4/fRKT4uLrD1xU1b2CsvfQIq7LdHfW4ZEyZEHAVix1tcRCAyspsIKo0vUrX
t8x0JWwoRxCiMqhskZx2Z88TksdYIk/q8Z1dJ7y1uukegtDtksMis9BaiCdjMEubRNsTLvxVT+9O
QIMzofWfXxoEYkjLBTgGk39/ncn2L4jF5q4Yg73j3nh2QHBnQxPxfpEgCTCzTxrtTPN9x915tPTx
zfdKbo+mT0niTnU/ohL2xCAwNs+Js9ID95x5IDgfBPlB+zrk4FwsFiNqni848jZeWfqBz/Cu36i5
wJHGr0Rb4ykcS6DXkGDFo0qUp3oG4pDX98czedY0Uv5nVzpthQffJMEJr7pYqYOw406UB/Rp0M3x
GzwZLlZdB+SlbUDLZtpYjOrkiKFZnBWkEF/dsxzwY82Glxf0Tdf0+dZwW3mh6Cwh7mmKAKQTcqdy
hxShlDLhkm8pTCal8K0I2fILfG400TL1VpGhTCPohVrJx/RNEHkNEQS1rP9puIs/y6us+Izo147Q
H0vMS1PqpXmN02JdBMyWO507t6fNDNxo+zPUuBuO2g5Ldvu7I0kx74aJ53O8fFx9rKsVBFMcazvP
ny9p4GcEvLXvBEdxdRU9TS391/4GR9sudImtc+prouwtF+DHYTSbgLrxoWQOB6Q/cBQtuhAGl0G3
A6bbWKkAMHfZRve8GzhWaEeakwNGyJZRmtBa0FzDo8R1vcj2biQeCZHjj+m5DUU7s0rAfYya2U91
bgAssM4RmeMUqB7yhbBfSCLn9VEA4pQ3EDoedcHLb5FrISHIbxScFJ2xpiqcyE5IT/hqbOK3MPbs
+uV0UDqmG9dJoCkTQxhYKSu7/qT1/+0W3qp9VYQa2Ki2HJ0CeusIL5f8mtkhNUyRntG7JxVSJJz+
VoT3btko7U6aXJSOWY5RqloXotxYBg5ZUoe0/axrahdpBpD/gaVTY8VT2McMiXudSc9ImpGqBYX+
yO71PzyBeWuDNPTogLQHfGVlV2emQPy0MnOHR/yJbEuI4QBQMeQJTBMqO0guHB3nkutSfiZRrz44
Spv43eNINHTTjpEVfc1WMJ7OMMfBeD7LCGJPkcMa1Cp/l/MkaZ6EQT6+O2Kz0+EioskDY4179P12
mqwyLDWIHSIS1LxSR7h8wNTN7PGsKC+WzMJDrFq1Q+mE8zHRrj9X913c9Bsr9cJ+1XNORtauIkA1
ydsoBFFL/dDDeUC1aFfkQ9sVD57uf9gtAulC/RYPch87DLBoaDBLNK/rdLyYMK7lrJ7axaMe3FMu
X4e7W/Tm6xekgkehAMNoVoGO/DzfbAJRbStznHES9r+S2xQrvG1NTHzr6weygztiEoLFTDpqLncS
aGnckpXjQ/PxKEx8qwlTRIokWsCWS3pdtoVmOr8YCF/Q9DgzheajEMAZ+hg0WbSG2EdM7m1gwId7
46SoOZsSTk6IpJu7i61I32ZgtdwgAIDiBww8DDVka9fMR+rUOPnMyiU7N5q6RlILobWVmbiv7/6D
9zrZ5TslW8M7HybYvWvN7mLm4F/hQ3DREBcmdG5BhmAs+B8PqjscwsCl5Pta1iUsg7DWI4WQHGnt
mwR5t8NFuYGwey8JdaOcqCJ3FwP7bKX7oDEpEeOzuSBlNMl35WcO/CZAJ102+o62tuO24BFpHtFf
NhBG7vKaUrCzs7mdKFER3san2VQaXfhU06FKwmkDYNRDZduQxqe4iVNnDWo2c+khMSM1Ng9Z3uGU
19wbKnaFR2jIRYbi1SG3HQb/j1VY0L0hXwGTl+CUG+FJjXb3FXwULiMjA2r5OKzEVrHrTMn59b/p
u8wn4p0emhnRfaHbZYr6e0kRSx0bkU+8yE25UTdmTozEySieytzQrgUR1AB1L7KSJYS/wxihZi5b
KJF/fY6Euv6p88j+5qPud+8FBsBL5fIDF2ZSSfufQH7Hb8Mv3DNdTb/o3zf2owIa9AnIm6q0A1lO
fGVLdmNcQSfESPF6ea8e5AiH1CN6KNbGQw3Wklk/qsbaTLLTUuLHNsNV2HeJ5BNU/k21EVv6dX0+
9laF2i1WyqL3A3DC36+Cv7wEyPPpbSj7MqJCSj0OTl50hEBJH+Xui7NzCKIXa6OuJYwh6rAXwDjR
/Zz/eZNNqQR9YMHTEkfpfm3mhRsyh3ipvpZeqZwETwICpIaIco9SzQ5LRKjR3wuQnmkNkBe1UmXH
js5/hOg/OXX/MjDxYV2qm95xhUNSxRoRDRG1TB+fEdry6+Bs27rWoPBa4B0yzou1dKgjIjv7okUR
md5KGOJ1VynMEpTI5K+FLzkQRRN55nE+J9XRGO+hSCX0nos3V97nE7SK51ofiNsQEgUtvdGnGnVB
UWpnhE/m3CGtVnlK+O7h5FIq+TVsjj6ZxAcVkEE1FvzFFalxFEWukSI1oB9T43HYyvwDHhAgOf8G
7Vm9s7dokvknnyvhCJY+4G2JEnnP31iy6ckbeDncMGU0w2qylTVSD1eDBybQCoPvCUDpmKpD7fag
RyLr+wcdymgRbGK79CNjXZ+5NOkNSAbya66WADBwBQ+wcrBjWmdd1fk6vOPeC2Hb2XtFYDFegdjX
Q+lSvTZ8sU/Ovarl6m3vthUh3mtotrx/Jw/ZjhGmuYLoX8i8/CdRi4BtCwMExm4zBLbCbmsD7mQi
qtg1P7ZPRsW4z91o3h6YSRadT0LiVvh/xNQq3xGeHB0VDmPH8lJgDEIeGoo4s78184ViD8hU+ihJ
BEnocdHUgOlCYLDbOqZPWaDC00wzmzTu/f1+HIWYKm+q7T/FOpY+8d6ZYZcMb2YEWGyMfFzZMZe1
e3tpYHl+lHUtqwFzPXSu7WoFAbZos4/GDqyry2VAXY42Zirejg1peu+EmF1sdnZ+It25VBhlKhAP
Z2t1dX4RB6uNGgIxcYuU9M3BhrYeogLJbFyvgD+hnIG8qo53EdW9gmjvdToFpXt4uZ6rOseqjO+D
xaiBld6dvKEbyIvhBhgagc630vc5rXLfzNIDeMloJtcH61m3vBvGgy94bPjbqGEEPcCXJjLFseyk
DAzz2/sLiuZb41+TyTzzl/gZzk9TaHq7nN2epZ1hjwODNswj8hjKaDH6jXKDN/1oQFcQoM4490Gx
mR4BWD638E2pmTXqgVh74ZrZlw0THf3J/ZFMdFKS8ff87qBQwSiyHXDaA+6+vvJQMS3t75G73kiN
J5gS9tdZUOroPYv6THcUTjZ62zKvKMnMnraS98EcQ2m9hOOzY1qSEroSzr5FLiPaLB0ITBoc/aMi
zldxcu4rqEDkb2Coc9yuCLv/ej1tWgZZVtgdzytysNX86VC9TgQTNSckVojJGSjAVdtrNWtR20u5
o3AlXuh5y3mwSKtdQ4uclpnIQKoH1yqtwHQ+/IIKsPsAfyM/e9aB6X6zPX9C+QRCZaKJLeCnxbEg
qof/+h1LGy8BfCl20I/lDtq5Crem0zbRaQ0QmLH+ua+nwAja+yqLeP//SwAqmv8Gxs1BRavU0/0S
t8iwZ7ubvi5v7xQq/+va24p6/Td+j9FHu4z95rwsSPRbG6SZaUieXXavJ2gTPu6fNZI2XkSAhk3+
O2jyXB6SpPHeNr2SScmgdpb++Ova5k2g3R9228WhSKj415onDImm96GB6S0gZVL1M//iV+8HHdwu
oVaGFccjMIhhMeX/P0ad1ebMhQ479ILhJTiVnnQwT8fc7Jka2zKY6rXczY7sjcLiucbYg7zIBUzw
kNk3Ms4UgXyJUW1JAeEGPs4gredAVreS/WZd+C/pVktn1EUmBNIbEdMcqkqe8qtzmj3GwJ/2HYCL
aWDp4cEFwESlIxiQoCj8489mOaE69zqVqVaNuWBsl1iakYg5N/+Q3fnB0uMcQ+fsKG0+0oC3cpgU
YNBl2oqaojx5uxKv/q09m+RPzCBPVSzV5C/tuvCmBvJ7g5EuU0KWNBckUBwapSHxOzcTZWwaViQx
W/jnBaoBF0+u8ey1S6tsB3K/mBQ7PXvL2In69ed6PTT0pel/KuQjn3fnVER99Af7wDoQD6JgCjlX
i1WcJ7jHoKZd4658u4B0DvHIxcBdkm5KnlvTwk+fZvejNiAgIhKsfFOdH1xlz5oI89om9jGCm51v
roolWNoLDFQhXdfjkraqMwiQ2X8zpRXbSiYHMoP+FijaN+/wFQwseGi5XRr6CzAMmsEEOcsslWHb
98yjTQOrAIVd3nHepqYfp9yrkG04VpjmSCwRRp7n1csZsbw0p2VIb/kqaWFcHMNJoz9bjfV2EfhP
CtBN16doD+HPYl7aDjCEhhaX2mov0Ln8/DGq/48rvHfUKJstMWkqsXzEV+6w3XJqCW9PjnxIoeNl
kr0lP4kU773rQEYzdJ3v0bF/xLSHeqM9X18YrRDdNE2FKr+WQZd+HKoBiPYM1zpqgiGOMIn3KhIh
Txc5/z//eP1bSEUnFr6mFk1DrGT+H08ypXTmsmPlgv1vCCTR3pWVNP7kC+RJdhmyxgGBhJB9Ze0B
dXyy71jEk28WbxzYBHLrdvij96BcOOWdpyUhtsz2/CV0hvM28oZJXqG/qSxRV0G/cmCdrU08EzBQ
eiM4ZdWDJVca7k1BPWRIcKSE0fPYJZ5/QlB66asBxM7egU2aeXLCD6B99YhamTRCjNgylXg+meur
P0jsPNBUsNbV0WkAgdh5CGVTud0hX4t9ngCfEu1oAfQQC7fr0Ij8zNhYd81Doxm9+QQF63puVa3V
EsGxiVqef59WsvbtNQ9HsnwPfiqnKfNxxdIIFduq8bZc6/XsbQ8z8cnGp7UMwLNrFxA8TJnKUpFZ
JyVLNk6+3UQ8we08BsPGyrfxWW3jcsRWZCC1Uhgtnv1+hKEYvVKje+mlio5UHms0fbzpvBwec9nA
BJVgpHIihi+wMLa0pMLx/RRGtUUB0Nl/hOZEwRgPY5DufNSJWaF5HQ9oYaP2isEk0AC5Ct8wXgpS
CsH3NRCJsbYCVTfsF9sVGjZXqez+PQo/WHxkzad5H34OQ4y7zOD8pTBsq4hTLD31yyTeW0F5cXoX
nleaQLR39DTaqB0vyxBiEwIKaU/UYFWkHErX2pEciR1vjPTdG7z4qMvnLPxR5SNcb0PpTRoHpxyC
FUaBHy83Qj3nXcB9R++MxEsu6O/sPWvhC41yVkUrIFSoj2QqEp5Ea94ttSj7VI6/1CP7tEpzhIp+
T4hjt3rnOx6uOOhO47bDn0ofZmiGrezLyT8Xt7shuqM3kv42FTWOK+3TgqYv8/4xnzEuAPP/7mOd
rgqXJLQ6KZTih8I7QX2G8zaPd4umPhzmipf4bNIeqEX/WaReTz2x0vjD+iUzWIsgGDXcDLZemR7K
G24X3T4Tfv8uSYU0rhgH9Ysewx2YQBVbRHGQxkro6WtVsAwcM5o4i5f8+EgR0m52l8T+8sLiRpiV
A3g9b61dHHvGtuP2Rq2E/TKSa5wQbeui7tu8PQOiADCdO8JjAVKBae/clh/PfdrIXmU98a5dlkt4
gEgeFOEY4T/MTrei8Tt8Sj8y+Q/f/kxi/yuYPz4/w/uaKzxWkn9/CoQQETN+VqrQX43wXQtW5v7O
o8KpNUMwZ8EXV/w1GSMkfoUvAhB/7oSzJd6mKVi8F9rwMoIRhr1yWNSbRhSqQSuMXKooI2mUehdf
4hRFQUCe1CVL3+Ungbuxert+BcS4Zh4/SFAc/aMXw2MpZKekrt/066kQZ5zS1MJ4SzAhfd3MY9kN
5uuPo1dig+ixpA/hBoBq4x+paBrRolaxI8/EAxYRQp4EuPPF+uLXDZTvA1yf53C96dvZ/Njz+lX9
x0g1QX9xiOLYsdhUY3nLxv0EtW1akIw3sEUmQsoeoJvf3BIFsANfsfkdiKjn1oSBl3rw8KeR1ufX
bjFIXM9RlbrN31xTAiBoWPpdafnZBbG+UMaubd4Lu65Pbd/mCBQXvozBwjOf+lz2zDcNRXahIZWW
bKHS/uIUDgihlvmWvZptuwy0EJ974wzeXGVWTv0RnMtF8CMrApD0adWHz/GPKThWEsONHj9Dem8l
PDhtsxvKyefQKGzH+bzDvLCTN0r94Ivqx05iqo+SrF7fGT4tLB65Ukt/jUFgPHi8I3kxyl4PcByu
Vqh567rtDge4Bjwo/4vZ6oIDKr+fDdhJ/GfppOPhiaScGCkXJfRWHxqSnkmNqnM5gZs1rDP5XnMo
h6udYkxeCA6e8jeAPpPjhh2E6afYo+O4l+0dxvUv658QFZJCB/VJxst9SyAieJXh3szdyWmiN6zg
NW6OH2SSvjK9+kw15o+++IEY36MO45166quBTc46g9k+PQuJiRj7hoklq3Ut2/ZspfG9U2x0MJHs
3jMraGc3SXSJ8qW5eqd/brZQ20y6e0LU6f0MGBDz7zVsIIIknlIqBd0wEgjpE7kvvV5eokn47iy7
wJAV+C5VuuD06yuqUszBcZPWQ8Tg2C81ON51TAV1JmKB0gmDtWmxLXaL43n5PigGZ0OK0ApwKpC2
2l0HuEkhtIkiUWVfYOCBXom6vtCy1bfDdYmIu6YxiHXjaWHgZofF6K05DcvcXEaCZ90SchZcwsQF
b9QST8vC8guaAtKGymobimOsvCge7/BJ7EF4xq5FsOd3V1AQbw8pdn6vDOMdO+ESS2X/jMX++Inq
iq08p3OEqAH19uUYOz7NCNo02BLE0AAKGnk43OFMsBFdLq+HBdcny6iBb3zRkYJGFlM0w8AQ7/ER
o+f06/Ob0EOOGIfyNNwnjQ+H2WHojwWOywFV58vCCIKUvOlPfoaksgVMXlB1yw4Omk57l5rf630n
+X7imJ0dc90dWQoTh/GrBGwpAXXHlbzed9zeNUVC1nPu+bTqSDXrZMq2vuxnGuxIo+YndWCPwbum
dnoJjLetpwC8Qisdbc+hwjrmtzY+r2aHbGMotP7w5ScHt28WwEd1I7VX2USRw8V1atBzHrbEtr6j
KVHRGZWrx6l9L7Xz2QXluRhUCoj+DWQmPtMK4pT9DuOakvvd2VibRvxubOD5vHgSblMUB8ZtteFj
W/ZPTqaTR03Fv4xh0BbYKhuLS97ehBdZ+kI29g3hsZK2PtrqZ4c1cSEm83iSGJ9lmHs4yU2o65nA
4xWN5dGgYzGJTWhO/oPOLKDxzUj2irKzLMJ+ZRT5gqSPa3CtoxRDRrfUa3SzYb9D6T9+riZ529c+
c4FPpdgvggOqiPaWAMRvkxp945HS1jAU/295M7W/9/Gjlto6YD6ceav1/Vc5sOVy4pD1J/kPjPGV
dw8XC6v20NA+r/8b1CVgu27JUSPgYiMgkxYeIdIqjZ4vA2myrNtvUIVUyrJ9ibjD+usBfVjpC+3t
CZnvnOMGR9qUuSNE1jufePvs4hwyjrFECSrz4B32ztCeAwsUL2HAq0e0+Oatz4TH+2Sd8B0Qjox6
UlrccWZNBxKu+lOXHrwgJnriSj0vy/UPBRwIzCe3bNY+xi5TLf8z7hZbqetPem0jGj1kNF7l29/f
G6I5LTq5xM9vWh64gAXdSBlvp9LMFj/FgVCcyZJZ+nRfNZxtBg+IMnhSSXAhZS8oPUGmN35jIjCQ
zt/T5vbHi/2k8VBi7SzmDdys2MTWpvzv2nAH/cIZaSCXESzbeERlnLU4l4ZRAzMDCU9PklFsmQxW
hjDMIx1rjtHPQTzenKtC3aRGyRyioNOVimTtVXNnZlLC08qelTWMjMAw26N2RoKMKIXEq9jvNDPA
L6ysqCIhNLIja4iTh1bZzq7p7KczgscUaGN/hJKwmBcIPNQB9kzAPb0LPfOMXl8MLGyz7zouWP8h
mBj0fGTHQhA0zZ6/Ny3w0HarEvfGDuFpn9s5JgiS/aYiKSVPP1jAH9iOZUOTi5A6NTfcYZFQHDzU
FgRMZrZtV34vjP+iusB3ZYjsgQND58KZT5PCui4utygA0Tt3+ZR/gLrBwB0MMfHU1qn8isKLPSHB
GJWzg6LZL20JRCvDHf9g5dg+B+eq1rU+m018NGvs0g7tGSdw2//Wqigx0VmBH63L8HBglvFDOF27
hX3x3G3g5wAOX5X46QhzQaSs1X+wsUHX4lxZtI0cGwiHncrwpl9yjVs2LmuUS1TuqDDI4M8qgzKv
mjJ51O9XrGIky7MLbbsK01ZwraSpQwjXPXbndbc6TCxCww/7brBFVovP1/El64ug9jlaitH9m6/K
QdJ3qR4CzatumUyuFTMUd+klz98+tmbmBqAJ4AoMXO9ZdPzgUqpySdxkK7bzQt6Sc1NNp6VxYg+z
oKTwH9PKR0m4FbJjZOVNA2sgYbiYOgR/N9d9/QFUhvwGZp3yExEOLzvG34Z9gLwn3MMaR3ptYlQC
NbSbpLKiFpJvxOO4NHNaXl8oe09VC0LDVHcyvXixvjEMKlgDD9FrXhX5iKKN7ZBXWEaf0D+fyUkB
FEPlxGNTOuUEZZhXF4HBcFqT5VJ3g24poOZiZMHRm3Lul7+m2nxsGfh3rjEH3H0F0j2xaSR5cy8X
8m7i0utaLQ+2QeCaxG16K31l/FAX2WS6KTv58q2muHe5KHz5OmdRIgl2Qh9gNtYp8niPLj6WaPI7
UI5vzYWJHRH/Ou0rWzNNwWdTvY1NBIbviWCk7IqhKoTi8LyQR+VOdWEs9N7NbBz9HqinAID/Rfid
oLO8cM+g40bSBSeWv91D5Pd/DN8PkR8BcED+zoz9DbHW0AXJTfheBJ2xSLqRux9s77dMIQR4GY14
ddTVU4bWjMbPrCtTcOfBBkQIUj4tw1h81++IrR+E/0uAcS2ioy9pV5JFKB6Dc1xnVYZjq25PP4hp
pXwS5hVQSU0qBz4Ite4h0agee5TsvKiUfvpfqea6zAF13CZCgMm6EqDOPsAjjfb+L88tF3esLnKE
zwu+/39eoIFHY13ukl7ya//Ytf+xFBSHH4wCLySyoWfnG53heSrVyg+Ejs6soFSurTxyDQcEG0lI
Z6gbW2tOW057gic7RlVGjbFODbR+BJO2zCkJVIivK7SKC1j8pRhAdV0phQ0PlaV+T+QrL+Py8FP1
0BiKniRNHNWQdrD/BLNcgkSUrTzY6KVpRweve+ixM5f0VF5ZQ+Z7w1qd4tcXV+wop/G4fz6pw/aN
+S2xBlbMauHXIMWXe4zRZAP+vDq1zNpx8H5xXjve4AlDxHMWo4TGh04oVEHg00ZWqNt9gQQ9oskD
jqLexRbyMfUaZlo4lXnQvOBMqC6zlVylC38Jt2me2gpP3qck5imepu9b/me/YmSq8U6EPKu1tBEW
yHV88aUGsgM9S1/P4tq26zx3RUXDTvW7cij4huUIeE6lOn8iHNjZ+uWEwEKvR1I/HoxzQR5VfqaY
TLp/Fnos82UPfFcvTTDlYMlg4PWwV8yCPlHcPk3wUOOCNBX+c/yjaxpYpZrnX19qDkEacLlJ3w+6
3wF2GgqJoR8I9i+0CxqzMSQAgDQqld5pO+aN7W+SnWoG9hnMyxs7DX//0CzdiIWj3yUX1aJhhK97
fnL93229RYDwUGMKR3YrKCtMCtqSP5ql4AU7iw4HbjIqOtVYwagEjWKf9UapO71mHVkWzRLFqPad
KgjsX5o4PK+KgRrCz9koZ/s/s8T7po2rcZRsivfxSJ65wwaJueMyj+YyLJMAS+j/6E7DdMeQ2dCV
CcayESM8DxkOd9R/9t8BJIz5kaYQ/CsZMAV1Y8w87CZ8X0Xq9e5sFlUD7CSn0Q0B3U2Nztz+DWHx
41ffvaoNpmP0PHhy+HEDlNzDgS9iXiPerGQbTCSrr/xU4CCVElGIFvpmOwunwCHrhx4AXvNNbKb2
IC9JXYINuw2lH/YTj48xhyQ/oX05SVQ0K3sPn7eUm0DAuNkjKvuy6JMv+jnTQhS+OVHgZdukqJ47
pK8veo+H+hFxLjufWiCRxx9U/Q/Y+yxW4nbAlsxQSKyHQhsKlQR2VDXwSFowq9wUjP/o1xoUs6rH
GdNI52CzwJLFxWRZARsnqZss5C1w5/WJUCmt5Pp7qNiNG5igSQBCQsO/9U54jDNC3ZaggCZoa67D
EZDKT4H1HjN0x5Dgw2KDwPPYeygfq89QpooVkELl7LgzNoapgZM29saDHA03PmtyCE3a3iqEwAFD
CEBvwH3ohYsxVjUgR2cwHryDcOjXavk7z4wLrkvBklbAO6JvLJAn3Bxunw/LcICVTzrkr/Gi2eZb
4jfICmXTTbSjreIYyFY3HLvG74d7dBPVSfeZH3OXLUUmfJ4xJRD/gLJ//vh0eWm2XWI2E3UVFJ26
4ByaPqPjX2XMljD+c4akeKFU+QBaLEcgmVRCOlHM9EO9EjhpsW8oFj4ITm6ih6+U7aVW7BVrIE/P
aQQlmeaNoCOGxqi35T6HdZ3mavGxzZlrkvzOYG0zL/FPaUofHmqEMZCnvj9+3JVXCl0BQ5KRi1Ns
1eGt9BxUDTPzktEWRLZTIJEWKMNm9Ya6AAs0sA1tS+8fgjXv+RRyn9RTPTNQEUSWgOyiVbyWR82K
qZZFninEFPGz5hR81vUFDrRgSNZT7SL5Cgr7p232p9k6bdQI9XgYwWYvLnkW+cUG+VqArSRJwooe
H1KwZMllFXIx0bG/maOYJsGurYCuLisaHoNRzO/c57JZKqNpZy7/soOQKMXQuR0s5Yrl6JFcEX3J
WtvZMTMdbMMtYTD+8CkZ/ebiehyN7YPdWQtBXf4aU18lpV3H6xdNuT3kRKOO3RJRxTnjvsHajKsD
YZOQHoeIAyPigZ2Q+nUS4C8BEzcQF2eNBQ39YvNPAoIoqIjv09FzwHWt9IzJFHlbo3FmC39Olyjw
N1OQRdeT0No3wBaNOdqTAq1rQCTUAw+zFrjYep4xXK/o2L8/EnUGkHTMQ+9/zctyQ4q/3VZcqnVD
w2bsQFy9n8aInJ7VCwzvQpD3cCoFyFT8ZXiQ05i5U7I8zpXy5o4xAymZ/ma5mvvxaVlfY6xJ2uqs
opkP+/HbPs5MsOe1/TrEwl3vogyXatPNjEvPxUEeED0ZON84Gfq/rXYJH331rJ0pPaZkCCTJnBNV
a69G3X88DKYa+xm4KxaCFMBb7mijh77SOgAx7d01jsul9XpPbACVSck5LFYKgukbLc+CwvL7w6dP
A8BbuzdhO4mRu2WkmPAqnFg9fjWn8SymopSUmlNa4so8Jp83TxMeImg5/b0GLo0XvNEqVnq7ZG6b
KVY7Qqn+1wH7Ha8SdCfjCqqHc87jdZ6LIVp2i8KiH+aXIIhJpfICgbqnb/wTJ6os/qxW8hZEWzJ9
3SpOeL0VHfo2eLMZ7Lxhpz4cl5b3QdfWJ8iPPtJ4J/8/0z+S5BarW37zU0q+udgvU5uw3KWfhd/Z
jgNZdMVxTIUBKNKQSF+8t2gI/OV8qW6d9PClwsQ9pa2I3Ksxavygs9fDsfg6IkvZhHhc8zAFImvx
o3XGsg/tS33AkrAHm0tLAENhfTWwk40o2/QOt/KQrlFD8wqwuvviAsFU+SfeIA9r7abWsW9LwlEg
Qt3iFYPMK1MXWjfp0v1BNhM7juJ51NEob8+ROVDd4LZOXf1lVo/6qlFwM160jJDpFoDEtGVhiMYf
hgmfPNYYy7OLfmR/jqUXZw8o52a3JcwsXPLXAq+bO1ivm5IXNIOqN3CKukFT/Po9YtUGC4UdH+cQ
YC21VvGOuF1I4EAIOjX2yxNJMfkJsKq/44OyqOzVxIbREZ048BGLCEAYhfMfIwp9MATGWpWQipt5
IxbpH4qNnlD8329XBjlxGS8cheBWlfvEkfyFXmAEYDDTIPpdHWK9Ps+om/ZsplKc7USUU2o00FhN
H23vQq42fkZTs/iPrRtVBbR/G77RQoV0hucx738kMI23grcuBNA9YBRBF9u4bbIvv/XlTZicoz2i
GY4jSa/WExp28+HnlnBpcgYLj1sVIVAik+9zM8Ty6XL08KPUHfTwhm4HeY4/cGzWuD/HBVZ2Gqsm
sI7gfmZUJmRYoR+LXGZbPTLYAQ31jW27wBfQHPm/MXWlZg7oXg8gIs4MYpeesCSIHIJeOqCkn1Jj
yTXE2DWzPTYHPDHYWJ7jq1rK4ehCItJNISkatZuq2/88H+1y/D5PVFmkfw00KpjurJC0Hbm5TGm7
VRY1DBo9ry0abkvX/tEKAQxcMyxg6Q+zovF2sVjYbXGMZuH0/pW8e8oDSB2AOsmRBU3dz9HTHSpz
s3/JcLBjCnvTQxKCd384mVT4eLXAqhpxNsY6i6UfWcu8Z1TpN8JZgMKsq3HR/oJbly4BzxzPplKz
HspNXNZKVkenBPTVlWwnhU5FgLuvotrKaLga0tgoMuxt5Twt11QHORlHlRE7BIZ6+YXUU0sEXyqq
iUYAaYli6rq/WLOd2wxo2Sd1QRbedWhCyrw6ST8JA4jAYdMYaVKPBEUlBb2i3L/7+wdKtka38bte
YJtqHc5TRfYIK72HORo/s3TEsQzESSZuJbsYMz+WUSNZwf4xkKikfrwhfHENkRS6snfH8DaZDOXZ
G8INhCYHOAOhDO9rjzi0pT8HPUS9njiqJpLwghP0CTkS1i7pDThEQqwuMhM0e6Ui3YthE3BAKekB
WGa+z7hLWsxgt8PwMJJQ7P0bpqD6oLlgM3QY6+uuWwv+qsHkDehcSc38wXx+ExvM7stETS1sY1FZ
/xMLfMzSmfVwpwh42jUCfokIjjpJbQV0NEvPq+93kq06vPA81w+Gt15ZNuqCTgeA128XyxQkr6AC
HHPpd1AFjkNuKH3ePwG85EINduIH1eownyN4fX+qSYE0qbTzAovwC4X9faHz5FxaQE0n+KynMjMf
3LA01mCsWySsYdFWnhnCAtwkfIVhfb34WqTleKzOaF1lHzuy7CVE9t9F6aTIpv/e77UC9AbnICrP
Qcyy4YTpLtphfZ2o8esUbviiUvDs3PXHZPLo4z9wt8tlizWM3mpV8zBqFnP0mgyRmeMYFl6zCvsf
b4ZL5Cz2M4d0vFDTZYmVBu2q3lGScKyjYdUK8MCWjCHc4lCosxeljQOeHd1xBK+bFJ5XZR6UhQhX
kv/79TBcC06Qh/I5mA5H7gbruf+0jyjVvQfAu1utrsc7gH6BWhLA37Y40InRwGpRT/R9IP0cTnog
wXX/WNc95OChjm9ki1dlOuhhXg7+pRkWgwgM8jpUB4F8TAILWbYcrZrnN2Vvby6S7TvRSY2q9Awc
w+ea2f4pod0EgRzWByf1N5Jgy4sjjy5DmO7rkC1aC2F0LB6R9qlfCBKQmzaYFP0X1X9tK/sfpvTq
odddmZ7cudatIokUwL74VAgcyxbG2Nj5r+O89FUC97iE1BMDDDrrG9c84sUD2NsO+KDQJCkCiXij
G/6BIJ4Q5Bzz/zc+ltJ5A3mQqqd614izWK3MLhKkAJF9X66wCfxsea982EPnNCB++fKfS9e2OKr7
yHVHk4k2OELudp/fnKc2NHEfl2QejYu7lI20RJBYLsATSHLRYhDBcTRM7DXZ+J05jYPdI6mSd3w7
yq7eiTEQpyn0/eAeruolHMSvWWVBcUMK2Lf4X73pbQVtcv8h/u+EhXivxo0fwEyvEXVMzybyOBwM
sUzb0rxCqurOgAcbTdsxJgfiqIaM5C48Ye4JDtEnDH1H/BAJd61A4aa77AWyvf+DvKsu3sMs4qOv
UEZTFk+6Slg6I0fbyMUiadV5E5midnMw2QJ6ifC83R89b3qFYJ9lucK9Tauh1zqQi9olYVbv3SzC
ZjuBegzHkNOQNSEJJ35GJhcCglCJ9OyA7PuTLw/9sVk9vCMbU86nQNVpzt51xWCRenjau4H7mIln
UyYCrCLmLwsgH5mVgVJfsrjTGpUHvx5sSm65HXgFwnBjYrSze8cZnG/EeOafuJZ6yV+v/Pa+o2vZ
zA8NUnLFTKQZqmzS1hIG7cNJ9pl0gfvml1bEuFQeCdTSO/EZZay3pySWCT8MuhZ4EEB5i6nA73je
HSgtSDMwNaSqsTTas3qnfpCOY643f+kB/RtyKTMKxHaVL+HExjXmdJvswEX3rYHDhcHqCpvY3LqN
HvpLdb28TvLenrBVi5WagEOR3XNSbOySYDSZEhtbiUDOKCujbO8S1YS5AzOt329kYrE0uo4CBm8n
bCuYMOVbVWuDf0zzLO8lL8B2pw2JpEDir+i84WTbs0gvzTzIFICJkO0YYytmtp7iEwwWHt80MNcV
gYN0XLP1jLmB7j0CVgVJJXWTQecyjlt5A2VejzE0lbEaN7cqdhnCoNKS23MHniHvi1otXkf5H/wS
/OEiqZ3ZZU7mScurcKnGj/bBZF6a9bISmbL8pF0WfmtNHElm4PaAaUdQU6imnOYWcpZFhxPdqNXO
QatC1/uopZQWv3krgQKfu/qYG28YTKsURmV9G0se2EX7sKM4mh6JXZ27iX9y/dvdTe4DlsYgzvHO
7/8/Fs84qD4JL04AWVwFgNH+f4HucHGP8sP0NlruZqfLfbJ/L/Y/a1jphsO8ph96QXOp4nGfGBxr
vjLPMtOGH67wBqnqgF2CzUIg/U4yjB6XC/6oq9sje67JBlYn4tJRIuoTI4q78Qi6agrWjEfSdg4/
wb6jghPKB12KOkzdSw45DESiSMzM3O85SOKqv1QdnbcogWDQ0Yg+PDNNa3PaM2SKI6em6ByA3fwJ
m4W2PcCtPj5K+s+usk+HDmTtIJklBSoGocVSsu5YaZJEbVhwIgZ7CCdzQAjopFo33Zgm5hru6lXf
yKC0EZqAzr/2T9EGg97zGx6vn9wNF3JlmqoDB6LerHapzEq2B6bRbYkbf5tpB9rGhG41CfY/uJ6K
WCvNPJt2ZeC2RKxa/p8dQU6BPniAWKj+OK0LJ2lqpBnazC6ReF0NDeoZPdMc0dLbPX5gxfu4A7M3
hHsWsotyXC1S0A3kEzPAsnWKF5/z8tDldb+1kSk/T3XGZNtS35/tgpfygu4Mzr0q1JfPHPJ0AUSM
zuV3UzWjPKWaIZUnWaPGjTZpQXncdqmABluAOjzgp4huKJcRer88PmAPlKR4GGFrR9QVJA3EXW0k
i6mVuW5O91JA/iFnXuUvY98KVL74v3ImTooz7mAfPJBS0QN8zIOgkF7GLAoRk9wBUNkM2F0BQUEn
Hmxk0haS4niXIkZRbGmXdYaXSpmJdoCbRKzZKqvD4k+U8zZQ9K/dunBEF4jXnwMkmuaveCzz+oO9
bt9bflibaDS7UUPNmvpLtWCSI3hbmaxP19kJrVvSKHTyjCzU60i9FgUy4Daf/LWJmC728QdMVTJD
7e/suZeicfkHFkMSaugnhLOSp8jURrSUfXfqwK9dSVeJVZfHvfJHkAd7ZkaVOptmBUhlvl2Q8Uh/
SikNAxLujWyAKxl00zgMZIgbevyyiVWbj7Zky8DfQgiq4fBaxTjR4LQ9vYZYE9Sepvfl0FJ6PUlo
UGHIOwPQCcrZZE90izwBCR1udtotGGRNzJJobSKfNREwXxg3r5NmGtADxnDcZle0FdFMScjYOVwj
xpmYlu5CF8yIB2W4OMn/pVJ7OyqlOUh5WVlsEKPzZibbvcBtDpOOCczrNU7o1yz3CkAlATWjRuNs
yLPKQEFXvsCCfVWuq8EsSoY0B+f1K5DBjaHiV4BTQvvXtzAyQPujetok4lyA0enbzmCijqKIE5zY
j2VDnlY2lNJmRd2NbCIecjQaOqGRtwYFtFJVwAZn8ldUx4+buGW2sIJ3T/LzaSYIe7TLBg2/FRFu
R4l3I2yVSfyDLAj9z5Bfh2gzC7Z+gkPdyczM9+EjrEdWRJsV4U8LJijuQ2QEpoPsQlA32cd3iUry
G0Mk3EXeDJ82mP02KaJzC8BVxizBrXUDlOJDVzuKFHhTWrE6mobzqQzeajHvq16opzTgbH7QvMiX
kKs2LcN8NmdHP1okkYrRll1rUfyk9+FfUAxczJ6nz+MADwsBJNFBYB6ZApBy+Erek5CKcarRbo7x
zgvynIDDtIXafIY6kljvPjtb+zCv7b3zoQihXxoW4smOdzofiggPqhO0NPslclCKjqLY9f3AWIwH
wHfN/27BSh19sLE5ZOuN+JsD/i1fxKesUleqiQNCCirkGRAGZRP79GhnVDcDZF5ktG0MWXyxxqm2
pQKvKR9Ic1xw+qcK/VAv6ym6ZHzfYCBRQEQyf3rRSciP2tLPuavlMav7V4mTBINqC9t/Rlgm3day
GT8wPGNR86gZ5+WL3p/H7fu42ySbhqghu3mL9BdX9Xe3msOgwvXpDvQM0dhJkanO4beqy7eOtTyp
Rrr5AHWSMbrYq3AYALgKTYTM2QQw336T5dsQQXzjsHZnR4tiUEAw0iwc06I3TOmbFJWi3eYrKx0a
Vhjncm1PapF/cHvfrzm1fgTTGWup0EMBR+ff0ddFHGAc5oKVfwpSZY/FYE8PfXCLNuZw5GiYJ3EJ
MIjL3EQCMs7rO1roFQlzPUlN1g2ki0r3M/KnrYYepltS2+UXm2fkMymeNxe13gXJ5s1/cznX4t5a
gK7YibAlymKSYZjGgRJGIrj30JGNzNJg3E94ox1490nlMuxapraqSg9pvqqihNqCyPeII0RgUola
8bAPYPeQpS+NJMof3kVbvs8mnHUJUcvcnMTdXEonmjMo35hWzRVgMip+bUzMDia5Rkr0m9f7NlHe
QPze9CIOUr7EmIgigDtmi+sOxfTWXb+iwVwkbXBVEErPtp7p3I1tzXgP+fxyWS7kzzeEXCQKLVfz
HpeH9ge3SJDS0QDO9C4L0ydEx/iFXxloPPf6NOo8oZdmXuwpZLOja4L9I8M5kTPBij5wNlCsHhVg
jO0YG5XTpPtA8259bznQW76oSfBEKBfxd45qU1qtqGkSKhwN9a977q/9MaJeVV/elUjvOSfUXLhh
y2c5UHFLmeR0E3hMLEA2Ufu2A9dfdfgRikhvFvbwO2vljgOmVAPF0BW5WT9+aw6Qd89YfnDBbckR
VfKoxttuD158KWPs+TRHMslqd9u6DZEu/C/vN6yMFMnjxWUDK7B1e2ewiZd2vcD8LNDsAzHanMhF
/TEyiIBCsG1HCSam/mZLMa1BJM+XHPh3w3J72187qp0MwIRZO7g8qdWJjKW+QOTzDuhmR/6Opj+I
bF/GAL/snJF69nwuu0L+Hyg5DjHUMXmwhc7xZ10QdnOHspWME/c8qQX/n1UzER/gJZUGOxkYkQQM
rMrN3K8Oh+HN4OIbDbEPxXi8oVCgcOFY1nVXDZlSDNdEkgjIxUQAMRceoyLPHRgA37juUWjjKI8o
tVuVdhA/c3uS4EKIJyFbG9CZfbLfNkehaIhr3VbSgPQHuBka7jwG/SYOoTs/HsChfL0CENeSgDo7
FMM7ltkg17jfEnyRXncmLhPGpObYj4KVth9YI7OQc6QNzWXru6aVfP/sRriIHYQfrLbQGw9egBYK
R4o0r739+lQEldeMIt9/SjzhhkOYfe+hF2mmzwMmSk5MRVnZqmpH5UN/vr4DoAla/GfqyKb4gexr
vbzFP0cYcuLFumpaYv2PDikMGI670Dwwx3m01LM4IvApGk+shp1pCdCqUv+6XZxi4Y3r5TvPN4pX
qiRAPl+bbBmFGSr4TzYyw1mcVci8pRGA8mn66VSN+SRO6R1eewk21qllbyAn8yYEdpxSXcwgQ2yV
Kvi/cMAFHxeDZ9c71SJ1RdBGi8ff8WdIpcpG/1mgY6F6kc7xv+HuEVluOnbY32h6t5TQpgi1N6tb
630/HMpkHTm/IHc8w7mX0MnI16JhcjFRG//O2UkLbBwDDf0T1kxPnZXTSfdZNsIaIPEcC8Rj0V6e
r7wx7SrgDOIbnEwTbmRd66cM5+fZZNc9hjSxrYUvY8wIodbJ0phzGvwAzjbAnbcHjXOKuJHR0bXs
aixYktq4l1sP2y09gwUbINBNmEYdk5SVmKs+qzsM+ehuDBnU4uhF32QE/LcWiLqIlnKn2WNIUjaB
+GnGQ9GPrPX1EtIWelys7XQRaZ5eZuHegyyU2V5Sds8KgeVheytZb9tF5iqeiwWXKVqvy04kW/Mh
EFsIpse+Z4afWkmEhh9zO0PTQTyK7VrX5W230JCmr/DFHQZg/hGYtEa+2jgNsFGZesuert0k/5Fc
WKHCO8WBW4d+ohv5VxpLVwXzRK85fObEOq+klYETUI28AUr5bW2vmxYOEKJWuJNW2T6sGXEvXrLf
VydLMnA3weYu0I+z+gIs6odW4JypCUXQB+3RIWAiraO0VFfPW6Qx95jybqf/moY3SlGZghBwuEpH
FOndR5bm104RHYP/eB2a3cm0R/O286810knatKMaIBpT8P0iOIlWhfM601efJOycn+Frm0DdJlov
MHwJGoOEtTenohG2MKi3M+215ap7td5hlcGgHz773qmyAb0O2RdGQWTva2Ui6HofjHwZOQGLeWXg
+JvHOuPnftQR5jkIXF9T7ljAUH6kYBdQXkFIXjafGaU4DoozWYuIug4KVkN2YRmid6MdRiFuGu7l
26dITnguk84j5IVXLpU1x5sa4nzSnY18MhwRWLVTqYGxM42MJ/lHKUBV6JE19xd4B30R5vfH7y+b
lj2fiLk7asklj2VI9Q6rDu4x3L46RQux4uLg4INWXbdh1EVIFqYQ7WZMFzXNPHvd6PuZzYdDk9As
5miIoWPtbFC05fQTBuSz9wUy3LpUyFD2Q6iAfT751Vrl0BshGi735v9mKJjITpl7eswPOxJDLwhQ
i2YLvUg/2M4xCoF3KOHIQdWFS5vjQQ3eFdcz4Jvth+LR58Gt0MtsBRAlmjVqGc79OLZVs6Zh+tFx
hLOgSSGk4IC2AfNNPaAShrzgSS/lQW8SmbReEF9svYF8rSCjlP2RfXnIb2I4RzaImzXIUg2uRhqr
QFFxYCH6pdoNtjEX8xq5/tI6kUI4e1kkM0NVtjGkUsr15ZU3WEat7wNlWO0GdKyvxsh43VA2fO9U
uCT8Nzy7C1GixBGdotuVp0Yy8GOMg+f+ec/kMeUH5/1gsCbbeEUVzxu64HYDBUxiITmZ+F2kk4gI
zJNQr2cgnOlktdNwXjA/kr2FrGrpTF2GjFSPJP455NS7YgpIuFFyyGj3Ozej44kgEddNJUbUCgbp
s3SarbUrukBbrwlVIovFFay0hAvtRvz0LZA37CQAy4vwubatN1sjFa6pYmfdMFdoSDyNE1u6hndk
9OnEWfYm9gWzzlnKIvc6dH5jw5w2+b1ID2IW6506pBSDB5a/vuc6T/Fbva6r764+9mKm3wA6QMdu
eoOsqWuaVXtnLPlqHJ/eiL3Zz0tzmtsAKia6/F3Jae3AuKt61N/9O7EDF0HQeTQV7NRaFK7p1E1h
iifzA6016MOUmq5YfEDLQJDU7g9CnZHt5Ev6wQeYyW7WulGnJUPWJS02F2vLao8mw0qxezbAJNkP
ytJVXdsh2c+EJ77o8DuTtb6RPKkkkQytqt1lxiv0LpuDnigbWZSLmYWGTPburg7c/LVAxNZT0iOO
Ho77m5vLgb6YbQlyXXmvxIps+ZUV3b4Va2etJG4DBnGLp5mSYNyC9vGs1SxUH4cZTmogXtkHYIq/
0I3o4+LRAxBW1nLmZl3PUaiZnZ69fh4khuRam4TsESsyy6t/A3CPGRxv/tSerrEisUSoPVs//1Wc
XrI9dIKG7QPC799eiikHyfXqRoeZf5gMJg34sdf8xzytDuayMnqSMc66FnYuJeF7rj3SHSDO8F07
B7U9sjO2Mt9wb8SJrnJ9lKOdS8RbYE9TCItLV8sVFoEV/fpqStpNFo5ETaffs73qoZMJGT+VFxrE
RaXZtXmKB1yQu27XfCNTskhhEaanh4nCv+mlL2IcZX+/RYXI8UQkEaeY8AgftQrWK0lHkNvziW6M
Qof5KTxwZjtU7IPizMv2JwhXN7CKuUVDMKEhsiGksAAFQJ8mSOurNNCjEpVX7l1+0qhOQXCK3ouQ
FqcBd4hoBN9LJgm9rW3E0xdNlhCuHgah8su6rOqlR3uOyxuXNeDSGrHGmOB+mUcSMzkVmG50Dfr8
SY3JeH4MdAITAANN5L3rS9iOmcQ0+M2wPZYH3vbqB9h57DhI38LNi4yPijLn/b9HIJmqjAiCdcMB
ifxPJOlFWj+e8lc+0KHLHENo0VT0Tbdc3VVb9GnBL3cfBksAh48ExnLMgmNkSk7BgirbnmjmyOBa
P7DFLWJKiYgtP9nm5JVmAL+OiOXXOXDGcGtm60sUQHXWAJQGCcyxBp3wga/trgcHOZDoBH+24TnP
FJwmPvD8SirrTkQiT3KttCLQQYkGDt6frTtsjXrGYWNv5kemf0gVa+HtnuJZU1qrOEHLbvtOABhN
z1Ls1ZfNP3NHURrSoJ24DgLgIzNEo34S2AKAxeAdgAuDNDcHmOGUC7TQHFbn84ljzdB53xgMMxDY
4mGkhNf1wSK4VvPR62grVYm0Wh2/xTbSpoGSNK1ep7Y5vvkgz8T3ekbZDr5F51QTMQSTyPdncEim
ryKBOmduPdCtfAUSLZsU3rHJhbDEhGjXE0UecVpiO+V/qIF0zs/InWhV1B+9yMUtb07D8El8Z1SB
xezPKBsixzYEGfQPI7jiXXEgwfywXoMJwnX5DK/B6kM5S+iWqpkc/rapfETStDPGNvV8E1/UKuM+
LaaqQYMX1S9yCZoangcuyQERygGUFefrFoJgspJq7X/o31QAgthcechAN4FXi7H+ILWrVgM1cNa1
FmI26BJzCmhcAwZdGCwJ5ngFSbU7fMkZXGLXfYhXz5F50dB/sMCnBFm4X5cGEaEhNjmkBxsDUZ44
+t1J4HrVLYwTQSfZZCj7CnkghmrqRRhyoEyvcfKskmDuOmTwnLc0dAaOz3jpEPEks0GFX06goybl
2ksLKNdXg9Px7YLDgkhu1F5/1r9Ff5AwwhdOcH1Mw9JtGI+p74GQpL9AdvKO2LogqTXfVQrslzpB
DvyLYM2CU9cbjOqZYwo+9sFpV26/TgV4NF9+VLHZR6PhFMup1VRG2/EasX5wOygrDPFyqUTIIzFs
TLBw9NN+uzzaUtHWoAoBADg5sfKwkOwz4GPnY/hwUnDcU+R2rPzRKw7a3yQQzZ2u2tMJeh7Xvsfr
LSIOfIuaikqSChQ/sQnwEGrocmJw3fEzBBwW72gLXQ2NanOkl6LkKxZYhL3k+x4JzkroKYrQW6oa
6jB6NBbkkSlQ2EACanoFw3QPQplm+RcMAhIXeVMHwE4oqbVbT/je7nrVkeEnhGfm8eYRSRvJPymk
MPkGnpUebpBmRTvqMA0VaGjMFgpUO5XxhTUio424HHlP+L2sP3LpXezWoINP9LmiHy+b6/3hrfF8
aCKAqL3LDSHGrUA74OVpr5+abv3NPHDr3KaIB2hJ1zsvlx1gb/RcJTGyBacEm4+/oyB0BbvtRxGF
NEUmr9lBjulpPUmya7LJlCtjfgov994god2S9eRlyvNCtodSMtdebttkm9ZaVYemuvfwmYtqI0mw
EEEw3zAVorV0PXM/vZzLgMq1AiswwVxZC+3jUxa5k2oCebiX0ZyV10uDwwOQTKnrEiskK0RpY6cB
WwtrOxHuAmW7aWDL+REYLoEt/lQD6SXkJrqKsMBU4rDpjjn0PZBlPnINXHudz1SSnvagO7LIKtIa
2R+BQPRVle8LTcOZXZVD8X9ohZ+fEnTLKT3XSQ33zBXoUpXsLiyEnsTy6UkKsWhMQQtq0HqkbGzx
lxB84LJzu0jF9gyJbwsMFhnJ0ltCVJnMBwarfceCIApZQMvbZv4WB2d2cnTxLAcK2Yyv9Xp8r/xS
J9WTDu3utmrn8QuphMkxOAFazj9bOs25Crv8lx7d2psyRY8YaccTyQpUkmqS2t1Axj36HppfLuZb
2r8+DBAtjkNU2GNZcOsoY6/HVBLYouGSQm4JIySWTFHfHo4tsgUJ+2tAERT42brvgyQ80bpxFbZ5
JDcKroVyRKRpChUcGOvJkSjzj3Ayf1iU9G3/Q1p/PU6Ju3hnUz9x0wDFT23gfISxutoF92RIl07C
JwCEmnBwEnbZVQ47M+d9M+Q70g/DTFTHBPNhvY/OCyTFdU7yrdFmTqTwq/5xYTNT8Fq/8YMg+bw9
wtkGkNCkrCznQWCjWztxw3syisc+umKwSGTYa7lU/sZvtstvNCNI3u8w0JzIkwcT9FBxt+WYA4R8
G68UrUBRqJLvtQaetZT67f8WNrDAAATLqcOEdq5XMYzkzIyF0M/WBfZjyMN1abXTnhAk+H+shgAA
IytZrOJgaJkyS/3GqCrX1khc3XaJge9/HzwTOmIL0kDX7imdU5SUBXjI6WwQMd40RG3TQbr9E8tN
cSOZqctyV0KqzFS5CmIaV/xeGwONaaIumJH/kTypvJsC8BhIDoRAn/BAMqBEECnyxAd9oXuon4FS
lkUMqAqOBqkShvnpCoDeRu5ScFiLYho2b7K7Y/gPysI2bNHauX9ca1jNv7/obtbv1u+WQnLP+M5F
vAbRus09k1IN8mRZSsz1PUHDKyFaU5T6cOS9X8GfUTf8Q8ZnkcvPfChbYV1PDOGtuDDHjnMVptsj
UCVs9wcug7aHJBB/NgrsGTJjjq3WDqOhGy7f9NBdN2ccvZJTmfZ8RcLl/llU7bEu3WfRbTr4U0fd
/ezRq6AJJ5kSPfNSjyrpMky4CPdTiBumL3Ba8qKfK5rW8Lco2ylJ0T5WXx1Z5QjOsEKuh3jpHiBA
iCIGVDM02HmKdb9GSzkHW6Qh+GVSl8dwWiZ3kevUmeujPv3hlJw/c73JCe5HDj6gAJp5uw0eVVLo
eJcZmAgwBNzjNG9oalhjmUezDKRK67yV6nKHCKA+H6MIXvDUxj3klX6nZt+u6MnVdUx9UwvhUnp+
Iit9/W5W46kY5tDltWC5g1wgbIbSTJpMBhlEpAXjoEJ2E4mKr8mhVPSeuNH8YO4woETmCwLoFePm
CXuGV2BBCdgsBLvhOwiHcVMlfjBLi+YjQHyE19fB1pRSdeSqPrpGe+4j1c7bsuDSIh2qQ5c+mbTV
NKsfmfKaYqOwdyJ6tGhW+GESS6ZD4WaMKgkgELZzMcNBa8oh4fL9iWdonmrjK9oRWC8QrMkf58xn
fz5sph9vP4rsCD6vh4nlYXvIS0zpaV1ZKQiXSNjJ813sNG1+t1Gg/JbZz/1xvvZ3ejsNJciUjHXq
Gld3POlPCqEe33Xy43/xR/d36F4OyrC5Zf6MndD5p7JxKCPrxyUsGhJQg761g8qnXb8V1tPz2edc
xrWaB0XXgF7MKwHRpjRH7cDMDp1xCDzRDrl8Bdj8BJZmbgwqibC45/iKfvbQ3kg8IGp3CmnAiSsk
LtlhG6lNsShKXU/5x/PQgLQrJsKN0R4dB2rCljdNZCONlR6yNTOr26iCsNmBJ1cCbH6/sIZYR1Xa
+dGHuGwREj1lpdMz4vWsdZQzQGVNIuhUc7MwPYeh3AxdOZJEqvf8x4nwZLDr/rMf18aNF8EO7YUj
Sk4t3YfJIBgVBwo48SrsLRvgBv8rzOotDYJ9NjtKiUtQa7rk2GcpuoxCgKw0X7JHvr2TTTaiRV31
6jjkSzblNKxl4WCiOO7r2r2z08xo1ThCpcvjWKgEdoKlaH0tJThxbv9dicsOLlRa0etPUPDhQgvw
zJyzZuJqPvTtPH6nboY7Yc5YgN/J/A/XEZ2KfKM+bey6xQ/et6wLcQi2Py5KU5gzGqo0xp0LXf79
6ElJPbXo7OqYsCrAFkrfXYAagCBDqlSQkKXY7aqWtEnhclJyozSxY8WWpx4qN5xGQa/ozDBizUht
eh9cx5wLe1WDlzqZ6fb++L4bIj/3YKgkGo+Xy6QCeURijBVd76jC84EA4v9fPN5QY1R3/K+2Ary6
lda38omOkojHmpXPhfKWGFRQzW3qcXsSync/UWzrsQ2QjqJR+llUA/S1fRICTWe3cbfgrVqb7VwC
QGPuLiwPkN3WLT2C6UaVXxb1FhlNRlMVOZni2/vaoUh8xIO5j92ZAk6YdtK68ikJfe6giErEUQNG
20Rovulmk3Q2lbx3ZqxigF8FLRNmieUGqN9jIdZcD25nhZCbXlgc53KIDTCZsuI7ewYQAAG6Ol3g
3ji5UW/u2n25Gm1BKvFPBuS7nwii3RkB5CgSOonTFjemH5mGDuco20+KTdXS59Kh+qcZFmim26OY
6ZbpsVMi9XsY5ryswOsbYrCQhX5L6O2PoLyBOcn+65taUd/SN9xY1dF8LlyPl3ofYDIOJWaPNnVN
e7DJ4T3L+Vub3Qri45rhLMTqkWCSqHwy0vzXSxK3/3QA33nhGyca8eK3gCdqlYOu1equqZJ4zzEC
GkGcBdCmcw3oLsx+KLuh+Fabsmo5W1A6GUk6f3wREbmFo263JjejnO0xM05GUVA+BTonvODn9Dak
Rv1eOBwapBakTrk19QFs3q9116JUSty+K+MwR5QNbcMf7S7uChjKOFZO7b5X3LqBxrf7cQsqGLc7
9fKAODXRUxwV3I14XhTUUlvaJoL5xw/K7XOCzIsCg6QrrP4O3cj5lK+MkAMAeMpi5t1YqCqcxtVB
Kgjj1lu2OIpuHcASSlxgSw8r2B5D5m3EmHJBVNTUxP2E2oXkp/CMpDgpRY+4wfV+iaHohbad75WW
RHOCmpnC5aBfbE6h56x6wFtUvnWYdLjVz0IQpQstsliE4vLKV7pqxQBYyDrji/DLafINAbBjUs+w
mytTmJU0EIYna3yqLI3D4FW1H0LYBqdTVfNlknbulidDrfODfzs32zdIo9mxXGAkCQlkB3akqkxm
b6LXar8o1siNTuX6YnHD4PBnj5jIultKyJqPESBZb7S4mOGKgBVUo7htbd4jk9Rijpy5oRlcwiAZ
/9RH8cz9AD6ZAzT2+5YGOMJu+OqmBG/ITNYUvFs6mdciOnMVAeQMhLQiQLYqO+6+Ib8fTSed7fa0
s9dZkhjdPt7+hE0r9YCN1SDU+Esp0PUpHr0puQIjstdfobqpCTYpAT7/OIUZrQ0Ofpg7KXa7nLd3
Itscni7HqqPqEJnx/LEo00JOur1ZU22+iSoTCccTdHC/rF7/v4mAQtpGum7tYGY1aH4fVf3y7rKY
E4HvEKyLqaogOZ3UhJw/bREAI2T9c+qIOcjuIwbOpnyW1IxN8mBMlp3TVCNdDcEGtfndOiYUtL+d
0T+w9oAJIPHBgaqEwIzJdvWLrnCtcK9M4ifHC2OqGux0nerWs2aaNkwWQ2Vmqfu1fmKVuIbHWYoM
2fq1ZjCniviL9fQdDo/EJ6/DlkFWDmD44W6xnzD/8gwehTBSyJEqAJnMFFy5+O5qALPireXe0oZq
eOOY8iCmJ7qeA0nZSE1bSwqqy6zyLjjQ6iOfYqmA5EDmndYKBChII3Gw/svSq1/x7EcY/kU+an78
uAUOaDmH4MzlU4Q3oOeMNFJCt3RtLKhLmOlnGV+Q4cQNvtveyvQmA3hJOdHeCGqT3o9TN9WA39r2
4j3+fzbJCnmrMS09/0fxVwo4e4QpWPzt70l+W5Uqaj7qatgS2LZLdzT60yZfZ7zgrZ9axuFkFeFo
fjvKc6rrGNHIjHe/rk3vcKaPc6AE7XIEO6+5eU+7hsdLrwYclX1GoldP4GVdjQK2m5AdGTnV+4sg
jI38reeHrhth9zn0wnaRxABdW7b/27Ij9OMYMnP56PWs0PCkID25kBLkY+j5TRzB3fONDbqbq/zW
m9Z/nUV1VZohGY5wvFU1Lxz+mouiH3Ek5nicBDLn+LnwTugmCxIgh5Dh/wEXxsRUROwGyaiRzyCs
cVEVXmQkRzPf6UfrC27srQDNThrg5Gpdz10AFl95zA18tHkR3z4uMn5yBMvCQPUhgOuqN9R5VkfA
0C0EuVHOqa8Jn5pG9mLHYfP9DlhocCL2kapgeTp4wgrsTdhe9zSsXt/o91PwN0u6ruGFYxO2iHAG
gPxpCNX96U2hSBLpl/PPEVqgqE8gMToVHhdxeQIk6bfBTr4Q6TmusSGB7ClDyYlgjZtalqwqu5D3
VYX9urFvlELKyX4W3xszYEaZbEvItno3hq63F9B6M1CcZrZJm7o7v7/IhCpqW6zM0bv+6hK0ywKy
1CleaOQj3XW+OX4euUX5mHG8F8qtaPwPkMuCtOZZG9a3pttBV0b2pvzfwVFZPj3pORBOdR/kGG8Z
L5C8nTL1KAVvrMi9nGGoQ5Vt6afiIbfZLMUjCr7TsTpItn9KIIIHpviAG44IXdzhvZyfk11suYma
6RT6Ur1Vo5U8rD7ZsPIL+cFSEDBNmw+X/kOp67Hujxs9WqdFNPhTx1CdKT0NBN18ZtFi7Jthn7z9
2dYtWzyJVxerO4c8XaLnJ9qlA+SrvKe//BZkZGJAJRLZl2H7CuNq4SZuTZF26yAYzzZ1l0MnwPwS
hfUZfq/sADay5sV4tNBiWHZfk+7jh+e5s3DaRaa7UAS3RYogju4zToYKiKEl2gC7SJU1J4q421Il
Jv0LUDcROx0BuHAG1I5vtVnKaOo8CfMgcsureMcv2tMAL4yYmXMYAGa4SYuwVsb3gR7A0bEaLP9k
ukTYEuusyC+XjzPrsnMdK/EcuEhORll5hhtiKxndh0QVlSMJx8u1dnNfvx//jr0hQO2tzvcj4c/z
s96ZiaykN2cnXuD7xICYrtgTs80Y0DCCQyJr2hDGQXjCaNGDhQfAVh9aqxa1YjuKZoMr1NyRJAYP
tbLA9+kVKiq4y3+jy+tw/gabmEQiP/zX2wiR9BCM98SXNBdLfazTk03R7/hGRhM5nMyX0uSfVv/k
g5rjmzAC6PYz5a5AKnU2j7l+RuVTh+KgOk6Cg86w+oucCIC6C5mAveeu4ScXIqpyg4xoe3m6YpRp
KCkmOK2jym7UmdfMwsZXQKvwhmlSULlF3Ol9cO35lKqUXHrLwuY+aoqdVfFUcruXDhLg5gERsijn
nivE6cQeRk8rhCgzr2hNFrwKnDPQLM/kyVstTDImDNz8eSVNcnuqKgUFZahWqVbcIeqpxmuRs/n+
eLtAOHW4T2sds/XjD1oGvqFHN9Dka4+5PU7Ov79lY3rYHjtPOPb4c4bL9WL4EEanYiM1PTIo61W7
Z+BXKvuaMlCM4yR1qiXI4bGEzfnZkAFqVwzUuRAGmx3SG5mkb7x/TtB9TnK8w1BJ1VMkB1Mgsa+r
U94Q/qRt4j4MURh+CDjgd2H9JmqTOfstol8qaLL3BudK30Lr2smY0LaPYR1AzW0e1rfp0/IuZr3f
asWvLwDu+hk8Cs+1jtYOCvDe10YZsDGlkGxz/4FzNc3R6YziJ5YiTxFiLR+9Qkn9lyfIMECIm22c
lO+lAeCsKLULpjzUNa4cL2uEHqVd1lfN00PmIs1x48uNWoGtoWm63y6CNonrqDLXZ8MIA1zshcc3
I7mPHb6tJdJKEt0seeoFtWIh2vxznHiUJMssFq11bWmC02wz71Q91XJIM+2OkVQNndiqx5qlzl1E
a1jOlogaeCWUpR93NMY54DSgF3bImW3hhgr+G43gvZGlxgQRRNOEiL+CmdLLboydxV/ZFcHSKZBS
sQ2DO19IxDFUIzfpcq2W4sNq7ZnhYFrIULqXLrk233uxb5M96iFjZsHaIISKKlHxNMy/ch/WRyRH
b+x4pvnx7HLxgmpyrE8TqRkhhTDSeuujkkqbEoBG1m1+rUd5Z2yDEksHXfd6BjWUcU+bSVL38KMZ
qG7S1eugJMkpdc3Y1crf8GQ+YjClKvMTIVoF9E+AHZTls2ga+aAcCaZujza750m3Y19Zd4LMeWyL
+waiDJyfhf/KLF5dyWZBDRHTr9rfici6h/k9HVp3xx8OOStQeRdVPCz011wdH4JLiyBygrlkO10h
ZCW526z5vhxTEeLrDUpsEG42I93K3Ak0JelPl81lgUnpF9jhxaJrFiBGvI2kZBsakXAcIGx7OxfQ
1z4qi4kNuiEMppkoRFqPDTQ/6TkifM4gitbBdz2QHjMDBgMP7dP5JPDuqowqJW1hMddtKsNfWKbd
hOIrmkxhQjKbr9p/1CkoAPp1+Nexhgt3Mek4fXRXH4//fJ30L2aizMuVGznbAnPTJF7im29q5V63
ZCsDHwL19gLjDpevaDRXXIF2P0TrXawZY/CPJ5PdnSSKAgcr6her/GbO3jfM4BCdawkCZV1gxSNq
NYCriWPx41cKSj84rwlus6WGjUlsDasGBTt1wyPt/LiK9XkyEmlt1qgRSh4W7cP+DXopa89JP7Gs
e3ryNnb9cvbFepgUXewr9EyaqS89jP98j9wQV1tF3ChBtB+BQddO7M2CefUsS8vojDIUBn/CSPIH
tOKUpQCknEOdGezo61MHW14goiOySDIfvZHALdVPTPwy/L4udkmYYtHpELxNWEXQlLcOerrgmb85
dQghp7ceKt77HDmsd+ILGPaqUQ1ZjaWLSRkxgOJN9XBz4IF8RRjErJ/qpxgsUVTszX5zMw/CcIyC
k1BqaA0OTdxMco5XtMhfnrUaGh1WeArl9u9qpL67GndqqHhDwTUhO4CL9h0w/L5RwZdN2w8r981y
lT3w6UAabjEQWJcygki7CWzwIwlJmNoDxKeu5h5zIn9ol9VGB/j4AWU1UDr8LzBQzx+mpgQjPAUm
qOlDKH5mh/yBUfOSaH0Ey+7TQqSJgGUuGzFk/pnVKfoX1Z7iDjro56HkmFs09wt4E/yrKh8hC5fm
u78VxJtYoS4VDfOh3ypIl9tqYDZd3rLldZVoK06ZykHNcmZ/6UeNSZvuqbaA0Lj4wwetqzUwkjUo
y5b0RcfuxxU3mskfn7atLerbrL3CpA+pkqaCDjyC/xczmkBITImBDPQDQqDruOIjss4uOjl34ODB
ViToU3umdSyMw7e1oL122Wh//mWDUOJu4VrEoPthqfUKcBk2bwIkRWjRr4xbLlBfMBPKUd0LvSyD
gRH1I256rCWS52ejCMBdbGD8VWUqdD4TA+HJpcTd19UthACYKPCTbl6p0eWH+A5GsVsttgLmT7qG
GWq1WoeKIatpMbfdqXGnsffGRxOUjolYzDYEScfDE6VookAtteXcIfLOdmBwqVFi1yvQOAtfH44R
Bh5V5VpU95TZq+EknyUWE5OMz7x9om7Wn7AX3+HqJuA/mL/a0+T/aQgyLiRXKkvpJzQ4JXOB44R8
vkNezbgZS5tY8q7e0lSXapv4DyeXtYM8b2ayoMXveCeEOzWLodkTl+bTXAhzzdrcELUbRXPgT4Mx
ioNgfGdciXZArzjoXYeeym/CmjBycCRxg1FFmYbMSXDF5Z6zHF+LGX6mktuMtpxS1WS+31/T1nBU
3FpcdX/K2koEuCcGFv3/u4RFJ82sh0HSFsQcDbv72IUqze8hbMFYJGuqkQQnvzUBfwxPGNQOH0AD
NuX6mdztgOtx0kA3+4rXD5ZCNtAO/dRnYEX3/6Vf6OLtP2jY4U7yymPl0LUNG+5mtlPrw5MGpPiI
o7k7ze9e5MvLcTfb4crUCm7GFbL5yNO1oxJlDXAJZmrMFbyHlQx4zoJyoOevTrsiqmcZ+otiB9BP
Tn0o8G+7Gr7H07NDMdvFUQ+sGtEFJM1lENSPR5tYQ7s0as3c7VL4fefF0Rrdb1/8Ocj6Lo+tSkQp
xP6iuP68UKXCS/6DqVigeGDFnTXcZhw8j0vIhiEftD0fO3SzUniwBi8dktifgZmk+MeU5K3BKzqb
ZjThVWfMrapiy8/LkOK0FYeIc5oR4KKr7iJ9nF+Tanjs5T17mjmws60Ou80qJosvjv2wdctuDUTw
hVTcwjd7EesY4aTY6b5OUF9dFLJbvTMoEwYJ28uu8AZu6b3YTZz9P09xiZLhsUSs8+alDUg5pYXn
qUwiGFmki8BEyg8ANEaRP8Hpv9BsakPY6lfQPrwAsrdriyPpEnLjgX3oxYAhGeKsqS2f3NHquTGL
Twv27eWoLjyK65xpPvuADyR/+hmpRMC0IXSgNChhLwayaC7pDBnz+tgNvzeAkL9iu96YgCWg2Myp
PV27g0/Wb2wSqRmiiHmb+X+lsic4RypwRovj3G1vSJguG1F6VEYygatJIeXPxDQEFU+c+nIiiorq
7PoLtEUhSu9GNCslUvnycy6yGG3ZFdrBGgrh8ceYB8/MUsfJTKujscCS9i5NZ1NPoIOdMDBZ/2vF
nyVQQZQb9C1qGphS93oV+bvpP7t7Q5pqznvKS4XFxqHIpZ7KDhosJitJPW1jfdJs4KIjVLKopTuv
cSMdENBfFfVC3X+y1CRrbRlIoZKo9Zkpdw9aCTyYLTBTlNiH46k77HKJnHMFgR2IWBiQwL/0Zyu6
D4TwhDdeKuIUg1idnZkHY4SxuhNfP6OcaSSVRn7ssXMfy7CAXeF2AKmV6xxKMRWjy27NlglSOIff
Z1cpBXRpLWj0EHQ0qAC7FPpcj5dhSgo7OJr4G9j3dLxfhZfNc0UHD8KUqNUvxsz43fcPMeyP/0N7
/THb5R/e1X4yyS0KfUOmnqdFX/Gn0vVg5kqDjwLaUEii+OYaFiit5IdPbwzqrmAPfgIRh1ZYg2/p
WvMlgMAXxAKfl2+KXRmoRDtlGREy5BROK2JPlNf+F0RlLXK309YjPBPaQ8ku3VzQJIk8HgODL3r1
WEsiywurVC9Y31hKRYe5+5bWXiPJJ70ZWRLbJIWHK78wxbXeQlNobYgTicIEvK7cj5Gh8RE9GOPO
mJNHClW7Z1aEVSBxFo3/cGnIbyohbCELSHzaGEaUxrhy8LpXu7dJr4ZjHSQGyN2rFOlJ8y/or3Zy
2GfeAl4SuVfh1Jd7VmmdJRFsRB8Xym/mb1F0i6swcW9eVJJsYKwys3J/iWrAVN2oL1T7B5XE+cPg
UY/XWC+XCEd5PV4RhWooR9z3d3Pnr3D/cxGvHBIV7t+8WAwwYU3p48E3uzZLl5dlEv83ae+lkpIh
hb+WImmjGLgzV3IbCeA/1TIj2zwSLxoB0sM0AwJawO8dmJ0PG3Jy8sGLGGzVCrMAfgmAZ20HTb1g
lMI+aB222afcDuG7kU30Y8mBEe1BYzZaI3JozrDIWTKwMihJyhMpvn0ss+UmUUK3QdfJwBzzGIB8
HyaB65/HWC8Ch2BM3tyBKTi0vdz55kJN4CvE9E9wbKgxFAgGDypytBaHcCzKgZKIMaSCAuOLA38b
o11EWzxyWVqociHqi+AkGciuFylEx7t8W2qV9zUPxdSLl5fzng9Pu2HsZisuahKUNSoNU8SbKMSV
DmMAo3/Kg3w4MGDyGHBc/qzARR1PYuzppXCUdQX29d+rE2VJPS2/s5ydgT+oktnc/GiHCNHstm+G
VO9skFBCcqtOVfB8J/eTaCSkRl6Sce1UzrtE/L7an5oHmxgUxJ0VCFizO77lPpAUsq/EI/Kfz4tn
r98ReAAmEUtnc9mGt2Z8fuU2fGiLh0zm9UyoaXHy7OnyR4Ib+d+0mdWJDh+jq8Cl3WGzQH4EIF86
H2HoPcBm8aVaxQ/o423/i5Pp2DpIHUtUlwoC2qaGhnyGwhWzTkm9IJURDQO5bH4Yhjj7D0b7inX9
hZf8tI+DY9f/CgYYL1F/TgwBHvKGjRlNli1GAdIXpKGdXi1QWwfoS3qiLhoQIa94C2+jKTDAZoRd
a8xpjLVeN176t3SsF6rzBMUgW/60Pvo3jbfiRra4LfMN664AB7yMkbPKby3uIL1mKCHegfJ/CnD8
3er3AwGayfzu0fgFDi4vV2bfJpCGOFB/+SSxU+GW2IlleYFuVGHfHLahw8y1UDPvBbKFBR9oTDDb
TVXUHb7mM+e49jkR/V4q3Yo7FeyTm3NI6JHhVirTXoceWQ2rH2IDMLLgqWk5GWj42d34hNunFdNC
pbP3Lqx+NHwSBY1aSAzKhp9IbGwnjVAxij3eb2J6xoD+KqG8xahgFHRVimolTjmqTIveikY2z4c/
EnMozreoQBBTpXruzHmoBktNA639t+7/220A43Gg8wFRDHhZARy8Bkj/8/Fp/woIGJfsfg23b6ZP
p5hn0pdMBBMOFOrby2FFLXwnJiHwzivR7UofeyHDctHnlU9Z26sC1C1yyDNUgbEAu/49Y3niOTIq
PEdCLElq75onn1E+u8qr64VOmhdpUQuDxAHZeT3u0siwczxDhRsrA7hdXdKwddzrzDq6v2jxvut9
+CEInqpT0F1EOUkGbAs7oJFF/8I6zJ54gaaTreaoPYBd7ew5WRf57hgqIxCIEmjNUxRdGL+63B08
l+DAxovRvESdj4XGuQeWNJPENAdzOmPYYnpET0EmHQChGURRes30IOkNJtA0AnxKDd4ldAPiwz7z
L1+lxpSF6b5D8kxBRpp2RwkrhPwwL0+WtN4f8oiqj9Aziu9sMbs4pT07/OX794xlDbI7NvceAzBM
V4d6eHO/dulB6BRaB8uQwwcDs5UcdBqzLTuvE04yX5y/OMOdwK6yIHAUXkphJO07aQMxrAj3+cn/
NzTpPXeEiXVUuFRl70Yd4Z8/IwMl+LK5bcFfG5/k2hLcOYStF0qz9BZ2p/eUWVOa2h46dzv/uAYY
BA62jDJuMo13xyccvV+Q88JKMrEyFhQlXeoOGdXZWmM1fTH06OnhBNfkhUiyRGt5LcAMFJTJi5hc
AWmll7uPiEX5krLr1MEGCMemZ3RkNwDRLEVr3ZS+MVylwKyW9gDQNL8JHSXPOhXrJO4NNLkXc1II
qu9W4Jj++k2YUq7j1ygUan/woMJXewum6eRGP/u/a68WpV7cq4WroCaoBOoziFI6NGcGgCdW3ZaE
WygaEWXlEsUdsH9hZw4sNuVS8fMczGbJ6n3/lr/ON1GYpvytADKvSbAAH7py/MFb6xxyZOhbyZW5
tOP9q3uZUXcSIG6/EhsTVZxm+f7nitdh7j9GxryLyiPolaNct/cI2zJ56I3D+8EvW7S7BVMXvkYe
xVc4NY/Zn+FphOv+D2bpsO+EbNtKPLD13C5m0d5oCdbwu5SRoOUCFFE0nt7CoLfeacvGAl9QC8zC
qjcaBuRR3ywraFAH1ceaXaMah8q0R/UMM1BmyTGMS7IGP5Xw8q1s2me9z0zLYmk+MKZc5cRtvKmJ
ss6EpK6Rpnxvj1CFG3U+wrr7J45WOOmewFdgwpLLPIY74B0ALaT3V04RBX5BN+bu4RggSPImHOyK
GWpZLIb6T3h0ymsafx2kiU7Lhf6qoWi/AYZnkQWqEkzWp5QBdpdEQpAV6vCqwQpBTvG/yWij3R+1
NcCTnUaIc6UcufMHgEa/wulen7bu2218PnpC7ZKWS0yrbT8+U3MCgOG5dg2tBzbhYg8HFnTxKPcZ
8u4yAjP4TjMdb5w2WroyonDdiDtAEadkRVmkZ03smk3/HFde4zm7ChZZtLl0vVgw2zNgbdI/oGsA
hhQ6BYNvSHJWWYPs9/VvQ+0hXip1ShoPqGdhwonn6Kv61Q1SFc4vVL1uk30/6psvBCvbNJDH1it/
AVSgJZMphneKqCV/YljWhgG8mB/v08JFlJWTBY6+j1EZDG2QyAaok6ImSAolCstrO5jImmzliEx/
evBZelfzhRybdDQDp19qQ7XFNnABIfe3EH7OW/dQi2UiBmNZEhrwC0fMi+38cCLFW8teqzWIzbr2
W+uqlLRDJzwQB5UXDFQUKX81vOaLVc9TwiOzJWKzii2Z+O9p2c+sEPC2UrvNZzd2nvv8qa0t91U7
d8gqkq2ZWZdKj91kJ9I8xqGi7nLOSexiZKQN2/QWuQ5irSgByZ6MM43bIRmFqf4+WiWxxebeGT96
nl9HwMqucfvzRctBqJbZuTTy+KXVn/NKBIWxMcdKD2jXgcA82pmorfLGSjS7AALlNkVqIpBygvAp
FWQes9vyaC+EOiv2ZPs1kTFWo2PbQD6ucYS5/X22Jykc3CGQGlPHCLbCcVzJ25Scktl87eIHxdHd
XAmlf8t3gJfQHBO0VV5Da0MRGfb74qdUNjZFdetGKXUIQn2xQv9BwZ+mU2nnJ/af4Z81QMR1EiYP
dzxKmkH1vHKN4bX1THeQd5532nzbSJyMzK71CpzKSiqUmO6szqP46adi1DV/DZhJYEtonF2RRKKj
kgYnTiqgvpeGgUqZPkGwJKZP1qu/dpxAAvLW/hGfosvMLt+jFbbmAmq85oa15nV+drDvNVt68jWB
LGd/ZqMUTyl8IbspxxvLt3r7urBB6rpwAQ5cemAdP3mXgvAoFmt2TeU1YRlMaSRYXsL6JUnsHAub
j7q6vjVZ1z06vVFLa5N0ND4Jq+VV32dLdfn+s92ftBVr9Q7cbm7WPUH7DF0mZQkyC0ww3Fhfbygh
6NVzL0vG6BLnFjDUMuL7TOqbRwuJJgb/wsMe1JC0gF71jO2reGBfAe3G+VpgEJF5SpOlPONA1/25
9BMmXZqfAgDOpFeleBGifG3dEgPRrYHLa+6JRhRy/IjETbqYjw8yIKBeSCFDXgIwotAlgNvk1Y20
vQkT7IqZh2MdJF/8U8Hhof4DD/o9i4Y09MMgN0DLFu3Ib7m3wCpVP2o8F1h7mU2gNLsdaNY5RwMQ
/pdw79X2zPagBD+bfhyQoefoQ1VLFE6ED9fSJgOsPn5sAAQx2/NpNsoxXG+bAJGf66le2e6Bi/VS
Bx190wXssogNB9sQcl2HF5EKPzzBI1IO+NJovVxznZFRajFJFR+BHOJMD3OSGKqBVgMVk5gL39mX
SvzdTdv5FGVes2r8TkK+RHOVmTDQFICP2Vl0StnEzvVSxHEByA7Q43+3eg8O48+V2A68lOOvW2hv
Xu+z648XFgGovFapYtihUiqwetNzbUpi+KzDp2DuJGLKaIykektablNXR/Z+SYSPBBaRa7rN6N4n
ycN1fpVYcc+kL0RLjcUREtCievlH/OqCwyc+Pv3WHlgOHnjKGSoAhqv1fazkWWr+Tq53NRTKipvv
Xhz+e/rh2n2PZGGaEG+9K74Ob8JmuRb+KIJd9gL/jNBFqjd//tqjGwreZYo19h1OM1IU4IfgnNZn
PBqC5bVafxeszOUzqiYQXh8tzlCMiqNF12hIewqKrXy7YHfQ+iLXVm5CUhNEo/eAGHDC2+PHBVX4
npjLZZ/NVpTkRLedcFQwj5mS5m1oCGAktB2hpBjJ9b5PaTEVPBu9bz0nDVHcM7yY1aAy288YuKOn
HL5k1P/VQqJrC0l8A7GLRixutAkg6BatbHndESFQl1u6cBoTs4fCISuoEXZ4HEe9BG2ljpOrth2q
RqCYHudBP6G67ESi+yiv102MBqPMIF5U3trQHLtaRVwkxp6eEQ+rWHA6QOSLHXp+VmKMH+zirk2a
T7BNrZN6nR1QroLsYUfFa2kIZPWgDaFQkaGg142gTaprl/jQOF2nOcyIvak6gLIVUwsgX9/gf5K5
b5khTkjjE7a9F2NyhmfXuwJaNoqjI3sdhWqcNhFICSPDeU8z6SXAAi6biupkdHubpbLmMeppNvJv
rhDI124NVqceRG2MP1nSTTEvRjhosHvvKM0x970I36Yili7QbsRCRFgg3K7tACggZJMY3f8xWial
iFfJgAtjtYT9GNHo1B8qeEeOBRJGCcjjshbU0s7vs40YTE2oEnX8UtTew7WSXbrTGIE6WAZjiBLa
1CEiMsW8N4dk2asWymX1WtLCYe+OHAqz3v69UAcnEXORkeBAMt7SwjzIsYD0NJKkBTD0wR1FiuyG
wyCCnLW4/cLxqOBjxmkrK2gc58gBKV0tqkT66jhYT2LCuxFxgT2RmkFcbhjUrIlaG/h+HP3mMMAW
oebJ8niVg5yeX+fLDNyhFJDLSLd4LPWP/Oe2ty+qKqQ1uAE3VIcr5Hfu8CaIOeGj/dEmEp6uqLNb
xe16tNjbTxnmDCJd5+jBYtEmgcqFD4k1BDYeB7H/jc2anzsbqbXYN1Z2SwxPiC5L37WLhEQC6uB1
OOy0Za+lxdRucBaFaXzYiNx+RHUA+5Rr9ZdKuZA9up9hdCpCXvi6RYVmc/gKfFdxtkGkE3Kf69rq
mo/P9LTA4dgT0SPzEPnkEzT2DOobW+4Dqy0n7x6aNx3ri6ydW9pdStvFvShzFAKIYWkVwHZNGgiN
/6dT8+ZuEMc8pTBil2Pr9Hf6gsPmEmMGElwLH4g6m/ZkPTufaKAWdqtp9iKhvRXJzkbLPjPmegyM
/UiKIFTqGL0r8DsWD9h3o00UlyACnooVt/0IDlsr24cMg5BDdzjTAgp/qQZNKV28EJ723sLjQNuf
lgUOAFg5wLZuIcYFSBYLrZKATwTwjQHN+SBlORqP22EjrdaL7hxkYI5Dis0pBp5XGeQqkJ6eDzM3
DVa0KfwYKQFJqKaCFI1jfl8MlQ2LPalLNdmqKTmN+mYOMrIFz/4OoFo63kxsHQjIhVU/JyvpYgpU
4IBhNS57b09QQ6R10eTVnpeNu8jR9l+NkEjudqb6Co0W9N4lUFfzgKcvAuFECpXv//uK7bGwJUFL
k0nmBuaeqsj6WUBTjWK9wXv7vQ1nANfGxIVg6Ag0V9i3PIYywoH6VrWS/TD8r1k2Yte/aGV1+63e
1g9PrMKYT+JadZ9XIkglbcXzDO5tm1QIg6TFIicbdaLexw8inEl5aM+dEevSUs2ZvbkCH99LQrmA
F6Q4GywLfjNEdPY1droGHlp4E3OihlM3lIYqGw/RPe8+bzc2BkSzig8QsfUV/LParfzOY/fuYcPr
iVuRArdIXaNirBFpWaZC9nxhk9k0vHBHHSDM/kNLOur2lhwr9Hp9swyKWrYwpR+ZaMtTAS/RoP3J
BKFkqjKDnJ50DkcAuE/CRn7bgF7xTGAG+q236vxm++ZbvhsCAnLsJpd63pbmfDLVLvKj0Mabz3tP
+Qp3Uirp7/JC0VAbhLP+mkVfpdDB1XSMvE3yRiwAZr0iiFDq4LEJXcgf8EKgrvYJAq82MiM7+TqJ
OuhE8JN9KKT1JsERvYSh0ZIPHDeHhDU1+67QVduNS92YgInnoAzZFTXhsiv51N526Sn+v4UGgl3Q
GFWmiIrptFaOrGPxPGQZf/sP5gLheVTE5Xq/qQJhjL13Ddue1sXwzc0D4MHKv6iwNL0A5riNHfVb
gqjXiM7QJrvgREGUsPfMb+IEZ6jXBd9NhQbKMzeNBE4K5tGx8sqUfz+8JzcKe+XECVOJwaYfuNpY
LxBYzfImLwuy80dY5SQU7XCb7//jD3cxcSnlcF9KeAqMOT6kB9lEaEWqKf0Y8u4ipR2M+zLRRYfn
Ps3YEXsGUeh1co5D1MN1JkXsd5R2FFTm6XEE/JReYA6oT1LHHq8suNM/gSSMCV6PzoxXi+WcaB3O
SBHzsJBu8X0AImCzocmTFRL5ksG+sy2/lDjb6Ll9UJeZNVUDvu/eUJ+eGQmkrjfPS8dkIpi99mAM
BXXRPGqPvedRusRLTEf3MfkHUAbdeqy1vyqfG16uxVIu86GFSi36YMR8D4o9ZgtnL7jEUFLSLJVl
1R0TwXDyYieKVp3ml9gIDyxM0sDVn25oDgQYWSX99QucMIWa8nNdrBUhxtMv8J/3SjD38mA2eD3a
aMtDwTdey5jIwthkMU5vQTo/2XcOU+yemnS7Um7enRaxZsHSzAhFfBhHte+G9HEpvbLdE83WtNxN
UT0qK1yY88iRKTpwbmz2tPKHkGgxC1p2YxnpKFilhn2OgInnFpuXwanaHx7505BMDAFMQrSf56wf
v6DsVc7w/AawDaDgU43az/+5UUmAwJV04FYE2GopSOBcz6TQe0w8Op47Pf5fEWgJvTxVIIGpxyTC
PEb5qcbl1YLvrMQ2O0EOAhczK53Lc/6r2hzsh8Xpy5FS89qL1q0KtQeG7/2b2/LJCj0pDLODfn0v
SdTyzhY8XNjod9prKqZkyrE9L4gMCLqndoWm4ZEUfgg+z/ROUAcsynMjdVx/1WpX0MrGwTUEv83j
GSrnCJOUhEFfx203DVoee1s4mKAe8JTC/UNddi1gAgY7BpXwwcvE6ultIigpbFDis5pqJT9102cE
T3LtZ/SGJTbdVO7LrFSEWDSDiJSOS07LzKqb2YHjiqu66OvN0/ga7fFQx/z/+csVUyBhRQaSEq1V
jLW7knamtoGnqoVEwD5vPpO+PNDjbjaZA3Do3TpsUaAQEJIfa8n7YABeDAK9A9tRUpGKrU9BvOQN
UOAv6+vDDfHaLbOvpy82nLNctwRA6GxUxRA7y+9sgB3rFDGE5iXLZAYfvqaJ74DlGzuMQdHK1+IG
HSukgSBpqfgvGpqd41CPQTviJNoHgBw1F3uK8Zw2pYcrijzLI4slHVS7eYot1fFOwnki0vt5/BFb
4PSval82vlw+Iz25dTKidzbt3Mi9M0Ez9pw0HO4Z4N6ZPNa0UCFcabbsuOVngpEvRn3vCa/Y4+vD
PLtZhmKcgzhdamSG+RvTL3F+s64iOnSVADeOKVBe8TntMn+1Hi3/i+fPqlzBMYciJgIlSKBHv/j2
7ndLall3fI/xqDUbCV7y+2cwXsY1GGRs37pAciQu7p/1wYJb4ey0bx2domFIqemhdELdjTd+Nhfs
1Y+7XJUEfhTo5Z9C2OWXKx30c48Pg7KaHMTknZeFTzBRbnTgBp2AqE6v1zzVq1/pTOe7m1Z+o7C1
LWvtnzC/qKUZLQcvXf3y4TevSlrZPFrHHfhdk5ZQykPueFXsb/8IhS6bYdbPDTQnGdjLqE9CnbF6
pC5a6+/b9m2mKbv7ExzorlihiWef4bnWWjnD/yCAQFXVRLWT4Bza19PiguTCMUxIg+7LJmTkKUCM
CgU/E5InfBWVHGs9ADaUf6daP3KyAVYmHKdVLPblZojOHFRDgkfYszllJsHybhUq0ZGCqUAgVmwK
vv59HPMAImzvQZ1zEYmYa7HG9+tboKQoyBW5oK4FT6MGMwgs5GtGPDMLvUaUlcL+w4KjBqENqZ87
HDvxD/r0f6sH5WBWWsVeRAr+69C17+dvx0aYTuwCeGvW5YOgk4gIg8W/uliafjUwgg3dadvWIZrt
WYmL0tEJQQNA5Dy1itC4YvfPZvcS8nxdNvjI5rmdT18ofYkpaX0poL+y6sbIgzso0g7+6zpDUtHr
HhcjVSHcVjXDuvCg1DUkAd/ItTbJadk/KPpzUlfuqfl5F9aHPNPoQ5H2KT8b72Q8ZyfY1ytjyF90
iDoqSMqDFXzQ3wFFc0vtNCm7azK7pnmiwtyKNQ4fF0LvEow9+APPlbHNcCwcpOpk8RzyXAnQVO0/
+exD4Ps1/2L4CBHrA/tzm7K3LT+B/CzO7l1L3QElTIGH8+XAapdXDu0820D+jjnw6zhYlo/AjX2f
a57tuNCQiwVfu+CQBin7fFF+9az9UmSVndplwVs0BPIMtH7hbT5e6f5FcYQ/bne/SjzKQ025k6A6
noWZDTKMHEUb8Pj1EMbBaauTwNKIR514CAho9i7jKQ827cMNVKEKoLmvGSCmFKO9RXGcgy3J1bJP
psc69JGdvSZMnQUnRbSd1zebzQzGkW6kQl6T4E+8Bnluiz+tTpiKxvsS7T7XM94NgpM2oenWTvZN
WS96vGXJwvlw/9DA5+1c8+5WF0dOLH+8h/mKWD543j4GaFnAyN7dV4ng1R8KXkw26Xbx10lSp3UQ
rtZAMJAmNZlIAXgfL59hjIGSzxBoUPAQVUvwihA2PwIKAs8O1V51j1RBqC8+epJJuo0NHFMnCdxr
xvqRpogleFEVPwopDLkb76S3TLK+uJUXhPSpONJAiP+uHY/Gg9HzANITkOEYXnPPxL6prIMkgFb8
V3Ycm+6Z3D/UDkTleNJygRZ7JN3BVLGL76aSszqBhaxrLiFFUMzGmqKpvABcU22SwqoimyYGtMcN
ys3kVMqSXwzVLfvvlxBYWvtSKjui5ZDu151g1AN+5fVydt+/7UKCpUgDX++LnpTnrGPF3OnNV+KE
ohLjC3+VNo0JKFJ5wVWt/l8HPQ4V/OWcm9/CgKS86EnfVTG0QKzSlz4qd8B+WGI4TTW+nA6jQHVa
G/+GwqSiBLceltAEmqawmZdXqIckZfD07cQ5ALmcxTIPps09nLK2djNb1NRSUK/4rOlCM+1Vj3J8
NppesfTDmI2V2KyWSlSL1NrxIjxMwslxsGjmnxS/8Z57tE+ttaoDJm4iqenMJpRXnbWF1qXxv+Rk
zVJq60F4qibYyVgFBfcC7IorBswWYEffU+tqv2UqFTGyatSu8CqVgCnlx7dURkGFsrDsw0GzFIqo
EBh35gb0V3henw1IzN93HkqmPqoW+KGuHTHGUjziWGgmjYL8ewMkExjupsU3ACQLJCdzGbdnentr
h9mQ3BzXWnbPiuMPwFXT1R4czkhHM4UZUsTOaBYKvpkzhSuh8LJJ9fAfpQCy4Ka+qHHGBD0brYBw
Iz5+dxL7vzv/QDw9nf3nAh4KEwLQ73mOuJVR9qGLQnAMkSzL4A4FMO/loT6OvrSU87NZBmNSG60G
RtOUmGBMQ/QfOsXCBLgbvaum5PflxHDYt9aJugYjbqFPdAksFDP2gXR07RP/qS9Zc2VUbWGFnyIK
eetDI9CCMUuzJiiDcAJcX8EYjhTAIOcvk8On7PncXZ0/pmdLzAc7LCJMKdRgiWV5kGMTJA0m+nla
IUMRL6PaglchKcYA/enQ6mipmNxHPbctHsD9PpXJETFofWhWqxvb1+4KUIE6x10yYM28bjv8rh+m
6rxl0edEB+YIFssiSD8HZlG69gXR7pdRUhsLv2EbLWfdJlTtlHE+L99gZzwtsYIjxJP5bg2QqitU
HM6NcGhGc0qLJo5Ljo9n/mJTbkHeWgVS19utZmMhGRzM7l3DPW8/ogCjzkAeTdhvPvDWOUA9gtbA
uwZDLueyOYX5c6+WPzQQJm5NjkB6tsgijfDCFe5dw74qD2AKV1BVLWaJANcRVgf/I9kjFEaY7G9e
vbCSWLOeYt+o0HP2e/2by3HOnwcc52yW214otEj9t00zcxnJHwwkiQURlsqtqEWeQTjc2CBjy75r
S/JKVGuAGYkwY+jqS5D0lvUSuuqo0BRJMmDkC2eXTAdNeDJ+9qMg/1TmY8Ja4p84tcu5d730piga
/oS2Sz9TA4Y1uRVNR1Df7SNzv8D080VAvhG6TGc1ns0e1R7zJTEqImDwsSX6J/Q8tIIKrJgaMsPo
tzIfDW5N/KarbuLblJiHJmxUSQsOzB4W517SA0IH0AeZA2v2H1El4WJOAmIjOECPgjua0Fp4yFbE
g4bb8QAS2XvGsHX3c7U6gbcFpwHpQRMN9mbcyU42MB+syt5iU/0qSihi2yObIcDZHDrQydpI/b0f
XUCiQh+OQHA9KZARZbpaMj97YDLN6sMvQP8HyzJNhg0kVTR7bPj6N8Mf68QejE2bWQCBMOTkFyi8
jS3i+sLmoloZ3oGxQsfthUAXv81gTVijRZAdWvueJEY8bXMP8T6c31eHppb7Eyr1uNmTfmHwOueg
6krc6sPc5dfqxqrGXJw0rHFBfoWsUdSK7c9GeFy8WTS63JGUN5Qhjt2B+5jyTH2epG1mw8AjJ804
y7DFQpsjbyFl54Ra7DFKXpnRSzgrnpCMZNYT24i1S10TnurQkOEVzYWlChFAXYxp335cPFr+3iCn
foNTl/y8vMVkzNpQmso9LSUBVZHvt7czDZNLQ9QGSe7fcoLti9uk+4JPSRadre+aHti3oKZEY0sN
y1MbszS7MJywizXzPNPN19pAQKKQgYLfXxFqp0ZE5o23HbSTWLmMUsclqKpw6jD+FahRmrcZjmyE
sHWke5mcVSM+mdSfgWk9mgAhJLuWJnwEuxJG8BL5MgpBwCyBG1hhHhhDnV4x6woJSEIb8iR/wuFT
8uxpVCHssON0Ov2C9AJ4Q/Kx45uaaoB7H2QUaZvcO8xYRbmHi1tT9H5sTZCFmS/+6dWXWtvBog1q
Y7cm859BF+V4R18IKVQvtB5Pvee1Sqtp3YKlQGXmosCLz1sQmuMxpXX8TiVH1n/jjMFZf6Psi+WY
mQYmxFvpxpTiZZEWdoq+rsWhEWvBUjim5QiPgMh8dIax2hjSjjBV5Y0znDaEO857lMJWi17FJfYC
wOWXgIdG1iQVF1cDw6Knr+CErHpnaJ9jLmm3EvEIkNm12wzNHRxrHwA2P6hX9Pw8hE3i6Eq2lcGh
/LD9k53BSJRmV/k7NMx1OOUyu8SjA0WwuNxCMSKVH3n6Yu9Y+XV8ofjsWPqEk+X+Uxid4wr2fR0r
aA5w8oXVK4dj1rm1gmPJWijpFf4xKbCZMF26+KNB2laKSSBwGGIQ4z6Esukl3c66Oh11ZcUO+DG7
p7t/KKxB4eTY8zn57tTXaJef63TbIInyryGA2RfeJP12glidX3lZ1CEA1j2iD6OIXyOIwRKcjgpR
Ww1TC6tC+BKME4cogjsPiP/+Dkev6AxTTkqy7x1+HiK0/99zXwHoscA7IMGGMuR4xGd305xBHvSS
++PfkIS3hEcW1trGRUzMDmdSzGP179E3XYrpaPnV5+JimUxY9kcFER8ENgNetetAK6QjS4kh19CE
DS4/YXa3g4k/XsvDlQ6S7oOgA3R3F95797w0kGjKioTd6hGvGsy9xLNMilBXIs/aXcY9MhAhb0r6
M1EHeRSLgDAf1RB2sWBaA3zKZuFVAmdCYOpVcFqhJj5aJONH82jY4derU2+5AyNdb1htiCncgh3K
kQiP/xohQIqsko/DgeRXmeEgBR8mMZBbh8OmqdbLEBrT/BJFBYpRkONA2aTd8vY+p1vowUEUjOij
4MD/haeNwhT8J7zl+iBWcyqv5mq3CerpKwY4+JkopSH2t5Hq8/oQtfeyb0APVeZxxdraVph3yX/c
19EP/9BYmNgMYr41SwKXddKqm39G4C1vxl3M69GI1T1H37WYxuHfTb2llWhDBaH4+Izr7Qp+ROno
O0+vi8dp+mzn65ooKH+cE7MZ1EV0GLaC5nZ0fMfHt8UYAHhm/xTwAfbMJQC8gwEjVBrM56LZ3S8G
9JaS8+u2n1QepNC7gj4ce70dt+Sa9YY1WN+kumqK4wMf9BRlb1EKpgmTXkalJlrVtMieRvka6KXz
AjgLQ06o/UdGOEj0Q1MJ6zf9jOW5xe26xpsWg2etFbVx0INvBzoGPAcHFRD9J5rX5fyZAETLu/i7
mu1CPsx3NtiM8xAp2/5t2AmOgnThDtGNFb7qUerV7u0G/9UxJpgSrXBLWTYt7ymEerbkPXfQLq3G
bHDiDrhaa+l1KhNCpRDa7Mc4yUlL+hoNPd/qu5h8k1pWnhU7LBrVc3oUBBtGqDl7HTsGvgF6uL4q
RwGOgQyeUbnDVV5Ak6vXdtlzn5vh3c1KVA/0G45NIcO11D+ObjZHPqIhtVruH8tG49K0k3ScVjaG
I23C5KzOMvCFfimidKc/aNWAqa7ClBqRiBJveE8XcF5i8em94Xp5EA3cagsc5/+lSbaCA5nHvVm7
mtRBEYgMqq+3GzSsgmcgzYMh95pPeOGV/iwKFHHc9uDbv7H6BGjSgO1yIBdfddQ4CfVvDlBrUTae
mV8yO7OTWcdvZ8nr9+pbSGo7SggjuFgwA0a8v0Yw/DtY2gvCqo1TqxyNhoZ8LETux5jfbIQ6wyo9
EdHKId093NUAjae/iV9+rsa5UG2WsrMu46c423jWY67AqjNUCjr3L5MsvY5IcG9QNJ57rDcedY9f
gaTydL9eRxDk2RzmQ7VOoaQXhS7dU6hvw2HdLbgPpWwpj9aAmldETHsQXPVH1DlOAlwN38O1aaKv
+V0IdmSsptrtw+AON6ZkklXtFtkNf+o99SmdIRMgJtHqMvZzYOKPXngxJrE1IbITdiiesytuIxJ0
itsGcP7kKJSYCBhRGrlN2UpumaikcjGiq2j29aKtsyBV5x2c2vxgmZU8f/O5GizpbwToWgPQ0Aaq
PHrH+pjNTYsFDpmxooXaQsMaDKqpUOF2x5xemmAB+dHmbi9awjiXcclzjROE2xJLp9nKHBhXKlbI
0dvNG1oCP2wslwHZIe+Ou8wH4vISrz0kFjrf9gOu6J/XKO+CxDEMhKq2nrw5uXveh7i6ZRKER4Lv
NBmxID2zggkPRI6HxLU0+FHEwyXiqCtwyuUASXW6B8ltCtmVw4yDUO9ScMCqyZsUUGpr8yjaty/t
s0uQh2726wPAE10cY9FNm52kSsPzjvBrT7lEoE4y3Dqx9e7Rqj1cbBOcStZtf3TyOTGstVOadJWL
zX/Lk7Fs3IFkHG5+YBYEeMlPo+oiViR0fWIXsigg6wdZ8wKacJ2n6krtL0Fors7dp6+baWcCBCbQ
yeLvljzc+z6bx/2CSKc3IBtcl95y4UVwo6oOWDsJSTCedl/A4IvQndEobjpvst5dQkjTIo0hB+8/
GgVAYzSGkgQGJBROs/JfMJC9Oqh08lwhPcnFUPvOQlqEBK8foyy/pa2+gKCTTLf/XmAEIOokpfDc
KFB1VnZV9C2JzRx17Tht+xSfcTwD5RR5nhnMNJe4f9iP0FM2Rv8cLNv0XBbUWh2jmc6fewrEOnt9
nlfkrNsL+ZbMo8yEaRkD3Q3D4AWpK+zL6/i/pOMCcbg5Vh0VR80s1ZCJ0lWAU/oKJoRc/9YcI1ua
43HHf10GvGhDs3jpWD8BkttChX1+nrpf5RMzw2Kj+SL2AHKmrbWtgcMTC9QHYD7C6wtzAOCcEtTf
a1GJqNEgYWK8b3kmH6UFk1Tfki7ng07/jOP2yMX9qqtreUS9PeEnI08w661sBSr3+v860Bv6cbBB
sQcqlxkpTaF6n7dPYHafFWnH2u7KzyL0igHXh1br0uSehBIiy5l2mq8V44tUpp2VKve21Wb4VR8s
Igz40zqsUt0USVM5Qt26T0Iqao8mtxpfL5K0FGG0AJ750EKq07ZJhC+cwoMqUVbg5sXcNeQzN1rM
NGHqR2rhRC4Z3q3H1OKD12iwawodAEuqU51S1OXuP3dPBt12U2VAHr6kk3mljKQX3dPLfp8QE08o
scHlsBNLlHhLBVcgDlrPTWCbzgPtv0jy4tE1/g5chwtKeD3oFrstLKBHmQxnxjsBaULH1/wAd2Iv
ZojJP+sRD2osjpBvfNhWtBfbbPSS4NDxjM7QpY72WtRLgEyTOzgbNZHup5AIOsVw0qlSeevnNQfF
EQQfmB9uiTS+s5n0Bq++N+qIGqVOGoks72b6omzaV9wfUtWSyYGAsBSfMCEWOqegqfoZDETD6wfH
7Fv/g2SA1l2iCt+b0NzyzlbYdghW3UD4ZuZ/kx/gBaG0GDqNRKPp+jMz5kt/+N/ykOwZIYa++yeP
dw3PuqyueUBoOqRFV5QrCuSCUNip2vou9D7BL1IwMUz+A8oerd/ki6O0A24hg2ThlrLJnkzML9HH
pR6YGLnEIoV1TAVnHMCEE66FkocVdI7cAwpKSYFbVd++wV5+kFTfVejQdLtxYvSzkK3FWMXZXIoY
kjxWJaR/vBdYbdJTASZJe0//Pp9grQOKW5t7FjlePigsUB7LQjXUaT9uxvHXH/BJjCQ4TlyEMcqU
jp54csc9nHw1yFGSSyohocG/KilmFHqUTo4QUKdC6z1hh86Vh2e2liCaWyvFAsd9Wi1G0hQjYUJS
cW5gYHUi/DT+x7ICW5rXnPmj+vn2DZxCeU4gSuJiZVbObUk8Up9iTpYo6kYe6ESSA3fkwU4aspNn
OgftJQGEGILZK8nJ5IXOFoRCbmiQgr0P5fq9+JkbcOHVlc94J3Cohug7nzMkg3xtM25DfVhU09ks
FHAG3esLpuMmoL70n3j7DMsuyJh7NL8fzSRSEs46uSZtwBNvwSeQO5kFAZvenC50p6Kj9oJ+2Jdd
XtXxldgJ9DufVwzFFZT9FAFhnDlj6larOC269DWlIbwX1fsg36FJi475oZu+b80KvqICpOKrPBbO
yiCFgAEZKyE+QXexNdjNy67nTJREGAk1+qyd/2ldeTrKMgBDEknhbpWdb0XJXPGEUM+/z2kVmWbs
p6R7cHMpUOaqNWJs1rDf4is2h1m6ySRNQKZpHuVfWaQaaVQcVQpb3kX8Wp6pmt4+y816KSb4nq53
Rr3hh84V1v7nugLmL+z9uXilx/89OpH/mYdAQkZNwYywbQ28HdHhm2BPkaiFBQN84DBdBjc8o16Y
0p2YWwTME9efv8IsOJffllc/Tr+I808Lj+Mq+2tH0LiRFhqfA1ifCS7ZizgOvq4eH/GtVGdGss3T
+4ps1PphWLEwgfSFnqelxvTSJlfuMrOGFVJ1VyOgnPQ8XP8vW31CNF8VC0hLMKkGd0ThtQqvsV0s
TV+G236L9D78z8gbnfc3iGadCFg2g4mUDnKWBR8Pa17b13zlikmkj5uhXcrp0BwnoJimJ4E26tF/
o8qW3O770xkmkXt8JTpt4rq6FvQy0VI0D8RMewKbKuESHmU5x9kM4P0FZERF27Baom4nMMtDZ+E1
29mGakF4ZP2e/DpPnvnjQtkm2/KVKv62aVFcjf69kgFZgrnTC0PyCMr4s+NgyrnTPFoQ6TgcHTLT
JB1iq3Yyew9KcPOQ8SM1SGyeckzd3mpcRlJyTSZ0aZtwPbU1WYNQuBDJRykgQ1et9jXguZdv7MlY
g8KSxMmk3k7FelvgB8P+4YgsGNoUI5i3/Pt8Jf9NswusRsOOjs12I/CykIDhnALXmv4qFzOzrk+o
bOXnPoGVhKexQfAq5juTSsgfWL67J6Z7ms14193Dsp6ysiVnJ4ZFtbO2nB5T9N5GvMc6jyM4ojwY
cOfFZcFK4mUPD6XihRV8An8lcvCL1tdPHzxppHNCJYDh3kzGwmF2CJxSNKPIBMtRigKmurs2F5u0
ND+TiVjLTVrGztkrKBVz1vH1L6Mo4baL04A+MjEONwMECeUgyLZ+nHHMZJeKSKiG9x3MZdS787Ez
Q4nLZcuBSaGCWEF/87X+tl/DkM8WrYUyol9yeh4npghco9Kk+S79cNAxsX6dRV6S9YZBObYk9NPJ
ozD9GPFWPVpTUe1sLIqJ+AeXVbZbxBcnlzDIIhsmB5SSS+Y3WaJJtrRbBDCR95OGxXo8TVoS5JLv
BPulym3yHBWlJVXWj09LdXBtbxU9nLHHKKKCJGu72sFrs81XzRL4Y//UT5vD8TVzWGT4VBcZEgRm
/RHlxpug23gLmdK4E2SF1B1UZHCwQ4p/Wfu2XzcsERx2L/dxNq4lZaTA6m9AQFZsJc8XjoUkoku8
2L96+DhmydFrjLtVC/MNrFeBdwdGCIBaXrNls7r/aSC470TLict6xTPUSGKNiMkQiEUJE1s8g9Tn
HUo01+LJQ29tzHh9a34EwzOomsuD6TjIFiUi9hqylOrViE+9i+Fj0NYfkfTLbLbpu4wp+tub04TM
wbrpI6939Ka8pSJTjMNTKksE583+m4SnzwcIdFjer4kp5p2K1UZWfCFI0T3EHoPE2GSmaHHGY2sE
BUkDGw4ziXV8kemTAV697OdET+h+yMUyEXt4ODjimROMBxGy4pZFbkPM/ZBJvyFkzjEny8uwwV5P
M+X7eCpx414UiyeJ0rq+5wiSW40UqMuV61Co5nqNhNCXhVOCmnYchDUnzudHJB5l+zDdYr16bVQ2
O5T9JlwzvIdK2bWVZXXY88JwfPwuboWyJnwAVKuhaXOwBZyXBGuV49F4wTm2jI76ZJ/KiHMY0MN8
3K9JzFSKotYcRzvncK4xLpr0m3d8qr3WnZcyitVUGLcTO1+cCFojJwkXQSR8mc2gwS2IPVAOJSl4
snd/AQ8JQDipHUoMH3C6q2m9Rn7EYEwU/CAEJhcR90TXOvqgp4c0aRYsN0cIDmJ0cqk2xvlet2dM
gJMprV3oT4A7av1s1/dJFFNb1pEm6AqMjtUWC3ssm+ld2AKeuHVSVZtfCMTcqVD40IBpaet24mxI
0BhRfDk2BzPYM8nwHIXTvr8K9HFSJ1k9VZW7D8tV7SfZ2UcPFpyUu42You/sS8WQ2GDV19cndqTS
fvMmE1I72thPUR3GFmmkeI0htjQHp5rI8GWe6zLt5b8OppJZGhLOuKf+383w0cdTvcXT+VEPyu9N
kLbumeQycvdzapwCVllKmp3se5Wh4B/cNtgqbtXrX9bTto9n0190RSbddCQlQnqkPcEkCQKBF4g3
b7QaCz8USxwbakoRLjPjxGJnuJ2C6/Rfq3ynYkE3/YnKQepW0NPmkNV8wQxyrs1Gp6aQgTgDSKzf
Bci0kXYyyiuKBh9cPRkLKbpsoZN5bW56oqrcXgyw7U38gr6lF//9DLHC7OD8I59VR9/K/MVjYjEv
SCnZLpZkrwjZ1Buan9wzL39i5+zpO0CXpeCaLgjQ8JaADCJZEY+5H9Aj7s0EpFwDwpGIDuyEaEeA
OG3tC1aviRZWMKmf9VeNFCKweO7A11KKUmIRJ2OZpUMwaVpdNYQ21+h+/eyDZJ/ZsSf8zP3UxFrr
0HIr3B/3t4J60pVUGtPztT8do4T3XZne+TB8eERlDkavDEW31hfaKq4nXqokGWPtr0uNzorZ4sL6
vCFp64krmlxA55f60oao12/9evCWBkPkh7P3+VbQ4JaekB8TUlz5QZaPEx+yw9EfU0X9z0aHAQ6m
mPklgGz3+O814harjIfftExknqoyblsjHahqhS/VR0qlWq2bMisIuv3NQw6fbnajubbr50hwdhPN
lzkxgN2KYq3o74RDqXHJeLM/ZrFi3wi3ZzQ/dzlyk2mmid8Mx/4iAy5uZlUkCx01DNI5w8J3PJ75
hirLLiULp0biV8vOkisk4elwucehDLYowtpCCX1v5jfrNylUoHK/G/WoktMUYLydV2oyC/lUb3A3
Sw4UKMevvb/gdNL+7UqrAlpaOhTOYAQuwvUp/IZ0mvTKUl1Q1c4TBcD4GFcNNTFxN7bB3bYAlLDF
cQh1NJYOuNjSGKhBGaznmAzjTo0Rmq/OaXZG6neNB5EvOc9yhfdApiKFB0udYDnCB7KPgb6S3wTT
P3/anJdPK1JMWHqjNx75U5lr3tndwKjbkIl/niDI/bNDDTW/7TAog8DmHifWJxOCnQznhArW9E+s
JU1dxCAFZlKCS37DKA5h2ujeS2JaRG4ydFBibTT39OLWXFxu2F9H36BJbZzuMG1mFEmFmIo1XukD
j1ksP3FOnjIv4zyC6s/SldYGLCTA3+khXgV7B0VGopQMsgvLLGnx39Iz5u+1E6i05CmA15WRjXgE
WBTEXEl5mW68CQu59VOPtJo9BolRf/i46IJDq8b56YrvQbL7FZ7kEDJCzLfpnFa/Mo9Z6ZwhutGO
q+AFoLoYS/JUfe2FpLMwkUzv4PvNDZ7iJU0j/iMEu1OhxzkIWCKKBhwg1lrnFYYeis+Yq0r7FSGu
2fpjY60S2tCgjVAvxBb8llsYslAbFIInDTzJxHg0EhPde7QEcwfmvE4nSJlY38TB/HLsvhdKP57Z
SAGDjWsY1e9BLJFh+ZzLi+nH/WZNbZKDLZNs0uQklfOYgBEuF8qaor2p3ic/Q6c/ZpkaKeg6WqNH
FYboenzrgCOtwQe8ZcnkMhVFNaWX3zlsC39XfKkDOXDA6Qs/slmoVycclRP153QzxvB0NYmN/tMK
Zut9TEUfxKfPKUzNC+2deag+jaPk2evp/1KKCDaBiaKoKMJOnMIchuAQCyuaSGDQ/gJb/yXFTG61
kNw8S2Hi89/HxIthNtUhzgBeGzmUgaVKB7W1VqeZjjThXWXE2dvEB7UQ1KKTBg7ZMW4mMowUMGpb
Rinv7FPJgxXMyhzCSY8ApmL+6WZyRfSIybX5/BSgk3ZEMlFF3JLvYjPgAWaFfYXupTqvCy17QKcJ
AO75Wjk7Bu8Zk/K1rwA1DZGuiHSg2CfGUnDig1gFl/+GmkwCfD/VTnP73wuOIVAzGmj4wZqacAzl
CuEI9/7Td/XGtB+kqwrAIa3fiMtAIr9KvlihyK7GCGsnOZbLTAtgb+YrFoUEx/kWcW5v0HvUhSyH
7Imz22g8imUD8wmwy/ZcTMEhkOl4Jettk7ZGmDUO2PyaMrgUPMiphKxSL+PGSb/Wxz3nwu8WOyjL
xGMJhmGbrO5qWTC/SoEw52XoVXcOIllheiRZs8rhQOs3QKIrcjjsAUq8SMcNbBaGu02Nk5Yjgt5s
n9CJhOPJbD5Kf+lGVOWulIjX/uCmvhVMVMtMaQj6ZBv5L70tbUkP2wV5IrPpeTPH8kxx6rx0OCfI
adgi55IvVFjHAtTXC1TeFhUfPhZpgNFanyCLUBv8vsO81r3lUwSpVDKIKxW+2rF8ZIvIMqk5X2m0
05fBS9DlJ/c2ZLgizWISaSNcMQOD9myxbQ4L8xQ2Bpe7gtd1B0dcV473qDz+7bnbazOXGXlbuFRv
VL882FhCgh1pbaxCYBY2O/I2BkBsezXhY601rOpskSSwtiDxMiShldVHcOTuc8fXJF4yZt47/Mvw
rXk6rlqzVrbVeSzO9oi4wI+Vmw9qoIGSmSDigd7XFlH7GqYeTR0niJP3f9VaPBLprLg/zdU/yRZT
ER9CItrwy6yuwJR6MZrD8dMkIvLNXvWH+plyB5vBqYbECi1kQWkyGDFZOhQf44bC8YNZD6fz3vyL
i4kdS/rlzBHudIIkEEqJAsDZ/nNxIZ4ImLG6wxWeGnG/MB/BTsJWE6ce+5uvT0X3wl9pRbgYdURs
g1tAsLsgI3cRpV9fbKn1myR5LYRudgjhjGiCvMnz/mHlJxNm+g3BARtRooXZ3h43hF8flSBXKmzl
BLjuM2Y/WD5juBHfh6GKxP91DUVfVK7UERhSDo1g+xvzTYvAGD8bjGPnYM8yuFYR3GYVUbeeBo4J
D93B676QuJC00bU6YAhOPANZWm20957+Vssnfcd3e0R9Do0EuOxmvHsSzliiemaedDNJKaQIn9l6
d9CIfn6Dblx8pCg6rGcSptjjmNrF5mmOHFq/ZhHzzPOe/wntgwYrEiyge5o61kN/JM/EOPUI7vQm
rr2YSvbsVJnyJ65nzeSQdipkAdUJtBizNrlWS0B8cQHPkB6xElND9pyUo8jG5hBfNtr6UaV+O4eu
Z7cPN5bzrDlWS0miPZV27vnFeS7py3ksG8W4dKYWl9RjmgmOngfoqtCWfCeoWcJ3+Bu0y20aITjU
YFYfukpJN+FIaS84MjMKRIS412a7eA7LbgSFvWV32K1x4/zd0MqBJLup8EQOKSTIbkkhNLjsr4jz
z1VukjEAP8UA5pYN+mosguLS+Ji8K1utfa0I2sKkBONw338tgcAPYryzOy7wrIUqVO1JtbZnfu5K
yIGtwZTxoOUPBUTwqWozxLc3A6UzEt06YYRwdi38lMBzUFHa/assmLEPTAgPfSRlrBWq3S8Q6tKO
yRk3MNT5QFRMVVi7+Vy8/ggSQI2qeu82/vjJxKJc2z1lqWbnxVZ9BBO6PXZaTHRh3UGKWIabjyyz
AazNTTg3D3Y7nq4A5adoJ98JjOGdQP/irV/f/4JO+yvSD+4BRFjHrUgrpfPyj7C46cGDvtrdoKSP
qJXKdq96QUM62s6f9le0ZBAsbVo70+43/TERDlVaLxBlThQjf7trXUNFlvC/SLZceqXZdTGXi3W8
tkgXQNiShYbUZPaLJRGUI3M4XwxVNrZ+r4aYoVg7crwLmIDtDIEx72YF/qz/euKf3/AdcG+Cgudk
W1GrjKUVjjdv+gOu+7qYX6i7qJS4XtQb/j0J9QSIiz2dhJ8KHcLAeMleneSUlcTCVWokp77Vlmn8
Wjmn8lD9i8h9qPsbme80lh/VBtaCAtA3Qb33bzrjIf2yjgtLQOzvVb7VAQ12G9D6dWngoWbBtfu4
osiSDmEeL5XFMf6u13spK0t80N9uqTJZrqRTtGjCY60WXyzv49lIuzyeXztmAtlwc/M26IfnSu+w
ZFPyfEjwEE0EHQzv1AcpJ1IE+4LtfvjTNDD4RnRuioXz700RIQuRpZsMgNACMKU14vk+bAaNNNGa
iOtUL/a7WU8EsGaF7QLJtmTdPFJYn6QAyJOSA9gtg9l2QCqCNdA8e79Y2GKfnC4Oemuk2TPs7Fhe
i4Ie2/CTcqZyVvjPYB9d+mWtwrkGbTRn7E7WVIcEOJVexahUZiK/z5su6Vgu5rhhlBr9ngqkZpoE
wqy/E80mHcPycQ1/yxhHZ7/M6yRLOw2Z7RN/rqWgxChfWxTUMejVbq6TRxjBWVDvW9fJ1f2Oe0B0
fcadZP7hY+ykn9sPOstIZ9YkRz0gXYaxhn8Qn14UUadAcqccQum+giiHoAQZaGgVpFzT63C7GU5l
PPdWllm8/Hi1QT4R0lNUAV/6heKaZhPkPUqGP2WYgudw7pjXqXHRdN1QFtGZSnFX5I83FX2ncb8t
bBnwFBdPwEpwvF1OwetKZTFo2YOSsYLGVtU14DyyGyTePBXLjrJ7FTYuEq2OuXsagfzjh5i0Ahjt
8O81GG4mFfP10mhmp35id+A6gkSHj0Qw58p20zaJmUxCB6xvG4d9p/TMowpRPJB8zQHP4QEQBZvU
wasTMVKapwMYlDt8PldiKI8Y7ItZU0i1nYZBcxce+8AYAILC5O7LuEkkMf+ZSSg433U9Ll2QSzqh
da0gxZ7wPAVRZxhMLG2IWV2w3A75Znq9Bg91+xY+lFMNiPoNXTGX/DPzEmJm1Y8bxVGRAJcM/hk7
YqrPbckQCYayBT1G7bovVMR56+RV37HTFcDNkuU04ye1ZxrevZjTl1TZGdqCYyNDJyo5mqlBOXdy
U/szrCPWk+Qoj9bTnPVgu6aqYgKiOcYvx7K8+uH+RarQb53m58dZDZCuPJV9HYPWLZZt6bKC0Phl
6RoHC2Yr+xzacpnXQ71tlHdLDMawhTXw1BN5tdqi2J81US1ooIV9PYdCagDklMdR1Nprmt7tzE8U
1vkNUjtbSeamEQTNAe2b0GAfTrow48NpNYtJBooackDAsG4NeLJSKOG09v7GeDmo7tFNuuaDzsi/
PJSwo+ecls5JWtK6VAdIhTtXYfN2fS8qIDCISqEBRx5oGYKhyn1Ipn9YOzsnRo90WJGkmknsDnbR
aYrHbjph6KSuT5VMAS9ZslEpuC15n5Xt0e+8r/tdZAw96AiNJCTDTFdISUp34+ECtF0V72lMivzt
4kTxquGQ10BjHbU/v3R8rHdctvPqSJ804G2GtqpPPoPqUau1LTrzB0ek3dQDoCOYboclCs7qLknJ
2Ebym2vIpW7WmwiTn0xMy2ppxgG8gNFspjCEV1DxIyQm9t5hCCJCopCabVd1EhEK3LymCRoLbrni
o0MO63U/PGdKkjrvHh4LgyeQiu4tUbwpTcDD/Eo+ICAPDmhoeIMGkGEdOuaBTsH3VS99BxsFl+2E
S/agf2M0SPRlnwX7UfT3H5aImwLocO/wieX+kKJkdK2ahkiWFruR6G8/8Zl40oL/kuZeUDRsLBIx
vTkxgDQdD7ZzNg1VNuHdHWXxlOeusDjMfakPa2gzPqtoBzezVmtJUmU9wjOdJVcuTKKKyru5Dy0D
hI4X/KiBScT5sr45dJECZBQjiCGk0YVhsBpRFggoFZ205MVQ0xZkYSH5ifjOqch7qBO+GUnzkC+d
ek76jdgn9am+XtdibGpstEqzRrWOfvrPf+cgS+olZFAKp5YrbrTEmJFvyMZOFdprsLViST/qesUW
hirEMkzmV/7zt47LDxy5ZDWAj7r/fOiQzbnLuxWRNMw+dpxafKbARdvciZGLPb4qpewXXBOPSCNR
QoV+tfD9PMqMfokcoqh4N1lwwO12ApK11lFGRKcNirTwrpQ9axjDC+Ul5+hlgYr7XtmiE2n7kktn
4cWS7vvoP5Qb2UXF2/t8pvN4PredQGykLwoTttIcCR140bVX9eUjNiRPh5MCae+SqQ/rqlzVfTMT
yjO/SlWy2cG8a13A7UKOEDsmCRKUDn8a7sxOAtVfVP0g+DdEucvrKsmeOF+a9ua5xGLmnCb2YAsa
P/5Q5D0x8QBV78Gqf0x2/t5mtaMF6L+452s26ur7M8ImKHdDhTY+6qN2YTnK8V7kdhwrcpKCSBP0
q0RmqBxAz9uPWajA8+rZw/aP71i21FVb4RvnAm30VwDg75RKoDrKyGI4haNSMMt3i8ptyzOKGzdJ
tHVF1ACO0X5kBVwzgDRnkKK51uWzaX3kJAT7RZCTSvHEV3EYJl13EkuqFR7VEmQbgshoS0lbBIfD
KTAvUEFiOj0A2n4D3Q8/Le7T80fTLrhYlDeOojI6+iN6wZUBkh9BDauo9FhJRE3DyQLGL/YahfdH
peDjlfSgPEB2pvy3+DVCn1jccEcW9+tUU8yNRKh3fzWY56DzNKmvcJhxPcnlc3uwXn6ynijmIM6n
mgjuHNoEOqouNey+GKGJ9/cE7OiOY2kdGwX8u+NHBT+lotOtxjAHOeNT9uSQm95oh27M1KcDWFLV
f+h+YxzdKHEd6qX2xTqB5fhmvdJBgBAC6CVDuXbGmN+1it8QHUSlYZ9KQCXocDUmLHj4LqSi3uZA
Js4zXSTHZLMRgsumg8O0TUSk3bDX4sppJmXE5KK2iITFQACVeeRCpO3NTX8GR8DFFpu1wu3tRXxu
RvWJYPogRYjq/pbQ7VJzUF76byOLVUSCAXpgihxuZy1VyRNFIbeGDHMraRAV1Rd1H/dp623Hrr63
sLEF89c18klSfGlDb6IiIJU+7cvxmqGDZlYIFETjWjNFdQE3DrbC4s+hED0DkVpHmpjTl84xUWGR
HEIha/lj2d1ykscHncr678yyx1XlJ/yPbJ2ZbYLPNkubIo2j1rWKwbIBoQSCnOefXJHO6OK29Wwx
tk10fp36UfiM8VjiE3sBxDWnNimlTmqW8K3tgXR3VDIPA+/d23QWT3ShZ50fhfr9mYEpjdy+oyLT
x8lc0UJfI1wFNkWJBwz+FLuk/LXdeHaxDB5/v9SJx6ZJwzsp6yNdPMGataz8DRSwvv4/+qtHwOvU
m6dwbFrzFlTOcGiS9qjVQWDkCf3HOKxWPhnhEDRbOCGR9tiNRHkAB+qFaDU2Iz1Tbb+mfKcWmuLx
HmDmUX2Yi2agXlS/jqHaH+E7mwzv+5nf7gM/VutQLGjGdv7vh5TB14YYvgQkW5mRTDER2M3yHOK6
B3M33yx8lgah1Y4Ma3UEjtgweeRLFaKTgth3HP2GwR44iKT3e3daFFbYuUC3fdc4sGT/BwAlnUKw
KcFGihNSW7Uj+ys23RmOkTA3pzYR5/T3dsJU/2b/n05m2MZO3TydUlZzHyPK1zSVi6PuKqgUDjzp
P+7h9q9sGGMzpmqVZpsbN6SGrstWQFzn8kQriN712XJdN/61cy3NJOGfZk45YX8HApBSSnx9+2hf
Ekq5Dwdu2bYrxEQnY670kl1yjT+ENFwkRqcAV5nEWOvM3W2Kjbs3ECkD1DOW7l+//CaNL/NONuTJ
ZLSTktvp0a5v5kU3J1NszpkQqxSgxRrCsn+T+ya65Wn+CChF0vsUdFftw9Q81b7kvCPhH1H/efa7
4XmD3v0NOAAIA5XUoX0GPQpSYLT79zAI9PIH9KbFapR9nb66v0Nk2lTMPCt9tseCt6kKdsSGFGNx
YNd30VyDOc+S6HFp9dT/kOi7fLMty2UJTUvYqK4B7yt+7BL246/TIrdtOccNml0yPIEpFSW7BvlW
fB0UYkXiVowMi4Ta66JKg45I5QyooD2zKM3IzxeAmhiSLlIxKqMNSdd1iLnlpGJrS3wcC9Xq+zcZ
d2qOuTYK2kF1eykSIyD7J6Rok9pwxoAVLskYe3ooyAhkygeg6+UWHNqPckHY3zGegCY4Mbpu3IHb
iuy+pls1/il/H98MiSe7QM/JdT7ph28oGw6finzcsUNF6SgaPxNSGYHUaL6/P+kkCBin402m/1Jw
BQ1Hhskvb+3En0qHeQ4Ovrhgh8hJ8WHkRYtNfXB8odiczBdnny/aQzMDNQGJZl6oghx4OYNLbRjm
bvmS+2jywYu+neiPGPbx2/9ZwmlFHkpJxJZ2PxUKayqZ8HkDTQ1PUCOSecw/1Y3KSFYMyW5J2Vhd
GgirhPoh3PpILiqrl9cnCI5gk2SNUMLiNQyDFTRaRyRdoO1T9p6S1IY8+Brvm9uvdjgH2NOIbdoQ
mM6gmWdyHCR6TasUfyqIZfRmv8W3rJRhJ6sOUKePma3M55I1soJP7hyn3jfX/a01tVqqvrEFDiOq
gOsaCaQDd54hbwXYx8JUVf8Gms+Z1bDMYkVPn0i5EByiHd91jfguhYsThXkP83pa6Qm48c3IixAj
Hnp4cM1Y7TZr+pMnyf7kyUJlrDgmxtO4V2VO9mpxWKKO1yWGtUZnEe0BsO/ch4Yq/mvgk8fjFK3O
sEgmPoaDtLfR9sJF9i0ZdCBID41C91wIc7g/APAtAu4EEFfNXCf96ByY8DyDboX7dDnduVM1ZMKS
kE9hP0gcXIaYe3lC013SHQ8VxFFi04whYlylYuDcHEjPTBMI+MWp6q69Qe3CHgVfp8dgAigaDDAk
R/ZbmMQhOr6JKZcvzs7lKRfA87lY34rTvRs9xX5a4Wo3poaEuxsulgRcO5TB9gp0SloTRTxnlRpF
ntbYprs7lnmKtdyY3GqAk4hIy9StiOZ0oYjmGWiKhefH9q3zZngjCC257GMojObAWferd7A+kePW
Wz+lLFmJi9Vgn/M1q5NYlvg8LxGTsm3nSdGkpGwDxiUcnn8CJgQ5Ozba4d4biXqRrdwmGMmHm0WW
M72eqa0UQt9nECwXzlbTsz0qFhGsJL6h+IMKwVKB3YJN84kYC1WBVtUHDNv4tW6UBfqnQ0zN3fqv
BgvYUIw33D79Y1urCyJj9c2r4v6BPPuh8yuxqBu9UHVJ4Zu9cKe9PgYu9p1JNy54Q+jMwVYeN+c2
g+MPG/Z8hu5VUJwMENID3oV+KaFqp0IFrzLqXWn5mffMwaul+80x0Qih8B95jZ27PokJAn1lYpLs
HIAdGWrzgKsK2y2s97VUj0Wf0+LjgHP+wUH4fH5JbBZWcNGhNdiWrHkniCDrI1aIIydADIRBJ+nd
j9/cPzD4UMX9WOei67gIffszQrNLh1fFtRWBxQkyxB7MXOVFJPFFDi1DoG638pY1OM199rRj0kBb
1GdwPlhCKpLy9E773J5d5FgLTJVM0F3YmV6m1voywfvJ0Yv7nhjLn9w3Ce3bVGqhlTWTAYQIRwwJ
8ohj8ATDe3al3pspN5xFcxp4n/EWIXDtubYnx4pi93Nh0t1F3U1rl8ba2bnl3ZPYurTpEcFroSgO
x9/ole8Mafd52QjebPlPqBqagau8fUOPJJIRLKEJ+E16ZAC2HH8xK9wxX2v/Z7L8ghJDXHMyGfBv
4JhxKuFZwTiBSZgJvVquSXaWJvchRDbjtC4bBROt6j7Z/rKCwRCEwmVYo6DuFt0xMtZ9ofXihf9s
P8bAT6TmTyg8xwFVonKAGx4llDBMHXXLNmP03fPn29RngTjamHaoG6Cx0wwDSXHzhLFJD7bZnhD5
NXAayWNoIA3FY1HbDFnaRYEo6a19GoQH+Pc6QjAe0IsQskCE5gXQ/PxouP5a76Cdp9lQoc1MA//B
oTKSWNSrDpjHHlOMlo2wkuq3P9WDKArqJhAbAUkxqCo4j8jlx1zVQozKPPyd4FI6w5o46EYDke2w
ehqpx5ddhV0PN5xfQ9PNeg7siG+rQyOBs4fw001jPdNO0mKpQsryEjo8hxEuiwhiqEfvY3y288MJ
pSqF3UOQTJeD8N5Yt92flvJ5dei1uHuED0mYQnrUyjq6zyaeztMM5ILBKcyjJKdBIY6/axjP+hDS
767s7W+C9DJz1TXf3D27Ezl/KCkRSXkLYOeh6Sp4sVqP2/Ia/zwP6/qRmXsL0BByTaizY+TLgVVq
VR3qpQ85AEIqxdLHslb7JH+pRcwlo1/6dITKz/d5nb1UY3T97w8JvFxCPLb9vFyEIun3Z50J1wC2
D/JkXsI5UemdOdNOl1h77LT0UqWJU/XCKLYVJ+mUKquEdCzO0YJUvH3ws2jFYWyFdHhAfvfnHM1A
EFR9tsaniIHZH0zEDywSObIDHSZOwgsYvYKoLjf55ryybI0yMvI+XMLIIn12NgKgsBHsaXn0kWct
m54IOVzyuGzQnrXIhakokAEWGkYpWxSu0coDnM8a7W/iuUqcoPriVWO4kkQ2rKyjL2ghRiV0uE/S
/vKbD6g3epQlX6dfG/0fkbrACNFhf+1w85rlFyzgPcU8hwg2H/5OJuB+KPdg0b4XktY3mfa01PO9
qpsMblXQ4mdt4INYe5ZO5k68FjuvoDmxEfKISPC7mMjFDqjRkdqAbPfjbRJRdiFcHg1NtQzB/Fke
y4D6t+04/xkKipjmMZn43UZ0h6MJSUMrf8B+jlWScDEMrezizJsvVNO6iiAnN9xolV8y9h8ddPYR
ExouGIEg2OomjEZbj+bXcTHyN1LbJTIQmyJcDG9U13mCXmYMr/3nIGz1OObs4e2DQJJ7Ii/CzOVv
AdyBOt4CXhq7spPfNb+ubn+6l9ExE2PCRWm95Rsn96Ut+kA7k2BppKbTvSv7+OD0NMQwqLlrpwAI
Yhgivs8pCgbZxhZ6gWaURgxqfmIsWB/DHMvc2x86xAhF8unURcJ4CU1kOIwU15Fcj4FRHLtUY8BH
FgcqYzxHqhqulYoCuHtRgW3L64aQVFyvgIziT9FhOsMrePa5SlOpDheKbSppiyFJvFm+7rhs7brD
33qQ6ObD3Ve1nsjt+v5CrElhdVWB2QlFBcWRNnuktxtFeSk8kP/xWXcUhEvROwX68A52UAKP5Enz
i8MruRpMmuBD2VEUA3k1cmnebvNHeqJ3H1/zkl4/vg3YzCrXKRs2taFtgH34F7pO/B9KmswuJJim
7+nmf1wvM8NHmsxgnogbJYx6vVaLRFpIUBzYOIwPxG52y4zdmMrL0sui142Uz8J5G1Kcf4ShbFIk
YItVIoMepoDMSEsEKkJCWsFYgCOOXaLZX5/oVFDzzL8Kjz2W5RDHDxm+WSIRDdrVCNosCK6i6BAF
ltv6SxWhQJkdgwh7U6h0eh+BruaoAedjcKAEqyhjXps7Du3qc8gZcvclQjBpC8D/TEadZpuhZeGt
RxG/IC0oW4nZb0D4SH0ZlL7bZrztNk1+adE08PIqEOtV+PaOeRiqgbvQiXEWKtkg23L8LE1E9Fjx
uvQgImwXMG/EQ1qKuzNruQYYVN5p6SqXwernIFAPVhXke3Sb0D2NWSdsnIH1n2tRrRdyekomQ9uB
Dh1eJ1O+GGXsRuyMhtPDlPgGG+uH3YfVoqwE0nAfCYrhvOcC8gBR5raveDRtRplnVm3Eitwz8EZn
/avPi9jEA31MOV+qeXZTllZT6ajYrn+nhS6f4GdqQB5JPlwKlZMHboqzvMK+DJPYEt8wRQyuyR+5
YjuHLTFN0z3SwxJOXw9n2wtwE7LeH1bfPoSx+rBy+id/Rr1l18Kmuw2fImEvaojxxy0pKdOiVTNy
dQ6nxfKrg1g6NTx8Xjah6+SeYKGliimwm/C138NBaK1HUMa+mv1r1QnzZLaPRYY4vJGtSYHyq508
S7yX4MSZmoVo7nZeq0o2zBEi1STSdG/lDpYMtk6V1xcESjcrXUfK+gaOLRd7ywJezGUNDs7IHuLf
L3/gEabC7rAAOayMuR9VxsDmP0fsJS6xm+w0OI6JHp8WDKPT0+ycUg/pj1eEbt1TQRmw9QISahkB
wK13OrHlsQq+2vD9xxHHEKYg5vL29XAh3K6jXvVlkxIzru883EkdWvg62a42C4IIxu+2I29oBZiH
krFlqxsfoEEIRVoAQn7DFK0/OVIWTKLEyC9oSLeEjAYgFAZUH/WYmCzezhwVzquIbM4BjJV3Nw4S
RFt46NrY/G/GSo/JgBfmZC8HR6oVFIUCGrvD7/rEq+R0QYLBFIkISWNoGYC0CzMqOUagEETXlBCU
j4QDyYgJx4pXCEu+Ilv9KxqbCLIGevDmf14U994AFnphx9gwB3RPAfdQBl1CsqlAXeoNvcbwgFp9
eFoRdK5QlbyEn9Kjo9KI0Y4yDpx8BlNBDE9dl2CdkgqyfeGUR3/DLLExtXro884eaFuTy894HV9C
Hh7iCmQgrfOBJ13IjoqPNxTENfoLG0FiY/Dy69WXgGb6Xc41T/NKIXE6N+r469O36FUMkJ0moeKA
XiaTM2J0s5iQjqRvfvEI+rmfqj+8Z067YnbjJbHdFp4yPg/J/KkxleLcPjVaEepd3R3s98QzL+6s
7076Kc29v1uVYz8JhKSFkBhiWc2qgDczZaev8kxLsW8CVRZ/8DYqhxtizPTHMcWAVK8ur3UlpmcN
fSvrgZXHe0Y2T2BcyMeFQe+vPyecBBPrfLDe4ls3gi/OFfa4De7ishNNATVZLgol4y0i7sKHttiW
V/cPvfwD0/12nNjL4QEhD0hVO7KxHM3PkkEUoshCQdNnAqc9YQlExydpuqqdPHhvukbcOe1uI3+P
PhQNoxTCaVdbncBvwkOMyqM3mOlhXv1EXGQkDGhf7FO9eu7N/qTDZCLxM2tHZJndorBbs85S/mk+
n75mkLsmCNXjg9nvB3pCtfZupL1P3vqHD7i7Zz+PD3blZgLQQJ9ut5WfnIrfla8uv3VYoIPEAiKp
XuZaFy4brhceHL/Nh41HHsQZ+hkYOzI3RaWusiOwUrWTOnWOZqVajjWKRG8KZ6R8zzDO9wpwkkuS
BXAz2NgzJcCWckustDVbbulKqfRN1pzKxdrZnZRGMg9hGBOJ2WNc66m+0blKFAp/9KuXc4SjHQF4
CEbVDuu0PGfm2BW0n2WN2NU47Vm/xwaxhVUZYQxuyp16euVQwljhP67M/Fo0GVsyVNeIpEa8WIp4
Kf6bq/JcHypddIBbEdBkDQIO+OIfBzkm6jbvd8LMEFO26bgdGAxelbD0OwAgoOEvhhcscgMc2Bq3
+EykuPvF75H+2AHMEHDdBOztGIjS5rUvzDZTUonOGeCrnLaBr8DfzDKDar7BUpXjKwGUQxLNO5HD
xwu0LF9D+3P14PxRzi+f7Z4cdd1GKgVGCcINJr7605+Cn1EmzZ4GmRQDL/JnE7rJ1mCCd8SV3TJC
9+hJjk5e4tN3dy8WTyqoT/tJdfBnxT38Dm71Nq6S1dD3/7Iu8rjFS50Tlws5tCZDfTi44f3hNMDA
E+hDA8wVq+UBLXpM+Mg/4P9u7cvFLk42xHeUxfMZrDEMGWvaCK5nExVbPvg+a95zumHfn+sloJnD
KMdexzXHmkKwzcJBCG2A1JJMKtlwlxjaYmqxFWuntHuZX9XzH5xgsZqVrxDx8QvMllgV+5cE2Tb4
xJhDO30bsULOVpVPGeI2eZnuP03p/AYjUa/zxseoNvIVrr8lyzkmb+Eu+TiS0KPKKPa4KyohIcVt
hOI4X492Oo4TtpCd9JnsHV0LKQ8Vnx/hNGh97gAtaFkaUlt/DI4E5Nnv3dCZ2S8niQt53wYhk17Y
aXgHoThPU8xFjXOMK5u30/BpeRGXVQjwggHKvy+bEEKLL5GglNx6hGbMP0gV+kML1wJ3jSWWeUiY
9IJvmxognivKyWTNHQQ+wuLmeRNROx/O1+a5FME291+9pB8IIFC6iZAv23qh08D0hLPL8roXveoF
1lNDFj4d4eBhRI2s5ieub7Vogf6Lym0aMj8Y8I8oVqubdureh9hgEYci2nKpepn79xYCTXCevoYb
MeEIkK4Ksxz69AjXC43AB/BkmpNT4UUe1Ln55WXow3imLRL9LPZUK++ABSDVW73S6Xp9XSTaUXln
clR70ahqk+xnQ9WGL0rp/rkCXnIqTS/9JeFv9PiHveh8evLjKzHIKxbjDH9UezL1KZdDaU2w6WS0
48R8y0z8twmE7CWA9slynj5/2A/SNZrgzj/qtJBTu6Y7gslSX8JPHV5eUHH+JSa+q8/cMgU6mssb
TInZYMh+fkyBhdeqmS4E+Qc5IYtsxAyztw167xk7GTFIsa3H39Yjt8PRMU10cYNRxD/Ra6VSJ7E+
aA3sW0xthrLVKFE/bvuoGQd5RSPd3ch5zB96nNWK7W911clU15MNCh1Mi0bvxOYxoNva/qvGGu5s
ijeH+f1e0LZ5qgbZyPinLVsHqf3kOd9p1xaczU79VaTDe8GdwUv8nqnyZD2HWB0hb+N59pYe+Zk/
/Ub8ihq0upHOrXefLpdgiSO4mIbecI0pt3XJBW960GLB23R2m6d+FqWcXzBgEmQy6uPsNVV/w6fo
wmKXj0oMas4Fi3WOxOqUgJBudGalzn3nM7ImN340EX30unQEF03BvTVlltKOWOHN5VBUafoajRvj
ZT9O74K9r+MXe1ojtJnKe8hAWdVi22sfyCf2NuuM6SZc842dfABd+MWQEix+TaYzHwmhHlfiaAPS
pIyN15MG/+DpLlhtb93QZAnxRQrq09GdTl72QtRdG08VNEbormliIipxfKutqA/DXFe8Z6AUT+VW
ycELpio7c5x2l/syiDVAsvPLJGhQpna9z3Ww49irR7uEzCihpR6TVvS1ZNrvKQOwlfqSpQHYda9A
tkzvRiPW90QD2PY3FKOIbiYsH7MX8MC6qzt3mp9dVVWD33lxbskFNJnRQf1iW5/7md4gJEKYisDG
q4ZbHqDxljWTuLruAMLAICcJaRlAk+isXIEweXd7TxzR3QUPtmcP6DvxlSoIFH7BJIvJERdgf+MR
aBeKOhQqvh58Hntlll48FQOYbS6sdVTTnm5jGXHWtVSK2y2hfN3dAFF4B9YqZc9nk295jQjpejeB
s00QQLDscgev3nbWz/5P7r8xptrEx4hejuCDhxsQEHPluiXUz4Zabr+mMy0zt4iI6B8zeTv551qU
PlilNfn5q7OvPXN5iJknzeP+H52fKRB5mOdEgfjjTmG8lTs3qmhHtHtLAis7yD00Rwpptvur6roF
ad7PeeSpZUgz21JnK0LOxqYEzUsZYVA3ko/xgkUqh098j4etvWm8wvJpGJ5FwKjfAtRNI/lbaQcg
9ydDVfTJoo1Hn+Da1QKDVCOb5OpL5wMgPR3OHfi/amoe/4gk8/yvrwSMlZwJJljMnrWpi+mV4Myp
SQfg2UQdWK4jSZ00XvQwfmHiddQ0kQ5OH0ccwxfMUHcgvvw+nfxczCiHswjecdfkXpYWFn1I18GB
NgtCwzaJ28n3goW/0g+pw/lKidIG9uPMSb4mTB15Z3tRRDea5854xwygCP8TkHUmJHcrovflK/bR
U+6ADgDeKbPir3bwKvMLD7z0MboIW6qoOOXUZBeOb6Bl1LwVOIi80ZMaeq886qZ1cNS/tQwRSVDk
59+3JnsuCpjF74pIhaXPTDhlS2XJlP39ZqEhw8uoBKuZvYggNinnERzYoWZxDL8/wSUMMmgzEXox
RyjukeNquINSYXWhL6YU2/kDiXzngCwRSwFy0egt9yiOs3lCeWsMldBBhuoSRe2nKMgwMTqGhSqw
fiPjjBSHpviASQZqY4WhlgiO+unSeKlapm1biyVAzfbmGImw6JM8/OU6G0RPPsZxXNBHsX0ltJBC
UYTTQtjE8DMOBQBzXLPMhcAxK3zO/bb9vdoSODbdPmW+OnU3WrOC3IU7gvUi0W45uRSfFERB8pS6
eVysboHNfp+NGHFT0oRAXfbHTjSY37hYQkgLdn791xk5WlQrs353+ceQ6y72B+JAOw9eB8L5qpDv
Rr90tuclrYMoovsgQW+8O/lIKwttaI3YZfwBT+OzseJdwvEHxsze+yKv5yuV3CgY+gVhR5I8ezjt
cMBmQ7g8GXLSCuQMtCHInMccBwDKPp2iumC89mJlf5HiFhibcusGuXaPx/0xUi44Vpi+pgAaFOeW
u4Fjk8S7BNP/xWlQmyrhEPL4G4gRH1F5tJCPQkWT1IcwsJ6jY7Er1V3mWHuuVNuSqpvzvTqf7rbG
FtuPIp29ylxU0/pv0izXhKWVbxhYS9ul0X8ZSEQTzJ2zoO8++8I3zMLs3bgLr9ouMlwlCOvUmwWL
TZqvq4lZUuFX7SW6ZjVkBeZgm5a2ZADDqXPYgztJktba4al1qT4ppK/4eqlEZ7lyBuvt6I1nqLZT
u0q9/ZC9ZTdV8PRaHW2b3l4DSkx6YYkXM0XGLCpdXyE8ap/UwOL/Zdo1728wgQWsQkIUI7zvud3B
SVD+PM5EqXGOpl4NAxfj1jOA1YnS2RbG+bSMA66iSMsd9RTZkhvzqbSrjeZz4gU/5Jx4K5MXP0Rj
m70J6lqtT6lQBtTPDEAFouhTnUB2AOcDhR2gvUllnORcS4alyzLR2ncr7inhog8XRBW2LULX5Ua9
zP3KmlTvsFREgeREqo0sJOlvjgSleN0kRK/BXFfCv2Or37aJjAd5s6JnW+i2Yu03m5BfE5P7mYCN
2dG4VqYNW39Z4tRym6qtGbyZbGGWeJCtDrN+PcflDc8LUTt2kHwEiY6bfq4o+zuUm0Hcfsg3D4Kr
SdWv3eGpziTKF/U74Sj4aLf55Tu7AIJXHmANQm9MGNFtYhexE2EZ6q2v8DQQHIceTaZgeA6QZrWl
uPVN8GPvUjw/EVNR0Mje+fzoctTxV5P0Fc5G1/EARx0rKRXFXhS6NyiZmu+JeGi1zsEvFKxg0OoR
eKePvAiZLqabIDeFpRu58VzfZfrxEX9PaPpL/JjLIqEPqwUSBLF+r3kDW4Yw7JMB8Ktzf1Zr8xy2
bvGVoiYpTehDQ4yRhbvZNzE5aGhS7fpFOQtPX1oHSPpUEPVKYIw9x732Vur5moKfkUo9J+irzuCI
mUR1ZNHCx0nTfARybOW6ibzvhI/sRq2lnyFPGGJmFatr/OCau/Be0h4aBu0gONYptnnvDPQ20UlV
EkGPWpzxhSaw/C/9bT0Sye2wTHqzTdGV9UuAPBal/Uhe6Ii9klC1iLD2bi34Wx2ETto+k1pSuDYh
NJ6SEpREjnIERJ+laTAAcpel2xEz5cydc/kFu9MfeZQvDhVmu2lHerFwAv/D/3GgYGtaRkCrJ6F8
RXYpA7MWnyt5b8lL8w8Tz+gCvUvUiqXUM7ewKGF3YcHRF9YzPNL/tSbL+RYIEKVxriSJ/ZRiGdw1
zTxrvXDj36j+pjokTTDqJFqZeg0/OB2jMynLzf+PQYF96yi8IhbNhseDBq0+J3pdbSWsW29xCGuE
l1+cC1sIeOFVxXohRE+otI91fWtaLTvbpUwyHWhxmF09DNn+KyNOe1TsSLyxgmKe/11JnNw4DXyN
s1PaUMDwfU7DfmBm2G68nXDuvaLCjHrc3ayjcfPAeqsDD93fcEvyGXDSHrtzWBIwJu1/7Df8u4jw
6jgqbYaoqeObP4pPWFoJFINJlvMYgIghXmhB9tsindJwku0lWOoJQuwJgfsW9iqrchCnXcoU7e4x
0WZH2dyR9dTc25LR1vzxdQ8FaygErXxM2FXZXNYxkD4P2G5TYosPNfxwBS1W5P09IOywsvWUCfY0
0ABI1JvaArszk5GEYFqzZ4yR233c3TXx8py8kicumHcZC7LtR4Fz8XPMdpkRWGDfz0JAV+iZxSiZ
VrNx3vJiyZAfpRHXY8xJotbnLBIvxmWq3FFDwMAkeC0FONZnhDyeBXpI7w+69K0Xn7WF3TV4S131
gm4duTqKV1RjRkGtUw/y+FV60fSEMpipP+YDjVzf5hWl8gH/Uf7kXDFKd7h1KnliA5HwXHS3IqoC
vtmqBmk6ZwvmBrvOjfmy1tPmIzz1Ur8jn/AVMdZLMJTSUc9UXOowP/xUN9MFBbrKHnkElPF3gfJd
0DiChNNtBEqETy9YegN02a8oSry8FdFZ8FFvFvmcDkJGA1ViBbu6Q443uOElF6t0T75ob8JZLZho
aBCN6aNBJ2nXERVy7q5iJY1pAt//eslSn5GMco6WEa8AWVD/jBEbCrc9FizCSAejfKlfk34z+v0h
O+ZVsJb3fnfOCgPdrIGJ2Zs0QRBIBSWvbaEZ5N3jIOSfdZM2rClIIlhJjltTVWBJ8tEn2i75Qr28
Fpwynj+KAWjKP/1e8F6n1ERaoYPsK/oWgcEhKAVkCD6e9aIkr4mUmDAUCo3vd+s5dywtX3gTqtYN
8/jVYLG/Zkqre2dNoYrDOA+Pn1tfr8rUcEtBOUXq+mwJCmzo37SpXq03Mpls/nVpuPctmikwHNGr
vWuTqF+stFnKbl1Wy6jjKRXo+8ZophP+9bHcgV9WjcAsCsexe6Q32PXqoVbjKQgYopsY67JzCyrS
dV0WFQC7DHAw1VqeNxFrhTl0UkcGRG0HFO/FjEnG4ZnzOSlymEYNFYIXMXLituDDdG+V7/dPq+RZ
Yln/cAqivhhVsywtstSlmlrA1ML2lH3pBqO6woCyZ7I/gpgOxQCW9ZrS5qyBGxVJUt4CM+srk4VG
I9R2Ho44UANB/gTYL+aKsZZHRTBPr13URGn8ILvm1cYlaQtQ5MajxsCv1lqzYUAwt89UYZXWtJf5
xn3lTqwWV8Phpo5Y59ZFtoOklESBNXU4ylc50JbhHdPe7WdTBl0Za3kmseJLjr7X+4ZTwyeYXhf5
LhcFcAhRZZUzMrbeMsys1QHi1DHeiT7IEHTiC0BJS7lJNNHz6dLLj7KTVewBxgCTvxFOZOS2OzH0
e2GfyoS5f/gMxaqqM1Uhp1DqynnILVldVoGj6zezTvld4sPSPDauhVLauWjDEBGfntfaLQ/jnUoI
R2OJYprAJYChVBeuZA3uowP2Acl/jGrFRtRSgx91fPs/RZGr7zjPHBbknSsReoKNxj7XE2iNVlnD
BUsOs55nfxP71X3Tc38+6GKe8j06CPJaZTBD2ShiTWum23sQ5X3Ftfm+o4R2tum75LQuF6qaf2YP
ozWXYFy2Ymzj4SQ7sCMVO4E8FZ+i8nnvIYbLD2WzlMQt6b0CtsSwnfWoa2VrzfQXtNU8aLt76byN
bER0Y2PCUXaob2lLa+RDDqpH7XjQ+a+AxVWtPDCQw/fdTMmgK/2wK3Qv4Jv8JjpLPyH4CuzRjb3/
wBeouGYS7V1fjGlbCaXCkoJ3sy2mpTkRYLySdSrrS1NPh5b/6bF0f/6ceTlfB2W5HzLQ9K1252N7
D2sXZAL7oGBKEYYiXxa6hE/IVGBrTulP4lj5QrC0F7kpGxkKC1V5AOsDPyj79LK6c1tf3b3m3Pfq
sR2SfTopEwoG2rr6dnblz5vgFYeISsAFEdFmXcdw2Rir5eG4FbHxp5U6d2gH7SD479kcIvV0ttI8
acAhlDEFnAtDbNr8K+w1R8Aw/BJblulrKLYHGOI1cAruNHvOVHQHHSouAK6TTTvN8NbMR0SviZia
IOsGklhL/iBTsAoso6qePrKGcrdhscr+rGK983kzHmf3cLJdj9PwYr/KwaYFJwXf5ZF2BH/6pxr5
88Sm3Vzy+/Z+Y4FtyhL06YrJRKO0uZHzS3UxEQhFl4OhQ5zkn1/oXAr8lz1GUWRIbj0zRBkrP/SD
I8i8//ZrcmGvtRJcJIZilMY1EqwWYkGy2kXgS0H/kwPMX0SdkVHhsSjvBdfWs1Tju01nQxaL1Dp+
nE6dURmA/WKIGpoz7cFWnuANXPs3BoPj9xpPuoxPXOY9pB4LN9wd42uDMgGU068/yNFz2dhzJIE9
PMGIB/RR58zi1uTtn8NHDyemYwTcXgGEnexCmn5FYw5NXBrqrINB39en8S1MEe0YbmhcysEPssu8
Yubi5ACD0YzyY+ROmFMnb+mPgnNub1WNss+NOL/8JiCm6KJ8qrCIjEkV8XoK1ZOcYDUXvegp9Yj4
UzYqeCRvRajXvB5tLplLN3YK5Erot+G0+1A8CjAfGmbJT1SyJVdHiFaCC5xNupz900lXCDAIYn9y
YF3LixBbHQ+UqcFHM68P/ZHJ0jHqmy7vpKOkiCNCSMW9Wb3Q6TkdGN5oKXs00KvQSYKoZIQ3iajS
Blhh7mm+aL1UZPtdP62VBJdmKFKHHZxYwSNFFTDC+GPgDfTKVJ2l6au3czcUcA1XdDqQqtPaWFru
dleZFcFPH+zNZzGG6uYdMQLRgi+448aJ1hhRARjeBs4EnhRZQ2++A+Ie3hRIvYl0+B7kO74Rz5At
YDD5me3lmQt69P3nEAVFDC7Rl33q89/spmv+pc9TX24vPvyHa5B14gJ+k5En8dg+fjIHtSAmfHx1
sat/ZULjwh3zH+13kHtVBOzBpPyXF0/kjMIPXzMGBQLkGbzr/lahpKHNRTx1cG2ESO4vlSSUmzz4
sOJEdH+hsh2Tzyl5EUa2T988h+tbVb+Hefjd0QaGFZ7gkuAbc1HVS9isV/Ypgxn7Qb6/3obzTuvh
jn/8aJZFkEtf+Ugme3KWQM8n4OwQnp9M/vMKN4f0dc/Qg2qN4ELRD1S7/6rA33KUiPbgNHeWXNl+
HqVDPwN3zkIFNQ5rY8wggbOVG8aqoget6FQBN8b74RVPIl2Ry+Oyy+7suOv+ZaPFVDfCaF5YuADl
bSBuaJCqWCoeSsM+EoqIOhWxZIkNXpJcUnUqk+JTxFnLVYqiguT53q7CPP+ka8D9zsrE50VLSiK2
q3gqkle0qAfrgBFfzVbLvlc2rFnrCdGc3vdTNnJiM2Yj1M/OxoJJ/sEnMf0cLlUOKTevf5OGVO3D
F2n2BIP2zIZa91m4sqFwfHzjr8ReIcf5FPxk3j9hALiK+KacPP0tqJ5XhI0PSNRDLEIrhHN/zJvf
FB7A0qfk02XQvwG9XVOTxU2qupdEGcF9aXrhKFDaohm0xYIVZjN6L+FtQ5MkGFNzahdHIervcRQU
ptpv72kUJPcI6CiapbY7s/eUe7QWH/dDpxwx+ys53CkzR1BIc7ru5ANQeQV4/jjPg1KIWQfBJ8CW
NMaQRxMYnJMqX/3/Vrt47W1mw2keJ/ZuCHs0mvqnR3P64aXxOcH9vTjRKQVbWVgz6FxipecalIVN
KZ6+cQohk/a8W3BD9+Dcg0eC25Ub6KdVYnr3Qj9q7q4NIxxUEE0mqUdKW1n3btgTIY4yGcAdurCE
jYwzoRmFrwObHvZpmD6sI9z8NW60FKARZb6xINUyJ9UcagYYSwGSOdfdcGYeF3PuUfQF7MViNRmZ
EkA4aou1yg46D4d8XwO2pLusXpMrhepYRuvWRvSVbePTV4nTqhzBt2YR/VjlQ+JJrS4Ct5WIons+
kUPsiTlx5kt9zspItVFtbnrrP9SYtyPgwXPMl96u3yY9hO7Bo5/uo2KzUq9Ewr7xI2EQpvjrDW35
q7F4WSa2e5HaQmGbD6SBMWKGnu1WUhESpz0toDUcs26nBOWFx1iK97DyXah9bchOBi9taPUjNXyw
WClitHNLxTEg2EeBb9z2Z3NvEXASYAa8/reI1Ant1sNhb6NaGzV2jhKOH8+k050zE9C5fsLBGSUX
qXTkDo7qRbUlu6F+Wr0p9iohWWbvclme0aMIX6JjWGpXb9+qSibAC9jn2kREARmLLnYk8dZnldJu
ENcyRndCZUiTDdzZ4Fcznp7K9UykhDhHumSCshkTm3mpkveVMLtLsThiYdQir89HKHVCyTzHdAZ3
a5+UhElPst+L+N1HZruqdq1L9kN2a2SdYJU3qgmEX3TpH9NYWvNBwFyE0c80WP5raZ7xyxzMjQRQ
hXPd7DdO9BaGUGUVG0pskEOcpwjXHVcNeS2a+Pg3wUYrXz7wbLFNPuBaXaqlAG9Q1XdTPKDJQpJU
z5E91+SMNPCTIfl5cV9IqxET20EIJtMzhV8jeaVJuySynvoa6b4pxr6Guu0gmxg/ogWuNG02znxx
Di/hnO+T0pkwBCUp6mYSZAJWR2adfAAQ/mA4mAUxQnr0w+WLVyXKmtR8Kt4L2G5XuJ7kciJb2wwU
xijx2T8dp9UO7oR8CkCjspryRI8RxejzWpW/8lldEtgKgbeIULGix883NTpEGalQwiwUYcJDTb/p
NWwoKaMS3l0bl+u5Z5BvuMuOMdHQsLtmaFNOQSb3T37SSAB2J/IW/LzADeT0VeerACgxH9vouXRU
ncA77KqzRw4UdSxpE/ah71KRnPuuP8UPv4ZiYkiuYlwsxmpBxSn3+YEv+X6jNa3myY5KOkIcSSqm
qwPODONDTO9MHblrNaao2RF1EPtNIRKnix4xhOc363n5oBlPrEl0VzLEEn1AC+IYJrmSXVRFxPbr
9gRifriX9nHYHSt18OD0TSr+HCjKuMgLjcwNoF+yHmSoEYyeY/2BATJZb3FtfKBjd8ISwRNz3vhA
tuj6+h3iHf7Hkby8lstaIuTQj54wlicbrxp62+nmfmAqF0FS/pbyk21l90HyBLa8JyGav/6pXy5I
sMjknIjcnSP5lxyMEB1aBkb7cR0LlmCQSRns7GRjV4lsqHBHcPs1bvxtjgcSHrETAbKoyv+9wYU5
IWfqZV05UjZsz8u9b3ArSgbyRaF1/7CLu+/D62z8lWUoInvEgbufTDp0OFkOJPDWvxgccukkscf3
SNg/Yaqji3M+7FoXSXu5QGA4KSJxNGJAnIMH1DS+Kd27Dyyzf8oxhJM965wf7bkkSMwl1jP+8L8i
iZVJQybteohOwa0iZfwEgLcOtLRXHlTRx2lZtZqBc3VGxtt0kdSSsCipuwHO810MEHr7WuSDB2dD
uUrRAJ1lMwsTKRRQ5a4Ibun+oOF0iNdA1o47Ny8ZaQ467+iLFoiXuZWz+dp5GfMIgN3iSWDSshxS
4A4A+A56pi/hotGxbacX7JaUHwyoX212sK6u9zVB8wJQ2zAHhk4h/AcrIS01DE1DSU409I40XEEY
8YjYZ7gRs7BmURPcOjO+UaElVd8xxuqCHD93usG60thS/iQwrY5BLM1W4sjsbCSSjeUWbVViQ4BV
yagn24UIfOAEfgaSfNDY7mIVYziH1k43ympowUgvIEkxSomO0dYt020oQ4suz2ltC3FquNmWvuP/
/amSOOQSKNJ0cwtjX792+VWzzSjZNXB3c1XBEIGJmAiSWtenm/cJfLKGoGy8+xqeFU3QY2Ko2haq
xzn1NdMPW+WIhxgSPyrK6VYH9RyWJFT8EHnoIQqEJbp+fp0ewYIZMvDzF2tUnnqc1QzTT5Ta8ysT
Led6d9RafrWL5JdZHwCLcGtruUXvfk0BX/vm3vx6Om8W/7pe7P+MHwU43uYgrq5vS6l0J09ueOFv
iqByt0FKRVgbX0MoVPGrB37cl8NnzNpzMu/nSOuUDCuTf6iSocs0s6zzVLwSc5fQ/KSHticjbBNh
DynpytTwogczZNw7ZS2tVidZRhIU1c5eSYLh4sCzcDakEjU7X+DMssqhwERxBzUkS559R37fwkWS
bvtYqd4eT2SFDD9NAvgsjw9J0C9xTQLxst3+MZ8/tCQY6qk2VrKTR/OXTAlENiGcCjabpXo2kRa6
XZi5p7DwpCmQ0nZILB5EtuJIsKOxrfAMyrVakY71eS4T+vJHmm2MtGhZidSNQE9fUEqFhBr1UhvK
Y2dSr3+viw1Pnrdzdtm3atdtNEjZUwFrFEDdBp23AIvfWrk/a5sStjY/rhD5JA3hXj3/8KX7MQNZ
t6uyZsZlQpI9CIA0XP8BzbQIHdcx2KOiSDd/ia6DfiFS7wAd75f0iG7sYObmT1G41PUaFzDRoD4e
5iuSqAsGdpOsvvh6iH09hOBy8cx2HB23XksvyrNpWNf3SZvnMrSgClz4fEx5RMGPxbJyzPqkqcpW
+LQsztvxtiH0Pm3+o7vNvpPiTFHJm3+IHmANFBRVhP285Py5XebUg5KlLJc9GZUqgx4RHiaEjAAi
lyNFsktbfZFU3ZSRu3/KuBDlIuNGLxl+uQkz2KCPWDSHjPYLEWvX0AP7X0CwiXslndiHxK9j+U3i
eg3ODxEP837sX2L79ubcSw3abGsObdlluNQPMCg29qMuQ8C1E1Di16vCStb6Vt26heMq1HFrZrLQ
R/Ij4aiVPZUB4B04f+0D/cHcINA7BcKmi9+xrUUJTrdiSpwwyH7NpaDaquzjYmGSX5H1EQQAmPRb
YOvy0UNZm+drXsGIN6LPEYnvVPAaWNNxGTGuTwSZ2J9uCsTSWo69QNHPbzsHgvNzr6cYfeyzl1lZ
hiyGckhWPsiAZod+619p1gl1W2b9AXdK9vx1G3VWf3ztKeGqbV6Ix4Z5dW8mBurD0asxpKzELkE/
TEsaRCRdMIaAigw3qey9lkemUVKuBbQclCJccmWQ1gZheWnH/rE+g4wgUEUeDp459pBlPKVW839k
ntAPCB3Gn7nXvIL+dcg6MPvwzcIe43o76iuIBT90xCxpUDh5i3VJCI9ceaBToOUcaVL2I707XRbM
ZMaMRv2Lm+Ct4hMuy/YhvPHpEG8lcHatjXEblVYtnWk5wNVJTPNXNNvD6DDTwVPtiym46qdICrS/
DELoJ/NZNcOuIsF8meG9ZnIZvEGTG9HMaxt9Rqirq6jC9OBmFnF+j2BnHPYRvCWPucekQSQZ//v7
4y6zMbPdSDOk9WjH3xrM4Ix+xdlgvk2hrFs0yx4t8mKD/Qctwnfa1rXGFxjmb6/sFOvSssn9hftr
SM7DqW6pmgJATsyo4c032uokpEdzIVud6+BMBhogKzM9oUuSr5oyZpTblc53UG8wWj+fCN6K6YG3
ZzGfyUYEhbXBl1hr00N4ckKRL79DLsCaYBWQSsNNK6zhAEdzXVnv+4VklmGAIVdDMvqFzz9Z0A7y
ujSx9/XuV02i5ljI9WK4aFX9q2sy73M+0faIY9R5DnI6IKYfmtGjOOssQ0USlBvdTGPDFyTF0U8z
bbH6WGrZ+e2tntE+1h0GwKLwPc6cu/2eUCHXwiDD/rR+W9MSYR6wqQQPr18HzeqODpavnlq1+bwe
wTGv2B0/iVVx9hsH2T0dggzXIVVP3zQyvuVXaEaMCd8fYhAc9IPcMW9RMKyRv5M1uX69GHXhqtWI
F2jLvOIxIMT1qFM9fStlgwm/2xO974z6ME4chraASAREplMBr+8hFCsswuBv0lk5zikGX3CGarRA
dZ6Hhh7QbavBCprUvodLG2Sq9mbLsDf2SGTmSpR3t03xnYz7rVp/v5bRa3N6wnYdNe9dVDpSzXzF
hMswJm7n0q0Uf7zkcvxdyhlaZnfWCYxPQxc4DjGJM/f6DVi6qr6ttTcdrbg8e2JIonaZHIwKmvpO
6PJ3utnhJSm+2odaFufRljRpS5yXos3Hp2JCGW41AZIymmb5qq2ITFmy1CDGcEs+9uKqSA5LqeCt
9zq3Oep1lN5zXyaDhDCdW+BIGnxYD7PVMxmVC70qUFq6Fcxmr3wl1Sf9OIe+Vs3Kl5tDo57c/47/
vybED4CAtr889PtttAYa9VDmcxlnD8Qxqhq4SwSOvCq4dl3aJ8AGxruHbauxccwl0pQstepvVYt8
e0lPaDy+0FTSWLjJSgXuF0oijLkzaBsEmRtAFD+nB1aBSuWMQQzj9148wciAVZzu3HtAZFWhT7CW
Itc/Ij6bmwoZ4mKp0w2TAMa4PbPNtew+R701RcgkcKHjeuokiIhk3+Aa/92hOn6cUpXfqbDZX4l0
f3kWb7b1apdpqKgmLwMmr9N6gw9bgxH3owe/mE/ky5jKTe6J+S5Zpla7NNB8CJf3ry59zq9XN9+1
cMkl0+V4NFkZc6NP/8AZ+nrj089wN03qA0hwMSuBNGkVCUmXUs+Sksm1fv9rwaJ9v2Ll24DpwGlo
Yb6ewyNp/5GEnm/TFJwmjJgg8S50Z9YuRHDQ/0XVGuSebCy9Naz4IM0zxAB39Z9rDpWlYG8u0HIa
LpEEVh9FT0uJJz5wFr7NuLtQ3iJsXpJ5t6d7rZrEyFYUELiUbHaHaZv93NerSwckVdi/+Gm7Wg8b
U7HYt/9u9O3yLI7uRNBvZVAQUhgdU+I/+F8i78ahiiS6C41rvicaeJsBeHmqMbKKUv/9EOdBH0qp
GDvSt7dO/uxlLh+3Mv/JAFLddAgaEuvrJsbhNZA1IdntxXCklh1RGJ9q8yCeJRmXZsvzyabfAZqv
9YlthskvwDKGpx3sM76TWOwbxigq9GdhXizv3KrMLx68Leda5QobRPh6g4B4kZl3RJj/X536mklg
Yu+9z7Tqrx8f9WU2hnfWq/CXML9uqlY/UZj+ZKV1wcmxgcgTYF3aAbkO5Ib2yYxvNKRn35fF00p/
T/oDUJrBGBzBvyaPjNkZ6BLcmRR4OSMrj/iGALtxj186WKHwHDyFunrAAvarP7ucmw5zyPy4xMSI
ID5e9yBtnsiuzmSgRc7KfOIajmWjuoiUMMiNn0qpuiyNq0BRHSUkCZRZvJKXXlc4k0LKUvcqO4zi
H28LZPQNH7ezPEbEgUYb4CEIbJUorsTbtUBvOlIlqH91GR4Ko0cpl+Xr1FD34OhTmHB26LBsxi3Z
Tdb42jww868mh7oezHPhIjVjBQaEl4+DWNnHssYKb9yxpZHLlDOebCoL1w/fsNinTi2SRiLOCe+N
d7J+QlXRySajmVnuLzx8kT77l0sbS9QYj4o+p28D8sfAqhffMwr0JKGaLDvivkMNUgwip7JPlwpM
zxRVSTWn7FO4yglTx1EOauPn3Tq+RyEm93F3S2QFsHMpJTc2CcKAAk4sIIZfsPiIzMEyONCprTbF
H0/JcM40lrmgLkPe5s5Zk4WXfSD6VGlLSfQZZcYRKCzZkDbQ5CDjJP1/w91ZHzkUYTmIxNBMmd4v
b0JxsL/fJn2+kBC+PnX9bsN5ht918jdLckGCnv2dcd/yMGllvEemYnA7XPrgv11NCMeugvAAWPrG
jBLc7h7v21vy7rovHlliQH03gopCwHgG95hnpn6V1WUq1t8TW4NEHjqiPLUyBogQpZdpmR71X863
chTkVFuLAb7rZ6CAZzgpweq7mElmHDiZ7qL3NhcOo2o56jNIR1AUc+4hH264XrVteVCY/jv3CT0L
KXqOJvlFRtYslhOtcP3RUxKz/dUT+WvpHeRrY5qKDXDZWyGVJZUuzmDek/naAzGGO01zCnX4JGWZ
PgWraKnyystwIEtyGV3ZYhgEpD2Sm9UzvPZza1yxINZjF0XE6WqMX482lr9cGEiKYHwoVZp5hvd+
hT0PvXrHgZG/D/R9/2Ge/QTZDTulziEKaF0/jZUKE+ZxxWV/9877zny/aZexxev44OkIcrg2YfIA
jRXJjnPRxQaIcMXPJ3slRLzBxzc4rl419M7ozL3vrWDj5o/57E93yjry8BTXRcfA/6RFNe3pWxL5
BBkYmBPuWby00CxHlzWTs1zug2z62WV8/BR3fmgzFORsoGo+sRCXZHUWRXvZD33Unuv2Lf/M/MrT
YxaZ/CSvTYLDDMvRf8lZKOaSCp2+XZz71EaJWBNMIrx7dN0o6qk9MjN5fRhqpSJcihRjptwvYozF
3OoRUv47/ZLc8l9HDzvsMEUiEgBsMuGulzZdCy27cTtVfTzZ+l2vE3635CtV8w9c/dGttpkxt3wB
24tFp63EQmZUiJBEzAuiODaZuDD+X8rKN5P+2R2v3b8qThl8nwSiCRF7vNGnjsJM7LFauLgWeU5x
zqkZnkxmcmdcP29ZSUEuisndQ99FWYSNulkvzj1Fp9wDEVfucRTfg7L3m3/+EAPKE1113+fCDiZN
32NwpOsADnlhi9Jjr6c3CLDB1Y28YSSr52+YPnv9epGAdtBhSEjURp1w1wY0AWva6W2VuSqq9Cyl
Fy3aWKroGLFrljnUJ5IkrE27WwclHfF+9tKicPYwSVWvzj4gp6IYUZVGGDuGzLaO7ccfa4MMxwnL
7QNEQlhWqpOnbPU+ITmgKXFA7K9VhCi9PyKOn1M+k6ETmmNSDIA2CTZsqJSVV0jCZe3vU0vmTr56
xqIrrkUsCEO2pmdJcy15Msj0//GjtKeVFvpi07OBNB6OhaE4UWzhopGrwMsEgKMoFlIzKUTpir8y
Xif4XjBd0NQw4hiVRITjjOKoNnwySJYWEuoQTUYERxwP0jXfDNTB4geMIxpP0OqkaXrpWJZHNh4n
VPy4/aBtpJOcONZDLBAc/UQNBClAsvNqZJYuBN3k6jgQ5e/mNTCWwFQwA+NO6pHaO3EZaS9aR345
F+8tcJdson1NOGS/NCTMrOQajIyovSrC2tj7NjaO6JA85nJXMioHt22YkBMtacvD0m+j4jfKfuvN
X8A+levJ+WNBZVTiqjJ/5CaMGKDz83UtirXo2mDeahO73j/B6SPTikS4QbG4T//4EtNigZxL2n12
2sTvHqz8CEFMa97p3pMyZBuClCJP778GmkkGmbsKZ0T567TtfevZnre8aKLepC8wRgjdi5vf8WHl
fSdPfv3qLDgUc6voWzpdYkemnJmbODQiZtdw2iTWoRGNd1gJ6QPX80ntmyNERRsPmvP5ETzUjlUt
Uv6caY2tSoSrv0Qr3MN3fBYe8Ya7T6xanILisb7TYqQvWQHzD3FxbhG7JI/ox5nzRMTGU7ra2gKp
RTQoq0uPGeVg412KSr4JqS4LkIqYQx4lc4Uy8UUUtbSJeWoX56FPL16ycPjRJjp/OFslYj123c1o
i2MCQFvsOfvQgqP2SQ8lq/Ktou8YFZe81cR+YrY9oO4j9bp3hgO1Hm6sbAb/VfmOOrGFVRfvHD0p
ER/OlAZr//wGLo8JB9V+oJAam4Mn/FZqwYQHrMCEsYyat9sF/OfI+y7U75F5kAYSJJQZ4/QAiUFz
Ch58/zYzzBOwkStz/rADcOPjy/DvBTkDoFyb+W942kBgMzBM+nfJathMw83cek1QBuXsSRfvU/Wm
3SCZNyM4hT2o6/uBi+kqswoOPLiOekkYQM4FNWuIx/joY75vBTzSDuNRP0J6xZRFBsfTvTorB4HJ
HmmVx3lCfdAHpTQS++XLhHsPiehkrZaMC7vxnKAYKQ1nYxNdbIb+v8FMAwltMMtDvmnJO9guF6Zi
Bcy0K0MLOVd4BZfBnEIC2QUAJivp9S6JZVtd4BN4pDhM7ld53Gp66bJFVVRBzfBzswwq5DrpfN/P
gxFV0Qj2BE4ILo0nU3NtNBTotq771JYzrjPYV7pqwH2AYNerBSoR7wlfEQZW2PF6SaIR4WlPABac
vqXhyIkes1gpEGYDosS8Abyv8MnA0EYdY6yM7QywxwB1BDrOquq6GUEnnsD+qViCd5Ekb+utO1J7
D/pZZ/zKfNMdB9AehSR7UkIPizji/SVePqivy9IAoUcuT1xV6J9qxCX+espttQYRD2FusWvGMjAP
fk76H0qCLcvjBSQZBooYRNhoTL/UDgaUh6IEAxRg5TBcjvYwbAR4m11Qt5dZMGYhKXVHUDgcFy4M
CS4CWiMLcGQsvM35vVILDWAlwXxJk1rS2KygK5AVm1rjgoGnk2G8Rh379xdT00hnRGIvszEspBKe
Y/gA9XPh/YOZutCb12Ezsow/Y4c9uIz0YcyjxLIvI7AR7GpaWIYQIG3jbs5mC+I3zeA7esJzp1qh
kn/PBs3x65BuHc9heSLkM6A4C4HFS+5GFWmPKXLf9hk3rHzn1gl9mosC6yFX/QiGq3jigrrXuS5g
IzqUB+BdV3ngbY9f14QKC7W+F9Yge0AzEX6aVu1EwAHwz4L0wjnmOhUzZQO0yCtobhRRQSFdXp2W
6VVyHQumzxggA9SdpvAmYL2eRZzu1/IX7PsbSQlB8Qg9cZkmjWHLW+pjJvnrPVKYkOaUQ72uLyWT
LyQFKDzcOr2zzuExidOnHtsYM1WqocbPhdzdp8EAHXa0G7b5Sh9VcnYgtpPQoBr9Io4lN8Qezvcz
eiyakCRiXlrxpQGjO7mNt7ZYiXuILvMw7ZJF72R3TBIpXis4UY64Sv5un8ktHlMZ5r4d3qpGRaAV
3CLFoU/CO9mZVvdkpNnyd805wizR5BVhr67cknlFvceXFJkHifgZi60CG9VShik43js2COeKUqgY
bDRjCeTi8Te0fSvd5XNPXM1OYWy+eosz0WWzYY0WrFeXx0YYVCJXWY7o+PqWrbHmONy4iCe/sVS5
/42DOv0g1V/PqWkRTHIVCH3Wf42J0CRFq/yVIooIwQLb9iKX9apdpYOegbYpexfHg3ykpYi8072e
RKbOEjhnL4LoL6VOfcZZzkI//M/JGEmDQ2/6EUKNiRAgOPRE/Ypwa1OY9S4bOp78iJgdqQePtdwb
cro9Nl3OH7qDAn0k9cfwUeWhLzh81dX6w+Yv1a5PaRQGQjV5GmhZ23MNG+eS2BezRDUw6IKp/Sh3
ysO7TeQSUoQcRib/hcuNr24Dl9gDYVL11ltoad0BzbaK/sYhsiGgeYSoxU8paX5QBD63GIAmZPLy
7Z0Ihqa+eVRusmlqclIqWdwG5efGWotFlv8sJWnFeVjTQzhtLXgv48iZeQC39M1zGLIADntlB/I3
0+LWW8of7D221argTytnrSr8LcCjw/1YSvpwp3DzoIk6YfdMbDK7dQRncl3gznwmhCrHFJqxaZR7
ByEAD+Eqqu7Xw2n9lSBkoFjPK0dSQ0xR7RYtsF7PDkErQWouvy5CdEPi5/Aydcn7o1zMmtRc3BrI
DYjeTWi/NazlQX+d6vKxZNt3bVUqRcLnJnOmgSWEuykjWjT5gCaYt0hObY+JkbRoZJX1+B4MEnKJ
c1lAMu0MvAEhbW3EUsMGaZhd38z+vN5p047wAE+9CcrAmbCFIXd5kVh4cDnf/sKHuiJ8dwbE1a9j
7ke6WbVmGV78ojXFZ5IM7GU6cO40h2g7p93PzgVD60pO7ir7B3PlRdu7j2phIOwWjoblgmK21UIq
egokTXLBCd3xWwN9ySs8XqUb9EGXSObiHYM5gGHFkXi50w50W1LVTfYF3Ebe2ca8cGIIvb5/jQJD
dPSvDbUaRDJ+W5IrXHWn0aFPbLvWaMkrisyQyauqfkFVqJIy9h0NbVixnyIdIVVUf81yWZ5d6RVh
kteQdPflS40GXDJMiT1qv05s0ETt20BfBLNeP1kmURubzKpNbrhLyKemQc6u1FZ71qtK7O/+d7q3
RX/HDs6QgJbscW6neZ9MVSq3fivcz5csD9JVr8LJkXaWBxQeug5lxX1qsICf7I6maJR8pA5dilaF
224GQgN0SgiqIMU6qlc31Vy15DhR0fyGR+3rctICvoNg+WcK/5hpK4j8YvjrZYjFC4iIpwnFsyPb
+ZGa2g3fBYd3MMJPfZsQzbmjdpYOLJ3Ga8auF/AU7u1oRIzTBjGCRFWz/rhL+ttaJZnqUw/R7qYu
i8pUDBvUSExlexAjeSOGHcKqskraWzYvQJvp3ikVse6hWguGBgcVOBsO+YhMwRtag/oilx4KFmr4
ZtgpAM7Gso4IhRST7bDTnpkhutHYx2xoWypbQaMZuORsE+MeAnep/wcPhTLFgaQXJCxbZ6Ob1CS7
+3LnSzTwjKUracMOp+VGjva+QQVpt6X97RaJX6E7Kb8XqATozU0qGJQ6dOHnv4S0qX9aBtZpRj2f
ts5y7U7pNqnKbkd+qI5w4vteq/Nofp63rTw/w9iLnFenzHskr2daEDRKWnILn6GksCrgCkneZDKe
kbw1oX+0yF/ls0jlS+2WCxSXNoAD/iAV4KSwn7XP+a2abUQh/AknqABjr/Ur8suOOszxjwo4hPNH
aU7K2uXoKkvMAAVJZExk3d+RgCzwKjLUcfVMwAT+iml0T69xxl+/SMHZIE3XuCj9vsZe4IHyyvqG
BA5ukfGAolMIT0uMqwuNDFImcHdO/koZYJC1GvR+hq/VYkvRqIN1Ne3wsirUuUnhUpoXHuqAjIVT
7nBdeZ44Mo4kTes4mZ/glzMFVm0EFGtoZcPVgXcG7eAyFhjkGFpgy1b48ji0UIX3aQ6TzqtcxHmJ
9THXx5z6TpzOYfzVuPJC3t2NfLGhpw1j+HPKX1hah4dn/oodJLaZkQxOFSaJdzd0hPNHHuLmDEME
oecDjBELVBVombt3unMNXrbMnxTKgfIR6XK56tS/5oULtMPHna7TtjubiLGuwQCzg+LVtdjTlu6J
3ZnXKHf4RAzTfqjGdpEYs2zKZJ2Bb1OhBQFcVdjDRGVrh4MIjZeh/M+Kb9CZa1c0JTrj8awISAqf
xRxjIoFH91gjpjmwBstkwu06EtgkWkRPO+6Bynj+8FDkg5qdbDAY+YvEdi2VmBIJSIpp0PEcDTy8
C5OI2YwGuKy21hQx8za1pZa7AFCfyRAeNMmV0VFJazhHJhxCO5SSvBeZQw62EqlcwGYZimV2UvLT
groLuTgeimagFtcqNsHr8KRoHvUAfycJmHApTSZPZTu422uh13UcasP8ma29Plbjjr2DnVMU1mh9
n8TJVKFs8gO/8E1sOaVHjVahA7oKtiZ7hnINe97ezOVTAI0MFFUriWwaURq9ouke5blXqzEY5cSE
S4ADW7iwRXHySJpQTMBLtswJMp6Wl/cEa/tDQyHtrbscYsQPy1uJ3hvA6z+GouM+Z9Q0ZQ4mV3DF
o80g0CqLYJfRRecVYgZnk//29KKErCa+tQOZeChoxF9annEgySa8w/NRJRxJZk/S5VWpcKwJWBag
19ViPcMGrTngScbIPAaiu19T/9Se4d5oYPIbWOL4AiQ4HILN6OtIbpOaeb2sfVgcVXxNdeIgb5Xn
iBu1LKhXsnuAwme4WNJHDqHGYh6nx+xciVxaQuwVsQwMk0WKPM+ysvpWxEpyjjEwoB2qEndmVnO0
POes5rP2DnmtPLUhKHlSej1enp5yU492tPTdBbCg9UNqxNYEY4q/q+nGJpz8Zp3jH2InVmXZfwbV
csoytfs7FTD4ftFo3GzZxdNwZpHxaGDkvIOkT9+utGLbF0n6G6CUKLmwuAto6z1IyaxUwqMXAG2F
gXJ/d8UggXwkFydkyC04AjYwcbDkhS7Fvf+4Q2XcTeCwV3Xl3QsqVEedee8ckypcjopgu3qqrnAe
nxRXvF6QMi+ZsKXWNYqB3b8SCTdL0uWazLNnKWZbmuFnqW/hLLpfV6brK84zS4UnxS2m+u20OlPz
JBJWFw6ZHjZVaSfTupnPXpQeJfuQATsrSS/enzO3pJZje5Iy0/OJezkpv0QWJg0Q+QI2KVnQgAzR
VmwQo4uJNmEIrPofdExEDlpL5JcYg541zkubdIDcRzir0rWHbGbcFnchlUknsSqkaXdbdXV3EZ/U
MTlFwWbAJ37gB9Rn0AaUR1Y53xKYi0lsXMyTAoxmoLKmFmvpDRP24nKzFyZ1HCbryxP2nz7qsZcE
A6ABs4LxXRmwud4L2UbvAtlb8y9EW70LgD0kJpJmTV8R0tFt44Yk7I9HTNz9sQlO4LBF8NXfBIT/
7RmwqbMtD0O8WshlcYswsXN5npyP/2p1/6jolqFgIp3F/+gy9YUe5MNz5Q1uNhmYgIc8y+tZuDNz
a6CwsFHsphYExx5p9X9tQqVXTGaMSAbjLdvMx8VdTmJeIDiNUNTf/zC8a2/umFk8O/Xy9Yxd9qf2
WSpu0ZweOp+lmylIMT8n86Jbvu9GuyIScVIxdkJt7tzQP9+m6MoUHFS6ijnRnmobxQopw4tgT48z
1j5LoWx7HC5ILhJQBFiB9g2SYlowyfhNJD6xICL3woEgaDdCMIzO1jRkYDszuHqAai3p8ReaR1oL
wRAR3DC3BuUCFJTS6XGNhjdrrEL/VZpd3//0lu7SDG1vcMtCLP5aBCeFrDdsyo9JpIYr0Maldlp6
thTJS4WmWaUJuwu80roVRl570/AW3VRoI+hiQiJwv9yJ7eOxnMVaIVjs+scR0iybq0RdQwlFkXR+
888t0M1UEODWeQc7XGgqp7NStC1bFDcdHyYAlhdJw6UyDEpkbEqgpkyuLOobp5CCcI30A0uijg4B
LeHg6A15rPGm6EQEKjZ4UGg6DabiEHZamHEUgzNMVwRT6MHZWZQWb/RNPPeMbgLZylu4Uk6RwTc5
lgWNm405M3+vSszjexUFjRXZC0pX9H7fwdhzsGH6I4ra00OoxTwy7ADkfpuw6bG2Hwt16keV2lJE
eIwmFgC5t9cwj6n25Cg7sttW1BeEkA4Azm796BUbV7CjwKGQhVm7j222Cz95Fb1zVRfT+/RfY0OJ
rfDtrmRKOzoeMkk5vRyHbsvSMJIkcc2W+zCYuIwTobMFI3MgaYK3MpdvE+qtOWm5aqYR1/awlGSj
XkilhTOEAA+qzTOXUFbb70r7RG7tSN53VSM2a68f1HkoqsMah2z4h6ixYOTEuX4OWHqqhxB2MmFD
hzn210DElQmiHkDL/u3cd6FXBlLAqq9KNS+ecCvvkQq9dCoqf0FW/yyg9+3BNho+cup2AixHtaN5
qVgJQ5cgklTkfADneX4TX9VVGuAPE9ninUNu/OEAZBvsorsAXQJu5O5cjHavZnpCIfbQNtjfmW2f
0aGZBL6tsiLnX7hVjSiYeYVgdG1wvnz/9JYWljur149UomCJocjkOtAlAtiOXDtE2j9X9B0eRTdy
ODH2r5ZAbWAvxEQybG91yvF6vbRNqFwLwnbDJsIDkHjpAuMAnEL2LMoDrzMF0ifvKgLVfJxmHeWw
O758e7Ob0jjEIe0od4Gk3T3pygFYqTxyqoSSrEqETPoF7g1vubcInkTnFVcDl+9pPb5bOaNqTK+W
YiAJExOfaA2U1AO3lRM72z9Bmga7WJdcyJKfZOYriWtyFHuTowMCEGdaLusU2bp5IJLX5G2NjeiF
ZF9wOf11wVrAMF5Ipb9TOEgM95wqQFQtxV3w0oGoqe0/ntmwKOW+Q0K2woRI9JhEh/uwhbnHcQNR
egoTGKs043u878LeNsViO+T2QIBn0tOojyifwAY+3czQvhff6HZAb2GvIv9s3/sYS3Tc2kbEXEeJ
EVTdk1295Bok76dAMPUW4rJETGIXiwiodYjjnnQK4MBXG5flTXgKU/7OFRhSCzKBvuw+foMfoa4w
bIrvBESWpV4/SdkrxjOg2MEeVG1JasEOWrRnn/eNilSl43a28RryNtt4mcDJ0Tk6tglF4w+UCh7p
IpeX8YLxXGEq8noLJoCneYu37VngqCQ/A4coIERpAM3386l3RW78atvDvdPCOyo1aFAwC1uFnwle
02OTYZwY0gg6wXjiDShOq0iaTl/bXTtz8m4Clqgsz1z2T75/PGopi6cHlp35jraUDH2hc5xMlVQb
CN9toeP63/xA9j/fID8zmAQUBA+BAqDDiKPcSM1sy4hyG57lhew/+328Z/LsL6UG3T0tPRrrOCm3
lx7asIc/MFNGDYKYg8j53KWHHmu5Wpo0XaaS8VXa359wPOsDeOiVln8xL9mSqGiUIR277DCXwmYv
V4i8yeZYmzQ7oVfC74kmMsKdZyCtPPccXBTXPh3gHwTrYp6p9/FdcxZsuIASAQZ/6H2cr1m3E4qa
QrfvW8m3hRSKIczIS8RJoJt9vA389KX4k9XzHrRA5KdJFddEx7WY93dF8DP9KmgvnXuUtuFAwAWl
vXOR3kcIqnHIYEPn8F5iBi1/ZCDQOEcq6baTzw6TDdRipLKBQ6YzbH7fY+kbuxDcFRz7FEf6ueWh
o2NlxLzDx89b2dbtqCofSgelEe0/hi4hbVMq/OPY9+ud08T32x3dT2kmfOU8ggGUEdUqeJkzCckY
FHdAjGSx0eUbHLYMD7qensjQhwhNzNjCNM8jZ7Z90hbysFil8AEJpu0/48tg2Ic+62/VIdoPI9I0
p6CrItLOUD2gjdoln0APlmkhc25hAGkA0A4HjtLnLO1lJJd6iSyoA4d6Z4XL6/QTey3Gp7EhzErw
qdeA1SUl390bokV87kesQovlhu3bDLZUPwUbkBxWRC+1el28MMr0T6M4dXPd8yuZFekV0KebrYjP
RSYikzEVW0JN7+unNby9qc5j5uv/X0WibEsmq1SgMZjQJFS898PIHC0Csn9rowjKyTRZ6jch6iPr
C/pDhKt4PcDdNCKz8/vnkuY2Hj2PV8iaf0SC85oRlrtuWtwhzik3VffHaL2CPRZIAeIIPB6bnbZe
LJy9RctSNmCbXUOSj6CNkMVZePJkodBVpBDQmf+ZEs443CI/6nv9MHwLokD0v/FmnxiW6PF8/cbk
090tzWPiVSTQ/7Kpaujfw2AcchKNu6eqml3VSUhHZ9gaNhBU1jANM+R5ethILMefH3B9V86RkN/4
gc3F874sdervwBVUmW5gx1ja8ra6IPNcuWsrgN6TKnnRg78xE0IZpyHe0xdyXXjcT9snx+YStooa
1sKIbnQlTaEDH/yWvpUF31tRtSk4EunKxgcI46oK4uXlbi21CM6PA3FwSb9BtaynhOID5069Sj3e
xaeoj3AMeQACX2O400BJee74URbVUjTM4dUrjXn2YH45YQctDDLrEngSw7kkCETRY71sfGER7hoW
8Dt/udoT42v9zf0fr/soYsD5r/BOgJoasgZe2YfoaRV1oSTMzh5ZklZ8JlHRCyiqoDWkkWfBFrWZ
p5U0h3LUp98NYW+PHlUPi7TE9jCydJUN6RorRe/jszK0PAOhn4vsUjxk0t9GuXYH1W2aDe6j8QB1
wdCMjrVWqJ8JNhjbr3f0sRHS0cOytzKZwIBLyrzSBbM6Hf3wxu3sYrLMA3HvY27s/rQGE+r1BaCt
hdRqf0bh1J5a+JyMahLPKiujfXcAV/xR+tQNaSZqAZdCWDKO1hy+5qzZEsgHHnv9Itt/OCP6Boo7
bjoLFTnhUsfoGxzhCBftxv4cfF6iBu1qNuoupRfdXoZh++E2STVWtKUGvKBvB7JjA5L14WVwLPEY
ZpSRgtyjJxjosCX/bRmUdnmvjAkdlpx2erh1g1nFYw/uS1rjPVR1p9Bl6G+Z76xcTjBbY6XSK7Bh
EY+yB4sIsUViYHDwl7qqfaLXo6brp7/L6GgW85mVkPFoMaPqDVx3Z72pvHeKUeOZCGilHyfnbVQp
MmzbijfkqLWoCg6SNhMWTZpH58kLE0XDySEkjukub8tYoO7XTb+oOQiH4oPhzJxQyIHFqySUneqV
6ClsuPKLS3mo/E3/GCYuT5bZ6ggZzVwft3kdEuC9Loha46F7C5smRmWt3eRI/QOcXeL8RUl3231X
yoUXygOe+SP0VLDMUnmL+LBPRbfAU4LvhoUTN70nyOU/sfmMpqYIFkysHbuRP8Y80RYl86qYpRt+
bjGn52Er/6HEm0iCepP//MgDdKNxwLldY9oYmFTWDEovAxk8k7Kj4INEKds8x+e0x9tBFvxAWO5Q
7tRa0nRJgQn0xwdArLdcwqiwC41OyKJic6TgSkQ7t5QSYhRjXaqoaf1wkps94WqSBIGweePdvM8j
CPxgdThN9DUpfvUuO23xs+cFhzlmvEy3U2dfsbCp60+70ly+olTwPileBdezfn92p3dWIlEjuCv0
ZahX7iAilVFfeyg/L6j5GzaKaEr2bpnSFXAl7Znn+4HsG0//fLeaI7M6NjQIazNby2RTajR6GS0Z
BhY7h7XDHL1Z/4QaB+LaWzzrOArX88YUgn3fdIPS+nzgCpQ8N9QNiAnxsrDxyUfjbME9l8dsdY+I
o6bbAKzCTGYHNSBZKmXzu9VTW9X4AJaiG6OJY5olSQQCVNGzn8CCHQZ7Nx9DLIIcm7hVfqcNI0Yn
ZKX1m8cJK4eNkLtGRIemBd7jpBqo6YXE5oEfay7Xd04lexwKERCCGv0+EVvRoFTFqS+aZtBecK8c
bAWRCq/J2FlwjaQQifFOhIVEr2nRerrJZ9VeVxzdTXT8744Vk3CKKwzfIW+0xTHWztaRiTWhJhKe
6AaGfTnEq29pIgPzW2JzczY3ZBj0FkS4ZkuqgWEef+G0hNgaU2ArCjxOEqhCLI92sOik3k91d7r2
rX56sKrkAU8Fku8OpNwe+enBcOHMcsc9bTfqd1moDzo7rqpzk/EzOHxG0w+8x41rckyU2NauAS28
tHPHE5LcCvyNq40XMFyArcItznauK6kTdVA6eyK3ASsn9dTGTAg9htAeGd6LE/llrPqMekVAD8R5
wquaqg0u8L6bTUewn8bEeoz1fcy2E3o29L3D2FkvRs+yrh0hNmnndsRSnXgYyrokBGWsjeqx/inv
LMuKUMwaHW8sV30JlAZoDLT+NOmHkyAKT5SzTQsNoqaa7857vfPnFJmi66H4EBHukOcXyCbrRL6r
g4oU48ynB/3mBy3cj8InrD1JlJScYJE+aTRk3MYZB+lRF4bdSdHyK1Z6GunczpAVOyMGDE/nQuTe
Oco1F+HDCWzhtvO/2Y8goLbcG73nAsLSVRX4Z7Rxpx/oiYHzbLmUCwC49j+sKoP2pc4zHzMorlcA
FdLzByui0LMhG00o0lqK0Say3VzFeTGyh/hRn2lhc7zvEQ//gMEdSI11LZihG4EvB4f4tBVJDECB
46M6xWpClo5wlLRPm5B3+6F6gvR+4zYQVRU0jcVPfTngji7x9EnFlt8YL7LlKldYVmePKTVOTdh7
7Uhqw2pL9vKSANeLjwq3J0xDazyTN36JP+qw6IwIDnVspmgOa1+rSN4xlVD8lt2JegvKGCFytWxt
v5XicM8DC8eBZbMCT3KVIkY8H74NVgFBmrnKCbSfKCHt6IvDKvqx3buwFekM/SyGTT4lRimCJ3Pr
OvYPuh5yBkBipTdDg7VG700rfPdfSMk1k0X8j6+ACDDbAQ7gCSGXxDhp64tBBP6HF0oqVfYt6LqK
qEq8JM+qA8DucT9+MDFoCFZMYkw+FdJFqZvLl+1zR/lj/EYKQvMqm6H+8TcM0gpK0/DMTtytipkV
LvSihQ/1rV4Eu9tiA21Rxu604J/MsXyj6GMzxfAmMn5qElil1JARbXPDGrxZNnDtM7JIrWPA4ImR
HnNfkalTxN1EkBbqhKBUq0zOPyDZhDAkRpksgTkXHEpjWBDV7YEn4gheZe1eMWv0liH/hX+dcHx6
0pqTMsEVpyLt5xfxl78nhL4nEku+OFsaMm2hTnXZAmVdzckxEEP+nq1hk3tTwNulrSVEuGHoadjH
dW08owl9+BFZGfF+IypSeRloxHzRN8e8JQ21G21uzUUfPbhQ+ynY4Q0Oc2ZQUEXEBYcNYHWWeS6L
6srok9fpfOCfz1ql4PG2VjksLWMnT/gKYVCeKqVtEHBopvjoRnHC5RwG5bm9RtMHU5JgLhyGKf+s
cYZt8XvrApCPl3RoZV14AhY1bFdOHK5iN+NKx95GmMaAn0b3Fm09ejYQb2rwacHg2zjZ9RA2wkvg
pcM+tpTPJLvBemksGyztOmDr7m2fxQLeLBigw7p5HGwZdcew6qrgvvX/ZDBSW1jHC0qyv4gxVcI9
gNgqaUukw8ln/eUtVdqB7Sd/WDm0omNGf9YopSOI68mzEYyPG1rzSoGZKfty382SdQIH30tTJRZt
Xr7IpgnIOl+3Eli5ivRgkFsL7DD6izdqH0bRa681OMC8QaMIWxf85Fty3OxJqbUatCA7s4ydU/Ta
8uSNN41SlIAoSbnJU40ggC3kRajZ5YhzM4h8fyalHHaxrrDPXRurVXXyXHpcs7HHqVx9TAUfnIEQ
IU9BaWJ6j0QLs4FE5siVA90ogBOmq2d+H+zXPGnabedhf3EnTx89k3JuyTwLAwxY6rCmvWcbBWlb
w6NvXI+daYKMS5RmIT4FCx5rkgSrSD+RJXp+c6LhhF62iHzm7GRrYMFdJfDJv4VTNPe5CZ64U4/w
UFpJihTVDr+XmlFFwAapss6FEvv4YuirK8Zw4YM1G9m+T0kd/McUvsxbLvDzwhaOXjYIAWYURUzW
i33C/764U+zfrAj808SXH0gGPJ254byjmQAQqgkpsjsQngxl2vzPe6d1JdKNeEdSL+vd/xzQdqil
0MKaGU21cbxyKDGtUfpWmLE7I0DdeONGYkWJ6Mmo8fiw6ktwYNZG6D1jIhXjr77xLVOssy6Nru41
1AiTFQTAU8X4yUsbEb9Gm3jhBAdTREoP+ry7v3OhMnjNSW7ukld7A3fce+QX4ecBZ+/FMb9GL12M
fK9ic1Vq2cd60oS0XcC9jSm5eWkzJYSYzUbDTdKqFVWEis3yPfmk79mgwEJhs96xqbsKYgQQeEZT
szhl7vbXk610vzIM3fNMeHOLORT/m+tFJC+g+zPh0WbuEGQw9Vng1rEwcmCYYfRpiMLqtvTwtZ+S
gegTpFjsUwJZoynHhp8jV4YN0JQ3jvaSLF+wtT+6mUiIE6PTNyTWTeEe0j2tJrRm7X3AOHbtyXnL
COX6x2UXPIwiX1VdD1rpurXQ0ib3QRhlc12BNUzXmPCJtapEoWagF2+ZPOh5uM9LpatmucVIGxXm
6xWOfbQNJk98KxzCo/OFpQZGFiNhw2PeEWhlkZnrU07IHjOQv7+x8vj7fLkID9PrwoiBp3PR917y
ftChxD5pctnN3UEfm1tdzxWjyyqUkFY5f3j2VdwnbKqtmq6F+qHVF6D1jzWzD7ivc4MnTpNLuZnA
Jd3aPSODolPrjpaKPA6Tx0Y4j5k7FzygzP99NQyf2Sho3BmOEvnnC1QJrlhFhBe800DeGPo2lrCb
tjTgYdGaNRL3mE2n3mrhu/M4otM8gvBgK0wYRoJL4bC7Nec+0xk0ifEE1H7ar7Csdz7AV8Iaa5bv
YzebIBmU9HRzXHrNIOKYewavRakOU27g9bs0/n/yCFUFnAagf6FF0kg/Qp7jfLTW08pc+ggO/9k/
wBmV0yMo6QCkJ2g83eq2KkMs1HgGd2Z75i4f+6ZTHH0iaUIdN0jmsg1iHWUQYXQOQfRQ5XN9LgaY
bEkb5Ba4hcEquT47nuPu+MVaXTLrAuyHSpU27aI/1mB8xeGapYJYaw5TtSkrOYAv6ub0INOXPBVA
+nG+Lw0pLtQVRYI62FRRWliOYSATGAMUWAmKtNzt7cQpHLfstfFcoQjHxs5brFJRpscIb6U2e7j4
ihRKRlN8T55pEi/DuaDh2VGRXjrEuv3calLrXBvJMqRiGhuR/NhLIXHT/fFqPLPu/z1ELBfm4wAn
Z7OXbgZtz/JumA9qrub+D3NxRhlI69PyMbUV74Os1m3EGHX3O6+Y01A5CJwwD0ygdlYoxHgjKwo6
xrlcQiugdgoeo84qcsbPwQ6Sl0Fz+xeZciYOJtwfJrx6C7XC1/2iiCI0xX/efarvYFSVBfis+B65
zJFgnKd0Qck7inCv2XYmp20liWN82RHhVhc2BuzTww5kvKxPgS8j9eT485mTx/8mMua1Fuub6ka7
i/f/gi+HXzGUYjAbMdMlEMQbM7sgadXQy70VxwbzbIZORg8UHQy8IEb5Wu1CgE2V5ljWYVSPFuCR
KSScKHbFIA2HQSAxZllbp6iQo0+RfUvGGc4ohzKCPc67+yCrzCroy+Vc18SvF+g77sJIeWt9gt1C
ruS49iWF4nO+7OMX9fuTlAV9Fo1nQSn3bWAuY9azDN/iThjADhaq+lSSqxkqoVoCJ1MnJUcTs2x8
NK+uODANHQ2qsWHDfrsANeA2ksg45v14GkRwrBRXUTzCGJFUep+htuC5qGmn2kdD3LdEORKZCJnp
aXIVaYicaV08DfV/fq9fXGVNpEZh3DRl0FdPMBM67BBY72RtSfCKG8zjKuyRYDvxbHUS3nuqPTqW
UKmTuJIWbobA6gdl0xiddOK39cF+HCYGTHIoU2LPnIFy8hq+havd82rVLsajNFNkbpx1Q4GpzMmP
ElOrvN8MZIco/K6Cp9dny/QgfrVFdWhKwSOLyC0y0p/JB2snOj7jwcHI+bDMjRyE5BEjku8u0D92
JA4uvPyCZfyk0CVyftUOO1rHqXMLyJL1v4b5Wxt/Atcs/OpyfSQZFKszQl1VDByDs8hw6l3JBwR2
3g6f5/YwVsPJcowOhaWZcMb8XADgRwlBJIEwYH3PPwk5OW/uBXNmM0Rd6UQc+xzA1rzDpvJwWhuE
U6t26wyt9d/2Lv1T2sk7vzk+sjXJHmA3DYl/rPTx9eYu2iNu1pkmrOoOJOHASNajb1kOShrk3Ha5
tkRAI8EopjL1zZbSn0yyc5syS5fevbg4tcWErpi3YoTygoguFOlrDOtco9h9+tPczc2WTmaG/d5a
RO3gDCaC2bK9UfGH2FUK7QCKrk17ODe9PZZLwPfqJ5QgRXe4MoMrDEguk0ooXhrFoNBnELehCRBo
svmooYMpw8qcjvqCuuO8zo4hug2lPrD1+RspvhA5FC7yHvU2QBn6e9N6iU1e/LN7tCC7sh+vqOHE
7y6k7pvsa1GPUklxUCpT/uaUEF3PUs7bWENPoFvZq+TG68Z1jaJArMu42yuC7/zvRAVEyb+6fL3J
sa4Sr9lhRS6fUf3WdzxjZdfhIPV4spiJbAUCZp9VRxaR3kjGq1advVTxwJK1sV/g9eukQ3NtGeJu
uhcH1qqJOzLfwpydaV33BbDnm82cAbHca1wNi/S7iZ1BjWBCoc5vnSpp+ULt0GJBEXq9I9QP35UY
BMKrd/5CdvsKbZlDZaVZTS1OXrzwWLKU/M+PkI/6aH7fQQSepGENxT7Nk1fQK6PTa3iVVserV5zV
QKtElbQF5u13nrJYsjxSIFRBMDkeYUt7+9SRHSqtyKvnS231PhxMB3dhR/5MF/OSOnzb9xqB5O6i
wQ6JJTqKbRLRFlFn+eVBygs4lr5dVgftIeEnGjEmt/79zpgVGUexhJ/GUQHyi0cvF46N/m6SF0eD
NBJDAX7fIxQW9KaymYCJlSZcSHDxk7y+MSdXNjRbfPyTEZcFzEXKEPOI8Zt3OfQ0lYvUPWL34w5S
9gHbK61N6odkGyyacV4ChTGc0B8kayrfWLThuhj9Ikoe8D7bMo2a9uvz06Qp68jicdf/mvhmo1wr
a5B8YqJZS06pUiM9XzAHF8okb5keadYn4mPLFyodCrFHpb7xXHpXL1EKbRFEWdh2r+smrLULdwZP
vj0XyS+2QHu+iLvft3LPRKg0Atzw7OiMWCucE5eC1WJyJMoS+50H4aFbSzajuAyqInnOXc2Q4GYU
1nEuV8n7/sDHw9RwUik4LHjKzD72ztWEgxNCckLobmZSltOiYUGQsTUko0gBsz+87ZsgSKSw7Zr9
1V5yh6B1+hzVTTbvpumDUXiF+xZSnI6Qm9n/4gq/Xks45D1RMifY9YDm0/jtSCp/ilVwF3HT0E5g
FQV7KuqsgMc8yiR7rQ2A3PfpwufnIOUSC2v/btYkYWViqYxBlm5my63p4UTeHbgBp6R38XXhbxzu
+ao9tvE00pHDjms4Fap/QK0FFNh2T+uk8a+9T4OL48VHJUPapZZx1t8g/ER63+fAFs7/ZPIWb9G9
T9fWr35/7jrU2gQVvvndSDDLzWXdyN+RR98Nb5qoesKuFS74rA8lKK+wnM89iOgzEfIZBoYvTv3y
oxa4/lqOlg0gkS42biKZANBcIa71eIl5HMMHUms8xLKVM9wbBAkVghCb/AXSZFksWtpDnucgozMR
eaeph89UPWy3m+dhbH0iLDsdykvNqYG/TfuO+0LKW+CTO0FtexcZxaGr+hAe1IfpVYeS4JHMfark
+WqJXS4sDrJI6Ym6n9AjqFbxDvEqCJ1IOwYp7sLjhnLugtvXraV/w1O4knakusUI1nNDrdBPn1mI
1XChfg3FwQTW+l2FTNsW3ptdNqOrFIevP75j9LmpNtorJ/CJ1jLfV83ld2M/XOBLKpu12R/Tmm5s
AGsQeWXxNfouGEtbLNYObm8lEVYoGOrZefAJ7fN5eRPqtT6/cPayMWS5DRByF95XGvuzohKqtUZw
eC34dnZPuFFVAiHga1VYjpsBL9rcJ9EyH2xyLJMITv31toUh8YspUDQpfHmV1PoTgJjmeSTFUI4E
uKcHZitvTp7hreXPW6HNqpq7Yu1bqnG2bftmvzttiudiA63BGeKs4L1piJMZp22+FTmdFDrG+gR7
2QI3Zu1G4sHlSIJOHFYHkETpa/DQ8OGRHnswHsLt7yTSFG0dtcYTLw1Yx34GFloD9Xmbm1QPx9AU
2jISoGIOWsgoyc+phfRTkoVdGwpsGDnTYEu3vBGOaGsiea0zaOOAFNJYEwMIT3TSYTFeErJrGvDY
2z016QG/aAQYuBvzCiaGM6sZWXJyt8J5XjLGXa0wGOHLKcBCiAPw/fgIX86eIR8vnPDNsuESDnro
8Uv2LOvJqx+p9uYGHul4C1mgi8t2TyRY1RAj2/E2yOmVsESv17Z6UVx1Rsk8uvYM6xC81LK8udVn
mE8bmt7lylf8/97kErHwecK0gK9hSu1FotOwGQFLCQbZtcD4Uvx0LnvN8zzVeal9V5GetCBec+kN
PMKUzkD5bskvzwuWAegfVE/XhJt5z/pW4qeMWZvS9k7Ceq/mfczBknMX7jArzajv/vYGrV9FhGZG
jCZu/7ka/TWSdbmeUvRPVFLlzjk5Ybj0qyrOT1ai5Gm9CKf+bmN+WJL1cG3nKSCaGGJXgYjF9hUn
KKwdudW3ssCp62PoV+GqAdkkSzTxQhFXtQXx4Mto+jYftwRjNwXN0SKxKU66kMoXHDpHHobG63mf
VXkTzuN8mmsjYNBbh1cNsKGqbM+d257Q3NpE5twBE7U/bqp4HZ70R8hyELdAitB57j+A/KntHdsw
tMq0I1qVWtkBgVEg01e1u6tfqAOubtOl7AI0tM/Uu3KJ8DhX7sbo4dwDy7I47VulRbizdCWYhqta
MHJzsDT+1WXkNiUlC1aJevBvX4YuUP9IviqROdEZCpYrwlUi/uoP7Xa2cibmkzCoPqGI0XbkTrxJ
2OxBVL+AkQXv8+utHj50r+96Pm7Yf5ad2SwSJwdAhmG2W4059dMyOuilG5IijRGmIF86mRo+msMC
VU7TjgJ1ST/5D6/nO43OfCbNkP2NeMEgoi/d/KIOhLaAQVoGdWgyNa5AYX1xLOKkarC8wJil2+fQ
yGuKFqZITM9f5CflQrZGmDqpf/urPJp1UrLyhf1L/gkpDjR/oX1yLWIrknr8uWcM7vVXl4ez3sYl
W8yDJBdmbDLkOd6P83yxU5iIh1s3qnDWD8IzThBazaHHAaiHGi67Q0b0mY7MK5g2a5PwqWE+Q9RL
KK7hSEggCJLuqxYRc7VMlc0SJQoqkJZ5Aww6rFyZNUGFoBNObWGJ2G1+6unMHEvBoyW+O1VPttAF
2YKU9ZPFyeN8yQ/HW4so29UmttNJefzjrmdL5uRi1yApyLVC7cvb/JmM3hAl+fb3HC/3x2WntQk6
XycOpp9kp5c6qLwoEKxmqqHKxrWde0WNDdSNkBEMeTDRms4Oggil2gjdUoa6pGoKBvUQnQKHX+GM
Zpxwh5l1c+88sMyPcPir1ByRcj0/VGa8gzz32SE28aIuswnM63WAAieXP8rQ7E/Wuh8/FVEzXC09
jsqScgs+Do1yAdiODBJXHznGzSqzdI4yT1J079LGuua47y9+U0yc8ijfDAMNz93R72lAyx443j+f
MjBphuBcPPzoPhRTpHPBQffbsiJCvn9UuPjwa/gXAzql2Kc4cJM1W5wpB7AzqErEXRa4tPiQ+//Y
AHFrHUFB/S/Gu7J4Yv9sS4RwrOa89RdInR91TEo6fgrIAsBLGJvcLf4bjPbuxRrvGGj9+OrvV2oj
SmTT/MDlkIPbo9gSczJAzQulVL3f7GpbLmsgCznRGuL8U7QTAqYwB1Wy1/8qiRoGApPvO2S7SK8V
/sDva7v+HARhvGRoU7AVw1t1tgcvrylRqkn8G3T74Pbdr7YA+8I2wXoWH2h2xCJX5mc1xCv7R22w
0aRka1ZOzIwpS+JaZDabVa95Htg0Ypbh7IrSN6NcSBfjxLoewj7FYZ4RB+1VvydU0mgtKyn+2TSn
mwRGu1rwZvGXuprm4w7/hTYh5Zop62jYtCscRuaUV3MKFjcX9vlhJlNeMelnk0is4l+ZXuvVuwmg
7s9QZd8K1ZHcVElVfSRHfeMV+8bAx0cr85zSFH+xp1iIlrl8tR9c0uhhyKVEZvjfRMXIvEn/24jh
tdT9725cLOFzxtP5xnPIhKdPUjgLZUmFKTUYqb3021jRrYgqdkYHau4jRfeouMMRF77pBTDMVEcd
rhGFr/vLLZVIpqtcD0BW/jMJpGb+WtIUAThI5E3olbCJQp2UqtjVDLNOCD2xZ+9uOuUflL8ZgZfw
DpqzAwYz82UDE9lM9F2yHyXmVUIrl8ZJqT3gYzs5JRFEpnLjOB00b+kC3Ucx6qXdh6oISZW4qoiE
ZDFqMPrLzmlWor8nHE7dpk0KKdcf/wzTbi+l+eGHyZv9VhSAwUFRP6SfVyUFg7VMEcBu3EuQdOz3
9lMkg1/ErQg5vvbjTibj+ooeAtyVsWe+hhoSySU97EsDP5lP2A/9RngmZ9hUmyY6tB9PxdZtQULL
PoAtJ4+vAsu7RwmNsvYJjMzQqXkFk5b1ZUsFPWdidkRLpNjDeXwTx/22TZZ6aqkbbtMlCp7YwW5T
ZMtYc7nsbzT8kbuKzec08w49jBFE7AO24kGu4lJRpoacq+sUpWN3ou7vm/gjqVLDgr1e2lXo61+h
41ovpGfKDIEnmUOha+EPy7/0SNKn5GZjPKqq+4nxgGy8uC6vOq7KmB84MskqW8kZQN9QfEX9maeX
RbTs7V3HaEe0p+2gN57kA6QXJfCb5wF++v+7TVAPk3lBbFNS9mllN7DM1f5h5cDz0adwDVRn41hs
CJ1W4HA4fjAR1nwnnbp0PMVxDLecZj5+UqX8Gn6nMEYRhWNgzPWyP5QYIVY1zab82J6IJk3Aro6I
F2uDloIcKw9UYJ0y9uSvmUBqasSiRlQHRYQyKZek7AF42m2jmzrrJ9C5ykiU9E1P5JgSUEUln1ul
rqiivtzPnzxF5fn6ZUjFRSHuZ3Np1ksJx90fQ9uBxT3sSItLkNEvnMLgeVbbFGTjDqX6OoZKDvXt
AULkFSCopiSq0Z6m/BnxGuhpUVevgeD/4h8RqU2/jYehVQNCzd0F+zWU4OFGJvMDa4meSKsXr89e
u/WD6ac6CH2epCuIQkUAVIy+U82gG85iFWRkr11/Zc+0hnq2s13L27Yd+GUtv7wzcVFMfY9SIGFA
VZHblFVZN98+8g/sypJcMcoqpS9nKrU0XmdRtn8pnzGvDOR2SgY1zX9oIW4b5WV6LY6/jmgFLK/m
pl/fCy8EjmR0DRZro0ku/vUG2gXtUE/xrwtaIDIn/Yi3ztp6FK2U+Qz4SFCaV1jKdB/SVqe3Y1z0
DC3Y/8HuPY+bo/qOnHcG6A+Eqo7KPTkUFshD7xnqua4LmrIjmDlFVpQsQ0nVxwR0kkR6JdFP8V27
GiUQzMXZHXnoeuIPB2AUibuJCz9uJrcVInC3pPznk4oYhMVnZRFGst7azX0nObAkb8ZAflGT8Vc2
QAckEhmi9ma7SdnjizKPCSwScvGf4xRp/sX7wdCU59xl670VVIw3WlCkx2pYFVnfrK+zOBKe3p2p
OwntiEPefyT4I4tHc5dnpYlLs2YvfrvFtnH4nfQ/FrkmnXm8sVaZOf2VOftLvU2CGGUZHEKJdUWV
UNR48K1hL/TSk5qyPTXiNP50zDvwc4X1gqZU+OLOwUcTLz+F5lsgyM2jTP9Ca9T8A+XrPR1Y/Jgq
S9aVKPEExHq1nSfzSkyCKLMdKuv0NlBviaBo+jFf79auCLJ1RbXwxt3Y9jhPYk7+hAWiT/7Tma8u
wHrQJFIHBJaLE2/yBMNXT9/AxllG0/OvrSmQLrITevKam/txrcEsXxeEjOMG85w987rJ6appaaMX
1cPkuQF2fdGHaJwrZ0OcjoV/qaiEKcgTjiiA2IG75sGVtx/yDQks+Nx+vgIqZWei3kiRx4yiXR/x
G1xwecbCbyFMgHAF5WFSxkx5MhZD3XLwa0kaRP+bCoSSWQ9gTAQv5jQe0I/2bL3Ms9aa0mxVdplz
MNhxAt7UmNHkDvw3DswlHcsyZYIp8XaPn5Sb04JUN+wiL0dG7sug/csqGE2t40P7l+BLyugatDuU
VQSlXcCc0FLae6B3R3kYtNPhfOxoQrRMclCiskfjhbUAwgBT+VcdUbaANPtjHol/A5AAPjXNiR6h
+/xPvGc9KgrHyU7Hvs1BdfQdjNfK+dqdIJfCp//FEGi2om9ARVIqFNdNiYjLUeSab/rHRDUq0G0j
RHGb69zZSB4AU5K51aFnPOTRM/mthnMIjUnDXvIUArDvRyYgrd7iGcSgH8WzJfn3G2y0IVCMB5Yl
Ol+N2RZwUknGxv5lf+7wLLUWKt+J39JbmwAy/b2p3q3IKwgm46GlU9sP/28M4bHQgsARrycPv06v
3rQhyH/gxt0K9pKTZ9a63dXjLcy020JOfTpljp0W4p5YnQC7O9+YxKGsqF4xpDFK7SLQr3CLh4ZD
UItlAzU3q82DPX6/3ek7R2yPKxFHIJsldCgu1fWZHUenROVaTakHiARB7/JsP1nXCLw1+95L1fNq
ZpK5615AACR6XJFP7f2dcnx9oMTcAPaqioortIA8APXR8i3/2TYVJ1/MSTEyccOFjMKzPCgvDZtf
xtmKdHa0OuFwsR/FKAR+qIneOZ1wvoJ2iPSyyjCykygvhrSEoQ9ew+tdFUyr18OGzS9LUGn6xoaH
s1LRbTimCjGYg9FeZSKZAMDSNjogazD84UZqLNm4JVHYeiLHdw3lF3vpgIoQvVRP+7r+oF74yGP2
unWfbYisk/vepCvkzOoPnzCc0R4VSiOl/S4OXJt5dcHDf8vZKigd48Be5o/wqnfQ+wA1yPN6JATi
xi4bpMa85lmwF4OyxEQ4FGOJI8R4vPJ5F1PWheQV4T+i+7se8B4qa1XExJfs6iK0dx5b8oqMUKiD
6Pye/SvbROZ654/DQDx0kvfR0wmXlXHUW1koLZpNz5jLzegmudLj21XsgHFbcc99Lvq78I4pKRld
lYuBfHJqBFQ/19kSYhNNfzldig/LS6IUTPIKq+KlaqW/I3AhsFDfAxik3eTOROdRAeRzzCfIBn4T
/VhAErKvAHzZ6U77gTK/+OA0Dfk84azOT2g8suY/h6j/IYIu/3J6wsOr+ZPBAdRbFk4zSXE112LO
GRGq4+XVw+IRB+8HPZ98etNln7zC5sXZaM+DiaanOpTWBNMDsLQSUnKXsCPoI8HtAgdYKe8eF4YS
QUi2Y5xWqAZA33vQkG3IVpO0zcus2VTmSiI1i+OMFEgJ5oSCG0FzmEnnBMAdDzjj6zTKYeTwicaG
0Bld3myCNEhaQaP+75r/4Sioq18lfFSqV/JDDpMkYMKre48Ik7LkUkwUiSTtqkHi9i7LxosuZ9JT
lJ5uR3pBQRmowoZTrc5XtSFokJhm9gI2CWxXvIL5vlv6l4/DMX9JD+p1F1pskePKp3spCJY893oZ
iT4pKPxFCK3sJiUjzBPgbIQz8WpfC8AV1FHY1iL3TotZdufy9JIVWANmNV7xSIHToJc+QjHrDC6D
I+Z24+E/OskekTkj4HGvoH+nVaXIJoYbvPgGJlY2Q226bXU9VzOtgZtjQV26nEGzpX3ZYui4b+kx
dbLJWnqAxz0UQFWTb8SWZdYNcT1ICaH+GqCG7feh222mK2brnmDkr/lHotapvkAI6ARHMralwYa6
68cpExg6kTcRlwLXQijTfR+zoIZ1CNOZN9kETd6sbq7AR/ldd2RydTg783C9M0zVqBjQXlzc3PTa
U5yNpx+CRxPQoJ8hGf6le7IQNjVIE79qxyBn7/bmFvf3yhzgrSOKsbCBWW5851An2TqUEYQRgP9a
n9az8qPXAiWSD2sRNVJhNx1ESfnjua44288+Qcq0YgQXLkit+fpT8bbMeHT9xqtc5qBmJK0mhPT4
ag0VQxA/PC485FfWHmVwvKeuQyfo9WV9xRzxu64It+HOItVu4dqLI1QhGLqNFKjWgSw8jawFNDYh
YYoW9W8ScHbWvnYTDUhQtrkKWOttDLb/Q3AyC+Y3yhBPqbxQY3kBKe1m8oATyQlypLNa2mXDsaB4
XA+fu42jGuVnZ8+0JYB1aYQ7nqPMxFbJKjPfpJCuR9RBp0MtcmYC4FSiip/oYhL7KjMTxVIcFrPm
18FyVVzmE3Uw6qSnzUcY+4MX/NFev0hZ0ycs0rRPqevYgCtybNNleWHKFyj3wLuiGOtpaPNpjrUC
Vgx3sahbXN4PQGcH8EuNXvzCedkqt3i3J9s6HoEIxxBL4gxI3xxIXIGtOMW5/SvcgBZkJQTRCd1n
OmdLArku1jLQwU8Df9uVt8hnwHfOyKIpXyZJGyrzciJno6naHZHxDPiEMpcpV964R5z3wJUa9HJm
r/VpIvAI7uUD6CXbSxBPU/8kwQjAvzePsIdaY96EhTpRvLAl/ve09m74RTEqFhMJVNd6ZUutbacA
8fh4Ci/qwAFO//m6rpQAciTkTiXEnGNudWmbz5wvf7tBGXmifwAIdQbJEA/REzegHnCa9NYCVsIy
Lk61NDwtGzVs3IbzJo1yGJjZVW831aYwpmsoGaUq5sxsM/1/iXLxE/gsIZCyVxhYDNjONO46P3Wo
tYN2zqI9WfH9lhVepIiK31OZfuj9cPBj0mxtoyuLjmOp4DCKI0Q3//LQHKzvzfNjmwzrs9xfSIrS
AOTPSB80qRHr60k5u3jZ2ekFMNOP4jWjmhwdDpvRKurQ3zsKHGSR6l2bNWduhJbFvIe77nx9PeNG
oeqQ0NNtCu+3333ZX8NIa3JcIpAsdxV9GldSYXBOOJVqySXy8FMrNjbBR4nBPTUcOdAbKwYyM5pJ
q6weh9b3mrL7b0Ch4FmCuyo1up7sre+rdlqQpB+euTPOkXz1HJ+5bgLHUDjOgOL+Vr/V7NR70Lgs
faSwXhfulzGqUEMUHLI9qtKyeaT670Gf+HUWUtOJ8IGXTSI+M2i0yNj8kfsFnaxZJ0mfpxDZWjRK
ntUGzW9bWJhbiLpifjqiwSkrE6EiBhjUqIqmIdRof0FoIsHTwwtP+e9b/66MQjsarbClw44e8pBI
ivuOzRmF8y4V35LfN7XCaBFA9YnACzDn9xShyurUbuxOL4K2TSzfznCBNAk6JlwWIZlGET7rCkDt
K3aaDAAnERmkmRqr02xFgvDf0HCOq2tXxOhrBq5PvGCXwL9zKPZR3QeZn0L9M2ThD4XxhUZZoquq
io+ucwWywT913Imz/2UGaix6XPUzltZCo0uxwVQOyCFHgdCrLgvwfPZgsVVijKQXFQTXZjoSqSg4
X1sfCGvmfGnJC25aWr0C3tgv6BMC+pYEi23Su9hTr0xkg07ZOJGFsX08PLrNlvEuoupwPVQkq9dk
DyJ4moDcDTmN8uQAMBciXpXYahjjuecfUH3j1dMwkHFnDfKInRnKXiB2XdYu7fyRLy2VRRE6N4tJ
0LrgDohQTUTZcGsxRCsCOMwOE/X9JZjZJGiFlMotZai7QCl219DPFpdasWB9r1jnomx9ZDULcQh5
nvW0FmrwNk8v3ow7pPgqAKKfXaX33MKxUxNR146JOPdnEwFy7Pm2eS7N+UsEZlmePot4JKNAr8KR
RevEj7TsK0lhUt0weFwPf86QY9nH94rCV1Wci9K9S1gqxMCeahfpPGhKmkXd/TatH1ayJXAvav+D
R/i46kfkgQS+dtd8nguTX+468upOcSXfR7sHH9dGeNUERBIqsx2QebBsrfe3o3ZLO9jgBc3uex5C
RPug8k3SwZ3KCNGY01jY8qFgsc76RbHfPL+AoKM19v4y6uv/+nYJ1mOZVZ7kZb5By8TD90xDmdAG
HYuyHac4qbhOo/od13WXXJ5IvZm3X/YGiA703JUfRAFiyElGiOgULl+cQn7UeIPv2PQzSwxkJG1e
/D5NC7lA///qM8YsMqW5SNp6jHJ9yFfhMKB5XmgXTbF2VjVICQS+xBzAawHinFUjCk03Vq22jNuP
iqEUq+L+rWR5A1676MbIXIR8TzjOPTsrvDTnBzF1mLcKEU38DnqBbHBjnmqU65r5nPh4EafamnD9
pUo9YzpHT6JzjSWEE3QYvc8NTnX6W2t7KxcWTAO8LBd+vz5mR/uG5ZKwyL+8DDWcT6J25yjlVjgm
Q7txjaSVzvWMQnH7Eefj3L6HUiE9xz0a+Pjb/cLc/YASWvgXI6fszfNO4kQdp4HvjjEHG2fcQqv4
VYa8o94qKg8CQJXva1huKhx8rZll3I/fnp2GsQfsaYCT/dLyyonRei077yov3VZ1lqqrX0UbDmMz
ZZ/+h3xoYxC+iTvLXlaz7EVhenHVG+X+FSmUA1hGZwsfQx51u9ySm70YNKxfzz8tAt/43ObWsWth
kmuRDNHdYNRTisoe+/uoiY5fFCNj3zGG0n/k8GK5MHYE1NKBVwm25j/xgAeO8G735FisAisP5b4J
JMViJ4Yw/M1CS6npofRmKlVlFF75TbSl42X/6hDR0LP4MuxRkFuadsGUzAiASCr2s4lEa14pFtL0
urdORWzBAj7DYplRMmkbxNp+qQT9PL6ZZc3t4gWpqzeCB27aCp4Oml3AlMgjatIDlrVy431+mIrH
KHou3b7SrPHQrzsarb2M/fZAXTUY5ovqwdFp4TbU1FbvFpz8ctK1ahRCV6Gt50gTQsTUKzgRSIIk
sKMwc+hn/HAXZnUiHcm+Q8BeaLdzuY/q1ELoWazDGJwRc17WZgKigmmvTQjyc/v/4GANas74CGRY
7L7bCOicVINgGpw78ExQa4F3FPkRhFDVecPV8fsfmbM2+o27DRmNWgwQeJBPQrIIfdLIo6ize4iR
0objyIFK7cmTykKqIM5q/iCzirPNzzRWMgdZzrcxdXYXL+eiU29SxxEiG2ffCPB5lBUkGO+pehmU
3H9EN8O2NNd0BT6YDIXjIZEkimX1WZBZBvcp1fNEF5/VUN3t8/nh6sjjsx4ttPy6FgP8WRQfmb3C
jNosmk/LIXFBECS7PMpbJNEDzwnrZaPy+ykjmefOmlaNlrtZxaT3u+RmOHWzXvT3Nrel2ppE4yob
47YLVOu0txKZwKNQQWPi+raRZ9W01qXw9ucKAV6EF7pVNCopoewL5+RJW5P2fRyN9zuvTNLzkg8D
qw2Yd0uaCmn9D4pzm2/uXiJ+fV4QcPS8UHGzOaXDeDSm/pq0x+9J5XmTo8F4whbFVGbD/P1ZUtik
7rR82cos2KLkgUdzkK8zLCe9AMLFFRrjNHTNrmXx66Q4IzDxJZg2nyQyWLTHeXNPNWO+MQVN2yWT
WH9F9LfSEJRSjmexguFbLZtKZAaF8fTfQ+9oGNXbXa23A7sMtxVYZsBgipmXfIHGyrJpyk/ed1Hg
dahnvi+DDI40AKi4jg9eAkARAgHw52ODZ14qkYxp4xXbTn7empiiIOClgHPV8dyi8e6UHJ6zumG4
4QvqYx6vR5NMbkyq9icqhQO0lU5kKKQdo+LOPdn1xJjtq0Grg4p/aimTnY7z8ae8zNbyvDJAlgYa
z7JlxAQB9l//OqH7C9Cc5r2azYQnlmLQ+azDCFaJmm+mLQuW6WpAYh/OO0Qgfw3yqQgf7KmohBa0
3z39HYqrMHy9coEgRXB4YMzWJzcm0yL9IGfOKh0aUC0jUHyKyqzTlQzAqC0Fe8jZ9159NyTiE3vr
7vIEsMFUjx7WT6kzuPu4oDEIFLR+cToKYI9+Xw4mxnLXsZcj3coGoHCjQwTNmOuElVt4FDuo4phV
toQ4Myg8W6NLBq+C/VW4eCFdiYWkN1YIfnUqGgpohmTNvcKJjQuvuVe1M/fhc8q0Q7By5a2CLQHA
8zHtlthAgzem1ejiEgxnM1OS89PSVEAiis4C121xuWZEVLtJBaevGiKD2U5Q9gpqH96VR0ClvxII
n51UitiUQwCYS7XibantfZ8jfC89J/FpaWGDaWVZRqGztANsuj2JngTSl6IpZtISdatvyH50nq8N
Ni+VF6FpOwAmtzMRLTCjMnXA+4H7MJrL/QVq4uC+moXPY7C+bDGPLc1Ta7mxKRuU+8gE/gy5Mtrg
PoLcnm9m0jiisdPo9yL1rSchEX+lILlv0QVnkmlh84TE31GDsagaAis0ln8YEqDT6wQx6gpXtqeG
eznwgdIwoSvwvzeg4IQ0T2gdvf4DLWC4HPQtjVHbSwX/caPQn2gtWE+Q24RunGmA5COYa1wpIWyT
MPbIOPiQCj8hlidGihgkbPj0L+rcDAP3zJZ2C7HTc+hkA3lLKnOGP1GOoc+NxtZtyB1xRdgcnHwb
WrBaPal+9l8Cjk9m5lzcZkt3L8ucNwst/KILDJf6a/X3IkLkliQ3i7eRBPj0EwrRByHIfwQdDnDu
T9mE3Q7plQo0A1BX5j+XsHfAsk1bS/7336Ui3bp1GJzzZ0uHkR2gApeu+dI4gymCqDYE1+qKIWN4
04zRrxzYBYmFExzW692J3yLIbXhN58iIi+VOo8Ni3wMHFrxl1YHCxNyYL91t7HpPcyRP0Tuzyr5N
1A/X9dKcm2/wNrgLPGFAhaXzbH6aty5w/ZKmbU/mEuesexSeZ+HfgK5pPz0VE5au26n4hojeuGX/
+TEqGUectoPUThBwhfIKAy/ICor1GVlKD7EB++cvpF88zgxpJUEuuRzqp5USMMoSkDUPBDt1iSe2
yh+hgcKU+Q9lqrjE4eAXu9HrqvSB/qC6G6Ap9PjNq72pq1x8fQ1hFgDd7IAvQVflc6apYjoVuau/
DH1m7ob5AKz5clQsRxlEa7nGeMoElyZo7vH0k2zC3VgiE5lJPNMc/7xELtxEYkPrnrQ39RYQGYcw
VQvcchXCheQN2Cd35AapcKg37tPU2qqdRVBfMwrDJX4h6PHZ29IOHIPV/k625NiGXq2s/hg8e1P+
qaGBcCZsNPEcqbXG9P9gMcfm88wBCO5lVMXPe8BdXGZWomxGwlPstzBcK3pdauOtcNY3rXfpg+Q6
qamcFH4YdoK3oj50u4JRtKCRAPo4CbAK6FDXUSQv2NtykKc308b03/j+q9HxKGSbGjVEN9luoKPc
OSp0Jgiuw5AkklPmKiq7Nr4GMAGi3E9dJM4XUnO2Q59RYV/PeQN7Ml/akTkskvaJ3UAuA6lxuH8w
3u9YGXMYhzVqoP/v7j7Ce8dqe/wKlGHpVZfyRU3n8UkjKslo7/1PNcLt1oUetTZQAeeT0XN+80bs
0qBu3/YanX/CDinaWw4pmlw2QJNbQpCKU777/V5EOo4pB3l3hvfPg+RnfebenjT5tjcrIi/7Xq0s
UVxb1wrvo9nBAfHHOtHzsPR+Bn9JTdvBPrwj3ZCzDS1Y5FqEMFG2kIuprqE9I1Kv2VLESGs6GbsB
CntTy2rDv/LSmWFWEHlxYSzTr03COE1CHwhk85/NDbGo7pLzFOiF8y0WT9lEKwuMll+3NJiUta2H
cvHPrFFDNUH51KTtjjz/qc7Ni8mVIPsbDBO2C2hjJzA7p9Qqoyy5wYVhFv0J566LV9w40YkMgysC
vRVDWy99ojYvd41uCRfp0Nfx09puOmMzxfvCRyzwSd+Zjl7kir/C/7Jhsi8RDonzayvJn3ooQRIq
czOuuEqmuWCVgZP8BqhNdLRLpZzs+8jj85tshYD3I70c9/48iPNx45c8tRpUcLD0GJ954ERDgtJD
khwLGJGY0E5b0Utn0oCXTHD66OYbQcw+AdQdBarJwZbOIYFWh+Kc/yre1rvjQ8BrourYoX2r70cM
I1MclKQod99SJbjynNZU+bIZhFm/INzMY6/xosmmdSJyXDSRLFnYAspmbl2vm4JwL6e1Y0XZAS5n
yRS59lswPcqH6Z41NZ8Tmj7ksBnunyxStSFM8ZnlIma/vP00nri+FKTgkAo3jDm1wP3j8woceXGt
qc8iE3DaIGxJIjhAc0l/bEi/xWHtC/m/exXORBVoAaUFqzlsFB8ZCSnByzwjejWt8PX7oAbro5bh
J9nVRveETo359UdcIyrWgHZrXKI8WnYcbtTzxjucNrXfQPCCb83LJj2kwrFVAocayC4jaG19eDv0
ZoQB76QFvGmAI6jGQYRN2bGCoTUbXLm4hQ07Vu54rX5aLyBo2nslzU4IOQom+qUhAfA8dI1JKDNV
fU8OAi3oxc1Lx3B5BYTAu5m6JXr5vqBeYbDZLJO/31BCfM7EuWP0HJdGRuEPEF4iIe3tC+S+2Fro
HdsEI3Q+AGyT/vxP9ojK4NWXQAccvaK0p3UWNAJ8ZUFaGMdsivN2fwSdZpTJ+izOrGHGYteQcp8Q
DQD0aJ0yp2QNa5pGPf36VIRFn4NPosYf3LX6X1gsbx+VhosDKga1h0qMHEAAWbH8dUy19W0cR8ns
x5x/FNvj/AklBGLkyksPbT9Sowd+lO6rXd0oTcNNxAM/PV8h/w/SpGPXWJ5xRbJVpYt8y1TAEiZG
mjhxUjHrZv8u1I2G0IIm4vh3u8G0RqOoM1bNPcOyhik5cZD7fD9oZPZRn+WYWzyDlpIxKSyI2rn9
dq5k/4EvjE32kJBTHk5xCQhU6S7trsFAFwe4KUvrozmizmhAJJFLyUKm2xlFqKhlXiQ4wxns78eO
jlUF8qk7XYmjOT3mVkk5jogeKRhjbN5hne2kK8v0WCtHIqX/2qdRICIURnHYJ6fI05Ntxf9PgZPe
R4ykE1KeOa3smKlfrEwWYlW5axH/IyUhq9QSfYRTxgPeD9ojt9E+a6MfohJAuH66K6gLsmd+wABB
+tFgbimha0ZjHBqDj31nPfYjXbmZ004S74PEWaFSA3tBRFe913IWbMTCPDo7aTFvCWYGUzChrFNr
ovfrFSySb+ELpahGbm31k30Zovr5GgEwid6haDw1mCwZY1eYPRhPYuT/d9094gFWAknTJfx8v56K
XU7dvEbNA5aP692kTHr6vKYaLn5p5T4yZMVbs9xSrzLaglII69mRcrtTfhjm/waHbVgKUlxdXjfG
6YxCpTBb0sGUS01m8x/Cq6O65/5yhzoMF+1jyDbsfcLR5WnbHW/mR7mUKvv4HEe3o3qfLN17NFKp
6UOH8zcutExNes961+Cr6R3Fmfi3C/mzi0fOacWvdNeubk8k3qdYuR2qMkONnkxdD7nIEpVSKEql
wX+vQ32kJMr/XpNcIMmU/8ju1hTICmvUI99vG0SAu2tpAj/E0PXBrbBodomyCQA2mcMlG/ZEFOOg
nAIOmWv7TJ3mP4mpOypECztO2rLpWO1+kiTbOkPmN+WdEoYGN0Zkg5JK0IKIKKCcJWjS1tmb5sS3
J+mwiQVerFDhN309bZz6zOlE1bM7Qwk8Cg0hvH5aGRdDX3vCW0Yp2YIc523BUjYUL1VdnoYeqo5Y
j9tTSVRzIJLQ4iuCrIftdbQsJWJK9UvRWIZ23s/kwfhIrSsdbzqDmjmOK7MjdOxsMRrFBIY4/cGk
91ghPmsha0/fXEXUNDZbSK6gcL0GoKY79ZhmEKgFWiYyUSMtoiFebbhBLnyvit3tWosKYeSuE6Jt
K9YqXtpVcUt5F2zBLeaUWry1SBIvbZZRrwrtB3ouVuUXDuZTBml8e3n/hg5phvxvTaysuX7j9vMG
fWuAomIIYX+9eZ+rcJzQRnAMB0FjStaH9jEKT2utPilg/Qrgfmd0bxtS7d8uCJ4iUFrvXOj665IJ
pWq3nk+AzxShd+kas0i+O44usKqmVmjQVg5tXcoDQtSAE35ytkcOXWMyE+zkbvsfIhU5JUrvB8yl
nbMYnOQtQLExDQEg2xMzKehWfCrm1IluTOzW5suj8Qut5sQiY/j6st3V6RlLlUzQSttIdiubvhtp
HMyjruhQ30tTrr7fLrGZz3CYamkK7EI9l8wvd2lp14uK5utfLeUGGL9pX8n0sPdWcK6QGCbGf4sp
W4FOnMw+VM21s7EObvAdBzLqA++WQ1O2ErC1mcjttQy825PoUrmRGJUI9EaAslEzmCNwBVmqGRc6
pUpRd8I2esN3rIcAIGgTg2ENZj+WGo2yKFw2U/w4+J+vnMxIlHGXRKCKRdXYlpAn02iVxwgeA7It
EEuM5zuLhN7OTrHiNUngts/IYifcTSILfJ6pPDS8ka7HYqEJFgLhM0PiUWllqv7vv0Y5GU3EsEPT
vCgZchp0iMlpGc2o8Vxpmcqyp5/2HbuVKMSHB8/3BWYJ+i4t2urKfIR6jSAZ4wTWQBVlgsDeTarE
UqfdO0QkbRWS8A3TIGHEhah7UjJysfpMZjbEHVvfXxwbYcF40tN+7yAGLOpOhmNuUl/6ogoOFJYG
nJCoUj5doWIfBoSf2ZZMaCc7p4341YE4P4NS1f4Xc+8K+yhibOO0Gsm3S1QJBSLmN+Cha3WkjXvy
iSn+g87bVU9JbGK05hAgucHdE7/4TQtQhHIAlyGuDSzzNUeJN+Wl/QmjXS44AYHjXlcHyiMV45Hw
0LQVa+AKMvGfFvzzQsEBG8h3S0Nox9saz0MxPf1tAAAatzjSTnXRTLZhdSD7pGhuX/6+LDBeh/v7
2WduFZVtL/FHZ9jAmw9dasOOYHPYgB0JpNbj+r3ppcZEz6pQqHzWZqNqPd516xEsdcQBeS/bkaOz
ZvjtUPBCmvJsyglpjiBsNosAS+B+Y5IpgGny3zwEwCJze7ONeA8gG2Y7KMCMvP3MB3K8x1t4QICI
BQr8d6eBSx/wEeUHHZOekYSvzdWsRAo830TiiR0gtnX3nMSd8NsWRqChPFQ61VhODkasIdLgIHgC
XAA+Su1St+HetEatCfbZyurXRAEVX6AtLDTvw6xAdPKc4Uxj7awYrrJCyoXOphitNmZVXfTd1SoE
f0bWEVwWLQftlighqYSr8nx+6trg6hRCPmCMHzzhEsizMQrqy+k0if5tgP1CJVIQgVRfLcYeRUpy
ew0b4bdwP/vhd8W1qQSHhdau4psIM77rP0LYuzIikcu7ZIRvBGO+3jIMUu3hfbEme0GgSqeWtGvX
Sem1o9e99soiS6cmDtYU39pVONh7BMR3GpNYQJ0VtJwJ3utNiybyVPwh1aTwJnm9Jl0gMftllYhj
jBSo+4a/9sGbTkkakV4xH3Hl6SnVB4HmAmEBczr/w4QI6i6IzIbX/fWHkJEIYLJVtPJ00LyRbm1V
yKlYmgeHGhIwuBginHYl9Kh7ZMPHR5N2O9Cpqs9fteVdi89GXeIkHusBSBClrT1GCxETAyRqRzGh
HjuycRMGxpS2NTIPRQXxxvDWVoey6lLp/2YdGAdNfkoi2Z1DiaLLuxki6xS7wAw69xOsNgAVb3cl
Q0P+ZLhU/YLVQcVqL1Pna8M8PApRvwEmQIwuFIUFZCnoNDww1jA5B6eOC+8txdkLW2EDHROoaF0o
QOplirAy1TclSPQKv7incB9R6+M2ScggjXF//4VbkxVZDjWnOyV7LZf9lR7xk5n4X6oMKD6+n1vr
ZoGqmvMUkYLupFkwMYP33laOsjHznSqa2hWPrpzVhsK+sVL66FzQBcnstsXvIPt1u5mBq5AtBaYK
1Bz8rTzeMuyDyFMvs+0ioThb28niQB9wyU7iGQ7CIikGH/d4JgqpiwiLkx6tahb2EBy07I9Zfgug
4l7bRbfNzsSf/OggNLP2lTp8jbwtacv9Qoc/kqTDjArCGMttZECl7IIM1wU14mtx4xUXx3CWHwms
rPWB8p3h/1uUwjm75exhoydkZGTWG73YHu3tUggEIzDTm1vSq5zuxtY5BBXETkbbAqGHpll4I/Mx
/YBB/tqR2BGsxuQINq1c/YDSMnxH/nfJcpr9lJh1ap+7AUjKfeelY8RcogSEkj0Hvcn3CF+vuXgv
ZWibcWkYLZtP6rdt+3qWuLYjnpYgB5iGbe29CjnrLeZjropRdRh6o8oMTLIn9Fuq/Eyr0ml4TWbx
WrUoGXT+zq9MYWBFOo4AAksEArAW6tX63kLgyEom4eOfPFvJSf2WUG2x71SLmj1jnEDZClIzqXHv
crb3R0vj9V/ErmRQKbG3OhEesAVflXO7+iVzW2hTPNb/6+QgKAMlV5IkEkGXzw3/tgyzzRqhZV6W
yqqGnUi0QURXJ9Qh0fDn2XBebKVBFr4nX6Mx5wACeGM/8lrk/Hi9UB3U+mD+Tuxf9trDIidh71Jx
641UhE5GyFZpM+1LbaQSi1UytetW7XNRPW0hwds4b1DbEuxWEWN9dCpmREITxMA4o19a/JFmp/rS
zBbE1UzabtjcBVpLeYIA7XN+wQOAq4sklW+dMeN094+zgxAcZ82ZdvE1hujSnG6cFX2n2gggot5A
zlzY4tpXyTWR1C4akTAbkYcJBVSatEjje7qrN52Jyx2fpMEUing3qZ6h2AiobteSC0reDZWVrc5m
s0qatP0rP9uq3J6ZiZ0SPnc9XfRXR3ZC2DqE3PDN36htWss3yP7bJbULfB/xK5Z5C5+bPxrJHiE5
gYff+lDrgePkxt4NjIgqZ+FJ7HKAlsSkE0UHI/GO9sZmsNQtcDbMC+n9aMUHjCq/W5792QAJdvgr
RqiUNuQdS/FhNB1f48P7sg2ND4Op7Fdx8Cj1tS6zVA+/zf05A6pf6gtqgDpRbyM0bfk33TX1Or1i
kmBSDgLD4Mh5pyMOhHYQmwcX2cRWTzxCq+/YCqX771hI8XJrBpwYcGLCLCZmBQSPRBO6PX5bIHyM
qTTM7zXQzW8Wkgomsx32V//eNXLdAHpbm2k57T7JwEr2BS9JwiP1UO6IHHFlsH/NQ7l0dGTB2OUL
wUWXNn4FVwtxvNgyREjzUN2ItwTwO+D5gSjO4Wj3WbSy6jnoZSSEK0UmgJCI5scidWRdezp0dYwt
+rEbXOw60VlQVkgFWmBDN0VAB6O6xgLPgh57zznoEr3ZvhaFWJTeEC5UyljGhh4XUE6/o5yf548Y
QJ3S/V94AwIUx14c00XrltAAyER9eZW77QuIamtEoy3LFuNhFwq397nX1ry2qSWGqqRlh1l6yfZl
cZLdAwqK0pFDQENLwggHrKQJaO4dLMguCpfQnFntaXyOwrWPROuR7QoQYl90D0jntjuxD694lSRx
uwVvDt2a/sqeG0vop1d2jojXKQdq9Am3pwkRD+67r3oZ0JwDi3gGI02zvaLIz+NJIhxvm07ZEix1
pJ0NY64BaBOh2FmUUFxPS25Q6McGPoG/SVlt1LP+NSu1+D7Yy5plAEDiHfmOwjBUwsz2qcKM2LqS
tbskvs6driTNyzBwS+RMFqIhbYvBxx1CDgGZRkPvH5rqYgl2cTMqIxi2kYO+mJ7RNM75XhvZ+thJ
SYYTsf7mMf9g+ziwZNwKRo3QfLePaPuoSOBderkIBZLRWvhdYli5CT3ta1+9aLFO30tgPQb/vDXQ
nPyWLrFym3RLcjfwAsi3I/muIt610kh+Nj3NlqIlBBIHKGApBXA9qQylpc5XNY3elo8zmafDkLVZ
xkzki8emuBFfUZSahnBzqEo15pEecDwFnXyQYYrTUP9BAaMtm55pckQfKOtK3Y/CWvfJESEOGLAt
P9mriLN9FTAdU3z80jlo3aPGRjCXtFQsnDqRoNHuKuqJRPQN9eGBIHIF6frBLfnje5t3uWrzZfDx
vw4q7dMvissNqiGoZVakKCDjpKNTJ25HRDsmruhO84TqfaH2QLWCh/XJb87PSsiAAenxtkrEMO2l
tV9dtxiCM+wfnPE5ujaBXajevr2p563IUCCkRHNfm3UB1qCnxa4rVe73ARmU3EzFNRnx81uZmLNk
iXIltCE1dRfcSNRqlrc/K/6mLvcpEnhw6BXEa+ttWkaBG37VtEi+67gZv5c7e3SyILqCG6Sf5PWC
GzHITZbU9+xyqqeqbEVBrmXevbMdJpFlLU3FRI4yIP5cgcJKELCK4iRhnCmVh/1IZclkwTW/KtLe
vKC0EvLrw7I/LdPm8bPIOdB6+rk+FHuIsEewwjop6KELJpkuagG1sSa40TnAk+XEek1M7FXcqFvv
oGX9B/+7BpSNAWQDn0RBS95J7QZzKenyy/lJeaw1emDv9aJwNXFDBRgRI8hwJJfOUajEgOHii6QD
WG7pqnu0jF7H33euyr8xlj7izhqKko8n2ttOtIvzLtbCSw8WgkA21ysIbELdLNYksxOSaEWtsRZm
Ao96xkwZBYyyBn1OJhIPstwcft440wc4bmOGe7Xx2DvsSGr+1pCKSlRFerJJFZqz1jddoiEdNP7D
OwphAscTH4IE/V5Wguw/PTImWUgbgQsrexNcOFDjOKVrSXDoDXwuuTKCfuS30W4KvSxDcHinARdo
NqKyePAYhNxDLkvTLdtII8QFcXVxobvi6dKYF1kN+9ddswOaw3/3XoJH+Fv5Z4lw4ZJlpMo4areh
c8+7hNYRYXkX/NdstB368vnsTIO2i3blYnK2KPrPW1P8WgOJBbZ+woi2EtAGa3iVBbA27cu+n7W/
Ypq2Yn9Ti7aaOt4wFsnJxhvG9iJUSerOlJcxjOi1gRN8hMejXEmDSU8AAI8g3fVV0ZoHEYJXynIX
RT/ZJUqpjyS1vjlai2K6lw7iIC+emQAh5DPZDiDjuAv7mh141538yjLtvWQS2tIRHAEUw/34c4xS
kwDzkvlTASwV+ensKe4TC6hIBTkdrLAmv7U3WmT73Xsl0Q5ctQ4MW98fDRwOfhu86JlTojZRPWDE
H66foF9Rwh2VHz8MasqGrg3/0Y8dU+6+OBzB0dJe9TJtwkuDYPRHpLqa/ijq+ACLt8I3BUf5AXCQ
LQaqb32LJfjido7gXqQdkF4fs3DNrtiNSoGaKglF+7siYcbextY90PXFLLOlgKL0Epof+Xs4fUrt
/5z8JhCHxgSdNJc81SlvyG0Z4lW45ukLmYcyHgXzw97b0CGDAlfZYilbRKdSJgRNlAK37EBo6Hsw
rghQA2ZNr04UgFGOpgwK4DEi7rnIqTDEWaFY6BsHI1/hCWiIYC8YBp8VUauVE9bgaYHOkg8ocHsz
/lF0awfA4erTt7lE3EyEDpgrRwI2tZx2QXHZIsr7F+e4sF4lB3hhkOMPGCvE7fAl0fNxKy1wE+tI
ZvkF1w8tag90Bm2gjdVeTzzPx/AHFhC3wiUgqUAFWdqcKcdAWLdG2tmRs1ULaouz43iYq6UXfz4I
vxK4I7wTmztNO8ujbIqMBJkxaN/olbHizvjt3rfHgYrL5vE//fYQ5f0yyjfyv+SOnjM3yKVmFpBE
gu3iV9YOVC1opiRpA4cGthgRbA7bYdbUxXoXV9d8hXLH7JxIcbtiwWsrV/RBFogNdPpKCjGgdC20
hv53k2D5J8KVQRx7ylf4EuTOYJOT8Gf8QW6OUEOWXm/GrMTV/SHdbmjRJPha5c5jjXQPq9Uu0Pq7
/yJoMO3SEg12AFFmL/HZs/I5QSUCXMcjASYe77EEp26+tacZoKZaiT3kpB8MqgT7UPvq1rGCOW4K
dsLPZGn8lpez1J4eSZBlfOEyWkjFhxJpII88/u+LGlx/7yMHtJI11YJ2Pe8pDg3hWWtWNjI6iwVO
pFf8zWZVJtO1Q5ZLBwSycEbhh+wrvS7zgcp04lckDGacnoK4s5U+5RrLXwjD1Am2x3OVYBeCdVOz
LZ8O+1PQXYyhkXz8O5s/C1nnxkMM/9ioC4PxA30WpNM8E2u+I+AVFdkoEsJJjNi9eBdwFWQ+tdsT
oVoRewdFhnaw0Jnrr9DaNERS5zA5tcEoasBAH8Nwme0+XZZYKLlHFdZs/G/xxqb5gtAIMSJBZ8R+
nr+tH9ZlN3pjmIpGKrahb8hvF5dNASvNNlQJKjmTRgR6lXQp2qn6BjL1mxtiOXBa/xlpNn6uRRPa
MMCdPYg2pPKXENexMX+t4mkHDKmzvQSufyyE/vIW07Wj3boj985gxaNlDt+M5lJkFvb9wkUMGfqh
nrtYaulErdqnDmC/BWiPxW90C50TV8TwNhnUJ/+4CAL3KQgwK3ZphhPB9OzsqidDW/tvBl/1gYIN
7BTAiPDMNxeU/lbgBk2V+uclyBt0UG/TQG1aLYNZKNnpbxGsg/sNBKFhhPkqV7MPKQVYfBUFSEhx
1q0eH3oRmS8noBDbe3rw04tmVAGd59e8HOInqghjicrIIHoIlPnwA8D8cfHiULKUzegcU1kHtBO0
Tg3j8aj6c29VrhVPow3AhNiIU9470c6vmfzj97krkRNf+Sy0jDRSKv8JuPcRcQDOmc6ld08VOKDE
IZ72JD8hY1SVTidHGqQHGb1dhk0Ic6k/zhqxo2Trlu/1mfksQO5fiN9Z8Yl7GTnbOSzezhI55z13
nWV6H26NFSYEs9SyKhhJK+7v1bsAJWNRfMq3SnlVoAgbc70G3TuIq4p2zLDu4iqmspbH0ny+bCSS
3FQFdnE10F8tYk7FQLVU8vK6PM6UZVprV7Qty4VOYLvyb9Inv/CKzJ84Hq6/1YSzJMHeXueW8kor
cF+tM9mHIHceq6zcWK32QF5oX7DOdPFstxWKJv7Iaifjh6NtWAqTAY0g21X4Was3+Qy8DZouD+TG
X/KP5yTn7oJbQ7rEYHobLeRJhKXRtjDgOhApabU9ZW54eLEf1idmU9YIWHySzsXEbRSpqWFjvfX3
Z0GMjyY/QtaUP98Vb5SqP5MoBcGB3DZQpad8RKJknoreLfgD0ysfQlIdtsZpY8peAkOhDOFAMzWN
RX6ERv/73XLWP/5Zs19x4/+Uh+18GXg1el9GIEK9O/I8q5AndoAfVZia9Om6HwGoarsig5GS8OZi
gOiLgJoa/qVlqzrnZlFlDF18Re6365lyfLWXmoG/wEXauj1fnqeKIprnGn6mfkEVhR/KEnlEomb5
UV2vfmIpMmbfRYs17RT0TWz8ins++j/WAaEY/w+76LF7Ce3C7PBQMS9xQnArpo1aKh2Ezl8ndqc/
BVzEFTBAt01SQqS+c3Z4SVP2QM6uQEhsAuRegH3NjQ2C/Xyl2AOpQamoFIHB1LdNd0iAs/oYW+gL
hjNcNCgUZrRKzqIz4mig9GfHLJZ9yZgqIuZ6XqedRjeuTJ3/IbAHwHd1W0FunUL6HzDUgblbLu2y
YkGsRo1NkOUG4R1l/hof9rvowe3YfHnPzFZaRA2BpDqZRFjWTIxiWzzHp2nOHy+8yjGB3Hou2eir
N5KMUMyqqBDg0N0tOQT0hyxzbBfLeJrZ5KuzFSxXVKEPNtW6XhIXlRP/Aw+QJW7Kv1jZ+hO9Bj5o
G2bYlXenypcQ1v+TGgbCv1F52P8KZHIIbL95RHNE183ZpZHt0RB+95uKJpPiA6x4B5ywyHHGKvC7
M8QtSNqVZQDlsOY3e9Mjx0YzfIq55RC04TYeQ5KjL3BKglEiIL3ZlMZi+MiASFErY2t8vkOc8Hhu
rUiNtcUG7zbBYwFO9LtSCkHLocBSzFeJD7uI8lbemLn6QZWIf6N2rUrQ016F6tXVt5jfXPbtPeZ8
ChJV8VehBoYFxlPy3OR6JkDmZk/a7wy/+kH1QbpcjyNP7EE3iXOYX9qaNxc/tgeJ+8TuCall1E/M
UKzCvz277AESBHFNX4HGAicmVGBhBut+q2KZj2TB2cbJMJcm+S8M7UOaHKSYH6+ONxf4C7T2anMH
kKUfsPe1wp6tlzEZLOjoHlxwtmrMsBkya7mSJP2VE4QL/sVhlBVvfTCaO73CX/dWr5HbYO4wZNlz
q24vP4NTgqodOXx2vgonPk6sNZhNYSGItpKp4Ik4jHQvvgdHCjU0dbIIEfnukV1jpNmXmDq4rbhT
oWQmCqCmzsdYbNmORhxXtJbeqJgqUvSTA0WYqaC9FgVZeCccC0mlpWQPhEZjPu5xS7cBT0n2lPVk
z65WaROPoi9G9OZesCv9EdNXd0aDGsfsDowwHPUDmI8/naUqAZMkEAUnMq324s79kLaULYGT9N8C
SlHa0oLyhCo00eDXFG9ciizlMHjIcIFDGrr/votTbQJRtz1UfWoZ+HIwK1+GddpUM8sBgyRg9kR1
Icr3OkwehJIoDmfnsX665lScjLQg4Z5P34pHc0IaCcAT/DrzLSEQw5C5mMOUwS0jymWqCyIoRbBY
0wuK/WYvKL8bPWj4fZXdNxL1swV/krAVjQEMD5XhrbGtO0hx7tApdSIl7V1LU6SVwUxk66bEi1WM
Mh0MeWjugZYQcGpFTfl2jbGqeCVyopSr+MaVL6i8YoUSvOIrkAMh/y15s1j1C8GFbmRd9NTzQKhP
dIWBJviBUtGb0WtyIBKaDBDKaNtiIehr1kv7Vjpnz+KFwLaSye1diUDk+6S8Ey2FnU7pfcKJNB7L
H1FGzm9Ts3VdoKNPG74Cgto9g9g9dIUnURjtE5fXGscVDbRmmIceIW0y6ReEzQaAeC7/wxFznVi4
wLMgqKOnx1uf7zS66VjPzxbr88lfn3jHrwKzewjjorL59+p5Xwfz0et9nekeNgt0aOWo2kBxn8qv
Kecgbq8jrR7JbIg78hvAnCZ2AIKh1+LJ0++4+x6h3GR8lwJrG+w9ahWwt6SPtjPjN81ArOf4Qp4i
0i4Ygc2WjGHEO6Qlydff43t9iwH9F9wqXcAs75rJwNVLktJcffIPuQ8Qsb/S3FpW43ficRNRRMsp
r6XE0gsGGlP7Nh8CiXG9xkTWJ3cJeEn/XFRbOPhr0vdPxYjANmGoakH2GnWOMqEO6Uu8KOef+jyz
ihEaGGPOIcJkOSq1rtL856bvFpV+ur162CMt0m49ooKTrq5kNoxP5fjM++2LR0zgbiTOf/s6pSTD
JOMS9fokIryN5FvGOsSOlge02fysu2fMp89Q4qaiDrc9Q8fduxV5JKWVo3/pBRMmlBBMLOUB9r9W
xSXFIHVzeAQdzkeWws+PCQD/jzkLWm56AseWWumeAaC2YWleSNKaRodMUV+F8RnnV3rQGC58xLut
LWJldxUGWLzBRNKYWpmZJWv0yaneTWxeQ4uxX5wCJE8ffHblMvf28ciVoJgQ5ySIMV6XyStpMix1
pwfFJlBlMBsQSilVKQbC9CpKxxlqVt+Ujct1oIEwNrv66MuKVNY89Rs1spFw0S4q5i0XvZv4hjEO
IqWaOlOcTzR68BrkFkXrWitoeQcG87WuGfbatEP/1eOL42uY9HhsMQra+OP0unEV0sAW8OLjHBo6
zeBx0DwhcuVaQqBMwK9vTS4w6hP7A6NRGKfLRVdkBc5zK4Xyu3NytpfuAG+VyxcVVayXjhZIyTed
N6bdvXQf5V9S0k5XlafSrGDGYc4vAJ2CMTrbeEYJBKJLt8lXec1cTt54FXm+kqgUDwSHrfkGMY/m
qRVUCEAuIkss+ZbJ6Loa184wnfhVLclcmgFVC/ocVUlwG9dWBBPZPhx4Y/nUR0q1qhXO2qWhMTpC
3ePuN+n1ldIcqHSkC/iV/QZ8zkaftJyNj9d5sjPbI/XdpO/Gv7HZm0Je9/Dntmky/AJQc0700/5n
Md8PpgkOnvk73PqfdProvtW2t98sn+V/7sQmDkbypXjrDgFq2LfkoqJ0HKErzqeaaIJC0hUu7lLt
RH7LUdPtBoULnFW/1yRgpgJRu70+3I5bA9R8F7Y0yBLkDaoxU5WVbVi6li8bKDCNy2IYNuc69JoN
BKgt+iUCVYToVEt8ARXqYUIIhpoRzl5+8J2rBP4tP39MjCXukOkd7fUGqCFgmKH67X4WFey2QirY
BnZgssIga7UWw3wsa+0rnJBxqj54H7QkcFZHAtBh5Zp8MrEdG6wQF9RDGKfrXulMZGfWMwVMlKQD
BqVypuBqSVUOXEkprlmejvbA1L1XgMSm/ZXRrt9b/FQU0GnNkJOB1GXxsNi9P7Jvup7sxEY41iNv
kEbJsjQzmuZSC9VVOzTOsKRY9isKqQH2EtD2R02BdqDn/kUEM+ocfuyKgaQ1JEmEbQeOWQqqeBbw
dfLO60EnX6e7jSXkF4aCQIGb3iNDLx1sMp+fnGkc/cckgkPuzdb+NVmaaxMcmmHnnCu1n4STyBsI
pK9BdCjuG3mhTTcfOQugCktn23QvJzddGgcbX6SJBn+992iVJV8UN3atDgR+SdDHytVSAGbje23p
UIh1OuLGCM9CJTAFr23+FNaNBl3JbIb9WKFMkLf537sw6RNVg2xsqGx3Q5uQ37wEEgxGi/W0No1M
HLyJHl8BNdx2nzexworWa9aWs0qpxnrip0QK+Ss0BRMeY5kluE7JtdOWsNMU9lSsNnNyATkaFG+y
gNfa7D2AmxHpTsPktVyQaVAcm6+JBgKj7tcQAH96m3ssPPhkGYMaK/dLDGg7wmKsS1h/IBkJIFoR
Zf7A+ar/Q7GPQRM3PKrIVP640CCO8/rxUaTIeuSOsCT9LQeMyONfHI3o5RXec3ld9vIQLZUoDb2r
GObWKcAT0ttuqnM9npwBnI5+WPNt9pnDborXpvh98051OCHuqrRxYDNV2E68SDHA3u49UcSV8Ot/
gucNXrTt4vmiL544KsLBCsGpJQW9m3lQguXGYtEdi8roZbQvP13/Be1Sw77DWWSOYTDLPoN+Vew9
jeUQ4D5qwTIjxnC/wDi/ZBpLGCqPhLlYW3Beqky9snrym1cdoizXu7XtZABdqEe7TWkPdkIoP+Ti
Von+K1igph3Nuw1kbQg6CdPrBNYLBad/MLaQH82dY851m6OJyCUju8quBJ6aPbAVrjwse7GAuTmX
KDs3/iaKuM+ZgDAOH82iyu0dlAQNMU3wxy7pXqBCrsFtAUKimfVuyQwnMRydnZgNiWtK4cTbldmG
SMQFa+7LM0LSYQVbsCPsbN6yYohzlNOikBIv38T1RUAdEJm7byFZbKUYkVbmccxuwffv1Fkq1vM5
IfjbPIfkTYjcNyVovit++AqVJQbQvfZY2TWTwpcntN8LhyeSUCfMM04IJdJWr/wvQNYW5IQNQ+BJ
pIIc4AfVsLTPyKb/e+VUnqmMBojsEGzuFlkSMMnTCkk6MWrxP4Q5Usnz1GLbt3jtum6M1ff/WIJQ
YW1jLFEwlQoobFB3AXUwHGL3IhbZlnu1oryWvpcKX5fDpDz9SSlJT+RBXHwOgcmnukdWzjKNCylM
WXCIjURVaEcg16ff/zTC1BUmZpkdkF53h+oz95KzdZYAZf4cAB7PINvy3l6O7gJMzBTa/0AuMdo3
DfE3iZx1rI/jU/iOv87tjvK49/ybHmqCOEaJa7Z5OEF99ZDWXPOsn3pw+7sEKvI4I4o+K2aT7OLq
MdoBfjnX37/1cB8UBkcsJq9ifbx5cQr8EGAO7t7gNMoKY+GTSxnctWjwIY4mnFQ5WMIYduc9sXqh
OcQHbjeYtJERxLS42J59QPCQy6un/I2bR++FpCobPWhooaDhq7OE0U4JtgmWMErV5iaaDZ6d1VpD
FTxqfAaYq3w2OGsYVEBpHQodI51idZvx5y5dmJzup1nYofHHkXYPMvDgw8IX+qMw4sgfMhUK8M0L
cFLpQYI/tiuO7Zi6cLMRX0vyOWI/5CXTupB3hSs14ySGpqlIJ9F4U6RWz5DCp53cVkUsn6RAC5T8
hnv6c7TerWgKd1eR+cwR+0R5s76r/De3kbR+ER8ojBHRPyMaPXQShnLb7f+E0F8yOUG/Of+p3zpw
5ZwoVbCVTaxD/Sk4AD/YxSqO2ImWH3wxAmrvbh08xqCQj4jv08cqLRKmrz/DPQ0fh9RmUwJ9PcwF
QbH4gbIFOCCR0HAIqNoQDUQXIOjOOPqZbI51frOYpQ1PQQHSfOjh0akuqS5KOtxf+PIqGVtqeqHG
Py6C2Kot0oyWkWVrSAnoeEyPKL8A2qi3G4VVr/NaIp96ySR/5z5NfElBR6pwSLlXtXXf447t0PCa
IXUZQHdHV4NhVlXKTU7rICJ+7LIZHJI7QWVJUCYNMdbYp0E+tegOBVJfADT269u8rTaq2PxpP1ba
K8RcQqQAd162grEl3IBuayRKJ+IFGPobUaZdheRkqAWZWS3P/I6NGkDimb1rKYllx7jgFFumnvp6
SUi3SZn1cgFc/1+ZhFeMF7ngCA1LQOA/WM3h2PlrxGAQ6PbA9kUzYyEXIL+xTFp3dw0T7WBxSlkE
5qtMzl3VfiN6cjdapZ1V6H/EMNXXLzS8n0o3/kxKg2zRxf7CzPaaRj3vDFSPnR3zUkX3ZXYwnMWs
1mw54kxwvxI3Qn0xVVzXbrympkWbJen4hbUhaizjyzb5U7nqFBvJskYqVcil+dnyMnFn+Tiw5TZ5
HTYw/SIhnvGsPFf+TUEIBslYiHnoD9FpdLsu01eW9wF89jMgw5GlayxsnMj0pWYS8hyiKFJBO2i5
oEXJd23U4a8fi9yj4kEd8Fioyq5mVNomYjtwcE/5yhmHvdUYESrBRTi23+jaOsOb95lLE5KXH5Jk
oRJnkbRO7ymcZM5m6U64oB+RNVywUZGlcm2ME3HoZlyiTOn2vCdEQ0rNqoXnFpFlFw+4SN6ggZUI
k7aQ8owQWvKAg9S5rObbe2A29C/TsfuLm1dWEkPrk7ty8WPW0mv9ufc6jaOeOeBRg78+oITpZJ3n
3jQ5pkf3/W2Q8sllO6+JzafErXimWZ5kN4sfddW5PHh62IFcGmBrtABvsct8SFBPCeBNc7oC1OTo
m/MxY3mHta81yntEk2iCayFcJo3Ci2S3wXII7ujKkHjjei5CjmNaunL5d4A8rwYFK0dTfuCgDAbd
9qZnYV/tJNhoyZGgnTl7XEFyyjgSjpfZCLO600cHdNFHbXNCRhDYCMbwnIxEJTMQeGHAZDzpTBgk
SyljRzqs87Lph65O1/mnLjSARa3mI8sInzmp64EE/FNZcFgIF8j7hDZ0ARVTyxI73V5BxkSNy2KD
uIN5j8nEtDWjgyachx4ML7uHJTSAQG/EPNnitKr5umDZoBYbG4ed8FW/rnpHz7dfBGOFWbUmfABJ
bC1NabeXEHhut9HDmpcEKtofSHwn2PwAIvcgh4x2D+F4HZfszTBl0OrQMa+mg+dpbqHUlAtbpij7
Pxmejsd9ZjAVXgV3uDV4ZkmDJ73keJRuMvFcMO8qO9d7J/FifiXYQ+ftDrFise8jsoGiuTypGVpi
OwostAaznsI4jFsuenQ2zHwAtkuj1fvoyOFrlVaTcAnyIrnrxJrf6RTnY+3uWiwsL4q+wMjGBijV
zIxZabTgz46JhQyPHZiwCjOVa3aEN2aNRBekI5DWeFuuyJgZ90hL9YQGvApgZrG5A/+qZTm7fNa+
FFQbbHH+lijNyRRonDB+SkUnAQbCVH9GKH5Foq5WOS6WIViYwF1Wh9SI9GwjmiYfOCdEfzTIJKwj
anaqgzMcrTLPHmaDuvX0Z4ul0MoRm78KE5j9rQT3pu/kUTWSup9o1dD3H6zSDlNpdQLnZLZ+sswa
+aK575fpI+jMgis1e+faxwO3SvjHagxVXfdDr79gakQy6Ldm26JUufu7d5dpHWtYvjtd3Kq3BRgQ
FFbxOFZHPn1swufXFEvozG5F7RXCPkwFzwN4oXEoW21peUiwSwTlKbtyRpwFf1h2KuuGB7tKHfzh
pVMo9xM2ywN49Iwb+hvjP7m3DgIEN0mR1s3KByGElF2Y0NO0p4c9bKds8g7ykZqhzp2dhvJ7F40m
pRJfrcHasp6qWw2V8EDZK4zyNolULdU8ODgFjKpE1ksW0jMK+SOTvxO2tDzNycGSgmzg4PI7Vaml
GE+isvemAyiXSvHFRrOfmI+hQMiRhEgNNn5GX+3/t5tK44YL+Z+NBBKwmGYYFN8u1AbGQuXKq6PU
Tn639uyTcdN7TiH/rO/TWIYdlG6oLaxgPZqep1kP8wCvr0kKxRYzJ8FZdW9T19B8Cn+WVJZG605o
iuKGYLYXdnvg5PEYqQJo4dW7kiC6jpDiO6HXmVK87hcX0wDatS2rdECWCejvTdwXTuOd5mly7kDm
YHUBjGCPT+CLNz8butV7/iV+Ysmm9kzWQU6Kp4THaZlEshmGpA3Engqoi9HgTo7cQD38bFE80Hj+
kJaPKD8fCJOsPsbcvCJR185zQEP45Imw+qBkZbWo2mgwYE8CagGOkftozD/c3+JBWRzeiPk4q4xE
B6RiMnnHumqyYyH9sQsMPL/H3IPcN8VwgidBRP0qKhHuXfHLsVklOnLraaZN3y6Nc1TOtADPc6YA
gFfuMpaRXAsco44esgTLi/N0LPjYI4k6+EiZtWxaDVv8CZ9VK+J2lRzpdxtc0Vgjd8uCFVgglidC
7r3QVuQzfr7KTc3/udJ+VZ6DpGOzBZLwc0/PwElJ02HrdMvXVhIxxMFjwi2wbt9uOwRXp6fyc1+x
tS30E8eNMyUcdpyaG2NkDLZj+RCD97kRkUyCpHGrj9IEZG12Dx1zloeB4dcik6WPwtyRzZxtp2KA
cRywqAGqQj1S7UOvj2IJckrNCQS2+UrWSZFYOrcPxOAn14PIsH24grVr0Q5wrGCYseQxeANmVy4B
aDJ9C9FiAdB492z+rvLXRLHYXX97QUqUP+PCJBFS4fluElzTwOtW/mRsfKTP1Au5TkAcRSZjtPa2
OWoAa5iQ+5ZfEzi0SbgWRrRh4ELi/eC8VtLaCzJnxTvUTWktqbve5MRYS+H6jvgAwRoGLPbjuqGR
cw/YbseX5Mp6AKUKzLldRp1sI/CpCbuNtAHnC/mUrwXlfnqLdWE6UuxsbrusTzZMXzVRg4LH5RDn
Q59VX14eomKgKKOcGBTnI33kgAPeFYiw5ockqBP7/1sBaVfi+wJAw8oSZuqdmQIpl/nnSurlB6Qv
vXUgRT5eyV96uEeWrUidfWCy7VycyxZmZe714HRgvneWkEFN927tYO7Jto7hKe6ZeynOLrHtzajo
Rgr7cxCtRnHCkI8ruzLIsLfy3QMYv0y+SV6YsWe5tQP577v4JQGfi0SoOSCvDP3Eo+B+E4WJZMke
hvKuvEJy3pY1Y7vKa1GhIRBM0jcQkGOp0kjqCbSQvC21MHeUanGWBMXQHSVM9tti4UhgoQ2NH59Y
nWYYue9nhVAkM9bTmed3vip3zZlWEj/d90tpR0Qa24P8NA8c0YGBjqFMZyhtNBqJcsPff6ub/him
HYsp4ZHIT+yaq5mCI9ADBm4FS9F86UWRiP+bXYiLUDnjiawuDj/0dbTbusNkoDfYOJuxLoFGR8Sr
IIAPpnLfrxqdzfAg1DaDhqwOMBJrTiuqJ2sSwmUuYAJsmxioSmIHzaVHN48LmPycH+TgvnvbQM9K
botjanRKvi4IDGir2jGcqu68e9nTLfD/6fxzjELREUAEx9Wrv1OZhcSGSwFdF5pw/xoIi49m1O41
xNsDbKAXeZva7ZHVO4seGoUrp3M9ecw7vlHojO9UOkmARvzJRrPR+6GXbIbzECx8bNw7veMlD4fv
9ok67NVx5oDWxoG7hGG+y5rKBTeKG6P4CaisF2wxhsYaAug2nLWS4DPLZ+9MqXyKbSPm8OkOwPKG
D0xugVVf5W0tTfKW1AyYcB3asxqY4/AFD6UbBgten4ZPHlJoAOelrQayroXo9z39JIRKIdWmJaYM
eqXNI0imOzynhaiFYr1BK6O8Xy3/ChPI3a24byZXwkAl+GwQofI50PUz+spzu5bUXJLj/g2laWQd
FS7qEokYVnRuqrqa0KiFDfGBmFS4NZT+UdI9oE4EC0Pl4JmUSka+LpWrRWo1Ojw8ng0nFu3PeaIA
70jmu8HlSe2cm4KMERNqVXX7fP3KqB9aju/vZvlfyL1r2Pnv8LQideF6jYrJLgE2y4TlOFcMsFPV
dFxps1U/Fxx/wa6pVaAvP1KlaN15nuFlZYRdeWtOKTxBW7LZjgKjUvNEeBsqTZboTO8zDzrls+sK
uLqKDQ+yjV1bZOANtEtNWqTpToEKkoB0nmGNYAym4/yASo8k9j5OuUFZK89iyXBd36MMPaWR42ug
sogl6kDudFKUYfAiJkrVA2m4Y5lrGVjP9rJps6lnavXEvdc6XFucLB2xUKDhkYD6a27+/a2nS9Z3
5M4dJqvugUB19keFJbZ8McRcMPOA79CWMSW0sY7FPKDPI/FizNxm7XtIBa4oqyEangbrB85JZOh8
QBWoZJRg2PzhbUHtky4oetd7qXYHHZ/o1BxsMIG/NhaIF1TquKrTeNo3lw3RSnT39Jc2/69asJs+
2xfRIKtzC++R5L5+9ftMhwwmrawfV6iXRFyLWKIiILcjxWrhjkni8OUhI3ovo5sVYZPO9eMLKx9w
RLnAkAQCS//XLX4pk8lcLmaC/qg9o+uKv85njKzp8n4gV9jjhLawgOfrNNiu5CmAezy6ViLAn/c4
+XgtYwlgYYSxRhYx7c8fwDE3I89fUK3yXb4ZuENRF0OS0PYGCVaVEZCupcVQlNPHt+c7QUL7jfwe
rog4uxAopAUe7eLapR4tGTwGxS0ZTXtnm9h4HtORSNuzUpdZlq13jmL8WHRVGTIoW4Wa3uNxWRZi
hEwRyt8w+PQEu2NnFW9zzl+nhpIpgzrMkPyQjHpLC9nQfv0TnRtFCRPWa5+/1oM5SpMiFdHxv3p/
GvIvt1rDrr8FBsU+c+S2NPE2E/LuzpE40DLPj1RLPSdPCl/eQgeje/vVpscloq0RoF7HwEO/PIrq
XKg3cTr3avtjg08PF2M2T2Cnh2GmcECm23oDy6LyfMoIDI2dPqbQqHya76z468xqgCDrz037hux/
MbcZRUXPE5XDJrq4GRLiA6/le1TOTMUkT1zj+ERbiWpqsenKk4BEmHlMxtANQN9aZU34+f8Nrn5p
xGHor+12pRE9tpEo3vzOtv+RSdz2mg38CGxdazukzEKFnhVkDTd5g0FlC2a6pr/OT8Cym4tYWOMi
N3NrgvTzcHf4VUDg4amtpqEm2vlUaSXJ4633PCBp34d4qLgkDTlcRVeJOEKcF+BFwTeT5CZ7FE9j
ixK4FyMqnLBBNvK8pPsTOtcZ9HCGMAynvdoTuGyOxC4O+TCW3eqRxXpSBqOHRvfj4oa3XU8p5xGo
kvmKaSalxfqZ/zCNpSNjlugtPOXegtyBv/5gOzh0jpO3pYODFE4gtAKYGG8TfnPLGdzAJkc7NuFF
mjHqoK7wZbVRNy/j/Ya2lTSrTm6d+p7J3sTgG45f+Ftx9XXHch8dLr5f556bcQ+LmYkWG318z44b
pT/L57q2g127icNjECLQyR3iNpOBGtHKS2f97srvKzYNVBzto1uFKNkwM/NLGyeTn6g6T2wYpVko
nNkhtASmA8JRyKqcpmqjaU6N31zyhuYybyOBu8RSaWgVYf1CtZmfox3cNXa6dP+QmgOIadjmf2KX
L0QycIWrbGljqq8LUlm0gFDJoJSOFP4TZl7mVnRhbXWM7kfnSkexvkxS10EwZO3PRSjvFs+CkKc1
bg3tI/YbMryUTVtjoXioXs93+dlsDasG10UNo87WbUi+l3f0imr/0W8P1VeRxDiavleGJO2bHkNO
RIYT/6+f2MmRPbKwPL29xAzRhuDEB1qM+Moz4Avv8nXzPpUocPT/puLhtimSE4RYffS57TYiMRnb
6qKbstH72/KNTOSykFc4l5MZtty/3raD+nD5hw+mt/FQcTr3nFJztIafnDWUYd+WU9kISAeHiZEs
/XYIAqu2cRvn9iXzWMflhsyo2YwRccNeYCg1bFlxb0jqBFW+ADqUn4EeodLtEEscqckf7pV/wZg0
93bAPa7Fk3a2JUs66/OI9bniLp6dA3lvpJ0RYVRLfThwjt+FDX9zW1/wRsYo7+FO2atjWCSJyrd4
laByv31uRcCD7SyhrOFxapwyGi5CWJKObCD9Qcz01+Z2WYgUqHhj1uq5tbGoVaJhz/xpmlzq3eHG
9ddKORahjQtc6AxHAuakPVd1EutTSEm7ezx9NWTfD0Tm++g/LktH3ot2OaQqf96lcC0uY1X1dsI+
HrGpbgvi4v8+qH4svrXS4TCWkKYmvvMMbzKhxoL6YjmUWoAYTDC8SJf09+Z/nKmnYzEloxdqF16c
3C7AqAtiJRL07+/vI2vW0QRg5o2i1Z2hYt6lgmoTeNws/gb6VO3v4v7Zm+WPQQ5qlZ5qBllwLbQ2
anXEzyOTKbAbDzF9vnkUr0CveIjP2wQUoi4wAiUrOGIsXd+b5QZCH2ww/JozAYYRiDuekSLuSs8p
LZabh8xYLZUexarAkWkAtA5Gjgg5yeOzoJvLrYwLKDCp7mquIcNI5X2RWdroEHuezMsVmB9oxySJ
qM94MgpkN0JsY9j1IulWob0qsmdSMZxrQAxGtQqJ3zfO5zFdKinYVshIviVMt41YPMx0TUN4aQ6E
koFZqZiOqWL1uIs5Zjzmu8Eds2G1GdFYh54iMaq4bq/zEZroVd/IlQqPgtR6nugYsJPNJSz7u/kH
H9dp6fIga2Z4C48WA98rwJaWqchw7XTFcMp0QFox+fqti73DHlqOpZyJNG5v+49W8N0kfNWdVq4Q
BuO989Nmu0tDNyiRkZSn9jhldYmHMqkzgYReQocDC38VfYz+d50JPhWUHgpP0j5+l2krUfD6zxAT
a79n53AnZLGX1UGPrStROoBA17lzP43+XmLOYEww9ZjuHsgtY7sCrcft9vgRt7I+9HXhT+W59eF7
qGkDibDzPI3/gYmXY7qi2Je2gOyacNlkbxddGQVv3U33/UbN5/AkUlR3Fw5R+VwQI0Br5c8jZ1Z2
a0tQWOy+LvL3VJSzJl5D7P57HQTfkbKQHtgBadToYt3QS18JYgaN9e/udbF0QVmZm40LLIA2UGnZ
40u/k9JFYwMEX2obBqEfHhNCuSuh7rh48y+FuiRRUMQK2gX2Obv5r3SsXQnKS1AummwQVeLMp4Nn
YH8y3t2HRfAv8VSL67eOPm89a1tP2DTAHH5ZaciHbnfOuOPjjEKEmqFJrkIYPUxu6a8hO5BNs3EU
aeGxh4fxVDDvGz5+XYFO+sf2extQJgtJrahpizRSg+RSNOExvrQvp+po8KXYXlJnyEiXqEyWcQ4e
RpLrQh0kFcYOVlEoQ4RK5nkUwLC5oVI66t2e6EVOwZs5mgagyPMMqJUxgwh2nJudbVoO+GsqXwd+
G1tvzdOb0d8QGIN8CSP8cPUCiV5bhQeTPPbHivIpiqraFLDaN48C4FIjESOHR7GjqH7Qf+mBhcZf
2XPoPI6xvHguDq1EIY7qYoR3EoynF+UPiP5rjXoCIqQPmhUJtX+JU9soZ9mSwxuiStMTTvLBDYqy
QnnR3I2ILElhJqo1eDiRyrNDfeRVGkkbeSx3Gfp0zzdLoCkSkwP/zJe22zk4wwm2TIG11X4vWkCF
0stQRFWed/X+OVrfiI8ue8zpBmx4O77vDBKICdXn8O00NssHWH48a8GmlfZajrFZaBBGIyx/J2M0
esXjQvTrv54bKc2HLBQG8SNhVCH1aw/7T1MCHDJq4G/B3UPuy/6JNpHkMqCHWO2lOcpivs8ZeVr6
Yy9fxb4CxB+mgZxD5fvmNOsE5XPHq6sS+Q7C3ePm9AGTLkK4uTMToxzSnGJEBhF+YaP8tGg/Bp3L
AYC+xJ54CTBlesgEcUvmZj/UgiGT39LKIopVS8NbiKraGdhfUQNi6gTK8K64HMEl27/tirTriJD1
A9V1JHSnS0kRnDkfw8PbNSyFyPEm4RUZZpmFrO2wz7NXvnIMK5pA7R+7uPikrrsGxnlqqEHw4Fij
p8P+CDAHIKSheAUVguXGZc4o4gKOxnrtUzPb4kRoKdJ0adMauLdIKLUlJk1lIM25ccc7rRY8tvN9
Zwi7BCQYQBOTZgt85RkKukfsITFkD20BOI6Z+6zV/cJEz/Uyr67wyTC61x480AAIV2mREtZ3MfqG
4TRBFDoJx5uMtz9TXhc1zTl1YlQwFPLvJGaS4fMuHYYBXeXk+7TxWVnN1nQkShNgIILZ4+Hm1uVI
Rt+++FkZkSUCghXnTdipDxbWo79Xstl4wLSQBOS3LlnCF6lAiVuRjJQiLXmNoMqXSRS6vu3BSto/
2hjv6hwjVmrrXgCwJ9kevy1h2GNypgQ4IuS2JXHWlg+b8jzkWJwwy41vR8gAMFdo1ytnU/UKAG4f
FcbTPuQEyCQlnz0TOH1p3VUlGEvA9FsTBbDH2otlZc33VNizo+zHrTfS632Q31ro5GIpbf9GBpgN
zoPYcxW1HR0EyX9GkzqE5XjCekej46c7vP5MZ4Ub1D2DdyiCmqJzRuMKmxdAKxMlHsF40lnxfNHE
koJ7z8WRdDijrqRdijDQOGL3EbfIqz4AAsZYATMrAkmS5fP2EMRmpGfAuoYHx6XLt83CdHFxzvar
Xm/vRmcx78wSasui0B/NG7DtLe1S+CVCZ2X49inVbBMaVyT3d/webm3YkAuMc6BqzNv+AlSN/zQg
EXcf+IjCr81rS7fK4sihriNcCV2J3VP1PZ3kmx8w4xJ8PaRuIi0P3N+qTxPwfg7Y2l94y0Qg3kky
mo/fHL7H64UJ7xOkcaff9Wdsn7mTUGXg5IeFtNZr8DCE3M1VNk91LsVAKTykeKcKc3TniGsXbPaI
j86QjbPP6nPtZbNhMx2SWtDW+gaWbu+fdvD7HeqOLJ2g3ZIHtOBY32CozU8e/Rh2tEUGNCZlgOQt
wBiHKK8HCfuhY9iJhw4OGbQGU3/sGHLmW83kJ9jw7zrQ7oE0qyCWFBRVS+3LM9492xQBETh4TCuR
KTfUEP3rZM2jYwR25vdwKYD/wVxw28WjhgVODEe6sGP82xIFQWRnlzivSa+DRwNnQjJie1YCHZr4
tbJa7IpRWuB4k/RTLHKApPNktFsBCcR4/LssinYMkj3o1Q0qbIBLdixLybdSvRCW6nn3fZTK9MJC
RJ4IaJMJfZpJM0C/kCSppL/D8oTOONS9AavlPo93kBw2/8+awd3LqgwjufhDMcPtR5mkllmf3VdQ
zbqncUY4/GQtCxUWMY2jryzhdK5isC2VWeAt/n2NX1CV4xW70H+H5xI2W9mwR5aC8HUw5guD1p0L
AragK/cCGuEnEZSzy4xO0fibhW0ZVTpedF+1/waDC2sLHuc+qWWKY6U4CBZ4m3gZx6YNMo5i7ss0
V+ZNNk+5GI6zPeKg8yzmNdK7FTPjb4+dDgkq+xhm/8RiUQpzgtMs0JSc1o/eh5UFAHjDGpDh0PZ9
9zjbccEoMtfGg9Um4bsrysVPZ6Yv9+lxELEP2ebcZZ7VZybEAzgSDd9H2J2Du6nvY26aJT8xzptg
+4v0nHZUCv5c8NP83UIy1/z2CwZbPnstJR2tkvh5HzerMnjh6mRZonx5y5Ej6Gq9sk3ofY+i1qgT
adgtJwzHuUw5FITi6fKc+GoCPsGt6iuRBrDFVSEVwAwCj4kQhzneMHDXygC6oOHxYGdvH+voZQCr
Rj5qvYVmXURCuvR92c/hOprBFtiz/Bvc0+aj+8hbY0HTmb+1tnIcwAXtdbnHm2wXlTKrvGojjrvb
nuUWwsoYJfT5l8zJjqF/iCriPSDnHlNRMJpxTnOUWcxKNzrHBINb4pIf9CLaAErq7vlVXaH0AZlA
wRrJU7rgc1iTTzsW6ICHxlgm0VLdnqk2TSy6BxIXd3RLgH/sdKUF1TA6gLFpFlia2JFdNOpPNm1G
wQ4FRagsS+b+v+vO1EB2qOgS3qtKWxGYq8zCV1kX9+pS4Ai7uTPwgIAf2b9kSW6umPac5+uhZ5CC
/SiVt1hg3zb24xL4tKyNqnf/lPkNmLKlb1Cad7yiBJ/OMyXmeEQQpqYgHWyYpErN2SI0QFYQJo6k
lZ2nwDyvMt6xRVEBmevqebHbi4zJRf230Ul5CjQgD0L4sRxOnVSDvq6M37DmzqoVmyk8cHSpYWXR
CJ6LLNbCGTitFGxuawO9VCNCjGjyaeFF6E4jaPb0W7rvhvkwMjIW7aSK9HKxq90Ck0WS4e4X9oOv
xbwSH9dZOYKXrDxQ/0QG7nUjEUfVhqp/z9JwYy5GNHTCoSK9DomVvJCd+MlugQCEKcs/F61yJD3g
l0JlioL+vyEBjANHYYxsy/klb4PNT8tp1G58R0y1yKzmW6Su4WyIGL0D5Lne8CZay1Rw+L6ljFqg
Puk2MvNpUCGE79CEak8ELv7Y43FjXM8O3RJAizmVmv2mJizS8dCTIPV9k2ULqZXREwqC9HBCt9Yr
zZxr74INIAANf185Z1p8o/pR4Pc+eqlqyxkLALEEsvIyGAuDw6du9urZzmUZle3t8X0qSaFvZEgR
HCUBxo3j/11PR/2mWtTWz0jvY3PDm2+BEew10ekf/BTpJsQeX5mJkvbfVzyC55EW968j8CATsMYm
LRrATk0iISy8HiJLWV8YRicuHQaxGjH+aWYptblngxwFOistg9Lb3cWQLnj/rSmK/tXu8k5RGWRc
nUrjczrqwT1C2p21U9mQEb8FnPk1MaKAqhHZZsSY66xvJzoxe4qXKaus+76IFFlKTuBXQZAFCz6y
HCuCpj94jPk05MDDXbJ5kUHixtWtt4nl2HLh6OQMKg6ZUVIysnUWvpTLLsn/CXcK2ACiY1frRz6h
GKct1i015ZcEFmUQK/vpRragJ227soL46LmjFrItbWYSs3EEYjwKwPeIeNwIQfWfdEGU3SuGGU6/
DaKovWdyY3AO9toXNvaLQeJZ1cZ9eXImLbw9F3AzEf+/1ENueJZUtjfPVmWSxNl0Mfmag7U4NKAZ
z3lLWg7gOYkj5MJGsGeOGoSDFye+t2VY8JiCV+i8AgOonQyzvlKqpjEOKbTj4I9dP0kgoERRZmHg
7ndwcnZDcUoFIj/NUJ+GH2fjH9sZiarN4qF/RZi7Xs2musLZsPqbBnBlpkUA0h+7UG80Du/q9NfB
ztkSnB5EGTkASCTBUgx2VHpO/x8gDHqHBz1XAngunu2mjrzajPo/YC5CdSSi/SRmylqJy568Lz6A
kSZ5MTuk2pGjwnJtu7kjxS4L5el3x6Kb/iwBCcsAcZ/l7xTatZWz4Lv4wGQjchA/XxbYfqQJah/q
MfA8JpWIQ9ulDhxSBuCd64+/Qpf+dfkKHh4kNylQJqtsp6MC0da5ah3/D4uSqA20J7HXZ8jX6bqh
NadHD0MDjbFsbTPq7DQAWpUZ64AbnzvTmFq75l8KXs04cibiYyVAumubw0O7FmuV62uDsDtln/uF
qNE/k/XmvX2Qhkp0+5e+79PEIgZ9RY7ocyAq0UPQyZ3sLOD9SeTAR4p/og0Penv7jTNr0nlf1FYM
jojaFFJBqLZqdmxFiYVoi3pfKxp6NDVU1DwvUA2FPs20qib8vu9EfpVPk85X3JoLhecvnS7Zf55T
QWijaTQ4UGeN7PzJm9V+Zf5HxsvUoZqAeQznd71jMxchBZ9yGTBIpndwkDABgDewPwLYlPRxsHrn
8LdEOECZlBMy22pjfQ0LYJjnf63xzQNPyncVqar6TWwetgjvdjNAhv4fVqHG1k9I64Wo+WYoX6aK
aXvs4ZlSq+MSa/x6p2n3ynUXbsjxyIdI9WrHgTBR9sqO9DS7G18YrNm1Y8oh6tILidtQIVv49j5G
7MFwXqychqIaJpIUMa0KkpF/LeFVgKAP3irRWWC8SsyIj3V/m22Gy4n0PBapaDG6mCG6f1QdRS31
K+WGWgjUObTzHLhQHMHJ7w7qXzBLvKz2PU4f6qc2u4aZ3hOikDDKW4DVVj7/a6Wj0klj5+myyDSX
dFrH0pdpEhP9A7/sE8eGMmZmrvz/5y9HpqQHxGrOVSLWbOebwCCsmp/aEQGiTvaCcKN/NCzRCFQK
MaTj5vbMIVrTW4wCO9coh0F2vRRH/mdIFk67PV9NwnD+l11rPhEMlRacgs8U+6V3u2/AWGl9Hveg
3TxZBtbR4HKqAlHXZ0hME2imW4xDKqPsulN5zWjJhLuuoDw/f/sjT6l6GiIQ096Frorztek8bA8j
yUafaKx2XvZhKhj6afpv0lnd7CF/+Bx3UiRRkdl9LN5AtL+ps8LaZSiWn6lZSpVmLUlPnDonbrtu
8HFLCHVx5mLOZEq7qXuTdqtssUArfAVDQqhz6k6MiE67X1+Pj2Ctktf2FuQdq2Iyz+cq7/t4dyxA
07uqEWqXRTJxlObPBd22tYWJJDfig5LEHjUf7pRYe3V/erlzCi8oWwVU7vSPt/3fykxFIMeftiF6
5kKYLouoehuZ+w2v5Sc3u68Uo/XbI6d6N/uxNN+p8vad7OI+3cIcmpNrFE1SyLZwq60+/UcgT0HU
abvJ8vyNOQdXW8hhbTKg+DOtEZB5c4lz3flHbfXg0zeTeE9BOclW5uSYkPQ6uk754ZPuUcwKOCNX
/ZoHG8c+zmwgS9o4rHR+6unfonmdtq8quFhQc0iYZz7RVSjzEPpm9TVNzAoGNPllDtKvf+GLqJJ3
wuarc3LRIf9EUum2svKax1TxbebPD4+2ZnrwDORk9Z3w1H5/Ngwg+m6SCn2vB6lOYEH8tRqnDBOe
pno9RAqSOa6WTyfoRUA5nZctXTlxlYL+r2oTvdUqw0Crdw4oDtUX9MqO68JBn/iv+31hFeKt5Izc
bd5PFQzCeotYkqOJgcgRNnDAYduears4IFnIazGxls31vefs4TMuIWCL2MIirHknrRsomDOsBInF
y9opUSP5wv0rjr+kKXIVvmHGWwg3qQkADLKaTxoYUlYlVJi0Tyq2+QnWvKZff1ANelyKtqbjXh2v
ui0gViGODcVn1qxB52WRUYxF3+ABRDHOShK8W9II+0qhKgLV6LsnelqpFtf+0ZvYh1BLsJ8ERD8e
yyICvBzYSvpLOEHjbm84VKJrMGIfE4rGBgt0uWiIlgmAHoCAXWK7QxGw4rX40IUPB1fFcP7TzotW
obd9O3oT7KWrWbzV/K0FKtJ/cdserPZkmAuCliI2/I21I17s3TqzJXCcyFvU3SGaOzgYFeLNzq+G
fjoR0jcNmM3Rpku87j/FNx4QIcUSJl5ThFQ+JK2bfpYpBLK2NaDlO4oykn6xkbioT4eMlixc2uLN
yzlCrh+83TBXI6/w6UntG/c4AzJSOEVig8uDXtamUoQbxTxvm8VZyNbo0WiffFdqoZaimp1S0xSA
+Kh51cLGnYEn362YO032oqao//XSkU8/IhN+z4Z1l6VsjRjduLLM2fIEIS3cq1oqgW7C6q4UeP7T
7w652bY4Uzed2KINwq0ZItN6m13QryhgHPT+Qje1etG/U6S+21ZYi5CViP4NS8P5fkgCtCQBn4Mu
TJXYh+ZItKg+ptoO/Rr2a7XZhYptar26bNxQVVR5WdqFxi1B/UG6WJ2w5BkKQh35+CKzgM2VfBo3
6PDXiVD1zKWFfmmy0wpcXDMV6fxMEJo5bdT2N0isaBxEIsLknlXRpgs2q8WZI6PxN3FkKDRPyS4t
Z+lq1pTuk/rwWlujjRqCCddiBRL9iDR2UmC8XHYauXZ9fY3/KmqsT4egcVVPPxasCtN6QQeaNb99
tnaL5ydFxwFo8FQF6bQb/AoXujHqL5D8jwq2BmwrdXfzdZNPNo0m1LyMO0AeXAOM346olrdcOaxm
zvf1rTSwmcem0kUSre5e/e5rrEzlzRbLKdpRjAdpzFzwKYTUqRmHpCqlCPcC5ZPugyz74DeV4UVv
lzjXzkaCfgYbg73WeMQBPzw8nRII19u67nuVTrBPziWY3+l/Rau4Y8D8leLn1UzOdHEO6G88gtGz
0xmqsqSl02jWleD6m+SD0qrrBb1fRp4nep4UZssYjVZEYowiDQ/FaDiQIodwySY2iyR63n2EF3C1
qkKNsdbQQqnICuN4KheeJ85jzDHY+vGIbD9vCOm5Atg3t7QU6IvhaqGzc2R99kw15XvB2DjujTWH
qISz50RGNrokvJ67OMgWW8bH3Pe8wUAbgkK4WXz0BF/zPXg/IAFXZxNN09TxALwuNX52pPqxCep0
9asSMSfg0O03syG+j2Trmw2HtJQcopIP4CGERa/Zrv7lK62fbOqWNKju21ZkIHtCQfKiNMOnphsv
AdYsaKQhLYPECgHCLY+E9f03tXG3KyHEYm1WLnGDQYKjrivazcM8WlEcO+t9BR4GTz5HULsX1bVG
l3FHcGtcOMQZHD+2+LE2Zgxv3mbn995D776aLh8V/V6A6+JFaX3YWk6XvWqN7WFcH8peRgOJRHOW
dPqS/TfH3scnLboQzqos+QgALrmMNKpSRYBHu26SOAUj9y1YLe4YvHAvoGLemcKFSF6xZiMgHHCh
DPed82xf00iAoDuvsSU125fvfc/pmzRMFNLZA4gaD6Z22Cl9cUi7lzsQ98+OvZTjP08ArGAOgk39
HZgXkW8yaFjWU9ky0GnpTuIue9YfYuXDIaTBYnpKKgFnHD6/WASG4e2eZEoGlT+kvfamsRCLDhaS
vWGhMXXu/1F5V7H5r4QxqkUih34zSnzVnzCVWQLD27ZctvtULTjACxEiDkWGQVqy9L+D6AzJzWc6
wCKXhjPNqGmz5X0v3C5459sWsGwJWENKWH1ZqZCsw+lR7XdQAr9ab7rj/0S9qwCli3NVWDDUiXHE
6mWrtNmN8KPqfhJGjdVRsNy351toWxBVM7h497FDOYhzxV7dmBW1yuEmaW9lbglO7CEqkj1I7G8D
jIO6wb2T0rFSdcgolUT8zNJomSoQ4vKlDY73x/Lx9APBv78IvkgYikpnE5NvPiXL7BzNmozWCnBR
5fnQBxgVRsFr4d4Uq0hrF9acRDfiOZRSq5f1bcrRdmEHvCZ/bcRxzTt5aFAkxnpD0Ii282+/eYu6
hyEeGhWJ1s301hLBN+I4czLYtZm7J7colMY8sFKxCEYl3yAdabasdBcXmfBvp2kn8APVVkPcMCGZ
rBLgyfCUgcY+YfT4Y+o4fVZuvJWgJeB7QmZ8SvlCHYODNlHMiag1GrconhOp9PIueVGBLnOBQzfc
0llbVFXoEa5RMBhiSIhRhwCJk42p3/5CL8w+3hHHwTF7E/Fh7gkdOSnxhjfoXuKyUq/ndLtQWzSF
IsLyxD4UUrUFRISDkdn/ijsZQGv+LuqHIeyfQrIuBDibZR0i7KSSgkHmIQVVf1g+UYIlmIDb/Rrh
vlOSJT7X7rZnOu5haT0p0d5HgPxXu9RLZH9IwHXPuMrASzaX96JmAMXg+alYTU7IS4sqzqjTfRWr
qOrziDEcIDoaJu54Finnr37r02vfYJd5eR9iru9UImRdLW388qenn0LQUhlkdqdrgv2Scq0QgYzN
AuVmvSfhA5vxFa1UZ8pQg1HGxqlnuahieBHBf2NoWXD6I0NgRAmbdss2271T5VsmVfLHuVjQSG1I
Tv6Bwf/+O4fwJkAnQOEGyyrGIizOuEXeZdaYky9nTXWv9pE+HDEsLSuGxyhsr9og3KYbaMGw+oR6
d0iM+UlsTGPY3IILvjfYhk8Zi+YD5DMFoHiMH8ZmefI8V/9MClUBQuoyXOR3I/du5hQ9LoGFCQbJ
IGBlpTc+to06Yr9JnCMp1bxge+OrWT5Lvu0lCe4NSidDNAR6JVLSHSsFbEzBf3cphhdRnHHZNSLG
RbR/g9dGDjMZkCTIPu4qGeEXBgwYqKb151PHqFMTMKsf50rYm3xvZ7F8ilMA5mSgQTei9iEUazMZ
0sOESdMbnL8WGRwrRZz9X6gdXLv0GnEpouocIxcDrs2k7h7YvX7bTt4dhNKtpFvdl7T6oyE+0V2F
8i8HEgnQSDEMzscQdn3+IxOUZslth76C8h6X2NlO3IhdRCc7HhfG2udXvsWfzvhpvlT77MSIhbuD
06VV2mpb2RjXMey8s4H1QOVvTNn5oF6CchN/vMBo3U4mc8wosm5X9bHYV6yoVGlLr909J5RG+6LB
2dUSUCE2D6WOKvgpw8sQar0Zl/k8ADrSRI/6YI7HXA35egP9oKL256kAFDTX3StGxKDlGNG7/rEg
PsUrOn35qkNQKA3vqNooiUzxQ4nZ4ZhHrm9xoMTSAgdKsAh0aRGLlmisfJ1GFilPeUdS1kD+WkSv
Rg6Z8Z3KHvfgpWzyCmJefS0l0LagTA7nPNkpIWwo49/XERnTRvsJK9rRGhODtYh1/ZjAg44NOEeg
hHtkLGbLcydYMzaETVXfvm2QOOzLMqQQxF5R70aCKzzVFlaDa1HlFGo+VS0imRhGsk+mO/ExO3z0
OcAIeZytzpWPcIuKjgMN0O/ZRBKs0YV6S2QO5A3UvB8dGT75gPgV8Gc8QEbagc41WmyD4/Wm3VVe
ICn8hlGCrhkUwwB7UqQ/fHMxqf2W8ePPMtK0QC7RP5vXjUpmjYn+h9T0krGCiTy32g7GB8ztZSij
HEmPRx9CYhzGpSrdsAjSFHnmjK4CMqb0P7M6+chpdK79hPHqHxuataHMaTInePuVEmXkkv4hPX7g
LZ4PPDo+8OsjTTk0HeoKNl+FBVkMWJPxIHn93r7KwPBj12+koR6huvDvkrOAEWPHoUUdLgZ0PF+O
pVhe6bMCQ/GWsFTCL9Imp4iZvYO9sGlZyVLzR6e88e481xR0Nc5XJH5R59SvicDkpY8cIi9FK5XP
LGUfE5Ifz/xx4otQthaUj/JvyiaDBm2kshABKVVJrJb4//GBH4BjNkqF7sk/8outyRd9l/+JG6I8
ka+UxsqAhyeziK5OR0pVC8eHoGzX3k8H3sWFo+8iovz/5fUemZKScTzbz2scguFdUMzt3l7orv/b
W7D5h/z2Y7fMq7Gl35xZWCmZOyp5QPdEhf5NcPpwvp+1fotDm3ifCk3Oun3n30IbCAxVNIibBhfo
j6iiJ20Qy9cpooClXecm5hBDPYfOSlGBsv+3ATK2ALzUlvaUhEJO/IED70odC2nsfqiBbXJiot4M
2LJzXuUdMw2/Oziqx3XbMb95bWDGquu5H4CMAaH0LONbzXzda4TSsqc09Ano82BQB3q6bgfH0NDO
Xuw4mLp/xRTVZpI+M8PRC8x+0S0WkagAcQmWQSSdk1yXbWaoImuwT+QRr6kTndgbAr7RjCnuAyvb
f6adyggYHr7A3NAsWh24wtw2AMWWVMCsxKLC4sBF6vQkfp2JPmSePv+UgMUKWWLlJckuJ6v3zEAK
TojJuV1G9iDhRDdk4b9qyAOzg0Qy6G496ZvaFLdW4F+7FenyqqZcULhONH3BhW4bmJYhXXit091G
BLg2SP1yMfWa9DyGVJsLxh+hQdu8r5yoNd98z7w9kQpXD0uK+GWtE3PJpxpjo41AqAPdZHFEHElS
fT3dVzWLxv9/6g754sMGZ8pgZZbKRTImpnFvwg+7q8nGaaJ5ud9X65JMemgJozRGiubCHbrTumH8
ry+d4fq7fuBhHigo8KD6Kz++1zi+rM3NGUrR3mQFxwXj0xpqz5reZagCsACrt3e5XeVH/lTKsGRp
1ywyftv4vJWVRtCtnXWzQoWYXwkkJQf5SrgZDqOAJE98yS57QKFYKaDWgBLFLqxNFhCR/AeD5nhb
vSgsh4qsl+xYscMKSY6B42q3BLeeomzziTxYNfkPXNtZ5DRC73dU7tDdcyM7wSiEC7qd/y0g7xtR
5t7mv+AGR/MbmqN20LdVO3VNkNAhGG9DUlVC0S9bWbr3bt1ZRAxwqu43TL/1OvvzsLFg8et6GJAR
GVdBZDznda+Ft5PGHacjhQtiX262xBbHAy04Ryl2FIA5PJglEolKkFiM9oycy6WV/YHILW4NORdO
yprHpcY0aMHsNGXL0eCot8IUSQAmpwsW5nnZxCGDggzW+pEmmK7onz4qk5SNfEk99PqVDgfM2Ec2
/UeOI04rZIL0ikS6M1HiciABD59+oD5wgDppv+MbqL41uUruf9+DW/CgYgrPhcwJZH3JM+VlCUex
HwvY3XnnW+UaL4QiGOXsvVkNSYUTTX384F010y5D7eQHOfmwd/+YfqCZjCyJhpEMEKTmEdEdJHXw
NlOc5p6EWhtK92YJ9/F5oRTBXxGyuY2HBHDPSuCsR67Nn4U43a2s0oyn7EJqfeDbgoTWD/FmS/0c
Z7TkhNll9ddNNg356PMjv5nMzZDdtT5/YSRijaT3jB3shAmUPSHj7RdV629qCc2yq7J0BVLsmS+V
8Jl5TcUVEROxBFb5m6kdBSQRvCBezMgXUCn3WJNb1OVZReEkapXZwaR+HJ9hSbJtpw3yvrvfXjK5
pep/wcjSeZvZoV6lS82EqyWeelEQAMBecFyLgceuYUYCEzvdDdExVJeojk8d8+xQ8AymV0AHKKpz
FqNqt9YX4amKupLPyXGKKdOy5JQMy+jHVPIRQS9v7kb4Cl3ahCmyFzQFVyt8fIg1fDUAiK1OCzJr
GQzkgp3/Rz2MjEuE71EyplsKlaJZc+Hfxdqg/jrpxNXghYXsb/TGFYHFQoWPUjORrT1CEdb9KZJ2
VJ5jqMbnLztz3/rXuz1C+mjWvzgyfOhzG4TT29kD7sTL67mQICZ+Bf4B6VilvfFYZI4UShXkUbun
jDUK9zKgsHxVSqdiGr50KWsgzot6uOH+Q2bp4ddueO07GbVAGzVSvCYSst+58KxiDvFDpOqImmhX
VCuvoONg4nhsDOHdOlNPN2klTf7EM6w+iAUtaD3rUWUAfZDNMf+F4fRobwiwABdAJERKQ/0Oa+UI
73KHopbDFkxHCjd4Dr4iaiv69cEEuHMKVJfjGRhI1qSzbSFzNwEma5ziuZqk9+MJ7Mo+VrxAFsB7
7Kta8Eyh8ZEpvg1qst8M7ikG7spIKWT6hQXgIKX1GIsuMKR2BbYYtVdCdUIAPMlrbaWZBgiEm/0q
q5Do4QGKDaifhmO30PiTiI78Pm49KTwTQLttW32/rHIbaRP9iD4W2pUwr3KzS0r47M0LA4+Cb24h
JwWYqBdwOShDjLscfnp4ImC8MP03wAczHodcT6VxzuV9xkxoMnCSwHaArxa4g2HZP5ZBb3VdMHmI
pP0oX0SXwBGvihK2sTUmcwcKTgLeIziwbbspImaUYKyTmb8M+iFTY2YuqRpOgkcUIk2pnvGYdcIJ
SH9YuQ1TMoSgsRqc41o31u2YcvOPPu9k1Ma2rjerLuX3yFZIaEEsmuJHE0+ez77VX7HnHsf/lRyI
M0aaH12zawJqAnVMO4JhGlftKv06FEGxe8cG52EiHVb7yfENO689Wxf7666aQFEkOtjaSpmeQSvY
Q+eVh+sulnUU7I/jt3scja9SG0ct8RVOzbQ4NvZHDgHYADe+PyFCmyUPBqvYc9S+GUMx3+fv0ssO
2tpGqgw7KjR+7fgN9wMzMUVLUXpqFcGgx+yytjeLRn39+R6m7rgNBPVDQyvUeKsZC+NLrjamV4Vu
2M4pq9Wcr7xocUzbXAG4o/o3cxbRfr7fQCQ8YN/CPLK9pHQwof5Gk40EtmbGdQHiRTXHEt/gH8vO
jfNGXHjaXBStHHj3YmTwxYVlhuD0O2JjAzm3CHSloHuMvSGvQwALcucTIhuWK2gO85/mj+q9aaDm
wEKBLsKIFrnkVrOMKSnyYG8DbXgm/WJR0ORheK1D46qsPniCvtiGJFnJ5y1aMEyUVmSqHxI3O3K4
oAO5n1GreCImHSVHgZ9Sxd8PKERmD/6SVZ3wZFO4nCIynup5QyEzSZiGrDtK4JzdXHzcRE6jftP+
oUz0CSk99mWYq3OBeJLBwnLFAcluijD30oY5xZidK7Xm5SPEiXRa84ty0egTAe6cjLVWQY0dsmLP
2oQHnL8ymw6xoa6W4qNTCwxFtXLCwbymX+X0bhFp780+LcBl7a24vhAr6kbkNvO7NHAUNWNJXaMZ
I1R8pizZHFvUFis/4E+I7hejIzeuJFhEb2XenYjCki+whok+KEse50AYbaPb7offnyjOUWBHiu1k
ZEjsLAXzSyZvU3qS8FwTFfdbXR8wJjmvvuuT7eXIopF6JOpmMbKGD6XWmZH2gGFdZeq/4H8r5bZO
5YPPb1U/LrxpzYkvxj5g5uMLP+YOch4XyTnm/tE/ioyz7sMIxPDTluFcgvV++h05PQlFfxWgl1vT
pj6bpKjaQl+YWt7aKebdU9sOQ6/A5Y1JH7MKtX8pCjfkzEp8ns1nSHy6UtAMjAsQ9qsIzuSf+Avn
Mwt+mgI5SAKlFEgwDXSOp8nhE0hp8Wzm/pMi9VcP3wCUSZ4ljllw+oDmOXgHptVLiV9dSu/Y5nbW
wOnvXOpdg96o0AM8zu1mT7z99X9T3KS9nUZMVDQmiTqsZt8e4Xu6/tG9FCAH6+2lC2q20y29i6cp
/Pggj92/vO3wsUWqWvQlPzE53/rTEgJizFi2GH1jaRq+4GAY8mFOUFX19WjUm8HdjdwxYNCgpdR9
XPWh3KRBVTpr0/Jnxglswo+oNcCRNeqyFH6GAgWQRlKYIlLHOG5zxrYgrbDKM1q6RbmNa22Ha+rO
HjD81aBUIhDAZrDjiwhNIpLOv1KCB/+fvtGdpOwqbvy8CTEs9De3Q/IlTylgaBEqq2Jh6vIrVogr
vSzY+8XwmgTq6Cyf3HYgBJZeg4hhOQM4p0je4KRkSvQqRXeSyL1axKiRqkMmbT+WeuRVvbhUWTZp
0Oqgse8+zB/ftGpBxc8MC8YxJYT0J3BrzZvqW88Hf3aSizpW9HojIc4Wydh0UaAZ7dYe23P3YZiu
R9aA+tW61WeX3pGJkHXTu7BxPIQSz/lYR/+BTqvSX7Kdur3Er65L4Un+yMgbRFq53X/ZntzTUKtx
E4jZy4m4cuMOKOMi35IcIGAMVm5aI6BqO1o9sTqlIrr8iFF/UCnPHOTZXdEfrV2QrE/ATWGufJdt
41urHbOBvQj4DlJR0hppp2uhqEXnyup0SRp+kvyt+P9Fs8BLavTXWszdRJk5ZGSBPjw/Z7y9AfX1
L4mrgIsjfkBfcPQ8l7aUUy8ELlxvqgq9iIDe9wU2havUGoY8fSorV3zE6Os67llxSYeuJOdFH0PT
doTPnE5V8ZITxLz+gvWbB+Wrli20icw+J8eoPZ83IBt2wqnprfLuQVUmRD3cUt31idFLv4k9okIO
y74wd6h/DfiOlt+DUZDXSdCy2XGsiKMgdrQsrzLQBho6+eK9bmxnai9orK1yjvF3osJggmEDHk3y
M92Jh/BxwetDEO/rw17pYGEWU5ADwF0Q0Psz7gq5HP3YMQhG44Wjy9st6Skyi2szJ66p7wth4JsZ
0pgrk3tV3JBa9h+K8OWX5xA2Rc4+VezxR0XCcvk2EqChLCaeigI+tK2VqgBSm+MX3R5FVRi1qQI2
DuMxf10Wn1Tz8YgvjD4np+ZSQTpfCcGnTArwFJxXBKt87wyTJdBvqHgHkNpFFhJv2fo74UlAXTB2
AV3twrC10rqKqdbhISlDW9ng1AnuiYDuWMAe08JIqzmd4hblfa2R/8/rex4MBV2lJoDowGLTAC69
g2hQqK1b1Cinl9qzmSJ/mNmJtNxRnzU5Ei/ho6avUDLVKJK5tmZJaz+KpNshgUq7sVbvPxuTv1UZ
9954aRb92L9B4RUfYgpqHB/6Skr9yhlRor81H73ZCurDMDnboy9GGdGi9MN+O8bUtMirCUofux8z
bpzwFrMGO9G5wi84zmGf9F99gF+jprBU6S+DqewspfwCS8SJa5mrT8Ztkts8y9LdBVz4Ad8LGVvi
g8wDTsW8xSC9KgNWziyu/R7DPv2v/EL+LdU1sJqURaLcQZX3616y6aj6BVjTkH1HckPXn2FYHPQ8
o2yCAi34Ql4JuLLgDnnZxln3dKDrdSdZjIr9LpTJdGqRCDVFf1Gt1TmsdGWdp0rJWpoFIVomRHu2
lQB14fSN020iD0k8KXGvBdztSaEp1Tg0mGXR7rrssMr+4Kd9Njo0k4+7PYXVZcuYs50h/qxSEFkD
J3worYv90hG8dK6k/d46Lv1BoiDJVVwBkQs6Xbluy5B8svHNUoR9sFGFvG4jBAz1001jCCtwlhM+
CnLWQNZCffcjWCYGBVXfYyM8sVKln2LJ8BdcaoajGRYHnmJRn/ZS5I7cr3smzu4YLrLN4My6Tw7I
vIrYlC9NwXn+ByI9b/MjKMthMXM20xppRPlNY5WLDFb+jbrBEzUnBC+lrDlO+zh9z4CoLs/WQlTe
kTBWuVP6q1PvXS6ZID9UfHezuF0wOFUAJHRwvZuKZGKBvkcSHRnvTFfF8oDGC7dyO4rc5U0ig4el
g7w9ItyAonRT8yXD4Il2LUwktdIVVvJZwCrqqNN4PPrCO+tM1diVMlY9nG6IfbmpLGgqz7v7yWYm
RRvLpM8ApQxwua4wBPs2gVDdsbYliiQISmhvmPBMqUgLvlwHTGLey3gNR3BekNrXtbnuwHP2yv/N
E9UT4G02TJ36EnJUVgYjcb/p0Kz726cLGUBA6mzfBlkMY5U5GhHv6cu0OytYec78JRx+Dvfo+ziL
MbkBnQ85x8t8FglTQepwldHJMMRj9f+LQCGDAUdDF39unywkoGv22jd0vb5zG2fndOAyiaqIonUS
Qdj+Hg+4oBmQwy5ZGHeZSqjL/oGHUv3qDdsbfOcqaZpx+csTrVGXs2UiNW3P6rn+olY88eIdoDtl
LcCBDBUB+KqRoK8ZnAwBXNwVNiUxzXIbpWivwnko8za+Fsw3XMYsQNztoTTS20t3u608Ai4ehr+r
KpwsFCB74SE88KQmEThvzfafH02Be6jRG+LiUwMUS/GHViVMBEbUCJKlj9sQx6VjbFyD4zNCA04m
b1gYwPHHNSgXkq6dTpXGhFEhtElSQo0pJQINiH2+J5JzMm/rk1fPXAOSL0N1jGE000yB0Xg1fhYq
QLb0LLlV/JTHrl9LKDQTuBoBeAXrcjwK4i39iy+PMYVga1RhoH6eJhcinV9iB7bCE4ALH39ZhVUH
oabNM2/kcclyoIZAzAyooipztBn8oWdjRV9zkIbsbmp75o6+/5JXpMz3+zOxGtHJC09QIwgC6nAx
lEGD9gIL40C4S1dcJYZeXT95hpsYPPryoXj52Bc2sHxxzPbyfOvN6200U5GLplrjU4LPMoER4bln
GiKvbrN75qZ6h7UBR/cszLo6IuyMal4d2Z2yvHQG9OOaxy8tWoNwWpH63nFNT2iu6W23HQbEbsWb
n/Ruckgd07krsDDskSKdxLqS/s8aQF9JrFC69q2uvvuzdxHXMhpeHAsw3Cn4LeKRbkSAL7O9Hoh4
AvqUjlmv0o8hKRVvpXzfAOxx8cXsXxDK5R9n3ZiPgs/E041/4e4/smjM3ZCaYrQRfLsf+b4iCAFt
ZkPPupcp0i5KP3AMwJc7itqaRiP2UWTdxuEfMEGXpd7g5f6ZHDRTq+zblUTePcEAW5IncjCyxEB5
eP96FU9IpGRkwWw7saSsTtEgMHD7/24M5HK54ccje8ss3E7DWS81jyzpsZt+NGQkcaFcpHwmy+kE
j8KcJ3kKV7OT3wLV6+THVqHCL6r4x1o8fKHgti7pne91nDkAQUgjOr93XgLMw35PKEL/xm13wUn/
hRkClLE0r2uZRhukpu0I0IH/nEU4nGsmNppLpjMiL05kymKrK2IQxvL6dfg3n9HA/hR3Ex1UBDzG
vQwFU9k5rLP85NUq1fUgYkptHaKUH8FjxsQWOlaoKdg44AqAq2+DRzOiH4epzujvZw4vcubHTMYU
zSR59Eug0ahuQI5KxeKMs2aj6DvpPLMaTT9Pi7jm5ItvyiYLUZdhLnC1cEZEPPyZm1pvC0lW5dB4
5x3j2Gk5yaFoJxQDSu8PUIWue/krNUuwrM9d63acyIbrkzuAhwuKw/ozDm9Nkn3xhRDF8BhQHYg4
fNBSJTqEppaiDBE72xxovbS0nRlKmA55HZYjd/u526XNtasSBahmFmK7VH8pmUPQr9XXmHNo6K7/
+9BzE3y/IfpTomTwRph2JLv5UoXUkfEX4v+ZVo/dgtuE95LKc7I8Rr7CuhjfDt0h1SNZuy6RU65I
XdXZ30RYZZWHhLymFs99CqljXWUcaLI1BnxZNaYUDaNbBtso5nrZi+GZjqZ8SfUKlFzXKla22z93
dGBhwZB87GLM1wEPdJLGEThP0/P1YFNeV1q1DdigxYwBBNh/os6bEeweESoI9l20OYeblyOalMZ7
FPzZzDKEOWVAZJtujl07wUKXSzigPBa0D/BSokevhdPwIrAP6byqk9/IT57STzjJO2ZFlT6ZPKnD
wW42N7mXsnf/NBgkZHEY86GuwbElwWyVaHpvysAEt07WqSNNkOQs1hHnIQW73M4Okr5CWK8vLRG2
l4h0yVi1mS1LvnywPwBB8LIpdo46p25l6xOYPzq0dkw7+qYxBXmioxVe7TPIFkjYqjuVFCra/TLr
+/Nn2zzQwX/LLIQl0YUhHQC7jR+EOrcE8yabBVxmw+G4a7DXgMOkMMSOr8MzHqNjF/nZREy+Y438
8OJ5/fb+waQjaPbJFE+9o8YreRaYCun0npa1YEXIKj2ZAMKGDYD655SE11aB4ovfCKCCrmifMdt2
HmDdaJP80TB+ZfE/h28/Qf1J3vtIwX84HDSS9VqQs0XerpyGwOqFYeiDeW+vKUFuXTqn+qpMlLzX
IVsFufEJGpx31p0Z6Vg4L3j2zfZS7AX7vZq3iK/wWOHCqYI0mDN8BFvuAy7AZpm2pOIDxrfounLC
Vyp8WnKSBRj0/Bj/NQOcxRkBkMvHiSrlfNGwBp5uTn0ONiLpuUTI6DD3VbLiJ/m3JN1tIwLhqyX+
O+tSr86M6EqsL2ecDZAeH5O2/Jvn4dp8oU1EzxaC4n/wtt1VKwcJDZ123Au+YBG3PfMxsDNLDuV+
78kNKRS+yNRTTjAZlA7jbMS6ZsP+Jdf//RrPFqkiaNL/Q6bqgjkwB6Cx83bNejOs1VSIPkJallmQ
IE/2lR0agzn1r272yaJRvRmm/D/guSrIoyP2KbleEG58FvIdskiqGsGEuo82Kx75z5mlEAyu10G1
LMRqu0uIKJ5jBQM1xDb2jJ/Q/mFr1+uYKwGojq/obYV3Rwf2N/OhzwK/VJWuLHj5CvepGqaFPu0b
hY8RodjRzq/h2zu9HGEZv21DM7ouSnY/WVjiqv3DoAA3ZAuRep5ULAW8AMzs/JobRox3pD/d4MEP
Bl9dzAovd8qeujobILgAckmCsSr5RQNKegZwLOsScANRoQHxBe3FmI6Acmi+v+DPtcRT8BaiVmrJ
noRzcFgIh4R16iBJCHCZ7fj6jw98zkg6iiCNy/E5TGodJcKfGDKDzJZDyjF3z90r7NQovztC5vP4
ocDJeUDXehlcw3yu5tBTAnE7XSmPiu+0PDSrFBfhcH34i07ZZFPIElZg7ZznGNhXVCj7sFv92s8d
NLglnFqYrxYFFsV0XeLGjlBKKmddGKHgp6biPSgOHxW0KQGOs2Jn4DKsjxV7YiWnT6fBSv4/BYpp
loA94fa6xAAgJRkmkl3M9atr6e6+G8h0ohiIGxzx/drO7Wui+SEYQD7QJa8KYAK7kysUN6QbhqcT
mHJLtaM4y+flK/GVb/f3678BTRLaNH/ijF0Q0N///ZvQBDHoeTYZyujyTyV7MBGY2vtWsyXO635C
lRpaJTTEmcrO9HJr0pfaw4Fp/8gZyTtyR2WCQwt69ytFv40Pw04qSjuyIt02vDRs4ivEYOu+jZfI
YPcLLdPYiGMrtgbt3VcJYwuREtXvKLHI9J0cwvteWdSAQw2aOJx1mCNtsBFVyX2aBhdxYminSt9z
1R4EVvD31iwW2uxg81kABbbpsKAZwjt/dCipYWEOj1p5t1wG4FxncxY0Me4VCUKJIHpzUTHbJxQJ
IhCujkbkQnzNAO0UaXTFNtySwFXEuzmUv9LRXV4XoaETjsRi+ByI4iMtdAz2NdpUQw0azrRQK9Fp
zvZ4lIY9WSnbulDN88BFJRX8t3pFVfPwhTALPJSVP2ixB96goKHaFFoc51vGF8hpRvkvBJkSXg9h
Akw+GXnVIeHr67kCFztwnqqtJPvuN5Z89y034SnRe5pTGIjceThPFIbabLhRh4Ba77whhoUz6Z3x
dYhYHb75WMVk9VFWV8vPxUNWzsQit+LM7ZXoQB/7cd1MpgMsm3K/sVvS6BzUhVifX5CszTlHGGZC
GvH+HxXs3luEVdHtpwQ1n91ZNz392OfxHYtaWqBgRou8M3jiYQ5R0i5u0OUpMrRv0l6Pkz6MezK4
ZbiZB3z37lwNW6Qh9IHGWuIKMKiuxrVsBFrii06+Mk7DRM5vYAc10t8pjTtjoGcf9nf3kHOxkkGn
tbRJSmw7UHkJ7NTxOMF5UeJlLOdpttm9X7xO30od8cjtTxuWU/OntMD1P/4O+w3yXECFfG04bwc8
w+IlV84cUSnAe48k5/BQKxaeaTixcBYnB6/vq2x0GnZeLrirQBwxdJGW1BHK7+wH0/Hxd5GMgrxW
Lq9zarGX9IF87T+7sB49vbbCb8D7n60cJM5wobAbhhrUs2GPH9jtEXbMnhdIUXLeE2tBvnEO78T3
YGYB39OKhpHAODqgZnF+MXzXAvmB4nkFeEf0nplT362bI7RTXLBwx3clDzTsrTwb4gQWDJ/lXRDt
f4MJfrZxYeDQCbNBZFcpXizs64WaW5tYrz+BBEsuL2rzjej+OreGBIZXA4kGYUxmPUr+dw/jR82e
lSw5CtAwxodV0B9aYQZ8FO6v6v+9C3UerNWCAELhHtSWs6YdXiBT7qc0qmTYRyXUt4C2zkzepBla
3tjcIJenu1oi50No8oKiqGUf/9QHDeI0I2Oyxxwr4BUgtbMkzUQZlaW/CJ8nh54ML5Qh/pbGfST/
zqhlznI5buHwDuAD5k3TrR7Ypl+x601kKfhbUAEEWI2xqdY5UKM7RUpdYmz00gtB5FTuxZpEn12i
qaXRKD3RlOU2qsIxKSu6hAc+dOXS5HmeaXXO/j5syaqqdrTeFNu0Oe76jnrwAc1Mqz6iq2XS21aH
DCZxUoxLj+bbBfvB1NOwKyZI21GVEw2hz84++UN6wyKFG/hB9v2rBkkYpajOl9qFzjubhPUSquFe
YbbKR81LiZ4wxEyBE5/qXGZXhYMBGzSUjefiPhqxGlriAOhlqSgosuKVBOMvtynCQIcIaApUhzxX
p6GdvekGhQqDL4XvIepPHeZP4SG5anSBrosxJNZKotxtmuAI/GG4sDxeYMeZrzSiqx5RH77yHVkr
yCZx06sqMkGJ6hlkMnhJeoC4ct0xIo3oXK3csg7SZejIEiGaLrhQMe1dw5bg50WsH8eOEDHunMNQ
/UJsTBQJemXe84NkkUQTdX3ynEAExdwdV8pTU1jFN2JsJaf5NoTFTQqxE2em/FZ5gI6ZvuKLkENW
56gJiPduQAELTPPmcCka5Tmmb25F5n/pSi9/8ahTCfjun7WSO5MzrDy8YUb+wf/HOQ+E0G8UWMHs
AMl65BQ6CNgg1kUcqP7om1v+Bp6vjGNCVmItxUt8iX0XxZJs77LHRYgM9rvb6T0ejxoMTtuZtxYW
Qd+L0lBo/qxmN/VsQTD8yfHFZpiY+Jdc2MNAKDFjCfJvg2Dn4KgQ1M5iRI5P7pXpY04WMGQtpaJt
BnHuLJU0VFMS0BxJ0Fu3JjkRJQ8nEVGZmP+TfHdnta45pyDt73Gz4GwLiOCREyJxNTmimK4IaiM6
m8sWm+OafJZqds6qIYO+KDJmYM8Gd4qv4uqs3BWBCowyjyF7rea7OMz+j8VIof0lVxPd2BacWYzc
A20F57vUDAECI6jCtHAV3ddy8T7mKyP2+48WCcFI+LsGUvDXeCHr5msL6MmYTfwQMdybO2pXjI68
1PuLfriJ0tnvzkTvqx63mQ9LsxK+Bh3KV8EDj4DedFlP2HMf562H/ACduiLzQFCzoet5HGqUKkBj
7GnHCtXXox8Il1D5Tc5vS+G+Imw123yBv2Uqs/aivZMSkUxhRHO4t9YAX9mCDlLpRQcD5chtXjzR
GGZpWAYmS/JR9S1UTwXEGrNuQyDBcEFX8AjF+NKOg0Bja/aKxIGhH4uksqxgEeFl6SeJ/cTSCcUO
FfC95EpmpS5aLFDXGkzd1fIev+HYSQ8poGN3PKj/REDfhAijZIUSWtvwn6DNSh8LlsMZ3Wrtrz45
2YHdRIcEf5eVpmwjecej5RcnPgIKY3jqcebs7AZodGBvM6dZIDGRdTC5R8mjORFFf23t7+GLYLNX
KLpfRWX5fw+Zv6S6fCKqGRsBDVPVxxyhGbyRb2qEONFkKwHyaQuc7JWB+qtvg6Uf6RJWYH8W3zel
Da6UTX2OzzxWsWohh4si/89gqri0l4dH4hnDwaNdRtKIyJ60Q+s2OOPv/k9rB5UoO3cTpMimcJjS
Y4B8Qxxmpsb9Dr2biLvHOQmxchoyjb2ted21MMGAaEi/ynhrVmMtTU8pFVhNQKgSj1lX0TOFDoV9
fZ3AzV8HOq/LRHGtMowKMiSrbNrEa4GjSEfYy7EGySCzNVhCDOIYz//VEBGdrihzst/qN6Fs5stW
0pFGqC+8Gxq1hZ14ZYCFuS8PgcnoAjpQixthUaDndRyjtjsI1/aL3N7JaVuDGAJoNvQaDzlCvD8e
+fjf1tc8/sNOdXViHV/z5s2nY9KEBcXQtNOT5cbjilaaFHQ0Mvc00acRsH6yzSPoBfP0PfAzdR5L
SOBP6KAe/Mv9k6Q/c+T2+h/7a/HajfhWlxPRKqVp7kMyPsmG1529OUhNfHUeJJpKJ6JHURIcak3I
aSayATdqEHxWnEu5ex9LyIrdzscRPDtytFNIaN//OA26XwM7LOwbLXDn2XwHApe1X5kQAIuNoP75
pyaCr1N0elyxx571hecPsWGtDumYxNkJRSgDdGTdCFX4QpivWok1+fWAh4sXS8GHjIEpaT+H/usx
U58zCiPK2iD4kK7/7+03ITmGADlyY0fcNNXjDguuhZOVXUFSyYEKsrfFovXCrGJbTU5Mm+5Wd4uF
+f7yDbNGhm4x8j3eKqJTEfJuP3IviVMgaiZx3fsFveK3twZRNoZGnwixmmB0k3eG0XXNhlcDryQ7
plAqs1CS4ZyJZmZpSvp/Ub3k4YfW0RI/4crUx4qY+gUYufLTJbTU9qYNdNndp6fEeTCrAxhkRKMp
vBaJG+PW2SP8tN29AU4RVltETYATqk9hr9fFDUHDdDiwAhJFd50UnYZ7TOTKJbSQk+/Rc7PbDAQN
2Ou2aM4pO6lfTm8COuauqzC+0zeGiNAtWm0gb7QG/yvf6VUDrxRY5i1xym92mt8d2x6EmJDTEBb4
MHLZi91kzkmfyc7AUN4Xv7Fg4AC/PKG8k60IOFAY6RcLXqPT773iG6jU3/J3jnJrS2K+hlK0eZ65
KiCAOFLNw3MpnnR1MOL9Lg9SBS6mx9MzjJj6HVLT3YgraU441B1y7edFkUZn2YR7XzYlo16RFhG0
t/PJ6m8tUIV0XTsQ1R/eosbt319xPEeguvpBH7X4DeEqiQ7h10zqjMrRkqe3qb18PFUUIkLZQlyF
wxJ019gNiVldWuJmc8YrmSOP2VMbfXuCSl+j6NAYZUzmwh+Y/t5JspD3tiev/EnLXZEM3cawhpEF
RWdg9Ltgp6PPw73iCgbM6J7RU2W5o+tHC1EIrcQMsdEgmFw7AL8rc2ifpvEg00NVxNM9nY0S/PHT
EkL91WtYMMXzhqxr7lQjab5fj7dv/0GOVtEpICw+F2beOcsKhzJrH+Awf20Bfmc8/bJRgKyXwOn3
hzI2HHHpEMFSVSBSRjzo6wUbwNrn8MSAMDI4QhUURMTHKGE1mb7187mCIBHHfbAygQDUvm0HpsVJ
FW9OR4Pn7kmaQR2BO6d3Yf+knHOkiYGnjgDQvr92H3dGkwaEsL8MYa7PIkTS1k2LimTyMKq0Oy+R
X9/CoQpcKhNYg4GWbJLDHXYZwgLDqhsen+QPBhqV3oGUFNMoPe2fSDWWOOUc+3tTRcxcCTsORbvb
Thtm7l8O9GEEU+xUuQTBaYvtX+FDFYvLGrD8f/hjzvY2aA13r8wOB/SKUhEEMzZss4vr3/ZQc5ko
ljl4PVweU1kzffNhRLcsSKekpLr1kh399yYfHfMnXB+ksTeVPTLtA/eS7VL1kQP5JNRAh3yoxmkV
2VSZXbx88dEv57R0C7YWbiD7+PhGETXjEVtCM3vKutpRwSte18NgSWa7PJPYvjAwg5WPdNpgPCTD
Sai0h9/sYLHHkrHEdE3+GkII3uVuuDq2GQoWKmnUIGI5pWv/OirSnXYN9wMPrmidG5O0Sn/oKZKG
bXG5R+2g+L8Ov5wTlVnv/zW49+7COOfQJzI6IA7asor7RUeVRDuHvihc8aR68S9Uy7PyyraK8rR3
wJXhWMZhDyrRVTixdDLpFY8hXsr6ztmlz6mWb9h1MdgrTYD5YuM9Sn0XvJDSzVXCjrk6poib5hFj
gsx5eosvIvwuLyO97H+RABqj6Rtft6DHs2XrhNBic5136VcZ1bxoT3DNNVMhVvuAbRrPe3Un/TrQ
9bjymGas/jxNzrZqhXGIo1F/6sj1sewenC2XJ9QPzk3ik78bM+4YoF0siJKYEcR924Hj7/86Tqlm
rEX3u2DPANKCy5rwUJGP5oMZl6iiaq2RZFO9lA3AixU3ETWxVpZEcSN8kxAPC/IUCYfLGUmwF4DL
hkGqINOLazhrgedKPjoGI1KAuS8i9pUwdzJ3JfKJPoJkxRswJrS5eruVKTnoJOKMlhyeipdBfTkF
awVPH0PGe0FXY0bzLq7bIS9QMSUGmPFeh8vCm5mT0OLPvEDnnHDa1ems2kOBgBC37xqL6f/iHVWx
e1NU90dPFrMHjI5CK1KpImtAynD/K6XJXX3s6/X4an5lj9n6Mt66gklrbNWZvjJOx6zjI1EM9EKM
tJE2/EUsMtMQKECc4I6uHujhfkPCkmzrTmTheD3GZ46iSdNeHy7dL4nRI9MjxdahnF+hPGDcr0mi
DJZjv5by1MnNgmeZMqC+mSl1LEYq+gkTIBT+H85mlh3t4xCwZU+MjnrO1xt2XtwJgVCM1ojxfuhN
uoVnZ4uFRnE6ooLCII76bZ7mGYpPm/93pR+8COz8+mzYHTyd5r9h7w3Nf9R3ijExTu40S4m85NJq
2bCFheSrcjCK7vB8OwOMHCSTr5DTiJcsV7SwzE2DEkadvwlIT0oGOJtmYcKtMXQib+VNc56ENTpU
yVifCDMgdNMz6iqiL95QEg3sZ93q6GDTyZaNIdHqtb0ffHeDuU/xhefo/YHrQ4475XfnHPxi9+Kx
nXBGLBhYkxDc4//vIC6usZH6wAgU5zNAqOgP/cvxnCvUfj503TdUNKOuMYVGft8DjAsCleUs60Le
dgqoKd1ZDGAp5CrCepwSyOdQbcmq2v5TKKvbZoC1G7n1C6suz6keXxJhXSCSBs+iCTw6PWp7KVX2
VTkmkS2q5twvpE0l1NP+jRM0ejlfF+FtjzdaJRkpMbVHGjYIgtkZ0GF7CSWnt3gVB281RN7cekJb
i7FfE50Tk6go1t7roCZQpx1YjuYjVcm4e7PRfILcTGzVn42EWx8VwGPBrUee8vw21uRi2rpE7gFz
SsUUazYV81moEGHZZFzmXKA5xOyl5ilmxFyFD5FrX52snamYxNcW2OVjGpDPswJG3rwG9i2kaU5r
xW0vJ0HVOibz2ZXT2Nzv73TudRddg0EozrbUs8BTAjkJRrf0Oi+y+5yRtC4oXGt8WlctlLauPxTS
Ea5gaAscNxaFhtIVzmnZfu7j/e4ICsUQdb2QZKWXBz0vccbiM7NMqfICNx08t3mjh8MgwzLkeG+N
u1NpgdCdUSk/oHXF7Iil8E/QkQEvQW5Seg+HeTmV4k3EtFCXjIkjeSVJ7wNMlPHc06NzdcYxtvPC
19KjyeybFzmGgGKo+cFHPiFf++gK/KxAaQ16IUqAL8o0gjmiaendZ8bOCUlGlk9aOxwzuOxnEeGd
JfwHCfH3pLBvLEdTjkue/+n+qFJx2bm3Phk32oTIpfDoIS9vkSDx//jQs47pqOsDrOIEL4OLIBrW
EOuNRQ/MKEV2Eos6M8YMOYK6j+8plhz/wpsP/SLocThmx1bN7srlKIhsdoS4pctnP/JXQ8RuHmJO
3KFWQExnxgdsVtHEdYgqbpSaQCA0sVl0WVnnutTPrY9VXmtpcG6fmzB8bxNaE7WAly0GGe7RIaIZ
MpktyinL7QH6KR5aK4OXZ7EMhSp072x99337CFMejq78lnxP/AKi5oM3+MNIBSm4fGGyS7kD/tqV
X6sVCTVPU9p8fQjgthkRoF43FC/KZDAXx8T+UimCaphr3oHPKNDqteUfBmg+c/ztWphmpWjQKfO1
euDfeSfuZuC4hSWzvbKe1JFvZLQ+PHASmvxixDjCW89WfuJ8lTfy7TF+V+iRYi7xAE3zWSZufoKA
thlYzoVy/cH7kpp2yssukwmTtJkSu+EWoxkEijmwq5CdJaUxFHxgvqD3sVldohHXflm9EfPBAkne
jUngEXmZeO8RyvunUe6glYtarN1l9PA5j22e3piQRIRXxT79lZrWuyOG6EKKdPumnTf8H8dhKz7Q
nOS0kj3rNVBVVbNuJTblD118hDvKkj3fNl5gFnbdFhCcUgLJNQF8TUcmyTVhkGOY7iDWM/7erEOP
b8uxc6SLRtiRcQv6Hb3+Q+T+q40CD7+p46kQ9hx0zQSwMD/fERbI3JOizLhAdCU34WaJK/dCIZu0
IUu8IFhCHrAYgb0U/IUMUMub5KOwljspvLbNpysYEUXcw0l95KfqyekIGsrx4ZRHElqWKT6ZfE1m
9BY+iP5nmBnIpCipwPkyBPbvzyzkgtfMrqau/+ySR1TvwtouHfAgm3MORFSToDj4cCHJySxHiwu7
G2c5AysLe0022P246gJeXvzFsffWMSHxpkkDmxT7ibvjY1rNdDZ5tHHLnEk24Oj6tbjhbrz/qFtY
JMV/6CIoDPxlidaX6/UHAlRpHuCi7ot94MC9plTLp+8t9N6IWqSJ9r9ibFBqOofJ++eP8StCPsx5
CIumWjFrYGLcWgWjNKTVnisWlsMkFjgK3UhUw2Bs132va5iao6CJYK7z3n9cpv/oKgUB+MefMJLL
evazJiLvyZsloYD0sLfjff4UPdExhPm1gzBZRS5ZGWnxHNVeEfQkWdbXBz5Sn6345LBg4H372YkJ
woQZ9YdaNWPx4xxNZymFytcNbn1rw64Zv36nJcwekzKHMgL4iTGIjze4+kC4KltN3l+ucgryznZ7
wpg7qya80T282hTX0Lj/g7OjYkopG1fJlGUHYihermRjoTvvX0WWTDfs0ykudxMghdFYVYD7jO/d
WqQ6UryPXeUfKdpUWSPAoU2Ys0IaiI+ynEIQhtM5F4iJoevar5GbUHJ34Dvd72HxvoEVV2yWWnCZ
7iYl29exWKkkju8tJEevfZYs5wbcdTz8k7Br2+Lj+9dESy7ksnNczNvVqKpL2UA9sOpxvKJj8T6+
O+v0UEUC+yY+KXOLmOZYmjXq+6ndFYIlClKBqrGL2Er2W2vVChv+lD3zQ76sLiUA2Giqvu7DRNil
dVh+VgIeXjq9Dcdbus590zal0g3N5su1tatswWQsANdSPWNPpTQ0RKSO0F8L2gUAl4zBPTzUDGCE
16eD++xvgcI7JS14+TDwtOAAmH+npJ6UIUR8GYE+EPx3t01D4d8ZZ0K0SY54+14IvmD4J5Z21moT
kiRcC8gW7r20CcQNA/IyB2+JUj5g7hqxOxqSxuybdd45MOH4zm1QXCuQCYWYEuGgEvaAC8zgzWQ2
aAF4FbtNu2pyaz8H86keRShur8bFZIY/00yDl/8bEkNyR5RzWIUWKA2P7LC9se9hsjTT99aaRXP+
xnOQpi5ns8bY7rg/c6UtDOvDSJGP0BNniEtmBbUU/pxdNjbndHIOH4ImI4jO9tskXZFlrtIcuOH9
dz260VI/Int+UgBUwXO2KeuRrfs1DN+pn2CvcV8FTy0z83mvUPewSdbqVfOiTqYmdsY4J8/2DtE8
s1HkMQ9rY7HQIiMy6EwGUS50BXgRZuhGvqPaLRQfNXDS2LIlI5GWkD7RrEmqIsDNRS2U6ZyxlVNp
VWuvwdZdm1hfv/RKB5/t0HERtFipwV9h0yjKXw2GPciH2UFlPE3BQ+bbPqM/h7Qi5dlKaFo4MCEG
k/aaJp1OuBnAGNOY+k4beCvlTYMm0nati7SQzUXeXbb41oOojmb5EFxfnt+h1+b449Gb2ewrQwXh
9Ru0M2VuE9m3PK3nK6O6u7MA6OYaH7zBf5ateeIGUxjWbeV2zjRDNgFQCpiucodCyVDaJjUwROIj
0GmtlZ/sttFFowmkHUhWJx4oPjpjqe9cS/pSrm+7boJeUURrwPJ4iSkfw/xpfjmcuk297g97GDdz
qUwsw9ecKNbus/9lN5Y18t+qS1tz4nRbmISn6hw6HU3vuy3zbHrJyDn80RlFEYNjV81bYZYQIUFt
MVYq1BS+ab2KZv2RAnrosYg6TYx+WuqYC6lAWnkcERjD9QJ4YAdnbgHDy328lXll6SIQ1VHTewOZ
FXc9iCEnt5m9A8PwGiIwyesR/Ipirmys+AFAZv+nyqccmmbv2f7/ZIx8SEMHU2Aeheh/4XJ02Wld
Ugk+3Bxw8ErbYH1ggKeCurRapb4kl6/LoF9X48h9+pCWsV6ZF+Io2bT19/tAArvI6ePqAgshA8EJ
NeDFjPVzdAblDWLW7HRuR29gLV/wV4vCcqjDVVILODZEGD+IXUfwhsQk31IVI88Ony3JTdsJVMn/
IxyfftqKB63kbLb0HDEmtFz1WAAhgpHS112YAo1FqjO/sxahRCB5WS2D6v/ZrpzzSZh1z4hAt+gt
kOfo+BwGB4ZeGjFq4EhkAmoEyhf/hdNC2/AMK2EIwZ/69R3j/Te1RFzAu8lEzGtlF/BIqJ1/T8Yg
9hVmvqAGb2Z/04BDGByeKpM7Lkl1Ks00WIbGZdVYK3gzosttmmVq7hjVgVx9DM52uiu/imv7a6GT
6SB9vOu2ypSz0KGP0iCB1NX4+3jnxibDwC2x3t3mQIFzpcGRGO0P71VwRcju819Vz3PxQgzDy2TR
fUeTS0+b50Pw/dclXEjJ1JGxc3OhiQM1t2b/dSmbl7YNiCq+CeJ3CUO5qdh0fRNRn+vC6MnDCwyc
fhMiKlA0ave6tvaAkZHGKbE0aA4OTQ82hqw18baoEjrAtlwNwiUvEwPd3eWLMHiST4zTvtMiVLaf
Qg+Roca+J7WLWn8a1G7w6nPzJkuf3fnJzIqoob2CV2YqRvi/0j1UFBX0vZifLKIW53QbZWNICdM7
PEZZVhw6MoOO/6qdRCiGlx1exvF9qdfpokFMPTq/sg7w2Pzzv/zs5x9U7ILnkq3bElmmTGWA72wf
y8ZB5Fot8xJ8JvnlvUuPi1jRbOIZ73XP5H/w1zb33ziBknENFTGbqMr2x6gLgWcrEZGaRr3yybKf
JnKg6yORDqNsEidRSWOZFzJaIFuW27ZR54UGzVnirUwunbr8cIvvUZeWzuEhwfMbyDwm//d78Dzu
qd5dYMfWSsFgO9lZKc0IJbmwKIc6l0bbhvAD24wgG1alcUQAreqocIjGTziXzzncizf3G4mRRMg2
iJ6xKjijSL5lhuyGYfX7aTgTL8CCSObr0zBhZY60OSiUG4yIyW2E+aRtKHGjU1z2oMQhEM8Svq8T
QaoXbhha/H5d3uPld+1zzXoOwrmNs6jBX/UyaK4KhaeZmj3BVKcaAEmM2sd+hOGZtGZup/OCkIXH
qWMkxMGenlTYYupqwzhFKH0/kNb1b7cR4lAxDzU6ytHLzKx0xSgtEemogCALdGGX+jkLcjBFYdtn
S93R5qqPO0JQ7OCswlZ9P3l1lURjzzUK6jf91PUvmT5W2tdU+p90YMLKN0w1t7xLQrRjJo7SM3GF
sfOG6HxVURObWJRuAj3ehxy6mSPg6G0JT/q6ueB96lMa/H6oyI8zhtseYUbCFfLaqdXUG/Xt/m8n
OiSB7DHOnw9PQzNxogFc9h1ZXRMftoqM0q0fokZ3w82AbyvwvY1Yy+w8Yq5RPJrD2U+Mr/TffiF/
E3tfkUjE20I1wRnFuk7zpqttDukP47nZvEnEdvWMeQ1C/yE/Yq6+hp/QzYUOaHG1JDUyPC85rHq7
K1CdOqhYOIucSVswdykEk15VY0ugqi7Wg3aD8B7enQtparLJdNGXMUh+7zXJwWRNq/FlzsO7Rxiz
ncxhD7tCOo+I0wnhzfaaoqASkeD6Wj0sYoWyE6e+6hvf6Z5zYwJq9UyOAJdBOl/lmVOJRorsZWRH
4Z4OclDhVE6z7d/tmyqnuukRKWz01S4i5g2zLg4dVwf3lEAbGBvZwjNcQu9caCWyrnObCHpafzEL
EcbDAylcw2M/9iMZQHsUP7dljkN7JOZhf6C3gtEZQ9Y4ZGoSYgHBO2xNCqMqIDMWf5bhipV/xmz1
0XDGVANk7YyLXCkbwCKh1akMIyF1RxXy9/TamVujlGetNgIFoP9jQ7htK6xMQ+WPPgUdb1tZYohH
r+eDBkU2l6rRzEDrklxg7cPq5BlFDNvl9rBK09eU1gujcQv4aq/+8pMXoBzxqtR/E5O5yCAQ1v4y
ooZMO2epVww5l2PCkB4ewCHLhMEeizrIL0OPdziPw8vCoTkyGL2pkwR/1Gc0uAdz49RqjqQbFnct
AMcn2nqWBv+sEk+M8QjDUiu8uPTi+6LMRustFM8eZD1m5A/dM/vth6Ieub2BzSdSrZ/z64+gStyW
+1CEj7fU6U4ujyNVXQWbwVpVOFR3AkjiOM15MYbfFTxdfjMWbgIHAliF3l57Uzq1K6mbJLrzJXgI
erkVm4iv5pte/pWLpf/7qQWfw8u03CFrOe7hY1Be6GrNsWQ1e77a4W/QPM32v42xxSBftpy0GqWX
lzDYEdDfX65IzLJuhAMz6Yqp94yLX1+H+/Clc+9UKnDZw5ZSzgZD7TdRbxdlekvA/5R0Q1wlk6ve
tv+dEd512xoeBWev34aBa9bIef75B16WRtjJoQboHn/T+CttaoP0zxcJ7U+TwX9B4mi9YIYbOk1e
SITBSg+LnOPQLT161Su+1USAjsNoHHp68r30FZ/vrsShJJvp5VLU2cVXG7UIilG1K2+uTUywXUFe
54E5FJbnASoMYOi+rzRpyPBjA5gr/09wmeNRmo5fBBiOKWoExUsEpIP0Mpj4/MoyC88/H4RsvAMH
cXqLztDar48liW3CC5WrC56BXyD87hqHtkIqLarzHIBuDYU5FBg8R9cX0weyBXYlk3Yle8Fy+76L
mFdaXXKGXyH6RRPmTcM8RY8h5HvzS1HLpEtcDI7LVQhlKmk2qDBgJRgcTe5LbOTArjq41cRsOX2o
1tiX39htMdx4OtlFM+1oYC2THjaCMXY3+AVt6+p7iyauuLjLtz+e90uMB1Up5b4n078/IUkhDhFg
2gCAEltta+Ouu5eZYmMWZVoWb0EaARU9KcOQ+C/O53ELoG/4072iDYflEE9G4vi5fuuczDRLyIpz
i41fWMU1d0qa6FmI/5Klrj5z1ECTIuWEy6Xg9nB5w55pmEi8WQq4zI1aWYdzJJw1c/H/j3piaAIk
kma95WuUvO0/AfoGgIU2WlaGrmmIzjMdJoIT4tx765D48U432QoCrkz6vNIPTsJxKZ5qNSx5lHzg
7fM7H3vV3XF3VNSkweaURGhWk2gYH8ApORcM9okGOEHVHjGdm8tamuWLoSbot+zkcj7LltYadxTh
NJ7wWiVGc32J6N77sjJtoLsD4tYSZDZuKzOsWvWdP3Bgg8KKNDlGBiLR990XGAm7cR8tmrQbp6I1
OwE4dVN7mVjqoaxkNXDhiDcfL779zNCyp5YOzM0T/vk1Z6PO1Av615aXw9yS5dA5QKuoiUPv9UTR
qq6mXIktADhmT42opPePqGIEwQ3CtFuD/997xkMo9P8UqD/z9l8IEjLY+9O8cvAeWj75urjSaFiY
uHm3+LukVLN5c9WYmTbuYfbe8mFANOSj7jPkUwUKoJMtGTfi0GhJc/vO01wxzleA0HPTXWxQ4zOd
OF8Ugs+DNpSG/ia9iwLdyT4wW86k0zGyqI2J/VLe66BCgk59LGjRP7e7+uFNm+YcoGxPtWv0B5lf
XoUsrA8xGaxniW1Q0NRdEM8DxCyGJ+rkxJ4mxK5XMTvqZmCdYgN/gb3dEcpYFh0NVxzlFH8YOxCf
rgdfOUY7phr2RLYionkAG5TdfZdIGaNO6Bl3KGg4f5qAXSlcr+iLmwPFTT1MDQ+wSoDNRmx8SJXQ
qPzbs3RYrR1q+3hzL6TjQ4FY10j+SYjsUNlGxWksJAGeznHPgpurU3yWfKE3fMxD3KoGeMLfEFrg
of+dtT4YuuSYQrOIn+Bo5XWNxrnISqxiRbVK75rPc9HObejwoQTQ+wmbC1fT7w+9nt73fFisVyba
f4Eht/tgK7D0Wu1cqFw+PnBXkKQDhhEw+QyqVb56iUQV4agWi4iQcBngHjFeOSZ1ueRbRQBin9oI
fCV/ZcsrVjP1kx17ib9G3VDBBIQMJ7wNA8U+JbIvjHrbXQ5ikmgW7M375LCfWS8/K8sunuUroEof
MNydvH5+E1pRw2KckUfFhpa9xOKQyUrNHwKiaiP5h8pAcMHlmdn7ggTmRXjjLmhSY4QKUTbubnLg
ZQaX7/rbh2VUGQr706TBRs580mPjV/XnnVIL1cp3ObAQmxAqE0CA7apigdbpvVUa2MoBhOQ9RnAY
PAvTClBa3KUtdO6fhpZcc/5AAp668iuaknF0laE6vRnHcF/wF5ETVYcuO6bSrQLCB7dzgubkK+Oy
r86e0EOQuqx6eCeZk1Z/Er+IUPmgxnF3J4S4SLaGhz8UV49igGo6PsnV5QiI9RnMgK67IPWAm21L
xxxCxLAAIzVbCidXgXu/Ev2H2VdjHTzMf/1EEgDdw1gJZFR93OQspAH+hHn+ihd1Z9hLFytqh9Or
gP55kNgVbl8CdfmxW4l/i/eLPJV7/WXnHwt6po1/jvfZpflQGgA/LZb2Rf9lbRz97UQ2MWJPmw16
NOHIzxK8CiRjM5VVGsWItb2sBZlR/HJpT1IkJ9z4GRMWtw+99oHCMnV6e5w6wN9nZBvF6egW3rxh
eGgSzF4Py4GiC51/dTtAZuS845PXMRtwmnpTGqM2qBcW8jiBH91oOg+gQ5r1T13NoO6njH/iFK6U
HtuKkzJW+2IGe8M97sEbIZPnZ3T6c42SFYz9f/L6ADs+1+gkx17DLIGNBb22/YTmexhsA6BSZ8ps
1+OWZuPnkcf/BJDhC3iFUKnp8Q4RpIzx3SfsXccB1vc5Iyf8teE0gHUCt1R+i9vfvnTB7gDODg3r
qt8aEeMTf13jwH695/KYvwIJ21wjviW1I5xbHwfXAToQMN8fXCLQOQSzmpRN5WN1YduACM4QVJu2
SElEZv57JHGKeayICOirlPdvOHOXeyU55zrZqx70/+8GJa7J0TJYAqiXpA3fcgqJtjn5Y2gAvvtF
/lyHUD1gDc6UdXLsO9Dm8bl6tdvGBPxUXekNpg5ojIuohd7AmoQ32mRn/tXI9b6x1PgQVXbWV/t2
iv3hILubg4ka4XdukkU9vrGRMtGCeEL4yf35slkAD4jH4t+8lBc93g1BlG7XPOMEDfW0wIAIt4Qq
cdiUtLu/qmGkXrmPUkXR/+v/G2rxjEOifT3PI9BK188pTFQkMEFQXpaa/q1xkUUT3aRcZo0l5M9c
Oi7XJbxlLnTd7M6FNuL5LzwNA07xl+/DPz6E2c5Tj2B9fRiNKNQWJ6WfQxcirZ8U0xwS0EueGgwF
yaVgo9QHAKR2GmzINfPcticzQSMK5dYyXAHNHnXcrm8RDWJN5juhqelZOA3QUBr987C08tEsCtsV
GVuC6n2MQGwCimpCoK4NxYkwgDy1vRnjq3NTOznXXeIvbVS//duwjuXfj+GA9Xf1/KWU4DhtD5Mj
IlS2AOKfg40n+iOQld40prTU2xSjT9OryehhvD0olTij8ANHaFkFxb5ZynPpq8tDQtX8zoMYVOCv
py34ZvtDcmIqmQQmZNVDDl4EESLfcvB6N5cn/zWxisQrot/7H2xPJj0GZt/f/uELqpXVqaZith08
QQN+Ib/LL6rmVrzUB5EF3XG10t9BCffMVJ86sqU/2q6TMBrxn5D2ngMyN+ArGTHxB21j1vigRLE5
7zaoj6OW4g3A5TRV9BeCCVsIiKNJMLJa4RwBREPpXE5awyQYcyZ6czkKRHWpLLNPMfdl/5TVHkce
KSeiZBw+rQ86WubhnMCxodq2G+xwsqpEL+Ibo6AWULTc+Eb+Rr1vgco7veMwEqlcxwtoba3FyWsF
vrG0uBTTDdDlfVFalqyrdVeWXiF0SmP5T/dJ3a79NnCriUKY6RpQmyRba7VuwEsFbWfsiv5ygPnF
4n31Lmb5xAqXq8QxcmpzjQbDQ1Tbn/vxmIsaCIaBltke/1ENAZu6EsGfJXmCFATVAV6h2YtlTyYD
fUWt7t5Tyz2LOSXXA4KBoSCuUHoN8BHgJl+0/mEmB/TlYqeLa+q7RHZSAWD7TKp5D/XG95r/8Pau
BzeA5fzLwQcPOfkEWIX/p2TQPEjCdhUc1Hm9MtAyatVsTEJdmERQ+okxGzkWZX7mLB9XhMBaCfjE
AuaE6s5BBY6K0cenO096IewbTgWRLAeS43xJOM1Ipdhl+MnFY1xLLxC+sxeKCCnT0Wl9Y3lY71b2
fb+7l1f7qziTfsej9UE6V+43zpyuSVeJAb5ww3iGWRZ5Ckb6/92rLFUF8hZX/J192VtNx5sdo/w4
SulrUQp4o9pUDorgn1M5qO4rCkmK6CE4ANkm6nNaLaKppm2DzKzEjXFrFSnuq+cIVY/fPzE3/8hm
WROD2sfa2CeS0W6S9pGulaG1XfDkCWWn45UTyDZQOS1YLup2BjE79vKtjyKEgTzT2S1XMn89/koW
cbeFKFWcHI6N5hYk+ZZEM1eyskfGvaysozGgRd5N1hVN63l4zqD1EW4qdXCaGBge5vpqdim2wL6x
S46MszmFbLwt3IE3fJnK2934w9z81fpK8mGlBAOaEre4JMtzLS1sw9Uh7q8MzRBuExRLQ1S0Za38
mIk7gLBbT0g5nwXp5GN6K+byXYIVG16ZwhVnuW9CcLUv/K+znHYsAUerlN8TKhEQuwW+4eirX8nu
B0ZqU6o7iABWQDQMqpvHWrGriTopY5Hs8PtrtzzaAOc50MIel0ZjS0E6kHBm/oSyGhyyzmpilz3E
b7XZIGcTzRRk54fbdp6xBtqNZs/ThFs6Yv1BB7Pjr5JIWQdgDDSpfA5kSR/9nlvPADJU2SW9CszW
m+Hec2y4PRovApnj8hjKFZ2HOMeIambmf1sYo7zJvdBskEgbq3hy/hudhMq0qsyNXZRPcXUdwGJO
6Qa2JR13yzUNg/Dj18gH3Ru81Vi4ivzgUeMITRS2mHhFbRIYR/o9lR/Q2yWlixplXGsOl0iyNbyS
DE3u8VChgCNenXz0+eq+0L8j/+afnNd6UXhxvBH7u6/lBOZMgkiTinrnp5575RimF9nI31nH4OnN
fHT2Ey6yiM88mPwbGvsiDrViMn0FDhr5jW8npAb3sj9ynvoJwUf+MEGrXjMBkTaOdioLQ/Ocq8VQ
yXEejTgBxa0DpdqLtCf5XBdasB6kR69UBSLXYvffxIsi50ccRkDWZUshxKG/5rPYs007MYUL0h9y
HYE+NAqMggrAjX4QT5/VghD9xKP5rU7mMTWWLpin/ndtEe/UmLyV+zqsbRhkWI3tOl/uPnfLnZ5v
q9CFUnGmAP7SxAqQrCb409d5otQEomdexcY1W08+yoXdtCnI/ElG4kyz401pBOR0NBR7Po6Czz8I
r+e9Al9fS8k6+Yiz6Pc2YEWCQ0MJVwX1qE3qFcx+8QC6p9m8YBcc/Q8tDP0uMPrweUzvYvo7iJNH
kd4c0YtOYYd6DnANeNXchIGb5cCI6Q7aRQNDBfeCBnc2yOsZOojXjG4FfIPUEdMco2yG4lp9xdka
A7JpkO0BiMqmt2QbZTbDLMOVOFgSas3h6vkRfFdauFa3unKJ6hTeGT1Gj5b5i6VwjCWntxbPF5o/
0Lb38UiR/eIU8MbYxa2JknHIShojA4u/IB/9BSrDHKP3rxKLYetnCDLGO/jQ65ca87qrYdjFQHZG
g6NRX8jSaJfCn0CGI9YqGzyuvjcQBsd5l+8EAoMs9qHkhJjN4KAgXaWFqbf/uoN/tThgfHAsbknF
x2F7Hc7EWevKUFD3Auolajh/BURqySy9lY+11AjZ9VuYqDyzDbPdZeHSyGJG0WXqA5JOqr2mMr5M
IrEMp/ZqoR53mrRggkgv4z0TQEuCLKjbZzXefS/y8pmoZ4aFKFNaqCH1vg/BKM9pt4CarLAyJwRw
rSG3tSNXiIVzOiKUTIqa7BjWULSz5LPzIPyIBisr/qdKU7ojbhTGXNRJ4TMxg81MoJa6ZlOXStgg
X5Y+o2Lv0NjiagYy9jKf6IfwfSIUw8p/rws5iDzLAnf+hor19ZSGW0bCGY+Dt0fcprMhaUGEAIMk
Se226NoCt/cUAdWBpBhHhHNBAk5jAWcpo8SnHA31mWGMxM1OBLTitxx0qKPM2baEYR0hQ5aG2Ny0
6NN9nUIbfgWldSWTfiaOIq9/0PMFkaFYXdjNKYzJdgb915A/IWOo5slpD+ddS8mqJUerrnihOo3S
yaYVIzAqjmDXSli5hVafZ5D6vqC75pS89fzzBRvsBLUUloANnvhkbdJM6qOvFErmwkoi/j4R0OQz
QLyVD1rwLOkiapdYnCJxifWkzK/YeTWcXh0UuHOSfH3N+Nouqh49j5BmaRdNpvXgURF1RzGOlqqE
3zPeM/lSpEgjOjcEtULKqrjR4f3JEWEjUK0OYxKa/bS2O/w4SYS4RNQ0pau1QJJwmvuTfeGC+uOu
rq/BdKpOllkNCVMg+g8gW0DObPssogsLUdcmbrsF6BRxWrLJD3UItyF1DceIUuRO8lVsruaSOS5x
/INxCqvoxXar9IKa8TKuaSeXM3GvJnEsv6XCr6YnX0j0KDRvfIXok57G/Z6M1lwiNUQGLA4wwPMn
c4xFT4i35UtaJhzL6US+XYjefLyhIo31DAPE0GTFa4XeL2zc/Egp7Rdwbw5bADQRg6FVJ5t5iCPr
xCrbOEHIIw+AvgAc2rEMF8uGtb7EYVKWM/uN0ZzSKAhST58fw0v0htghQhz+anuRFfufpjqfCQ70
c9OFppLIOAa1PY9solmPDDRit/+Jv2Gmsu3HyIduunHjDpVDWrca0f7AWOruR39ENG8OhgnNn1qe
OJ/1xS7tcCCUCN7r8RxooIFDwFLFnXpBpwKUO94YQoWZGArLz9ehAyUZHX1ItK0rD8yVTlrSIrsR
pkL97PzKVi7kDj13PsC5edi1TRdgt8f2LihMH24AVWxId7IjzXEYbOBsfTrCnwngjZtlhEz2eANo
Q0xPLPwvutKuUSSbaTuVkGA1Pl4iceBOjAScAHipU1g5tTF2KSYB9HILUmCis0MOs2LpW3ucTRPJ
PSkm4qZ+6IymZx5B/903/yuAn5ZYNdGteKaVgiSN10Xqg8gcZt3B8qZXTPnLS5i45BQO5UJfc9lL
Q4m4IdidKcHNKXJkHleS54TWLPrgsx6rRGRUNXdM+NHD8NlJMaU5rrAhOxHWeW3bSUFD+0Kl7YG+
t6ddGA/UIp+be8t23RQaBhqEhDGkjETdxms+wBFmrj8yrGep/zEBEIMn+Kk6YifY4yuGDXcdWvtk
VNP1ZG45gwZTaOlK7UVa7JgkyRzx8ViouApLDJf6/nox7w0TQ29+QpF+eDJZkLTrFFsstjPirMiy
cbcljDXXTTaj42aGKXewUE+fE59VBAc58gZGJ9ig+BnbxJ2FMbdIAzAZDypw1KFmUFUuJm4QVHPN
KhtrSGTx/BPeclkFW1EXOnHbGB4jMVjymq+Qf/NHH0j0hqzUVOdbSDomfh31bMz6Hb1EcmM22fq6
70A3Ju1eRW0OBXtVy2teQVOzX4k/e65RmLAhNxZOeCb0uIb9/xQD0SBSbDE7fIhK8fktcrFswwW7
DoVxpungV5G0v7aAxwJyAG4KECccLo7Bt8/aFh3oKNAiJ60oGo9own3cRokS6qXXHmtQomfudUbK
g7a/GrDu52BrSFo/GssGqnqVKrcBS8LTawc5Dq8TJX+As+6S5gIIKJt3ba3A9OKu6BueSCSJvxuN
7E01Wav7bydSeYcicitmvjyHuwFeI0QOVT8dmuA+PqCBhpGEgKEHKFU+cjuLTDIECIj6kEU5uoow
0o7GV2llsBVCMWnxU2KsBH8PPE1fZ+nidiizl5HQeN12MNjNXW2wtYUNWdxsLW5PTf4G0IVYPuPp
vlXcUvkh5Y8fZCND1CQsZRKu96jVGG3d2EjSLSJK395XtpaR0dU58R8nBreLMX8pZnwF0CC7WBPs
Vj13guUc/ipfA2HrDNt9iN3rFCePtq2K1uaD50uFblGc5BnxMfgEb0AdghHcHIucRilgpzKmyNED
7KnY71SIfUrQczh/FPcS6fUz5q5cQbjyq6mup6GhlAm4mL93lGt7kH4ta+bfP+bzN1NuWYSZDZeT
jhLxegjecz6vUbHHwEn6w70L0rVl3hOwQaan1ac8A+iQqVbBNBItpFc+5tAl7sYp8j5f6nb359b5
CiG1sNsr5wigLQC3+jEUHy5LAhoh2tDyq3yA1Rh+LwyhU4c03EMry+WiGqFKySNQorEogfbDUD92
S0aDYaosbQl5EnHBzMHSwEUE4tGRYjHUeGUJvlpyZs0AKNBPhLmM1E9HouVK8nR4VD5Y1h4oKWeP
OkZ1kPvvid26BL80DxVMQ8SirYGk2JXWkrgwjWlMR6UNZ4A5zWZ5jhpCil0fmMLMkcMQ1bGKtEqb
60DtWwFK1W0/scsW/azBBaQuRm+8aj5BgEQOtAp5T7WqU5PClwHzJCHpK/di1MzIwnGRh07XMN5a
HZgkCbRehBTns/IhRyJHOPazRvIoDYiWg5ScL3jYDCZnbpy3uAy2WIr/AvgCyY0NxYVbGr/QkPjD
LIbRazoui7kbQkLGKMW40ljeQYqFkiPa9L4+6MPyVu5c7gqErb9uY7uiUD2OSP0+IH6lMjy4ydLw
hb8brkL7SZNLuCCcDU1Eh3X5DPFuvQsVBytyJx6Zy4aUiDeR8/NXIYE3PDfUQ33V6Y/a4blQjbRd
KHJHFSRzCFASq9APkrmw+jP/4cOEADHFG5XxFkoVAC+2XNSJY1CXzNzCo88XPjvDOjfJbaKYgXpT
G0HAO/+DP1c87IQij+lkWZXgiZZ7NNRr/DV72IOTojuXeYn5WNYphB4aUCGPWXexwt9wW3FupQy9
32kwa/TOxLb6ObK4wRVE8Kdrxh2nQyL9yjcJonJqNSn2y6qo3axaoOVHGubwaC8/jsOqTCE3AYVr
35brNXt7CXDW+bRui9b0LoMqs9nhWBYdIaSRuKKU2DwsGeOPQxAznzvKsOdJwFNTX8gtzjM5FwUl
PaTQmBUbM+WGLiqytaeP43/hdEMyLwNRu6PPFX/djFJshsgmXeyO2NZ7inwwBpl9+UpMMFQ4C5TB
PcZa/gWyOId9gIR+iBo4gg9fyMviFjjifiYzodR/n8lror3d5QPrzfFnjgrEIo5S+jssVLq6Ae98
PXzCyxpbJBg63TeAMGO/Yuwp+t4cES9Lks8pQCX849ap2TOV9ueaQEmC6X0Xn5+/qLb5k1BLSbxA
gN2sAU+0iY/iEQ067h2WiJiKMtLasH2FWS2IyAbWa64HsuVxBW3DgQ88MjcZD4L7Oo5fMZncWj+6
F7cxqvgYBK0zHilDUEw05v5EOMfDa1z9a+NagrbbcwGfJRWh9yaoPNxDp2KUQ3OKKcuUu1Htisnm
eDB8obYhL9vtko2PXFVz0Kg8A9YoCvk8vb4IePdPhdWiB21XeZE/bR9EXR/Zp0GGlFUgQWCnHVId
Nd2u7JHZoZXjJ2TeRWwlD0NBBagHmJE0hp1OHffgSmVkobSSha4huog0O6yWQFoJA+TZTsHS21Pd
Rtj0BpcktMh9KoWcbP3acUrYdzrb4rlG6zBYJVHHr7uJk3tpySh9hkCkbZTBD9YsXh/yT89JZoV5
zeoV7GOZYcGMsE7sIPycGcmgyiLW9bJgGDuQ2p1cX52hR2p2HGNWJ7L1IWY/Q5eYPoMUdzGLfrJc
Zdpc2ihfHRUDHhTNkt8TuNUqbqlnuUIxun3vgt8hUp3ZqWlTsj1RMOYWep4JuPQedII4PRRdS2yR
1BnvkaaqzkErD1ZK8q5xkReDwLWLxAVEiKSJG7xe/y2rdkWKvggsc7iSTamQCns2WR1juZCjaCc8
FDmeo2IBz77tYrlBjNIZ3UwMGSZ04VRVjyNUmeXsYbRUdiYvYYeBmJqgyIJu5EXebAUfXaYVqQOm
vEFHEcfz7F5r440MUZMQ3mwq5RM68Zm3BD1Hkvgt9ByKw2mQql341UyhDuWdywH6DEvSoKBfVMvA
iJZtjsSvTLYzzfcH09N2/xlncEUJ16dBeYDm8CHXaHOi0q9SoXll4ZAQjOFLvy9zQlIw2uaacKMq
mtnXMV7Wq8uS3lIFFEnJJJTgqW9IF7ONinlibaOd+7vy3jCjwPlH1UofA2Hexk0k4A5eM8w5G8IB
EiTeV4roNjXxz4BmIGuQbnhX9TrtDurHsvhZJe7Qv0XscYhExBCYqskHTkJeBI0qHq+R2dkZeddD
Dpb/1oAxWixr2PX0LP3shZ1zYO15u27BQe/nt6QIkXRFXdUgO88mwbRyiVaLRs8UPe99bhaE3TaE
jVB/7E7dvfrAwwHld/qDcH1ZZopXi/zcJvrxDlT07R+u54IhptHSTigVf1e9HtKITkEDIl1Hau0j
RWFtu8lGdlmQ9aHnB+myr4AVYvm6WQtuO7q2so8tGZXCginCDyZmhznA3o1L4GWA+ph5xg7HjxZe
28eKsSwnrAqJm5zqPe32BeDGLWfFO8rRUMVPtvBoEdHHfJfaTCVyqx8TUd1XsJjmVnS1NdhZBdKm
iOL79bcYtwG5Yf/A3hvrgl1JH37KxG4oBjrllUdBo7HF7I8vQbHeAQEQGJtg0mFCHh7/icGtOCTQ
EOs75djmOMSJKplxK5mKgsEgzuz2bo1UeaJurCGKxUJ5mdyBXPti8y3ifmTATz6eAOMJNEefQCJU
xLYVI+C8JvCwx9gLvjyUJPyY1t0xw80lyBOzerwQf4ZaPoANJFdsqZYSlu5l18U1WrjAm+3k9sjZ
I23Aqk3WA/+kvV8UjcLeU0rrBDmyyYmgGpdY6dSw00eOtujvuytQTKb0s6UvNAonNt/SOwBtIuZP
RJVkcCb4xSrggCDXmmHg+3Y2b7pfERSRd2mSGCM3KXe7XXT/cqxE2TczoawSlSriuDenfevSd6iR
bb7+hdcP12l1ll5nGlycGXizmp3xizfxN5sDHRie17xmeOI4J4a98HUugmCBvt3scAn+ac6LzHqz
T8BoRSWylI29fZWbEDzLe0PPB0utA00EONh57K4Kp2Wm5cGUjID98C37CHpEv3rStspUIq3jgEtj
ZwRK2Mr+vEsfir3eU0XGJRKymRL93layczU94wSI8e8YT7sWlXate+bumCMC2ks5A7m2cMrGZZzd
HgP3PTRkPQp/pRZgEP5DPu5OeckSGKbzCfK2mXWF4Se1cs1Ne2g2sKe3KG9AzXCcs0CmiTgFxuqQ
H8a305OCNxcayMzzQDhWd+6gDPuFd97/C+ojZOFljLlCQGclATOyaqaZT3ULU5j8+elAGbTZ2j06
O3kysc1e3bGRGjIXTDYiRIG3FOvoqvMW2W42srj9gYN9hPPY2OBKeVs5aRuqq35I0luI55RKoifj
BjKeJwIT/epI+0JTeXUOmikVk+Hgs549tnDO7M2pohs+cAEk2rvnmlHwHWIq/mwN6m1PKbpV1B9L
5tD9e4u3VS5kT+MqmGdsdiT7kRUhkH4pl5LcrXHnGAaQp9UUApcQ1pIE67v54gf8r0V6RPCNlGWs
kuFVK2ruDFahk9pK4spwZq9Y+LXFxbpbsOR8SVrbJXtcw2Xc7ddqcCITA69RTetgCkvCiaEp8xVs
ERlFUphuCFjO8tp08KLi0T/JZMDmRQV8LPlToQp40xTWcduNq64FishKOsKWbraQdu6sCg0mWunu
auG/1/LgAi0AhxZ2yuK2WBitgJ1EilNDnIdSshlYNL2ClJy53pIOaDlvBZUnabci79BPFrXrM92H
1aeTsRNpeqtmQ8KqfykgLuFOK8RO8xsSLNcMobR4/S7zLr0VzsTzgEbukb3TJI67YUthOp5YMCAk
u81PDohBlZF8JJHC7/+Nc5gvdlHwtVJUWsjK0ZmMjcpj7LYbDmixlQ7KVaE8y8Zm2u4zeTHuOOou
+SgIAKLRhwgvne65jD+ZoVWVA+gW4WV/K9ArIFhR+hKCQmVZIPpPBp7mY7aTAhS2AFiI2UeeSB05
xSkMajDPD0tH3T0h5KVe2rOxHDEslDUGzpLkVr0SxWXa0XqCmbCRpyntD6a/SiJf0610xIchWGYo
RPqT90w69eVPyOaINM0RGCdC0NAIUvNQqIvYfkFQL+wOc16m301aEhKkhmUYBq1wmJBXxNLFdxFH
+iETZhcHsSSfmIpoY/4YUOfs47yADhACCasvQmqiLEH0Vbmg9QbeSfIVO9QaUmjmDZ7h2zXgrNYO
hqOhA+s5HWQ0p0ie9Oa/POs/GVUtkvfhpPfSw5UxLX4y8mbOQ3DBZTiI6SAD4e+LRDXhju/ZXys6
3cYixymvbuZXkd79IULUieMoM6HE+rjuRoJPycppTB1vd9qMeZb07Ohd+pcPSo4axhwqVjr9qXRR
+qpRipUPHaoQYtfsP4toH+J9r0Av8rXg2P1VIuk8EEXsvPaMceHzKFtugMkE4ZBC2cHSQadIoe08
A5UDSa/3hY0Rdi6dFEm86bQ6zv6Kq0Rqpo2WiaXkwmZ/uAqYLmmN9mV/Gp48mnbZFk5Iq63AFP3R
XqkQYmIhp9W2AKf2YDYMqHI+LHsjfh21c2NeKDpVW6t+FT1PMN7FLRGfRXAs8kY6YrhosvWx3GVC
S6bCJ9xIyjdjZHVutqaNhDH/SnStHCLsLLpKCiNELfcgbpOu18m1rvUW5obBObF4VAfpc5RtkFKd
NwIWnrHPQ1/pFyapDJdrCtoDyn0b29XnTsZqgSsBAnrvLNZGTKVYcxIT8HPuKgNqhUkUp9EdmfKz
I0uQ68VV7XMUCRpcwYoAM6vl5yoM3B0Kyd+YGBDwBejNO7hHLFT7Bautpn1zpwhVz7G7oGUkbP+v
aP1AgPxWl/KvB4Q+l0asuD85MpWTbe0X+qbq0l9ngQTpYCc4rlOBPMhfmO1BUCnA4iM5KjfKtfxq
Q+SJ78K/Mqd9yzEiqY1hW0lcCoSLVeVOfpnV5VdVKxF5/SfZpLrNg7r2HVrldwZ70m9msTaT4/xc
uOkTW9XrImcgPuZMBDbc8sMk3uP3ZC0/0tgMFyn+xJ1SkDPgijdcqkitUDt8Pb7GiFvDtYtCOalC
RorvlnA8zNGmyAp8ViMIEccxp5j7FINjUPVzu71/lEp1fFI+KqHgz1rzzDpFP66eHbWe8hhczFLS
qJjTN4bwDE5CZMPbAiYJsH7F4IOrzlSnXuCcAIrrIXglrpIe+ROrZRZzYIqfdxt53XDQRNQ7eOIr
EqFW3Ua+IlHkCU8s+rzeQnfaQP2D8YBQFZTmidXbQxHv2ZsZrCd2jogaScKdTFB45sw0pyp7sOSq
29gRNOjByidEooJLRy4TTQjex2ENdxItlDugwsP6EYcYkmwt0BsjsqWJwgoCXeRCE9dXM4zEyksl
DJkfv7EOwUfAPB8rFdzmFMDag0qQQZ7mvE1APepp6R+fWWxc8esjE+rudKF4AIY5x6Iz3nN5gf7q
vE3jzJlV2mJqptUoVs4hmiVGvSH8dmIjWnj4Nm3JlQ6v32RxzTekuRwPfutSdvNjplAJ/tDVmKFu
aSaq0CG6o+NNRr6Qph+HDnxsac1T03XjEnT/ltJoVtQhXv3NqI5o7Z6cTcQgEzLEQtJ1dL+sS+17
7eRwpGcFxsfw09/ysJ19wnHR6TaifB3S4v3Y/InR/RCzT3GyW+0NfIBmRtVia0YLjEflgu2LXvc4
F0FOwsAAoSHZfZWCYmcB/IROmW3PG/+MDg24LQ2zY6Ty466mIu7KNsZoo8QQreaSZycET4FljRYO
oYnDsrJtCk6sW54QhjlhDrgudWkibtA87IL90huo7n8iPSNqO5sn4ynJIU+5I3y2xEES6eqOF0dY
6kGtqZsfPpc8fjKRTSE6r4xagYJNCvKObfYs1eNRIaGRmfBs5yKl2TUJC/mMgqdnSpuTEomvwYWV
m5840dvp54zxV6E0hdY0LiY5hZZLk21kglgr/mK17mZpEAMqCgcBolHgxX9pIQV3bcXgEjFptMh4
6EdkXUJBmHXQ81U42LTi6SdCYsGTProc4w8MlzdlzzhIU9DLCtVQsD8GdTySuhwA0RaoSos2WMLE
/lDu6N++mfrvQ8JaijgeUBDVo1BehvKnxeIUqFG3HlrM+slOMnivQeOTyAxJ3c1aMIyq80TG257L
VvLswNzqm+/ouu3rYaJqs+ePdG3omJ0VGtNDPx6RxJ1cziT1h8lxfKJS+HXZj6jS3RwIz6mIXNFG
J80KzU+gbv7qKhWZ/zbAygzASu8fvF/DNWpUgTzczi67rjwai8etLDmVrxj5hdZx0TdfaMm3WeXm
F548RYa2CdLSXIi1H9A9V67VxerwK1MYXkfWwMl2Pz/CqEtBodLus2BCxmBLT8GMZvkOwV0jFGXV
k/3SG1MKS+TmJ6x71tQZ38+eMUa9wmBt8j99SaCQJagSFeigrkp0aEUb+2MCY9TBrK4C6rHCar0M
fPJEtthJ/3pQNpsod73ASjxM1dHR5L84CDn4lqnpjuhCfgHyEvjtrTc937ZXKM3ALD0WDefIpKJO
hBMhZ1qERUtZvYdWPmlclX5pcKx2cK6E3wODrCxjOQTQVCzdaSaNs2KYIdOHikXNW8kwzwbG28OW
fnml1bTo+meK/MWvpp+qQ1qYozk3rPfQNbLixw97Z/bOLf7W28jn7Hui5mTgC38syLXoVGblnBMj
KsUbX2mCYXNMQwqOh6imbpCLH4IW543Tgcq7TxgJJwQYE8qaTGimz++IldJIYf2eTsGwD8X4OjOK
RBrOQXPfyVObEI6n8qTzYrBDfiZIDm0nkeshj5O8FRvvbPbk+ECKBEIG+UmpaS/DAXBAqEsq71Nz
xMeBxQ7+Q/f3UUDaU9cMLe6YT0ARalj/MbhlRvJSo76WxJzX00ezbCiFh6xWsiFCH1bTCmFdool3
XjOUtB907dcEG1P5zZWuWJAuVgidXf9leyYHiNDch9j6zXOlLW+u07LKyhusyCv3+Ql7rJqW/YDD
KosmVGWFaxWdBDu6F3HwF4AI6FhQM4Dm+w21jGVAYhYj2vW4k1pQPmD3z83MTc34Yogsgcid5gTl
yD/nBvc8Rk+ACV26eZaAFc9o8ST392eLU8ESXKrw142v7AbGNHbK0rd1rTtJ2cJ9Mo+G5cG77/0r
hh5GyZbAhClSnS4zMudFGO2QtKKrjTEvnAbd48PlisAUr7BuWTwfLmTB4zDCLWah9FOJU/RPAZNj
SLpEZysryKmAnYTOqO2GC+6x5e21ylnaUHwLHMzb9vlWXps9gbgcEupN6VYRITOujZNpXur5v1Wb
buCzvKphRPoIWxqvt3QSrq+QuaMj3UjQERsGybFGpeAt2GFiOqHhrt3nrjKwou8win+4svyRW1By
8RCV6FEee+RcW4M0g7f6AQpsKGpw9r2Niv3QtmvPbTBfIWRqF5Ssw1g4sszb8zRIO5NHwg1fx3Td
YiZJ/ESmXh2eGSWPLvir90H9uAErOtNtvBPZ3D/6F8KwD72Q5xOXzlWSecQsnGvkp+3lTPEAXjXU
M2GPhRJaYw8ih6m5HBlv3mKAt9f/M4fQUNMJIhVmkgu1PHr5qPglbREUTZJAGQsPVANQoc9aQ1sn
i6sAVanDeVgOhIN/21yhANQwGkneV1QREW6fcOXLLTusyIxKn3TZ2jacbYJgmvJqWG9l08QV/a5i
j5FVxQGLwf4EeMH5WQqetdnmRiQIm+KDs8NSeyKF3jlHPxTF4jS+HZ1IHEuybaOhMjq8bNeq2GHd
PMdYhPDRMfExCndKDmlbtkeW6h7WXGKABvejEX55FKbh+xxrD8sA/dJQwXL3JYkjLalbX18tHo/G
pw+0dDlSrrKDcyWVCJ36DRxJXy3GxWPStU/n5TwWZ51h1crQz5d2TBY/dFbUWn53Gzz0cb+B691g
MeNcjQkpdgTQxiLtMCKAUMJziH+9gq1h5Hg9AKsKqYsDWx6JaXS5MnqvWPbtzIByx0pbGJc6i2tu
2zonRu7nFlo2JUdIIP5kIbwS3iVGSuzf6mGeBESRR76hg9VG2BasRkvZQRSB4XLl4DwdJBVjUhE0
6Lr8FG9VeGiLbBfHE5sJXh8JEY57GhPOcld0OsNDg+3omSwjw84HkdV0vECmz7sbQ7zxyQwWlhKj
ifMyujQr2mnKgys5XhNxyWFdvSBWeTWBUclJNepIjFHj/O7YKTJIDszsbRuYpSFbW2rv7UHOWgfC
ftWRQ7cPF6ncuHR+TVBBynuQghDujrwkyqGVDyOU13m8PLVnxkt6yjD+boCAt1I+mgpI8ywMTSsf
AxUi5Y30Eo3nyJ/VPqNxU1TzazdImBtjQ0yRonYqtIWTPdkzwzAlYqmYAyQ5x5QG5/Xn6opURy2X
G9ng58gwzhX0ML/Gri3NQZhwGXwcnjGWQ5ND2jQR+WMvW17uVbt2UXRAQmu7RheJGyV9JjALRsA/
0iL6kLhiNayb8V0ggkwi/yh/U5sc4Tt+5MoPrMzjvvveaNYmammfUUGvHFdF6AYbAmk4tI70n51R
FhOGVN52leneVPFfBcpzNQlorHpMd3vzAtw3t7resUV/KvCzWqykiLjuoof7ANxiZClXXbIDg4Tt
KPVdSGPFgdFef8tpcqyxZ77vYVZ66FLF4n5sWRhwmo+Y0GNjcULqLxbiqZ4rMrHBZyqjJU/0moAB
iHFU36BgeCu0Dj//QQcI9v1wLtHjc1TPVypauUx8EPjzN2/FNg6z5HqFZ+fypwH8Y18WboZ+03Co
hIeDaokEFdnCggY9Xx6TVyPuBIOP33Sn8wTMY6ozUxskESTH/UHwud51Jc+eoRHSKhxwB7ACbYIP
qrOKdzwsl1zEtubXJNiKmONBgiqeTvTCdbd/qjUFaroRWFae3YqNX3JYjk7xc29vaQMIJKEozuGA
YaGmt5qs5TGblaHs/j4ogt/e5jevkXD3DaYbu0HXwTlGdv97ZWbAqKgDftuvZbqFvHtXcPdjc807
Weir49kn/FM70Q4hIh9nGbgnYM4xtW41yO9yxl19u3mvLRobhDcvhd0YPI4+UhxR2+bP6eqG4BW7
NfcFFjG6ZE23ISt5jIAQkCzBSx6x+7TUBiOJoclBzyVHPsvWJZkMqIdRVotCgyGt7CQWnxL5SZ/M
FwTSFQHt6rA6QnsQY4kWwWmiTUE3O5FgL9FRtNTlNzBAZn+u8eIrnww3/A2E0TdA00VeqhDwe6H6
2h9ucQTfbshXAQNkDKqQMiTm7K6M+I5FrkgH8RXdi3b3bzDARpRuNWtx8LQZnuq42D27xur2Xfb6
FHQQADvK6wUS+KrNxcbXXN0Ufx6Fk/pLZ80Uu433rTcAyNoOHTZyD6SuLFmT/bB5dR8BOrzvOOEC
IicWb94OamvjzUkQvksznB3MuvDCEDLnWXP2NQPx5A6bgNu0Er+XKJYZGos0k1r/Oi13T+v7MBIa
H8Ol4YrfDwvRhnbLw4ADo490W6tj81v6flHwWxpZJCnAfW4X+HM5D25fwH2Kqf5ZnF+iTfl3MmBp
Wh+ig+zruebyI0MZktuwjJ2cYsvKnObXdJJV1B9iWSlRRaic2ZF3KC4Fee741c2HI2wUva9cFCij
50sXQzaMlzn9pTBhmP27KTwzScUf8fUb9D8h9rgQm3WRiR6YAVVx3GIMu+rqbjA81H4oSPAmPVki
PYbTas9UCVWX2zUrzDbA20+/AoNQ/YMm6jXLy2CMB5gU1sBjXNt0kjOA2aFnwJOxXpCP7e8Vw8vR
8L912LS6ICN6WigwQZg2ZvmMBerf9D97Ffju/OuKq4sRh6HcBx9Xmq4h6Pr6i2EDRTyWSHbitRmN
Qo4UPDWy9VsnxgDYQe3o8w+kEL7FzXHux3VnEpUhXa7mG0PfZMYFv1rlg2fv778nJFOubz3LN9sh
aZOrkbM4cixp4RoZqa/am3a1BR/PZfN2aqj1fyeLUtBaCtDbo9pQ95k0X+o0eTDWv+A1NQACx45J
SMLySCim/Y+3My3DCAGX8WK0t2dfECFNHlmqrndqpNQS5rvDVVdISArmIEyESVhuQ02pvUzbdtkO
Hupjsrh4Q66unbAh9K5FcplzQ3rsLYQ0jusWDMBxT7o/L+cM9o73tobYW3CsiXuxoE6V7iLrq8x1
E+TrVv0S1mIch/oDHEhTWyyTnL8dsFjC4T226CLlPVvDKzBQ8buvrnJW21BbTwUzqBNbp7RMYbzj
j7Hd+J6aAH5SjyW32SoYd9b1Q1Fak5OW8gttHsEIxsXEfqoL6u43kAuoJH4rNoNzwY0D58XKb/0u
1Kvm7Y3CQgfzJBSb2mfZFkIySPFcGL9r6VUPkUchxiWelmjY0Sw/+/HcMaYuI/nCi8zh9GPQDyh4
SDeXPVik64O8z1zTj/w3MPgg1iRw73eEp5xzOtB2zO5zcno6tMdrPg4T0z5G6ry0Nvt5cHWyD+nH
CVNDL/vhnB01x3V+E/4+yDN0opDThQRBkEPjGZW8keP3Vg3YmXAay0wNK8qjcNdf5pY7vrlsR037
0nyHIgLriLoTv1Hjr6Ihxi/1aud5Ierc+RwHLtJ5b8MzJg1jqnA/GKzXE8wCRJj7VtOOz/ko4bBJ
nAZxg0e0aarvH+pZdReBxQTkBZ1HWpi/CKatU7rU3E3qWwSpkLHpDyvn7nwoYWW96Dyj81u5zkLN
FdymrclmOhZYzQ7kPcZMgsbIjyQFzZLlqdBoPB812XAjAuJDij3sjpyfwCDNwHIDPHMU7KiNNThb
qnYB2HDNkceughOaaPimZcYALqjHBkPdD/7zQ9nBWDFaZvLJx4TnHqyMHiE6liV2jyzBtGt0cZ5W
qwmR/6wq6h72B9L7QLxPZU75IRpqWNgmoysfHRgcyTCNk27SpTr10Ct9tfdpOIKNwYZYiOntXQFa
+TIhGGUOcW2Sn2JP0Dtjj08rzicWZTd8OJwIEG7qu0VSFr+6RThghwm1PsuEzDkWI5K0HrKU7rYI
rHptHfPQzKhNokx7BLWgzMO2Ljl/g1ISN6jiutas+hyvZHiZgZlhAJij8V0BHgYT3j3xq3VrOAxl
qI9bNu4k94GQqKLTzdoHBUZwh2+K7v4dOH9JXddIpe4nf8TR4S/VSNOccdhdBtV1wUEnnvF/Kn7e
a6d92YXCUbD88v0QKT3CRW9B+/vAX9OiHFVXAkWOTi5gzPkj1p2sRohJel62G9wK27SSbg/PJkPU
BzK1B4mMJD2yInAstw/8R6/JjYZrTNj9VrO58kW/D7kKB8piYNwe9B8yDoSYfG8SOnzQmu5ZVFiu
nTLt65nVXaJkfRSMkCJpDmTL9/BSlCsrLtrOWGMOshIcW2BB9VejM5TS3LZ8UxWHAdSoo/dRQLUA
vu4jjCfJFqd1+/N2el7QThroCyPHQSgasTZfBooIMDA9B9ZqlnX9lEsrpizJmdF8t+hpU0rnf2ro
RIajXMYvXUQQhiENi1fujqQTPxXj69OFV+CK11oL5JzQT9gRa+Vah8/JhSC5IN+zDsvBBK84toME
TNehmQW8T+dNYdWdpsUItL2ZmtFY0AcvBLGsA1xjhUyiT85P4T+Av9t6qCQCJS2KvXaFEHbYvEay
JS8emfERdPgfskUjCljjbhRM3B3npYDQUBHIzEeZTVik72cpVajkDJOoIMtHRXkIqYyLvCaOGT4s
EcUkXImfuc1S85RgC83rVYyI6LI1PWFdOFsJwYvc0aLoqyOB5xAmcphep6R1dZoQ0j1PYr2Bnfym
dflnoiPpOiNKqwuyvPgKk9WssnsVLnkRn5wvseBqDHjs56Bs/l+EInWqRcA+pETLvi4unoEmCgHf
4qzPZD/it4waGfO6K3MM/LyMZv40lZ3gfULSzyqJItnAFYQSiKR1YgVOs7db9pvqJfAbFaVWg2+0
AyzF4gm+oCLilEx08e49Qkt6jANMBF8YmChzc74zNjmB9SNTbO/LZxtx66zD0Zo1cb4sZd9to8Xa
/XREEhz/TpJ+E+6Ic0vAPV/LgHpgRgEePIJKMLFbtuywVGb9rQKq/awwhUdGIjBgLT+lwGQCPiVE
uSkGsDR7HU3nbLrKoZjEz1n6j5OlUAzX9QJrCrnh5Hg+X0iGjBlZt6O/xUqeW51lG0e6a4IoEYi3
MF1LgPN5kuXfqEABgkV9WClRg79u2u/QKmX0SQk6i7g6aqbRqwbKCbDhtxIhT/Xhi7ifnTJLK+Tr
YkGYHJG8SCiRKqgW6oiYbGKrAqa06BP3QSEr+UBtpHYeLbXlIGzGReOx58jN8g8ac01HQ59TIWew
csIeRqNpuucescuL7jUBcBkIMvGEFM1fezvVwMzAlvHDJ2UPTd4FdR1vdtdHjdzBdNR/JIopzKhM
B2O7hML8yTpQwSoQYmRxKFYNX1ICdxGTsT/CqQW3/7cdF9q/ngFkoX27RH9aEOHa1fFL5UrZHPRA
dVtKsZM6RL2CcO4ZKB2BCLO2vq42HnwJRe8qFKRnJaidzGC2lgCwV+gOAgmNjEQMQBR1o/sPlHi8
VgTrLiCmoHuobpsSqya1NaBfMk7mdrLjPWY3/xvBvOMye3NV00oJtHAznhxFE67znzOEcRcStQ7S
v0xFnQ01MeVy9SY6PliGt0Tv0tbWgMpVxy4fdobJjC57m51OjKCj53r65qoEbS8YxJ69PQuseYke
ZcHPMyuIRaaKHV4eOthXzOtAqRb+7oykkYb6tKHXGEt16fIHit96TIRAWD08qSF4og5g0RPjPJ2v
awBQxmfVR8Ln/9k6VWQKz39QFfjyWEPfAsNm0MRk5CUBwo3nmPzyqVNW2j1o+ZUC5PRe6iO1Iz4K
NGStCLCo0MTZENSxYVrjIRyvBP1ZGXx+PlgjcafbHYoY2Vl6rJhWCOD4kg4GdNXcdfEW6WsRR1/s
hypF0Mtpli38I6ECd9aSuIqL7jNC0dniX0gc7led4hanjW7soIEUYP1VLBHF7mVqq6C5l9rMWabI
CJPOHkpHrL2KnAYgHQFbSJCU48YN1JPWi4SlLd21GZXqVGyPRHFXatG978yijPPu9IdSdCXPyhBx
B6B5HWWJX02CAt0h40AQuJ6ryAoUzlTSX+FwS98f1UjrLRpr2PuJu8xZqe8MH6Vkco+wUKnOCirx
UOPXlWpDnK1mVei+kA/3RvG2kEhilKVcXQZS9CXGtTGGuUb8tMQdYqDNulkqJdfhnD3tPXph9GP9
O68xYa6Jg2Aj2+qqxaJHhseozFL193Qdn276XvIFnhUhw0gGoKGm3gwJN65qku7GwLiRqnK2aIz2
qChAGxwMqYLw00R82Z+1dPtNRljyrbpCcEmHEDeZU2tb1KanOTfdgM8epwJiK3D/2Fs0e2rxX0ci
xcOB6sZSt8x/NxIMd/+OV19ZKqA0AgDkM9lf3C1LDyl1GIUjdGKN8Q1vsGJ8VcoEsO6eJfVy2oC5
DOjCZNfnHn/NmAoiZI/uYmLFrBb+B2WFTeLa6j8G6LS2BOjG3r2ZwOWolP4mRmaxhZ9R1smlRMn0
Pc58/Zzx1sPFox4sgakbRafhRof/KTAQv+SfUAe/dUCQtI1tqN9c8wnR+6WG/tmDa+KwByqDKp1y
EDdoB3ODxnqjW16sRqqhIrEUE7bys6jHTrrkgfmy/NKgPgj7rrHaWNLU7woNqH07/pDNvs8s+Oxs
IkAWrymsEolJqLL1JZvl18reQO4ue8zpAp75laJWHPFvpBYtokIGU/V99qznC+a4TURjMHlD6Pg6
OuQcPo58Dq56o9M+21n7aRQi1UhxVtDsNuiokzOLwRW/mnmT52lL/acnZAfluhqwsxVCozQYg4T2
nY+taKSTm9PImcmd9Y+3AgFexTPvPFNbIlstNVxNtSLgIcKykJPQYddehl2Mvdp9cK5imq+E7zBW
XRAYNrGOQRYx4F2jkctcYZw2Fn3CxIkOC3b1WWovgD6ttjeZCkK8794LvWlNb4PLAlBpoUDuKCzM
tK8MtfzdnvTYrie57ntWZEbhoZ3WfRX6NsiSga7bvd6wOQbiYLNkax9XL8z+txO+m51upUW4cGbV
/WUnqqtAJoezIrgy48RtNBKS0XvUZc8oHiTz9+HCNFDIRfsuGqKCJQ231v/4i6C4vsT4Y/B/I77Q
EaVZty1Dihw6uOHwAafezh5AqLadlCQBsRwNA28Qn47/V7y9lchA0ETjmmkBo+A6HCPanjcM6r00
BAhbox6fnNsAJgYOjuxs/5yJmuVHXLmOBVkCgVZXkVhweXI9Uni9+Axk/cqRpNaHK20/wgj+XgFC
0Sp+6AHjXkBBuNXhzJy3cjFoSBVz1poSm4QDW6Y6Nq6A/1uZ8Ylg2PMd9mwnrvo0HSTAKUlx5+53
j8i/4m256moefP2MBhlcDz2bMVFhUI9h1df/qLvKPkOYDjwnYmhaArgASG03URpH5eUAdk92k9WZ
T7RR+nYqHfnTxzo6/RrjqlGnkexAX9G0kPxcDEsQkwhEeWBFlhImRo5HGjoXanAfCHGQtCou5aNJ
B9RSf8JJUurkBn/nZQ12lEhMp4xIBjYvStyti6rsHaqIX94gmYKubf5/fP/5QKKuraQ9g9JTBHt4
HrgZPVUOtpVXVr8IdqOagP2ZyXmKjFQ/DqtNuGgI5agcdS9H7gron4WoJxi3NXPmNLMSzs8URU81
oaZNUV1dCt0LhFv1J83p3PYwHzoDcgXTfLwfF8BTCbeZ5iDccTshtJNlb+maCTg1TsT1nnRcYSoV
vLmUZCqLfxE/Bo9V049sQ1GnDXc13JWQ7V5mPZEJzLyscl3aEw6olqEUZFqxD75B31E7gPh/dydq
Cz8R1Yu6VLIsxquP9OZO7CSShXpDRnHfwdHw7Uygx+h58RgGvpomS0uXpyaaNOh3ILdYUIbxqzs4
UlWcYTV0PTe1PafxgW/uVjYiAzjGEjt/wecOUj+kU76M9hMwT+lOW9IuSkflmwKDDHMl9A6cDNQl
z4kQH8u4ba0BULZ1+OdC3EhLpRrx8v1+SPpfeFZscX4bVL6bGWAmt7Kf0n0vB69Q4P6l96upBfcK
o0yfObleOYYOkXbT3EcXnjlHzfyN8ra5P5rVG5VHYzB27YHj4Z6X/BI5pq/dOKYQ1IFVj2EAAy22
d3y/uRnFnUGFl6dAG6TbwL+e3F2i/09z7+vsPqT8MVPBS04F25gj24hHF7yjji8X4ANDj72AnqWv
LxX2UMDm+9GAyaN0WW0tHzLPSiHmtZKHdKGCz5Ago//ulBneKNY6VgajwIe0zjqeQlGWAnxYX5pL
c/0SY5UPGzgDyUIwSHE/HT62V5v4dD4F0DOSy8WmgNV4PYJGpwM9S1kFWI1mfwmykJBBJpe7Bhj9
MmFriwnmpyxc//5DuFNwLozDKNpL+Oy8uTouu5sbdiOX9YfGlsn9YXJ+McURo+8KiB/j7NWAfPo9
hucBi9EqmcteLxJJSN5BdJluobO+aFRPaULDtFONahYDW8oGgB/b0fiYPOcT3jFyfH6DFPo8y9cy
UFKh/6mac66CpCpAO2eHbGM0ZLNpEyg61TYus9tXkkGqmGTa+4LIRG+QeenwOt5FivBxOYP/mjBs
kY2xCkCtNlZUoeWeIwepsmcpaRRh4P085zWV9oWyKNqf1q5tgMTU3VtVdjJxOxRABWRHjU17vpyI
dS2LZ5sY5fBoJUWXHBDQKfNSZ8n2XbyllGygnngTs5rM0axGz02ugbFkZ8GpUgt7odsgCDahDzQ/
XWJUSWuyTIY6YR+AVf7qYgbZ9mZp+als9vSqVue4WKYsBtytU+ErXU9WcmddnjbsZMVhXEZvBdaL
Wr/lo0Hiy27S2JKDmOxZdkyynppCga+FCN0U9aDYWo/C7UB50E/p7CzRzAlAYDDSF4iukl/1x5T9
AHGAi1qy0B7ysCSLiixXgrkQN5WB3UuXsV2IU21LKivTHTAjKfr9p1yGEH2cA+yoDbDvMUMDDSun
eKeq7xz3jEnXrRiy5xf878kjkO9ABxXLqdL4kle6kD8XO13riL5bt2ghMrp+72seCzbTlykrQ9ag
1gWIzm6vBtj0fA/IzivoQ2hMJl+Ser0XbdmN2/9En95cDiHSzQpHK9lFPMbuvVoQxsx5ahvJnptD
YNksgv2AS6OM5loKufMtZBdDglO00SO5MvHNPUS2YDLLrdy3NR0tvNUAIIKEjtw0QuSD8mSvhRRT
YzNhk8OCcGnU5TBaZdgpf+CzNNgREq+S6Vg/0u33j2LcUOzwmsM9B+YXZ7BRnQ4AZ15cj+WUT2RF
xtP0Qmq+zzmFtodUnVb7mimup84GMTWlvJjbje1nqbPpw/pcLUeJbifnjAFB7R8m/GHnW22nc2Gz
cEsQUOuupssXLsm3YrmWi4TlAPmwZ9yTC+iIDAENoDrOCh4hwQsonZUjL01MuAM/GXxpGAvrbMuc
y8U/jyckU+PhlB80A+e23m1akMPSxEZuVRGZD1sSBS8IPFKrrEq3nUUNzv9EE9jBT+26tEKWki/y
UwrjNj5nRF8gp3sVEJL0s9/u4BoLNUn5GjtJbBBtFpz3LHnkng6efTcW5k6VIz0P6cR+z8u7FhAn
T6F0Ucpv/y+RHgI8cHyfkJqAg7bBdIaJ6gdzj6omMs1S0MHzs6qTRH9YYaAKwFCKSX8aAo8hLsR6
lmLU3OUO1rRsR/I1BPc7V6zFMpBvbL4yZqxHFqAuPG0AKz7Tmqwe97nwIvQPtspxsBxrABfoyNfR
2wtGaFDgfxJOmXDErasWHqQYNDvEbWaTQpenuyeOJdMwjnsVqwqFLzqu5+WbaYoRZKCZ7SimJBd6
SXbK240ToRcdtdpwCY3HfoH4qq3WxmEM3tVkZkB8u55pubmq+2tEEe+E6hVGT3NS4KUfE/LZCbB2
Lo5VfknBXF0a6yNR1JPw9xcLaxGV9EFHaZngZSV1wq2jMj58RII99vmxwEkgF6gfPwEwt0k2Sst9
zgEYT4jx2EFHkn8tmtwfUtUygCc5O+BPQuRsAaG3Hxsw+7PVQ2BPWrokcXe4nTRvtN0OdKb3GEyc
dkRv9cqdiELIu3wRBLaZFgRFj03iDo0r5fxlq7YiBYeUVN5f82KQm+MbkwpoaihowLhE0BEuzftY
QFSrvE6SbkVLBQpWYPXVbeMonGBLY1tgrkz1bV4ZoIVId/pc+nb1tGYv4zLAQH2/AJ7rNYZuenm0
IVEHx+/J0IJEXJ4JqTB8oS/woWeZBhI37mxw3MO0+BNuWFobBhSmzjLGIrGSFA/uZAEM1n4DuQti
fr4IeruCCgTjTBFqv2Suks+ww3SHuxIzachpmA9F4b9wF60pcnbdOO0qpnsN57Ht5KaWI+ye94ay
uhYT44M3BiOCNgO8dxKmsczDQSdEAzPL54QCO1PosANdeL0oGDXxBSoQ9zH4fbONyLbfyEn0lEb6
GmXwUpf+BUwMh6vJTWJLAAoTR4yLatNhzDD1xIStFsPGnBowEQmm2jfRAImBCS8dmEn9lzmFOm/9
FTP4OdiyN/9wNldIcmBLDj2feoa8bNZMKVsVNRu8kxFePns/204UwxHAPmjFlvX/HdymrEmCCPpk
1d2bx45sht37cURtudJT874P2ZfN31VdPVKzILIszg0sgEV4DNzlGox8AngDP0lFtylDoOV5+qnC
0iQeqfAnvv+hPP72cqgmDsbZlKMCGrOsQ7Fwg+oZBeeWDRjgzN/PQGymZCcJHdyUuafvf8PsMCtL
Z4O/bSbbtBKycpe4T253OnLWjXF1nrGXGNOI6Cm37iNZWEmbi/2KPo8FhzQEr9auRRbC9I5m+L3D
9OEIsgqJIwzabw/MGRy02ZY7XAgKdj6VYBWixQpuKdXklSZ+KaoEvPzq22WDvTIoDIHGu+OQp4lE
bwxmr4a3MES2rDYYnDKfqimEJbKTnpKHJwT05oeQ8msHeqasXu6mjv9RGrgiTn70t/gFyQfO4qVG
JiNk1Kd30AG80gD+CCyjxgBao26ybKtg7/sLRtTmyBJFdHOX6hKHEgX1jW+bzKDeFfQc8m3x0xee
VHVOZJ2H6CU4fsnEMKzNbH1ltXNpwgeXZr0sI0FZyOi7rK7jkhag5LSXm8JaGdXSjGIhR0G7V9Sc
zPX9Wn19+vEv6+H1WkwOwNAaTFqiXA+lGqfZcI1by3jsYN7FTKQQ9Jk7JP5yEVaD9X47LTOC8UOd
n2rxBu4ZDXQQN4SYAxoSmjiFMrmMrnrb2OG0rvMC49YLwCr+cK0HmFbw0IJXJQOAVoD2W9/Pt/xe
4RRoDd7iXlMI+S4qm2CFtkx2uUSzHVXdNu3CljAfDpH9mlI+w5humlSXQrRUd3xx2MH4by0wPN6c
kI8A9nYroqomakM0QlCXD+Osm4hEi4ar0CMMCCEZbDIoAbt+vEVNvlnyuRzDqVvuYBGy1rf0HSZO
ukZAWK1ESDANMBVnHGp5/lJiagOPO9DN4L3Lot2pOR1g0WapkXCidOKfTtzrs4C9bdJ7q9+ckgwR
Ot5MmSm2Sio7J2cl/gMgUZF18MoUeZjbmKf7SRWUW68MAeeh2607+H8dACiEqsDA2WO5U8FFl4q1
zL8+DN9/5TEOuRcNBq+CpA4XI/ex9liaRiRYRNI5VnNfNzqWh/1vaSn2opKvcE9x6LLGrzQvX0W+
a0vMlHQDBsULE0PuFTQpiGxyWUrJKuZKNwn5owG9lQTJJOSMkG7WZBXdCd46F542kr9bis5x5ygH
6fjwH0PnqX7ncQElDJrjXe4apBxZQ6fRBB5SHj9v4jloXLrrtWDONEzcOS2jsMnS/g+S00vjW/Gs
6T/IffcdJbXQ8HVuSETugXVTqBGQ0b2kOC7qGbuPyP71fulQ3Nq9cF9jsakzC6Gz9U5lPeSoM8oX
ZQy7al4bBKiWVxFlaDyFTnRy9KF6D49M8k+wyhU/aDamd1NazvRr2a4MaX/AUoZMw/2hEk/yk9Jc
0Sr7uCtHp1rys8LRDXmkju+S6ES+KChzhrTWlMhX4E6izvZEXC+nDBZElLQGGcPtDcJYePKFNcs/
DJYwdSF848h53VE8GWOic6YQZMdDphGAFn2Bd7fe842mV3n6arUnD4P/uw+nGaKey0nBTX746ruk
/ebpvfggUQwhT0VdWTb5attS6Iy74lzrQ5WH1xBPfI0rN/PrJ6mfLdMuOnkmgb8qri8nrpVMx6x1
PZ69ytHpy0NxJMMmph/glA2+jpwHdeiy89AdlXc1j/UyuQMZJn6PRCw5O9HtqGe67ifJU5iCW2R6
Ne3ulUjCPVzDL5QpoLaykymy5+UHPibm4xRU8TybQ6edSI15DlmJmC8BE4TTlCwtrD7gXpQoXz7w
sLti966BLhba4V8MFA9a5eErJ/4wd/1EX18mqBJTIOaFY14C0h8p0CnEXBpe2QNAJ74ozXYS6whK
oAGjoorI9cET2htC+Z5jbnoR/wtj4Z2gXgUh8/Jl/XbKUh0wBRr+JInfTzAvQ9QZ6D8ihDljEdk/
KsRMudBFIVsTgUncnEqV2LybRmkLdmyHMzEE7nDWzNrsRSXke3U7EDQeOxE2jYh57fw17LRhLvkT
2Niqt6jbA8xXD6d4p0x2VLy1jMrLMZyOB4qnAH3io5qmZfRKaryn/EuS1SAF4i/Vd7NDWZejr1h0
BJ7mPktVOXp59wuqHb1PGNnQqFqaku+UW6pjftBVgMa+eTYBbWIMJzK+9WGFhb7ZqDJRsaDUr/TR
CyAQJ75TsWWPL9yBQ775TzZHgMPxX1pEvKjKr4Mn3NxA0j2ZlcvQ72FMNLh63q7ujsMrVQ272DIj
KbnOergjGf+mLd94eiynij9lXJImcGwa8DNhjxX/xNWC6KE1ONgTy4cUXvtzzzQrhrMbeBNbaU6u
9bNV5NgcJh7NoKw3qTPIOOX8Z4vNzljULwZsQ2OZLg9CFe6WpEVjQYVrid4eePs1X6fcajKBkme4
6JjY5Thsc6NTHnkRRYqyJ4RzsvMZNhltWWTCB66MYnKy3v18of6W8vkcy8sNSgQYJTONCQ/sV2PQ
t2hNh8PkUYxv+TXeTC2Za5WtCAVVKYmy3Ije04iFhj4Y8IgYuWJLOMjkhHoGwb0T4obcQ0e83Tjl
oUZsLv22CiN7rDvaWG/YiUMVFf1guhM2sxOYkW1X5O1+tqh+udu8vvS/CLJ333ovASGu1KngG7z8
8B5vKDAidEOp1GSo6HSq2hPN9j1WrB39+RWyBIgw9NME58unC/FaanArC/UatplGBfF39ODxAmjj
UZoU050whUEf1hwaXi8J6NYVKtXWp9k6M0o44EA+t6YuXBReC2+UAGTIu8Msz/+xM3zR2tUZrPqS
YMaaXNhVz6f4Tlum+OrzHTjZHATN5eWkL672/AFb91Ei8LnUpPmVwI6seDlThlg5hwiG6PSppVUj
PLFP5BcoF5OlGPwdpw3S2WtQPiHd4gd7Tx/DfdkTxgA/30aRGfI0DxKQNuvogccFQcEF7FgdoZW9
4Rr3seD22Tmt2nt0/kUU0Zk49VBrVyWJ1T3WrcKxrMw+/Rq4fzULj41Lko5EummUddVzRVmixRSs
MJggCffHqfp1uBA7fchA3k6aSF+57gtWDYgsoj7FaOEJccTaa0k+JeaHct7Ct9iNjCHJYJRoUrbw
c+aOesRjTl8Cc87vgKyRqjD1qepiGTTOHKYnzePwE7PBkGLU6N0kCQmgaRulXiU0kCpeVfC+jyK/
troRlMpaxxYUX8NJAoCtLdV+tCiawstkBscV71EOmek+1xbddsVxRbryqS5lwgBstTUDrfpfgCS9
bDM4q/OEBssT8d0Y+M+EPRvnIMd+Epa8/zSoFpvM65XIxVHIudl4fsvYrkb/AmEj0b6qeG/sKcfd
44RSTKz0TYBlt3ez+6Xt3UcpzNeWDf5niVEjGK5TllZ78Yv0Jd0RW9Hn668e5MmME0W6WWPw61er
Q5tyQZv2VxhkKbk7s22kOJoo1HtqHZBH8VQ+EGVuPF/Ow2UgU+TsGLJe4TK0Jnusfvvwaxut3Sl7
znBt9kzimdQJb6qCQu6SoGmo2xB3jYqkFbxG13iEB/xP2f4kHWc5VWNDlx0QE1r/TG6PVxlx1/BN
S31Q5PTkLtgJSycTqvzucs6TSgJfIbGJ6DlKOEVtEfjyneEfA2o8hjnUJgHEXIfwBExP6m0KUNcu
P4r6jbIynYqv+glDMrvJo5EG6nX+7X0Q05Hpa86QRtZYA+3qH5YC9leuQMdsUqhrDxVfEpTcIu4Z
3va9VDFQ0q5YT6oPZHT63Fvn7JFVM3fJdrOA7rporBjcDOVMd0Z8kd2z2jl2ATNhAlcWzYssNb0Z
bVEnzjzm22mPqxnCg01rHedlXXasDRc988PsZHFqhPdrGCl8Jxcxzzt3TLxL5qlNe/4mXbjSN1JP
dcwhVhpooeXd64B8lrtrpnafoMW+qNYFvfBla8/OFEUr0N1d3jmiEKhsB+na1xDh08KA7zhQJiK2
FmX1O9QtN59xM86ExhOPzrv0VTW4SPuaK+gPNYYqcnb96oswxJZWf2k6hW7a60MzHA2DTMEDcWOA
/gRX9T3mCSQEXxLyYkta3d2zAuTqtFzqpU3Xy7q4+uD0rEWJUIi8m3fS736uLn2XJKenDJwAiq6g
vzXmnBS0DkVmxyG5gme6Nk2CIBD9z5NpduDCnCjBZAh+I8hFFiFcmtRq1R4yrm2U5S4+hraVVsnR
SgqpAgcUtsgOhCiFl7HqOOgFkD+vwa85g+CI07ptn8awfBD0pcTUsaBs1XbK6PKawCgI38UPMUVj
A7mQCC5wD98LhURQY/iNQ0QWbMdFps7XtRRy59v1CWW1JZXJjjwSpmseF72qaoxS9qSX0qWBjiLW
6Jy2GYtdvYvVv0KrrvMj33PwTCC4tefzxCEabOkSa0YZAWTZn/CemlOcC1Y7nQSDgNqOQSyaSh3i
iGXW8VU5t0LtYrR0bEhCljzYghQxVimodfC8xUf8mwTIY+VEK6al2fHgbRRHItxjJKwHPlMLe4w3
rGL+b7iSBY7rhUNVAEdhw72IF2dgYBHqCylTTov6u90QvpaGO7NuMSQtqqXsHRzL0ljKGUCVroAu
6HItoEn5gbIO7O9cSH+Qq3BmTL6QIs8HXW5maM9H7Halz6vvP+avlGBQESceug+gcCzXWC9rEedi
8kw1Dn9tv80OH6EjmUOj7cff7lnDuojL4nWwmN7qc3YHVUoU/y7JZCGWgBX7+MCivgwfjlAZb0ne
Z5XdtnLNxJSUb+jTviYVsYNep0yCCKtcYY8I5ANe2Pm3SmjCsGtif78U+lEOxi+XLVXPTp+pBsy8
PVbm7MiaqnbL/izDkxh+qRSPduAQSaECv538CyJwUnLC3pHRSBHlbFktaN75LJg7r2tcmxGY9qHQ
hac+X22Dl/TjmS5XoAJasjmCsqWtUzVdDsXN35/hyYYfLPKuFgl68hEKOfGEoaRB+SV6l0fRO08i
glJdGcjPJKffFs3tA75xLh3BITiQI+DoeecO1UDMTpGvAiGQrya/N5yrzMxWkiDNW52McjB3JRNW
V99IVHJaazOajawY06z2GhbSZ0TLG5j9BJF0Rgb5wQGAnxp5sjTN/Ahkxp8yAlM7KLOzI46hK2ZO
giYowcMdSxlcskL7ckSWLcsr0JS0VENxqfSJ215cgm4iWOM3KBpeaEw3MSQCHoEzlrDKIveALOwR
DBkyoQUIWY1UYVMVrPHKHF7fzz8vCsYngWI0bPL3bWC0WOUyk7Lj37G00JnbMq7eTiKDiaVhD60y
sQoaUjNsAI0J6cyM7R4SMSCsj0tfVgd7Q3gbto1kfxQTG2kRLxJ42GRMWsHTcg9Ijg0Mbn4FgR1s
1H66TVZhPO8nanOPTN2L09h3yik+aBZ7hQRO1t7+FwZGgX/0YXyZ9reYQRdnYSvMTHwnb58g4uae
cus2nUYn93Q0RL/8AqFFpiVquTOoQqYHvX1i5NYjjRO5xcb9/Ci+UeX7/pFqBpKIqM7vfO3okPuf
fuGKI3hB4WmacIuy0/znk6xu2k+MzAPvfizoXSbIUsU95jxDQu4xTH3CQMDTEx66SizLD5mvwY7f
fnL6mDLvMcaFB8vQd9Kn9PJ9oAtxnBbhpIIiAKeIB5Tuwb6seVEONCg/rqNiGtsrKBJQu5H4yg0N
ADtU6inrEOruLzMSuU7gjGvZPCXI9X3J9el35tNsL0tHgFRAbJdLVAVjMk8HFMSaVeRqXY4Jwckp
E92eb8khTgpbkHn1xhRcJmk4bHlIKDtFG3cb4HddcrT0IHk6lGkbrM0+reslZ2qwSFtJqtVmgyhM
GJQmKqjZl40Ber4vYF5t7lnnZqf7nKIn2CIXDGo2Si6YWpG+aHYjseDjochf/exNsKXHcTnVQEB4
QHCAfHb6madtwxAn8X1KbZ4kOaA5IfsCsg8pTirwpVvSe9YO7fyj1hjab3o1DsKBRC+BZCSjHDiP
RXBtC6x5Pa2ktOqzbitzl9LGORJw6kiVhW9Aex6LgpPbP0Z9Mx9hIlZv462AR/IBCqmL6IvZKhtS
F0d9BYwLBnnm+qX0FJ58SAUh7bYh583Gj1wXDbvkPivMO+FG+Zl/gNuzDiaVaJOFEtBcD3MdQWv7
h5MgHDuVlfJvdH1J+zTzbejAW2ZZJIZPiUDDssACx0fItxwFuyf276P63wA6m/ZypBu4JTAnGY9a
QYHdvGFKWskp6sMxFSqXUFo/xUj9kzEIhBn13lKvNDZCW0+WVUtCGKBjTnhh0/g/c3tXLMFFV1m+
U/Y7uFN88jr3kIfp4y2ySK7z0A356sRmw6WRN+X5/M5C0U/9lwOLgXdSnIdDbMuk7gF70IdrM0NK
4lpWCYV+rQI2ckuqIAyUyo/TP2zv4uE0xBd3oF/A6bKAmX1r/iRPU8417dazc0Y5KEct9ZS4fxLb
gTFjGnmLGXxG/HtzfophcQ0kpXLF3yoRLeZNzr4EtWGjYPj/7zk37C3PrONH0N8SuqssbUHLpLqr
ScclKSThPMQbierpSGRV/hUFtPp0tDpEF7szu6d0pNGJdZ+q0wpez7iTqM+ObzR+qxNNON0DQd1f
vv+8xpBg9ndNEa4AtOEQ+4sSanFYvqkQFSmi7GcMDasQaNKgJ/Kn06a5EQz43oMq2yETxJ4jL4H5
zDeoASez6tPAK11bVk9xFKeS+xCLb7al6lVyxiebMlFZX4oR/KVuZE3Bxji94Rqaidg3apu5Szik
wOrX/PM0e3Z3jb15c6VusuPhx0VsWzoOGf/LrlwJTT86//Bmlr+NzA2F8ZAqFeZdCX5HaKqwwd0X
rGm3zoDwI4ePAZquqhvqp57wz2vmBOld2jJUdO48WQ8Js1q8slbFTTBp1C6w/DQijMVNb4G2RSwZ
gpucI48WKZAjfgNGbfQqYmfQPCzsFudzeVxniWtNEFV3yqjCBbK3pHgv212DEcrCBk1Of4VxHSqa
CuoOOGxAVb0gyueQW2zCDh+JWYitaB4GEeLT6O93pQyHpEN5cSiMGFgkpneu0ZRoB+ABewUENsIa
jaFCadxHGIvsi1LbIDJ+TiACvw7JS8NXXb8ruv6mtMzEpH8fwfIe52lDDjwPE8hg9EDXTLt28DPo
O7lYc+DxxE/dpH+nE4ON+g0Ef2JQE2NJlEHbm9/O3Xvr354K8RNIFVvatN7hKqwYgYEoREptGWm8
TnUSxpg0QVq3VseCDQRxQCK320BPRwVXzGfSUYCbcMiwjnKYQU7BVzOekmWIehB5YGF5In+T9q25
lOUCs4WNN7MgAMCMfsOAHgctaTEUuhIuTIHd2zt+6jAbbsmnwesPIz/KxVhc93Kd8w2ArxstmQyF
dSbRLBXyF/gZQrM8dM1eY0nf9FB6t91PGVjrseTCzM87Aa7Qmpn4gN2kM8bsocTUH90M+Asx783G
cw49Ep/o4EwAGznacteLa4LqkMSg7BO7upsU25IRLm5I70AHbBTnurv6k2LdWTbzjdFKiANNUACP
wNNemcFPTOVicorT+YxAEexfY0jxwiWmFTid5abYBaTPfpxkgJhuU9V2mBcpPuAgaZ/9zD1ZB5s2
gLkvKkGg9wNMrdCrR5toKdU091r8Fe5GeOMQr9Nk+SK4u+cYbtzqQXSbLNGwbNHB0nePPEPLkOIz
ZDHXYOWa56h7+VH09jNLwCUa+1awiyMsDxH8QFrZ2lhREd1UcVri/3nSNk0og7zRLk5Niod4ZvBG
hKkvJbgnPg4tTFLrKO71nWg4H5D0bR4Gtdpvz3MpfL768uwxX30EtbNBHcInQqaqCUemU5qEMtRl
/+FMpCKltPXnkDeBx18wH8m4Fu7EkP3Eo2uS+3ZOV+py72vUEPLH37shGCNw6SzYUeK7WP5nAcBq
5ZrC96QDiePljQ5iifJKdGrADGDqMx/qn3HVy+VlqDGtJJDSQ1b3GAbSU4TI1MqSPmGb81oFO24I
Yr4F9+Fv9DVcxwsW8JEKnx2RJD6Kyx6OAhypglDR+Trwp+GIki93yAeQKLiIwfVBI6dEVPy+Rvuv
EAicw52v/N6SWNMEMBeTbaux7Ww5LaQbM94j3CDKzPLiXUmrCZcyZT+VZs4f9BuwnOKRDMDMCoSD
8WTABR0csWSJNWmIFGpPz+ZK8FZ4Ar5KL12XYUumtSL0F9S0k/f0RdXF226N8Dfv3yKcujOgbuKQ
A+4EhDpWa7hEPtF3bNXwwdeRU9wpEnpXBTNI6MtsRjpS/YYfsZTZlJwUT/1Mkbgxv8Dbm/g4TKJ+
aM4LDh6epB5EAF5FGDTwCGKSrHPQRM4y/3HAByakgg+3e1zQzIIijHIG9pQLoJEynK3eONAAq1NB
LXxEDA+MPR24+ftHn72x7Ku3OPbP4frmnq/+OQLGFEGrONOe2+tkJKXYjbsDd7E27tOTK6JhKzaW
9seHxEfY5TXsJw6WI2ujdeUIUTtWiSJSekw7Imq3YN3xUtJfG1jtoTU/LVWteIk6ZO7HK0E5tPHS
AS5wxou1Z1q0UAm3snQ3GfBtQ50eeHV1/ZBUIfh9LW3vNUNUIN9t2cX7BM8EIuH435cc64tjAZ+q
fsV4snU5cWjs19eK9bpy58HYwSUWez9/JtZfflVfiEpayOR3rdJ3LmacmDrORRESFNiGEJjftHbJ
fFYRU8I3uVxxQpIAEyGGNjWDR7YDHhBw06BENaJ5VYmoxOl26Yc76fm5/ZZpsBLcU3hmfz/V8FTF
QAcPsANMqPGHaWjZLOGNwFNM3l6OX2kYQf5j0SzlDTY6wBtbKwW7EJJR1QCfddQLm8DCqjSbcNwc
NST34sWKY3DiFYhDJhwrhJc9I02E4wBw/0j4pNbLBKOh7hVLICI8gWEfx4uQqraTwIUbWSxvpXTS
OXUfMhRGTrpCtQk6eczJa2CiwWYgkvvy7GyqP5kJuTDnsQGrjEcPvR7NZR6VE2AGlayh/OVsJtJR
kvbmJn6BFrZVV3Bc28tGmghIGJ9WKdF9GoxpoJa4GVrlexkRvxeciIuxZZM6HsvOrGN5yY6pnocO
g8C+QjtvuLniJ2qsVE4DlXPREfBDApyWAmtdIr1f1pSRIqCf+eBzWn6YpeIax0OsCkO0gxWJGyQB
IQT/3i/XPEQCWxf6RkyMav0VBqpkZPhvU5BnC4AuhIGEbl0MPt+H1U48QVjuStePKV0fSZgWcO62
JyOOioPrLNa/SYwJzfu+dE4DMXLmN3vcsDJGuTICbwnUPZYpWmXotFO9FgkHsXBdMuWYMtMlQab9
SCKG8A+DEgWml1CnZa4AArXom8djnFCTWVbhiMMpwCiBWRqpC1d8fiGbvZrG4/RyMxs4qa+STRL9
iB8JlPwbjsocQWlgbQnWYe19cLzS/F//KtytEZfFhTqTEGcwpZOopadr3swkACE17JkAhk1Ba18O
u26OeGjGWG0STgsjYUew4QzPHVWWx/pw8oeQRoHJuGlnKmrwyYO6cKmbcgZ1qNuMAN0CrBH/kzX0
BznxdOYg8/CnkxyhCpgcZP9ePLNcIzAVFn0sQyrN+6OsfeGcMY4UHEXX2z8eBrAiuX5muxmFdaRD
ZgL/FiX7aokNInar+PR1JypQQR2WCYEzLTyFMstI4xQpB+YWJV6/i0orSORXDpqq81tmuv4MeqPS
6sFZRbPu5WIxzow8hBGkN8fsx24MSK1xGAKNW69/eMAP108+xoqOwtwVrh3gYdPhncCs65S5zEgV
VZu4tKkbueSi2qufcNMRjDb/hzUlMYqeFV0ngfklqsw5ZPJMUMGgR+bhc0OfQDX+Ioej5rzvs9cQ
Y2bp/d6PZ2BKBByrjl5uYv6wVPfAOffOowkY/q9civeouCa8WtuFCFmPtmGtDvHxyc6SqjtmczXZ
Ho/m4LpaVTHhlrTK4EkZx/N4N2Q0Ih51MzSHsJsmIkmdqeRh6aLnbASKRVkIz0upK//N0NUaQja0
PLjFtPZcp/6VbT0pFqkY3EC5M5UhLA+M5GS5WOPKBmWbWAMXasRwFDtncGiwv2fGgoMlO9coaL3o
rZqrQD8nAwp6tooTozrGyXARd0Yx2WOhP6qGsUK/DTNdeRTTCd/UcsjXnNZqKQh6JRHq8XT5vbuT
yIxm8OiSn3GG5QDkJAEP8LQ8Yn8iWhzJZzJsRkCgNkP7pRdJSk7GpVu+1/OTTykDzgZHustUhRAO
kjwAHYCWJT8vVund1uhVrc1mzRsCA80Xtvd08UVfHPsQ39CVQJ4vB0R4IJosIGUbB8KqPrpMBLoo
WKE9M4UQQEVJG4niY6noTMspK/KU65E5yxYZJE9BMeKdiHQJq8Hx2LzYA4xliaWh2qEkBe8GpzRe
f+fA2wYFk5VaGuvb93B7P/ml8/yV8MRZNFA9TQ4KFJhtSdM4VtsLLLa75h6YdV70vhEM1lMwYrxX
tb4sSMDcKFKOQQfOwwWaNRh1Co4FldbQXVnWx7Qto87AZAczPvCu+mu3TXN33CM89a9mCzgn8FSc
ngaMDLOOlAJtSrNtfd0xWp3iCRHYFajhz29ScQF+03uVsWoyh61Zsg5d5L69h+9Fv1t6OinxwAHS
59jbrO4jU7RBzYEhJn2ulQcn13Ab9hHzZdfkMPZeddAS3YoZY3JfwJ+xjZNud/X5uC0yDUUDnnlR
mSEDY3KJCW6roCurGR1n2sF/cw41AhyhrbcgKHvHThBcvlUc69RU/l9XMMZLbuJOgQf8sxCJxKJi
+y7ACh45AFSbHiDcMAiWI8PLX9pWVpZhcidcQABlNE1qZ+F489NaABT9X6OV/kwiDLvWlir2txI3
mPOtNfTFlhsv0OctXCVRYtksIzvjMxlo/oz3JVoB/5i+n9of6UPPnbe9+TomSYE1TndoWouCDV8q
d3Z/ehddBH4Nr4GOdgofn91iRwvPuuUc1FUt/iL1HXwkWITa33ywWeRGJPH6Hyy1uK8bGWH5Ixxt
CsVmL+JdaF/xi196WrQi+FLrtoWgVQhoSoxYlmfRfjamCny0K24uS63iJHfS18EvixTmiSHb3TL0
BEuCVTaWJWSQyNCfAf9CkJo9ZZCHzxx3KTiaySRWSs5qTGDzd33jaoLU1AxDFFBnFCQFyecCC/Kd
kjXDKx7E4ZO/vDGnnXMbc3cIoZJcikA0KVA3HKC9Lr/xt5KblENo1wZtyfIETZcJyuKwDNP+QHbl
rlO17kH1tk34Jc66jaFy9RzVcxsZcw9yyJe1Ph1KvCdreRKRoJK1UFrzOHeGAWaoDdFg8tutcjAH
DZ54gH5e7ZFRUD5neRmnXQ1eeyNBvjkE0ZH74tXMASaFmhCd2pF6IJUV2q7g4RI+jkWySc3gVH7u
1mkPX4CVCucDLEKxz9+FN2rrGdPh2D05PnYDZjbfaxRSn0QlCKUhV2qCAUQvMgKEjpAfdNMIWUen
ups/XG9Z4OcYEQQXPGYTHGFPQd1YHSG2YfHspeybq4jG3Ucq4E2MFPqevrL3cDBwVSgvg4oxfrQY
2ICQ8Up3sUAIS4j9MuCR0yGpKZ+QyiDtEzdF+IvLOL7tqr+sl6/VV63bB382gbofwvlcUdKvSZWy
msRSlzXoY5948diJdGXdBDuCeuPpFlWvkwWgXt/+N5lWjEahNuAyLhippE3lgzmaZYjpCb2MSvyW
NuczBOcynV7HDdI+WMftWfoAtN3kHGpfBVdKmaMXeqJdbq0WBLfjcVi1UeT8tekEpif2N2APHEWj
VI1gUpJwHogkJCDKb0p6iRaqaZ2tiuJgksgzgCeQCSFEEfIO84XnLjByhZ5QHQLiQuBYjWqGiV6c
F87zrfQar9FEeAWaCMa+/T+YsXR6TrqWDM11H7XagCvTvllbNQa9jhlG+affYK/z/+wfGjFu2ebQ
18JBm4E2Q94+3jN08RHSlMmveFMoTOAd0Mv4gZxzF28fY7wqTzt87zJ/QcPei5XlYqyJmWYlxQME
rY4wSQbf7CMq1x+uQF0vjhLSUygidvd3IgWn8QpLmIYCRmt3ADxVPD4MyYoEELAIJ2ertq74LneP
hokqI37EPXx5EHqY7Np4HLoXQBvJe2lM/j3eVTe9IO7Qaq+bsdDYjKDVTtiZfd4tqPRUl25LLP/Z
lzOR32GnjJze46K+fvDWg4aRT5FimNF1TnYA/L8nTq5TEMv8O41IIMHIOT0g0jMJf9xNb2S5Oec8
peNwO/Ctmc3p8t9fGEur4yyqDZan85YbrbQlsVa2YyXzOiDcVOe6RWLTiLF4J4BtjHWka7pcw5bF
h6bnDWRMabJHKB4qNZfESfMJMdEZ99mEk9bSVKPZMFE9Wk9QF7I4CsLoNrXmjtCRksVY/Y9YkYJm
Rmz1T6rnOCUZMnOTip5ozOkTIXoRdvqeMdozgsT+4LTkVrV9pndzRcsoNY/nq6/0YtjxjLRmvkec
QlCO3Wmh6QpIi2mEdnVyT+PiVerHBx6ud0eblck19eYUVXVpnobFgnNSCdZx5h11iZYw+sDfKiOu
wxjKctQBx+h/5KQjoXC6UOACyn5dAbSrexEk1f+DEnx3UK3u/K3mjiLqF0lqZ+WlBxLanM45O7ml
JLl4OKLfpmK6nF+TVoK/x9vEuCpS+R978r/0B6m4i6gheiFQ98lWBtYuNWWAYheRuZCkQhf4HtqA
x8MjJo533jMfYu7yQ713UsI09EFLNo20H1YYs514qU8QIteLz+DeUYnwO261ORMlKpca8pYJ7A+H
WS9STSceu88MICMwOlpGLx+dGivEXEVrhinspPb0kRf2tbar5NDHHC9NAvhmCwOCKgzg9TelrMK2
V85FCzwb2qRby5BT1+guUpg/RXfhR7mJiAS0XBRUFFq5UiZ7mz3QRAGRZ3ShE8ljmfAA2AE3wety
h9OC/VVBvT7br9wl/7J2mSOLND742CEc+1iSe3IGjzWlf4zpXTTAUkn+xJpOmFnZvuUaOgu4++W+
1Uu41qAupvo3I/Pa3uC3lSLh/JmBbicmskSCp3yt2EpIAWbJF6Q1tKhygsv6S08ITIVnkXsWOtfg
F/ZLsFbZewhtwL1tlrF9RnNtu2VMfrM47zGCB7hi+0hjjTXXA89A+Ft03ZNf5rpUvnSG87uxSCMK
hCvMy4uh1a44nMo8P199y4bLBpR2D/ZFGeFxrtcymN/zNclu/BGgLvbHXAczAWMi0EWls9tem+Uo
LhgB9kELJAPqVkmptPJuieq/eQvbmFHJQZk23Ji55e+Wn+nYUJRx4iE8afYSybsPYw1hE7evA20N
Ddvhcdie51gHtxjY5RO1o6zGHsQE1/OBGpNbxPOwPt2sbUKxStIHgGagtD6XzJ8G+qS+JZctjE7M
346uGv3p3cauW++/oiI3PDpVx525L/hrGybS4oToMQR7VYsY1QmNyRtCjckSVwof0qm4UsyfNqVD
zbubIXYW3jBCg2s3RdRbzlZ5GY/FQngUUBsb+SCVU6X36ZvGLeF2/gfTeoF8a2SIkJW+rMTm33q+
cFNn65UOzwiyJYrPC05EovyNH6cqshd0Yw67bDCqOTrrUUtNlXxrX0ptce7737im6qZPwaPaLBi7
cSV0rL1iufqN7gaEOsGA9f3kXNOH8841bNPUVlQXr4YnPPwRFD6X0BgQVoqB1iagmFR6pEVNxWXW
iRO5ZtasuzZLOA9nleOxil17WkuOGgbCnT0XvXOf1yi+Jh1OxGTLoH0ZDP0vSg6vXI8JKZkN1Wav
by4Fc0HTn3KoGnfFC32n8R97pZJyCej5OxkUmNr8akAIgBF317g6hr1Wb9kkIXCQe0QYKHnQCcJr
0wVCvrY9Qk3ETT0nkEGwLwTHrDh8yqEsXjOFzYCKerLaCqAmZh5rZXc+WBsMO1HrqN76tDaBsL5F
TbVGI5jFOm1+0kdH6tUtHYqa2B3jlSk24+Ek+weN7VeG+nbrv/G3qStqeTtD4hK3hpJgzr78arTZ
W5ELC1uYY0mJahrjnWVC8y7CXvhr97KRkrY6tl+Rkh82Oa0rfENXYylHQvCi9S5w5x19ACniitEV
IZyReriLeEAbfnx1QFZat3JxE3Mhn88NVTKklRJk24dNTex2Nbts7cslU4fKNdULiVmZbc68X8O9
xqrgk3IW5R1b3IgOA4uS1Z0YtYYcSayv25piPeFjPCNRxUB9PDPI5rXD/Mxs6qCxobdn9FZQV5+w
l1WjxNax0AgeKrvfTzRYezmYYZI9ud3J0s/qJ0mVulmpo7DIt1uxaV7S91GtGxBgG5uGyeBPPn86
mob6GHh3JV2FWJsVggE55F5qbiJkU45UFw71vI3NHI9aSoQiz+35hdEjWbzKpdBsjqWFJqLQtJwp
clp6KbvCnKdfFx4Ky1QJ/0BylMDZfy9oeLEHllgX+BspCPpWztaGL0n9HN0RpieB1E7EAC+R13s7
lCtzo/Qo44MSnmft+fXsIrESdhRCDsuFlsREOm7aG40u4zq4oveTnKuyCGTBIf/8KmlM+AguC0k4
oCZVUOtk9HB8P890RK7mM9FtUsG4Pqyg+rcFf1Ezy+MIOZUmF3edFhEBHQ6Hf62uRfaMFfXRxOWM
m9c66QPE9A4Dcl40UB89qsEZl4PV6X8PkKCMSai4irCKrA9O6lXZRa9dHLKmcrTvX5LvchTYHzGW
mYtu6pNvazX6XZaYabgXJt52THc/Nba7+4GqFsDfx7Q+XwHEJd9MimjZe6DtuVLWGM3tOvkKlkW3
cxgXbJCZmEKtZ4BjRAG4qWx5Fv/0OaiaZ7EnuoDQbq3HqeQ+rxtDSl8gOKObl1OX7ruIzgAhBJgl
lbdxv7XXMyiY6OnfEfbn0f9pqK2I7VUdtGxJY40f9Kk/F0QZOBKcvrS5Mrn7ddXzL6noWeKGxOuj
Am01KKuuRgfy+N7xMFUi9GwtdPUqzkvKgAH3sHhgA2xlFdQ3GXH6y4nuOW3mLrS5+5aib157Hk1s
1N9OzYgHyOWPmg++3I5/hiUfN0X+AFpswN9rW58TePT5QXnuxI0LL9SChO9TgvIXIsKE8NtN8if2
pOwpnZCt9fV1AVBbXGx5z656Q7kzuqIbriQVX3Lp0jea56sNhKyq9yVu4aUTJ0HrPrDxuPbOelwU
ZgcP426S1o3lgmY9aC1OJIw4Mf5NceexuYBxEVVfI+KTnGJNArhEVRlG63O1UEeLzfiAqmK+xqJv
0Mu5wQkQxwfKiseAcQ5YNgc3Lc+ZflqqYW4FOfOGuz3Xv8x3bKdXTydhg+XpfyQsawKMSgTF2cvM
UxoA8vHOSaxKZ3xirsM/ELh3jvWEpaHSLdquPIHDHWfoPc476+QjQYo5HiHw/l6lomqSNO5JiON3
6mqJg9UvGuEhYQTbrJ6yO9xbzusyY5LILgTqBFibp58p3pW6xNLoyimDQJPOAMwmQO2BxN0vFUTO
3o9yIaeQCz5NFTTNhL862VOC4X5NWgqBbaO3lfvSENsV1/3eng8jH1vdTXb371SEaerHoH8fHP6E
7qIPGDkBnq/joScluYgwe8kyEVgPWJ6D1CDuY43FSU0MMOurlj5IdoeGA7F9PBAHHD+pzSAVG5A7
xXQKYSyNKBNA+IhvGTgW7Ykzeo63Im5lTAJAA4MX065P3X/HecdXp0+aIUnVjdKReVSiCKjoUEyl
kQHBwngzqVj8ROGNFae6je9Q6khFatFntlGurOZ9YFIx4u23j4kukXUNmQUjYtea04/1i8397CsE
Rsg65Zf99mIARUXfch+ENindRdDFLEqzwUhGT8Gu0De/DFrf5BXVcWNUwkYdDbRlBBogdW/rVBKe
x724HUNEz4DfRZJ33ovVunvfCqndx0GxMte5T2A0jpieky8MjQQXzxEOR1ZrO7Fca6BQPVpjGhSb
5c5VPYVD2UO6d6HhQttHXP14L4ZqbjcNBCT+mbyHf1WkuTMrAJhzMjNdYU7K7YE4QKG6nYbnXEJt
jDUOYuaodF3XtnUWoedrraAGXtHzDfR5qYTCANvZ8NHnnK4NjXdfsbuhl64LnjPutcUrOkMlUXoT
QrkaE/drn0XhZ4PDywtx59xe3FL91VuUA6ttIOnhF8UPEd3VjCwU4g1poSTYwWHHq0Y4D0tLQXDF
4YG/NXDfipxtKh/Go45W4IcdE78Ew8imw12l+ekSo7WKJeNQ/XbNTiB6r9+C9479xIeq7Lsp0W5t
kBwNB9nQu1RQFl1UtmxAWxXUQKcSZP3zSjcy6RG1If5m3rJpSY0SaydVN+g5LuIwhRYV08Grc1JO
qzRtfsxXUrXhaOjb25SCKW6JSQSO1hEsaLQaDIo78r09CkNZquRsl1POl9CiKBqxlcWjaSkfOaqC
ASzgREQ19U7H8yLdpuA6vkOuH3gQrDIXq4W4ECvwsVdXgcDxUOZwmIHgaWnCWmVvOTdPNJSBDZa1
Kt9LQxF7OvFdEnhVeEZxfYOp+t5H2UDXCEj5FNBYmqXB0D+Se/Yy5Y0/g9aKKdyqY0z4KBfsb0xy
wVahla4jUIvzb7fXobcwl6KaQCy0UqbBkahRSK0xMPzm7+8ZL3qXS01/05MKQn1xp1PULXNqPyxL
8gz8VjreyRxP7AvVmHPcPKPnoBJ09oyo6kWmfnZ0IVXgoFLCYoxHGW4ZcNhYOmN6MARO0jC0QL7R
6v14opA2Xnsuhxca5NhSt4Y8Fmky+Ejnk6SXIgqRxmHAW0rgEK17kCWieSfH62VQMPWND/PeNIO0
pxuiFJ4b4ER8AOjVoD8fONozaBb8k0mkxk6U9QvoQx3nhDsWux/txxgtuqFIAEm2myG5Gvyg1RBA
xQMOCZAxAleFf/Q+Ds8D4mFaskSOnN5Tuwv6WS3qrcN8WXMguR+oil/oq6dBO1BaDW+KzFDIMUkk
E2H5as3VBxRfll2D+ZaSQDdTmLdXEn094GWsm6+vABaaQ7gCTpRB5DyjBJ6fvW0miiUqOWfewT/w
M4hqwkzUm6HAy7BfyGuM2yK9vxYq1JILd0A0cX/C+aj7P5nFJYv9kmG7tptPQSnY1jCpoVO9HvGp
wcX/Ti+gCp0uhmpvd0HHFil/i1z2nY56k8O0wkILrFZNJEyZcKHlhCiQd/tNKne6M9RdLj5M62T6
r1Vj6482fA23TZB/38nrA/Y8eiVYccZz2ziFCsChc1zFk02JaZEnF8REYLAfxGsXjXmAOcICCm24
WXisWRl9EVz/rKXbC9ejqevscUgPtFiSVr3OFA/ydrIoATSzcMx+vRyGnVrfrxXejCYejHse36/e
21L+xzvNhZ/meR0R65DWw4Lo6lD/Pb8MQnorVbIIvYnqIolP41Q2LNe3GiLFzfhKp0+2kYOACKbg
rgnNkxfqWbk08/MlSNkaP52Dx4s9VXWlPeL9WSGggaxmThQjceRaZAb4uFsMNIm7a949G2qPQ4RK
93J18zdJV3UCRa3ir/p3UZGYHplDcLFuxp3gdo66SSkCo4u/aenXusHE9PpCqhYuNfYp3kP8FeRq
8mQ+etmZz32anjsAqEGEHbaFXDE/l3Crvwn4df99DqYTUJ6iZu8iR9VNcatkYOUGI7JoPFRyE7R4
6jlbgDqKyRxSOyTbkNjlH3E5l6cJP1lyWqEmi7hvhl/kTw4S0Bw4Pp5eBlSSQD9/SZBJBWEFlleT
WJ9YVWqFdXPLR0KSDP0f48nINSXuTwXOv0lCDH4Ngb6p5X2wvs4flqNHz7PXglLBd8OIFWEt2U7S
ycLvFSJkGjgQ7vz9YWR7BA/qh1X/MXwY12K6QB6AXv8y7bL05r301tpkzaMk39lxvUzPgQKM+a1B
C/f27qqFbikH5yR472pFOEmfAmdtE3lgg86Ov+5vkloTfSuGSSHlLjuOpLTGXqvQB981MN/nfJOm
sBDKOznw4f95q+6+97Fen7vYig/sUa/wtaFpR6tYm6LsCxeLPRAJQg+Mw/FvZzBSZ5NepUDweI6E
TtQ0xRVg1SbtJn5mLs3F2x+jV8nlLfeya9PPU0y9GqHU03XMoxKKatPlarIZRdO012703QDZQVYA
N0G5u4xatvHFcWlP4+ooRFrEbWTYc//1LlMAdBSB4i34wC3JjKJh/nnGtqrHnmK1Y0zAYOM9FSPL
EGn/S0wJQpfXfsmxy9KAr4do9tvsFJwZryQDbB5qkU7h58lqflRrC1NL3sibyjJazn9pcfwSM091
4WSi9XQdo+Djtqi7BYiyg3/0PzDtlWtMi27FQMpFsptI0owi2jHnj+TOwql9Sy4i+ma8ciN4H+zi
RCQWY1JxkPD65QQl3R9oZTELRrDYGVqoOTVGGBf6mYk/UuRdwAbPsimR5DCWI4AsS6YZ5wKK+1nx
bMltVGMvbYdKQtMZltVY1p2jIatQe54m6qnXLSn/+DmHUCrkbhQa7aBDccuQfe81SMbrtHHtWB+l
JZ3Ou9sbvtp3DgZRB/c2OPzakvbO7tfA+F1sp6gB5T+Xa5VMHCf6w81RN3l0r3CG6IU7UMkMAPpW
7DSAVCgCjKuAIwIvVfnOBVzl9lq5xRcgH3Z2PzOQC3P4/um3yqAWj2Cx07MupUb52tWHUxQC/pFf
rN19zxmMYVpa0xSqk03iJk0DDoWdb8lpr0UPkWRrNlNY4jfKHhDL06NIprqIX3uqFAPjlzcrEJy6
yIonZa0/GwLSz+tVYNdCm1yKBrqRfL7oU8QR4Jqz/BfWA8M3qHb4LmDETR3WdE9461IMjzOsdiaf
LNEFbpfpzCw6/ck69ovJO03PkgpXgAsYeajXUXIc06b+Mt1gljZEHJUdhzPsGpIwJYJF92WalvY5
qIVSTIlKqMzRrQCEMBJ7HyOyC6NydhafAHYwqped7bmMyP8gC4dUOVGpj/c+fPgwBcBJQ2epDzlR
OgEkCVxUB0PcqxtFgp9J56UxQsNQLEh0zgpWtncCPwycvnmk1hn6hnghWjqrelo/xwLHYdQRPNxX
CMb6gZxHdkI3e75MJPw6uIAKa6pV4eKlv693B2DesEuqQiQqCDZWvmvsXJzTgmjyl9/woo2Nk6b0
7hTn/ccOPfD3DoT0rAjmxVOi6OsioCOAlEd2B4t29vX08flaIAItHsXqqTfZJkqfwXqQqK/1R17t
p5OSjMP8IJtpJjDG2EdiKwyTgNUJ4jb1pMoaGXJ15K6ZOExDf+o08etsMDBpJr5KqCJnGWQnDuwq
a0ZNIZ4GC4meWx35Oaze4CEcT0fWTNurKKsEXdjEFAbLF5AdEdUzjNkVdP7//m19dgwWFkUQUa40
KYhlszVkh3ASvqwLr6ZXyxvKQvf7wQsEBoQec26jyDfnTDuwYe5Lu8gtMC2wcM964SyDFDC6incO
LhqwNNY5od85WUkajJ/VK4+KYIuqVLs66086kSYL3viyRGqWLg2XvqpUb83WY/1Uy1WFDPEpGmtk
WBlQnDdYxujVGTbi41Iwgn6FapHE5ItckMATkXfPI4SAM7Dqq1LH0De7hGMJJh3aNNp/Jfo3Xhba
gfsAe2GrxniqGR2WDXd/v/OefunBgnYJBoSIY3YsgEw5J3qro+4z8FuYHmjtPIqH/Fh08JKbBVYP
3s+RxrSTFVoN2Ud1ZUq7len5zf4sfEnLrWIOn2Vh0W6xqbEhfXLjDruNhfWOyjjzB/EymDuP90uy
1wzK1ZYMLlOyifsg7eLY7+mztDMu3VOpcmSZKusgeYurOzM2YM4OPaCdwuzSIMyrzNGiuXiKP9O7
vn4rN/XZRIZPwwxfJYlmEM3c9CtTcZDiRh4+NJ/Tjp2kFq7yVc2GuAH90TJpSocnZPHKGY5AQke9
82LAXZIPEKvFzW+fG9Xr18u6yK41DKBjzu0JFlXcqahxjiU0sGaD1lZBdVVBUCU23ZnfNE7IDpAU
z9yFlkdkTZN8vAx2uZSBRcxj4FUqGFhIQ2GDr0q6jIRXoGlpZJXa3J9OXRedVZMkpLjr2mpTdhd/
G9UvN367c9BNDp1kkSDDtbGbZLanwjPUyframi+vrgiZTSugvkAZ/fN0b0/Hw68/NQ3owQRiU2Kc
Wlp42lbg+OXbh4GbrNMSm9O37aCl1GCdTVnVbpJsD+SVKKztTZOKrYV0dT4dQem9k16FoHk+anId
TNC6BlkNf2ZjVo5uv19ofdLOiClxzdq7yXcg1BNOLA/cvHm1e2wWzX4vcv57baa5ZbSisIosTKL1
e+T7jMePa1fbV/WsAkmlUi9hly8+5MTBr6KWNw7QsHdyBgW8Zt4EhB2WFYNyuCL8emdW9l9FCrKT
ZvhSmGRIlt3x2by/fn1K08xvVLZp6broiC5wOs4Xkm/FDhs5qz3jjBGOgJhrvuJjwWe4Y3BlUm7D
oF7glK/P0Ux9uX3oi/goGQbdWOhFekA/ERxyd74TTFef0qGiPWrIfvvmSFskOn03FNWZ4qjEws7g
lR7IMmAwqCRzVCfDNr3M62IInvhQvzPvVI/PZhWWlev00yKJkM9LhP1V6EYX5cuVSqvQZn+b0Vb/
5OJOD0wGSbaVsoWh/iz9oKquwmdDSu2o4XueHW8v20jgmv+7qkbW0AisOxqKOVspyCgJZ0yGRZ0y
R2TDmTuOeiO1p72Y7BxZrtSsLkzmlXBRmHpT9oyAu5WiINZHt9aqGuHqFSyyrENigPrveqhqdfWv
KBaO6F3RvT1prOBrwOIZ7jVTmR7Al9jOh8VVpEFPpRcZyu4OSbsVP/QL9apFvrlqD+USi4zjcR6p
3Tl3AZNMzRv7ryePDC/VBHVtmobfN9g6oZmnKBSCc4U1QUrG6f+5FPrU/K0Il+lUfJYRzdYzaDUj
4priGmB2Nh+5LwKmphSFPZR3oyziZ4Z6NrWnfz9zHZSB4Wgw/fNenRnUdjEzDNjWSAP4I7ovTG/7
nZI58lszfBc44NjMLqE1YoaPP4ymMfIeH/RLYfQt98Uh8AkFGrkJxLISii3WvGqHAsJWrfOiJ0k8
oMQnjbIeNKMaOckhjFKtt/JPspiNbpQAXetycgGfKYV6Qt7kXn2eZtsy+SZyD3UyJ9axN9LKVfN7
MQ1QkFscVMzoLwcM3eZwaauawFLJIPQnpI9zdXeAq0QpzZwdR2p4w3FqItHithSU7q3mTlZmOIzQ
xabpHY4oSybbqLR9kzSYkOFYX1fp71NChmuZd2ClzLipKhdZIwI+jCs5pAKBv7uXI7XE50Qm7zbc
MMkjYYD5YYcdFolp08LHLFQcBdvveYla10afO3Nxa0KY+SkN7aJVd/pNXnGbT2GI/GMPXRyZ36vd
tzAO/zl7dFEgGU78ultWxttNYHCpzYmMHt0MArp0XfLfMR3Qk+OFTQUU2sNt/qq2T6Om4jhqkxqa
SgU3WebMHK3NfgQvDEnsIMOEBGGdvuGJ6GCf+S8mfcNFxebLMqLXt/m4AARuT7AXyc5OZgprmTay
j8kRsS13T4UoCmV6XC00mgq0xrjnZpSW5MpPKx/HyTUByf7VVBCvVHBf56Jbr/W1A2xDrtSuiMzK
Wpq7OmjbscZjQirMR9YTe5vEJ7UsI2Sguit3ZmrGJCweZ8vDT9rFs7KyNA1jYf4IiO+vifEc/DUz
nJto1/qHBIbkh4lQN9JxREIowoVgmMsOm6qrqPFSWQLCgs1jFCs7i6JrT5/J8ITCAYDwKMojdCvr
9/2YCcBqqdAJ9PN0JGb2zB2gprPyMxGi+4dCHiA2D9dBYRWKxMpCilGwpQJ6YCGHBl5V+O/WD72F
p9aXsi5dnGS9eVAna/yM3vyYOxP8Tw7V+sdagXZWi6eUxLx7yBzFS0jLSX6uJlRmd/dvRvb0GmX+
UTulRRgvk257aGEcKzcwBJNZORvbFCiXbPzq5/Gqpm6YgkqPmJN+GuhOQzdSjFR4kgc0x7kS86N0
PDqCHsy7w2rAWTkv2TmhJSwoom65TFEo5viYqWpVk/Eev9gcQQP6F16Yf9EebpJaOkbCxfuabxNO
Q9fFmRnxuU362y8dsuIG4ZT6a4SJ1KSU2aqqqGNbNBYt+D9JgAs6ifd9+uh8KZqMHi6hfyZPd8UW
EzIq44NF3KGGm/6yo0SSlZsdDNrQO4NN9QdHHLwQKvMPNl2ARjoPzftcsOwxtHnce5uZ7bRgsIDk
tACi9DQrY99ZgTynv+DgsTcpl59kf/qniGkZ0TdOkYud6qfTKDQkgc19W7k9HzzJ8AK2ZHLiqaFw
oHySuOCRC9J4A0nqEFJh6n8aOquS7MwNNGnH/wDXQ1GKPMBiuN+78xI/417hv4WTS1aaYnltxlFN
xpi2Qb3+fwZxY3ZbWFKwbdWDdp6reK0tZxhujiclHRE1bWijAnOcJdzkJSFBDMPGJCKoKnX9RkC6
HPp2bmPrvBs9x4SYmEztGLCaGYur1Fc55be4m6ZqGZGR9UcN0/5bUOdBzr92bhY/6u/B49ZQ4BT9
egwITW61zwe+jhAIXmI1u9N4sHyL6OD0WoOwdGT5Wvd73IdoS2Izgqke7p8KSt8775xm6sLy05kS
5sl9Ja36Pj6k9TyFD40Ov89JwvTVi1uukFqkql3QHuFob5T2Vjer2r/VY2VQOY+Q5jb7+BpE+Cw9
I8jPob6SeRD6lJ9UhncSEzuHSxjSaxEZmwHVCrv7lv9WzgqLonCBmhlbBL6ElQiAGnF9shMcbu6m
/xAbw/obSGdQBoKbqRdvahqZ8ffvYkAyFGsh7CWSU7Qh9Iw9dd3q48eSNWmyC1Snt3oVgyGeRY5m
0AX0vrg+Br7B4SlkMBFKB4OOWjD1B8adbZx6x/0wCGsrvYd4PCegipX5eAZMSuNbXq8EXoNlwq5U
BjPWkVUwzXIoUFu2Otffp0enTKh8YG2+UaAAG2H7vWQ8Hf35Ku12YB3TypIjNfSgWNDC7C87KchV
HpVlBX49AN1WqsjW3JTl9WEGXWIKZKmIsL/jUOOAjO5V/MECimXlZzvnL+Yj1BtQqlhh4bwsIlVD
D2QEMGi2pUn+/WP3D4sP1aeltIspUR12vjJpTW82JjsljMrDnCQorPH73k8ThFqkzJYSg0QZEIRs
U/DnIGFvAUtx3p3X8HxQdAUN1/+6bzvE03joBt2eGNFOCMaG3LYk/Ru8/rVn0Co28m0/s4ewIexI
j+6jCGvMAVFyWCW8g+bbidxmpJwey4tkkp+5Rdoj6BNC8zFQZcsnsUw+zIC5Yp8L4XtC7PNAisqO
Kzpy5j5j/pFJ12puL4ZqrXry5Tq9SqB094ugVjUA3hYEUSBNOV89KS2Bpd3WlyPIVnW6urSPoIUi
Tf/RXhYzhl1IMANlANauw34MZ8Rp7VMSLiPtoeRMVC9UPXUd22iYN/BvMZdSPo/83XDAXe9pOVnE
708are+Htp3UWPSvH6w40kfAVoIzSMdlavs9fe8oC7FkMs5SOgrlJGUZ93p30ejYG0gB76L50Yrk
Xq1A4QQniXW/kFGbEoEh43uGZxqwgwNuYJRXod8BRJVN5ZWUHBK4GI3Z4TBHb02qEYdfX7F7SX7a
XG2Pe1jFkMzyFIYfU/zTeCdOsVeGJCuAvCKXXSNNfhFHYghfrFYVBtXdzF3C6gnNyxIqOpi2f46c
6bspH7hH/wr9JsQinlPP9DmUUiWaCZ+EbdBqyieM0jSpOcD1RcPMhm9C0hdAgLfytOQxUMr6dByW
xEuCQPVMTXwD318eNKGHXbWlCgywnYGey3TizKgBlFeBpCKOsZba+WBLSSIwER2KFMbYcKilfPh3
zTkMDi5s0HzJe+YpwSln9lWBnkNKOaMv7jAN01RI072gwLd3y6M3ezqgUHU8U4H8E0jT6oUBFMRL
d4TEMmWrV4fm0z3OZRcTFFRumVe6h9iPUBTLNPR+SL4Uym4bh7s9GuVYxB7RayPSvoDtlnUR9tik
G3YVHstHqqgCtKv3hSeXwFmECvTl/0LCHKKaAv7jf7//i9xa6jU9Jm6yggQ89WniMdOIc/aUurcZ
B4Xx7JvyLWfIysxFQ0y7eaW9B3uzOjZ3sTd6TfJM7+fEwMWUUeirKuDfHGoeGkRrkZLWEQCbIO5N
bZiY0rmqGIdnKm/SUf8tg9n8fKf/MkhKE8yFRPp+BKOfePoPExU64RYhusCIh9xpqOlpzzPtc07v
wu4a68LTt3g9K/foUhtpU/ekKtP/X5Pn9/ZPCELyp2CHqWeal344Q1zZJPxU4Q53Wa4Mz4Rt7VUi
koxqEjkLBJ3ztj6VWGxzjmycibpz2XECnfoACXwMkDR3GbYCS2aBxcCOz+ScY5YFwr7eXLwhH8DZ
S/aK2E+jWymTzUk75a7JUGcP4RWSZi5g9CzoPHCESl1Ys5piqzRg+yuTcgtIi4QRmK0ZdgUYcLCw
F2zliFz9fNxtqoirni+vuI1mLhtXyDD28mbhB5HCTRUozN/4KCmGuBr05qdFlofVyjEJWw6tsaNF
IndaQq8KJZwUPtyB1IncYbyIzss62JTxlLClYdeUObPxvvqjyk30g9F4Ogi+c0aExkzQiMKsLWjv
q4EObCi8ne5BFcG+xUajUjEarZDLaRR6/IIanPt9PVYbsk6zq+jCR3QT/kGzoqD8NNADlePJ+9ac
ECXJ1FuoZBs/vjP1LNeJWTFMEjvgIRSVF/9jVWR2IhiUulXXAXBatZM1dJuzYqF74eDCg1b1tW20
Ke3KcAKdiM7RUs97LMTO2lolYGLkCuM3nOsAkSU86TE8DhZDm7I38J4UjgSAA6G20iO+0XI3Cj0b
/+Jfzu2BWxNsAI5H/43tosQ/PXXRSS+LLL+CfSSt2kayQiXsK9X/TCD6ozS9qvsdQ7+rj1MZ9dYP
wZPADnZBl24Z3BhOKJ+sFPZ+WnXtV1gFvOZaJmF3C7A914uAK9H03ZeXUZC5kl8OnUoXhSAxUYTm
a6qnsbfzoaMhC4AkaGuWzHPRGuhRWPPqYDJHhYKLm47HAyFMTti7gmlXjedix+A5YWF38iY3ZHs3
GWjD/Wp5W0//KbG0FqDAaJqmu+pf5J8Js35/IHvgB1V3RujC3E5RKQHMUrEosAF8VHFwy9YL6vvo
3IubHZApSskP9tbP04x8Hf1N0rVO12rHQkJU7OcpyuqbsxjB5GEWcQbzbQbOpM3uyagy9uXNBQ54
ZZ5uMC5bH8xcn+B2vymhuhKZIC3D1//oWOfwcPdLOtchpzeX4KmnLpgD4zq/cQtJJJ9rbQdZph4g
TkpRVErOjP0HiWjtAAZ6XxD4IA/fyOlN0Nc7ec6jprbP+eZItepqKxRlcCZ+TI1Qb9eeYXIWB3NH
UdfrZQzwRfVfW8XFwLmzn/cTai9cqrYVm2hs75QdDjTg2riljCU/Lcf/+DgSh+OUYGreLJM0fJ+t
G7Ev+JuwzCiJVDgJUa2xJpzMz4k1WdSJ6DbvazIkE56KEjuVuSZMxqDmJrjCK3hZ9oMwnkkxevQL
p69LefRiCCeQdHJ/3z5ULIKX6uGRcHpAVwb2Zw2LzF9ZUUg499h8XQKTMbrHNQs1AMHctbnaykuU
hW24KAj+myfsPxvB/RJlSdGZvza2DzD054VvqbPpzDvRVka3euUXUhjCy4Dzfgf3naku2qgPkNfA
ZFWbNZHoyXSFvEJBOP8u0k+nxfdK/ogfTb9m6l5CxGMoJU7G7inBzpWcCru2RgVQ0YYB6pIyPTUY
LUbF3dVmboRU3mGllRhW2YH5U6e9cIoWvN1xkt9KzHOTXvnJvOVLFDoUGM5kjMt6v7wJFLZ/gWAR
xC+17zQZL8LHMcinkKnKZNy3SFgsRqWRyont8t500SuLQaycj9Ega9o1709oqOj9j4/4tC9LVoRc
SjKEUH/hFCyRn8lUs/fRej5SLy+aouZFPBiTuxPJDVjZWC/+brE+HRPTVCUrLPYKhT7orxwzI9pP
kdwBdNaaZAARqfVet0B/g4cwVMB5/NbcN9aq+qTwI5hNKr/JUXZa1syka4/rEJxkgA8kICjqKW7T
mDf458NJQTG/cgnQfloayaJM89y3rApTWaPLSgYhygItyF6+jNdWLnJRzALc8kpvDn6iBXMzAos0
UXBxxWNRfQ0C6GDpeuG6+E3d6/u03K8kCkky3iVemtEiZ1XkicZx9OonKzik5p6ne2r3TIPyMfV4
b7vVi7/1KR3s0pmB/y6UxGf32gw6FhbFqdyiUx4wVTkSx6QiRdP98rbb1/MtpmzBMkrAjITLcSaV
iUoD2LidfYR2z40YiwetQJEdSLFpblUxRLdpMrRe06b3ZfpLZ7FoHSC+4gXyBVjHbgHb3z35sV2h
2fTvW9+gRtzo+FDEIlQHGHDcEnEe5kzOc5X9lMnYHKxE5oeDp1d+Ovj2aTFiIMwvnSxJOUSdya8C
0O3ZZJIMfopQUHWl4n/n5aIm7uQC2fMsWVOD9WuKWkhspKVOH3mYB5+GC0ZbIMSltaZuRjFwYfJ0
8OPEGXkGjwPOxirr42uzmBptpYoZVK/ZcTv9HQ8/vlXmIk7Lq/9uzpI62wjNtDJQDaxrNPowogT7
Lu2cO4NOFmBXpY+sD+oeSzRAThmjKrOEmagVXjFSIEZdOFQkpYQUllipUb2x5MnEjk/AjB7Kl8g7
ywJE/qIkAFtev/wZuj3JktXu87v1ErMEVpxwFZu2MJM/Y6u0ytWCb/N1B1cxi1+seJTPRUfKOg8F
WOmZ32sd/AOao3pEETYP/nbusrSBtGUljO1MopIdEAK5RHhuYhq7xCa9nklyIhAvWorXj0f4JmG3
UyI3tB0/oh5yH6HMDs9mJamrD8exo/Ch4eplOI6QdxGkhIxxmt1jZUcmPDZSL+h8uk4OkVMbwu2N
OFGqeaxUdotA8JfVBsIXyTMD9im0+tBl7wx7b9wgsakDpi1fltc8VUHp2CBucLaAPGD4L64HStFs
adSn+kZ1qgn2OaFApX8s6ERqW8xv8YvYafiwMfs6epQLuqhaYYfqtZjgRNSJrqj3mCGl2j0B8qXv
0LetJZaE5aSnAJtF2pw9qmSUT9qCLyCAZm4+G2XT7znWYb0oGd22Yr+IZ8sEcV3uDMitgfaxy9m0
zhRuncvSj5ZXah588F2LNfswvCOwZtP1FpKErac8VHd1zSMUvXU34ipJggIbK5PhfuUWhRj6t+av
gKLDMeR5whqHUQGiO3vZADFNFDMUgSuFhIVM7m07n+kU1RTeC2gll4VqgPmdJ5Mcn/lIvdPFPKlM
LhZpps8+Afo8bmXMq0Q77U3p2ZzAMK0IF097tU8hkK9MHd+x5WQ62GXpowlmPe0Vx8t1ZyLL4zEg
bW2Ak5VGvNP2/P/7xwoFaIwfdSfr46w/CZ4ZngiRoLfs/pWGWHJ3x/fHDCU+FS/bOkcP+JtA2Erz
wcRDtBnVARroKgCTzIByhy6U+4SoXlcAhKSFj3WjPNu5RZDIG5f2+6Z2g9uVMxZa4yUAZzIvhoEd
OgNLC2U1mzjBC3hpFz+NJKeGV+tkWzQr+1LA2O2doKtSWPCnK+E5ubsDh7J9SyNSd9qNoq1rsgbl
JqwHzbFdKukmEch5n/SIg0xmoNRfIUlUmdfEo5cCQanRY8+Knrru3wfuIRAnFbjNo6Iy7iY8fKio
XzeYi41gpQaoPgdOaMJstBv8MXDwVQ9KJBtsmDFUTcBJYWlwtFumRjfMc6JYCBDRxLOW7FZ9ltSK
H6lX7OtGyeBK6EdzUWzUUt/3LvPq0qE981p19mLxMjoGcFJtygI6wJ0SUV+DQRvBws+yxCbc2q0t
3MUvXU66k1ENF5yanED6BbBSml3MZyOg8Cqfq1aphtKrxuOgNfhpmPzuVrzueCgEzyHy8kg5eng9
ZO96BUlhis9ULdvCjfMHLPQ/K/B79SWU98+iWZwpIXCEoHh6Odp3nkC8b1Vbc2CUeqf5M3qQs3tc
K98ikpVJda5zjeSeXDQVdVMMDnQ7E5Mc/JeLlf/HGZEdwsEkB1zl+bPlxpvlJryYNNY6sewsw4no
qkvfCVQGaasct4rj5hRaZJbOuGk98sss8tgLkyszblnhT0yBx7e2ZSOiS7VA8/RDxv+hfzysR+/+
CO5dcw/db4irkN3d6y+OU4PoNO6eRY7pF75JzGPjXa0dOIDCiIAUGbbUWmcuFMrOPII/Ca2D7G0U
DyTlam8mJ46c9QiXb8zU+Wf8bg6186XwByej5xIF+OsI8Z2cyLpQHEuZwvrLRq83FIgVZxLGaPpJ
Jlnv7qHghHYYOaivOtaf2hLo4HgeLj2uQpkxciQ6fVDWjB3c+J3Vu7RD6l9XT1NAxp8Z8r6yLGy/
K8CkOL6uLBB0P4DAJKTZyLF29FOMKG+nkAT7cm4vlprOlJPnJ4dVUvdu0ZtnHUmePhfUD6bd3M+X
8IhNg5dqbzCf/3TxJ4Nl4zbrvwJqY88EIW74D/vRwYzKHQFIyj33RY0lMjlaYJsZayHee9VzXfNM
FNTbr3o4naGMkiC//jtLxCni6NxQHfu+l5l2/4r0lL2LqjjwXmD3GY5cvNwN5TckfwYaTNCDBnXs
Ysi2ScmANOPAFp18jq9slB01DdJswpr+fi09+osAQcBNdMDHa1i//d/oQglM4jGy3LuOQ9TxLX2N
xNmGGcUmaqa9cN7e/lfODEijNsol9W3diwhrh9B4px6uWvx8wflxk/3K+/lu4Zi9v04G7wXhs4QT
OVqci3/VBxoHdupnanyYsUXKdtMxxeXHWy7PB2scINoXGNIx01xohIlvTK6vhbA1ECqVF4eB1MYs
izDQIdXPooHjmuPXfr82PrQZnRA0f8iSceXvmZQUq3da+VZhjI8MfPTqLgBUxUPPhfPLVn+1RBMn
+uUgjPQ51F7GbJa2LUNSeOGUrlYo3NJ51eeumzI/47Nr4mMgt2Wr2n4xSbFcavCGH2SWa6hrOIc3
SCJCvBxjcRIvIMwf/HbjimPIffUVdcZuKM2erCz6BOFQ71j7OFbDOA9Luoefj9S/EmrV9YdxWZHu
Nl2b9zJoE+ek8btW94WIuUapCPn5pNYS8PayEjfCt5lBMnC38sYjmjKoedMUeMmB9tk5f7i+si06
21DqBHvXQ6rpHa06FHHhvCXXdDUL2rixpmmd3e3JQA1xxsoPCAnKqwPwru37upikDkzklICn9kk0
SGwHcVnUKqmN4gnsRRhJX0+uXn39au2O6f+gXvUic/AcN9nP6NI5YSq0KTq+en2kTI0vDWeLEJrp
niUdfWyZjJaw5O9D9WwZwqkKy6W70fQhpqTIVJijgpCnpYVqdtCtbdBml5wYbcFyq77HceaDxN0A
zTDdVMh/iC4PEff/eQi5VbgSfvTCr53oEr4Y/HaF4rtG3g19/8huRhn3bcpm9KTPvQabKTihepIp
9ORHR1I3C1Id1wOVTjtgmRf8iR0bFySudCAZMbJlqcEbIzanYrWTn+Dzz/vQlGC54740cKiwfJdH
xiUHkxbGXR+x/Wlguh9T4Um0gJngtsFsDc4y2ClOyGe9HGIqFICV0Ei/kel9cnoiClRmlRyK+7Ly
ZF5K/Lt8/BHRhxtQUnDN2/NkLSA5CmNAONLp2bgJ26GwOK4Mi/+dXFd4ZoxHWahBCLP/qhDOdoXc
fpbLG7lpHrpK1bwu0kqfICoRReFPyIbm9avgriZ8MlCIAM99MXU6Nvb3rY0E96hRxTVjttdDaQYI
XCmScmvo7MX10AyKZQeTDW8SI87k19kK2u+Rnm5kPZZSZOelJy+NApJ0Xz5qk5Ku5I2uQCFZHPks
Emi9TLhaCWoGzT0++MG1K6sqYHezWApHm/JZWDhNAGTqrg+n0R3jPASEyHIkwCVvU13K0MtUKlsD
6DxkhtsDfsQ6kz+YHa5f8qGH+xkvrwjGUpgojfenc9xKOgwOHCzoM7mrAj9ZSuwxn21n0dBBjZAg
pA7b/ser8WIEMxi13bFzdzRBwkW6D9n3RQsZbJamm5uss775AhdBL3iPtTIEgY2vrYyigl9MWXx2
hyLd5xza9K3rkt8XNTAHZVAKL2QqndTEVkaSvSHgC2rT7oTF+DDPAAfcHFGy4faeLjrh6URmP0sQ
UGQx9mjE2tEPxwp8FV5nNEuxfprbMWQ4MLd6qkXzVQKYJvWdhzRg/FamVSNzrWxwJNgrcDhKhVzZ
11DIRhd4HRo4jfHkjzxmOQ/omkvgwXOttuHD8VELD/u/+zRIE2tqu/fa3o2Vno+0J7r+COBhB8PX
W3KNyB3+hmbagJMPxkXAC8dYMbx6B0QbvXGOEdq2XDzzl/gn9nwUqkIz+bX3m6zntBE43ji9MpVT
wV4k59QLzIU4ZPvRmkgRcA1H3IWbt68+7EgOK1OdkKRvHr9bsk4ht+Kmtdu90jJDGCNlSPsdX3iF
91q6a/Q58Srt/6ud6jvqLfbgpIA4EGkm0Y1CPoUNaXdsiFlbgdW5ssnqnadJIjxYu8/KHTXAnz9B
4YvS88vIGFefVkGYHgzBa97Dn+79ikG9NaqxAHaO8lMliyQWYR7tbWOilyf4sfNSUYa3n1mWYeKu
zbjlroG8jUdoHDkC3qVXMnSdMqoZqhEGKerQiXy7NyntkQElB203gfWkiKLq3OjwL+g9fA/oTwRg
mu9O51aCP6/2DDtRZLBr
`protect end_protected

