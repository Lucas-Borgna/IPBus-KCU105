`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SIpkYaJTZYuNRkk7P3FfZD3OEpyZbE8fXGxbM+d4C+oFzFHvnVq79GWar7FoKC6KRTRlo20wYhWw
jHt73De9Yg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
JakrkTjyUvpkepS3bNfAgnpvIJtFNdZf0l+qcBqQFvZA83VO2zLpNUzflXWn3dZ5RPdYc+GRodF4
PiZHiw7jbIWfiZvnVWJ+lZoof4urpjFuM9s9QGf8Fi7ZB2KxZy1I4tYYydn4FwiwXsj3ZfN53dLd
R1AuthRiifxTJ/jLXFo=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AQDVG2udr6kLYGWeIxLdV9AFdf55PTQUo7+oOMmD3oLbRhMfs1x/SPl0/XHXeecevCqnFWGbg739
VLuIbsD0S/K9w6VjvAuzDmBStmZkUo285UfRSok/+mfIiDvkA22M94LPygCdIdhlYTtEErgkSy0J
FxIVp5KcLVM3wjOanZfTX75dPQY0y2jKEoaOdt6RwIBkgJCg+9WSp0ZqqgSQsZdWAr59o060506Q
gcFwxh2mRbcgIgp4Y+x0YVotOI69Nyn7B/xsAfgXqgLR+LjHzl9sAfyiOGRfmXatcIS7OmNtrUfQ
Q5o9phH7HWW7GpjRnJKUBqmz8Tay7zKEhGOhKA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
daJdBBgJZ0Rlo3Jcmb0IcntCNF1DIB1jcoPulTCvxyFAFygegQFpyS6KarpXlTGBRrFRLiyMBMap
9S8ixR8a5Tl8tBsVDpOmSYnXLckto1HJex4ywkf5KIV5jDy95F1gvPJYet7IWpEV3xOSC1+SWDxc
Xzdn6HpcieSTkY7plXQVDzAr5ZJayfLIXDFv928/cYuQ7skpSghQIF1zpkGFpTXuWkoHq3ysbwRx
ZMpFkwLng8nHfpGZmPa7KDuCcJbXCf1E6kDMe+slPy5DviCo0HDzHqsYWuh5gUzjjzBNuMUwEKrc
LI2FHL0UoC4hj+3J22sQ3h0pcTxYWv0AyT6gOQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wa4klz/fsdmFCoP5E6c9CFladQQa+iMTS9sC8NSW7yJuBM3mdvFDFyefGP/iZLevm+IyNGn5fdUm
a59iEPEmBXkHzhV3yrxpx8Eos8xsT6w1oMIvGeiPUhuENIGQO+4MlkwtKZ7m5AC0RsvNcl/wQIBy
TWzsENX6wi98E2WzrelnparoxovdaoZHpPNVBl+hn1eqtr81FAQ6USguWNtz+MnXrJxroLVs/KX5
d15z5cqbk5jSuQJIi1tynwN4znBepJBTCSw9itkB9aw8D7K2nHPdDl2xGdOOAYROWanGbgMqRcye
g/T6cfmviR/Q2M7lkf23u9Vvkfd1RTP5AEAyGg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Wv+z04GW1y++JgPWgQxLk9+Ox9RU4u9nQV+lZjLjvfzcgrxd/TrU+vvDZlMLLXKBoaBc9oGwuP20
45Js9Mc3bB2RUL6zdvuDKHuP127/6pHE9neX9fvq2t+8TXQ4aSYRYFJIo/UrKHq8lSxDkYeJcD6O
wBpIBISZ2Mmw7BZChRk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O2H0B7Q1U/tX6c9BUn55xVnNoH+BecEM8LP0tgY6eoWdB+MScKNT5VttBIwK/eQd4NIa14cS1TwP
q50cCOUfkgkVa4DpYF+TCeLOK+K7M/3agp5leqbAHRgHcH6gM7shJ2QPOV7isdvyg/k7AaawJwUg
+pPFR71SuLE3FstS/B0ovlSZBr5+SbGN7yduezORDr+ZyBZqvR2++5gkAWfOBFM3n3cNuIZP8d56
3XR9frJl/GJU5gMNErRQFcmKo7YggNnJtztaGMluz3ZVQ9lM5KHh7ob3wutRpD7b5FtH+g1cUGH/
OZ93oAl2jJPN9zOLYkPV/M7KBJv1mvK1DKT/aA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 807360)
`protect data_block
8u42GVHWvtWaLmIN7Bb8QbxY83vG6oryPDv1dmRNz6K+TFvPvfNW/Y1TlK11+2mk7vESyrHwKdv/
gkVxhnfkMUlOeVPt3Li1KXJH0n5004rjszhbNcSZ+7kDc55UZbECcaUQaaWrYk436vqB14mmJD61
M/8vmpkR+Zk2XYDiL9JGkw1Go+D8gPcXVjJmzNHv6pXa6+/dcslCt+XsotoCdXQ0PD9QugvfRfN5
2nRhOho6JC8staMMA83tZkNJqoL8ZZptBFccmrNHoRruJNdm6ZJluBayTw+ULSpMA1VEQ7Uzf9BV
6avZCu+ZR2IhC9rZz0i+j5qCfdrNrie/sTXIeVgJA3qB4yeQqsWcpWmg0CWfT4pMaQCHUHnTXC8w
pnvmrdaC9RhMzqQrUbYHSmJUsR78s/59sBU/NXeNaqFX/reM9MunKwl6AbCvmQb46vildPr+MdG/
1TRDtk0Ye1CwYDZdaF3h4Mc8f84242J8SxluXtuooeIX7WVh6K3wCXjN60sTGCPOXsCmZtzohAjA
yjDgtCzYXJXyPWpwwvTvts6DcEVOWLccX68AwvhJh3lAQe0v9QshuZFhUugA9gNMf9TsStk9gAS4
WbkdU9acrjU/W2ycso9AwcCIxJMQgxVwudgAhMe8OFyEvuNH3k6VAiAOlVa3JW0lMuJpUp9uHn5M
PmW0x9km2vjOq4d/vtdr4AX1hS6/eV65dN1Mkby1qKkiwCSd2ivPRTAZYT6orc+36RTlM64EWCvb
nH6AIgLYnyDrUQWC4jBj2ChSJ5CGXo8Pi63VXI89YK35n7jjUyHgwoMWn1m3oA7+72g6M4M4RAhf
yxg7D0qDetKrKPobBbebiIAiwItPzreMYL6zZK5S0eNCj1uGGdyytYy3NpvVOqWVhE1alkDfpNXq
cGnJT+k7tPouQmkQVaLfdIheLUkWn4sD/q9PwQ5W0EEqwc38246Z1BzSU7jdFGYpEDiyIcgWpoM8
/48b7YqFJ6ri+ZORchuvzK4hLyCiJ+R07CxNGqwFi5SOnmg9Y2kskUnmbcoT5auh3q+pbqKPFnAa
YZyshXr8rxlZV6OK/C9Jhx/fUl4IdnAgB9wJNZ7hUsqlTUlCjPAPbUK2ZVCPUz6OKn9dXw2OeD1W
3P0QKE+jhmoQIwgQM+wQow33t21LVO5590CcKAVoqGYmbk6w83kPVyX8OXsUEbYm38lEMHQgAC8L
YcG5+L6IaFgqxH9p2GOZYN2blcEK/LYjjYBx8EuR0O7vVvujIymUma1nRg4mimw/667sqqWRBEEm
Fu2ZfOe5dFzukOtnvKhSSv7ygaV8DjT9XAmqKKUmjAkLMDU+LtJiIRXxPey6zUDTV9WHhs7O5HxH
eX810R1l4mvZ1PzwyNsmldTJOG0FsQYs5ZJFlzGF4Ybgy4vgXcFjN28tpvA36RaOn3cnfWgq/DmM
ehj6jSBEKnx4C4/uVGEB//ALBOR5+ppetyvoRnL2Gf7UtC8qtoXHCqNCUKNp+C4949dKLLEs9i0a
sktI2UDay/eqbqLTrKppVEgzq7raBl87x95g34zMqQpxydzBq56p2lZNGf+nBpsowFsNxNJ6iplI
YF6PP/V+pnNGo3/0C/NvU2RQk+vRQ9fl6k03sI8H7S+phYlrrBGqLGLw9Zq5XVzzubHJH8dK20VC
OcDuL5sJ0Qi1/PI92ky65XU28ygtl1hzGYL1DfjLh/5LRmwHbXfzzQkd75AfUdUskjhSZnFohmLv
bI9S73h7+IlFWmv6Q9veR6RExiUQ2Ktd5OK12sdVBy7QDm8nXyr/0R9JfSw/GJqLARqUp8i8oSKn
JfiFCB0vPC78yScLn8um5r45+vD3IHJh41Vuelakh4bhmCGGY1H+1tu37s+G4cXabGTQFv851tp1
CE5Ak+Lvq5iGgXQB2KW1E7z7zBWgGYh27bXkuYY9OAMJbGZyGcgpzxSX3gBLtR2OL3P3vOEOrJ6m
mxf5fmprPI+k3tuC1fUUFK77PFdkyVME4XuUHKS/GMi9gc8N4kYE6AhGVWLCqiSbJAalveUQUOlK
J+ZrMNBp7ltXVYT4uCTbVQZkPg1RzEYmc6oA8r1KEh/p8CRo6PSvOLUG0W09Gror5/LU+Bpyh3Wq
0xTiEK5n4WKMJJnlExNvpji+XI8THY1vt/nJ4cO3J5GLCLVJ3I2XHUe9waG2u7icP//xv4+anZAn
CQG+pa1lLn9WI9HYHA20SfgatUHBYXwn+MGutNEfqr3DTgjh0+JvWRKCnzXPXcPLXACizWKtlS7B
7z3CeoQlV6Q+02EDdpR+4nFl3qMDXfwRShLtA0zDTPEBIkQg6x2zIFeqZg0q5B937RmL/F80Jhfx
EgGgBy1md4gxcZUPtty4SJM6YQZl3izZu9jsnqqCbdSIvmpx5tOiktL0FRbU5ZBEEj1cfD6rpBIF
C5otPp++oSs+QHaUxB64964diNbBSOIhWVVDq7YHv7S6ueYVqkTAOnY2Ls12zArhqwf1fIWARIcB
HiYN8qtPvwHaJtMXEZN3XrD0E1O6/4UfXkd6Iap5z+37gGrqKntEgEWtM0/s9VZDjkQm+8KZrL4W
pVi9p63G4+xrmCpv+c2rvN13+cHEs09CtWm4MhLObhzvuIje9C4TixYrjPc5uWjQ4JK05rdnupmE
BC7ost+34/aH3XtD/Z9XVFNFKaG3M24fqXS+V7zjFVdQctGXb0S/rPmlhgqIurKPoI2z87kzvcRO
2S4W1642XBVNmxRPePW4HgpR04M+JrVJMudf40YLvvt8opAtYwNlic+8DaIe20ilW2ypaHDDj2TK
9QrGDrymfz76JkMjFPGPo0NX/mWSZNVKdMLAMkMMhjCsgMfHeNAzTfiSouz8QFftTvTTF9vJR5/4
3q+Dh/2mwzx1jVC3xGei55H2M61tndSfYwImVETTa2OZwV0aGQemUU9Ze/u3SiXpLLw87i45Tlbm
FA1s0S27qhn5E1PRFOuipIfLieDbJ0en1zqRYhXuXTdOs3Y97lSMAAKwPICsjpOYVwzXqab3csdJ
rxq5UzoF3sJTL7IoXgyXF6/FXS3t3diWmuFvjYToSMvSgPYITWAZOsIGo0haM33N0Wh8XQhEaeOW
+cmFSzFYTNwXQKtU4TKDlYjRE3+yh9uSv+PuC1GvNm1MQnOV7ZSzIB52yFGfbpg7fmLIzpeVXHZ8
e2HmFCPYn4VhHYMRERbIVoyche5K+a8Zs7UyrBt0ecDkMuxmLfv47YIGaGfNZ+VH0ODp1BNLQb+f
J8rqqjWS41msGeWRdG0WZ+NXuUueIeLad/hFu6HKLhq7NtmQniyQDLM44KuvY5xrG8IsK7cd0l1q
TvVwPLocmaGB6nk3qqAK4c5l7oR4GZS3xZxBO8osMWiuNoyQOnugp8WCU9WcB1eibDpfwVoHsRSh
5igMedyEUheobyTTtTh3VgvBhdkALJqWI+TBU50jxNOP2qOkxcyPymBv/thAjVrlmfkBApZAV2lH
XSPl+xR0YLCX8ZKow/Wi9IS7up6lYJJTfV9XoLCYLK+SrBxqQd9lpy1YA8bOAGNPxufLpw1E33ox
bE0Yz7G4qGphdFY8ksRy/Pa3LpAJ4UDU//xxG/MRG1TLYSRYEJd93grAxfKaL5oCacSZPuTUWCjC
gnH+nUSvF65u5T8zPAsnuYoujYsdLDfHSPloKoF9MhcQzfQnFo1bn7FJtdNhyaa7x54+QcoWGARO
3oPIMKc3j5NdNhLh68764EHnOvH8znYSl58grTyJTFix7xG6QXjFAxc3mOvunzO/tPbPxJdc1rBo
B2X2ULmaWcYXsR4SWbPiPmuPPvZl0j47Jij6SpmLw5Uv0hfwASOq+mPxJOKD8H7Prg8y1KdqqDt2
RUUpN9Cb4Ue5T0G7k2XDBZkNmdq1+kRqxb77/D70fWIHswQ6ORpnHSC7mS/G++OvN9/KyZBUxB99
mz+aJhIvNuY2+18wN9CgeFDAm7E2j43QoPXqhr33Fiz8Fv+cXl2JmPyLja8VuvA1kg6RQV8kd8y+
mYTv34b8gD8Cm04tEGkBgok1lzMJbp/zP92W8sjrjSVc8+yzhsBHpFZHYPBk+COj6xK7s1wci3ew
VNba2mWIPKBgSdHt8WVAur+3ozQ3Bh06zp3ajcYMuRg0rZN1Kw6Odq0nVrqlR8zMUUPd2GZ93d0A
QjhulPwJMWs8TYt4w7lo/JsyGJZvqwQR+Mg7nOzIz6sk5EIHVqHpY7y+XNiIDXxSVE9O9F3tu/6q
VtRyCiWm0eukh0vUxB5YL+/ulg1Sv6xKgdkz2o+liyEyiQ+WseWRFfH5YUs+BNPcBSG/pj3y3v2I
BnNGvl2a9xXk1sTSdPjfIH4Fpsrk7YgOBJCmz54u/ndWjWeyxcCn4742iSVt5tdJh/zjqGNR9Ifa
pLdpU44KYxbyxZ1TIIqoKR8Aw3BGYEJTUUYTvrFNOoPiS9qqxtIZHCAKX9DaRFQvit+h51yFmHJS
WAK1VfJdrkBkLeHjYoVb2h3GfOjTiJR9NFH/6xorSnAb58m2Uk550ZznZ741Qb4v5jknNgiEOV/I
c+rklbyV8vqa059LazAFsTYofMSvaphRL8mlsv1qHY7VU/McxqpTejX56Eu/L/S8OqjoXQzMswy+
NK9NIrqUh+BS735utstHHDmvf9BOZoJPOmTpDUBmBp6w4CWTMfaPuyV+djGKSgAA08FvdJTtF/Tk
6/idN3CIvlYqdHgg+YTRERuIMnfaXc1x2qlFYVi+PLH69juHtHMcemQXtDdh6JIoskiu9ePehW0Z
Mr8zm5/hiIype1z6EnqS9XR2N1MYPmtFlCn1G2DLg7lEIhK6PmUEi5+aXf2KO8kOLXGpaJVt2Lr5
rQrtB8h3zkkOsXGFTD3d1bmK5rWB8qJKHP0F/ea3LwljBoAZWGQITe6XydrX2S288vbfkrJtS66G
GzXuPREStt9hBbdoi2JiX83/H95pBHM6Sbsd8Pz0jZsFAwojCZQv5dKZsFuRO+QlzCHISMQYdasg
d6HilUpUlX+EGr9fNTLKwIFBrhHr8tvtZb8tJZ8PyKhT+HxY1gY8k4jkCqwMnyQQjkh8x6YtG92F
E7xA/5Lf8l4svmYxz1AqI8nnIcUWUYrZ3MwBu66dELc8mvYo2bdC0OQrvM+IvoJHZf9w1Jm6bRfK
l/AHay+tBHCrNGypRg07pOwNID8a6XT8/nRedVaUmCl3JiocxTMQShmHEzjHByQsOvAQuMnA6D42
WdtGU8yOFoRZnfFptsJcPTd/oubKOKqPklIk1c9h3TTUEvg5MRiJffrcYjZYyZ0BzLLYdP2w1Ns/
qnjCsj6nhSmHXvxEHOaJdYSjSuSdflDl9xdAyFkGBvkUvTt4CeZA2pSpcVpuIu7UaJFlHK0BljqD
9dNE3E7VNPDEp7W0/cLZ0hJfXSH3eJFvrckvFQELTGkJ+pqTDJWb5yQrV9HdOfVTs2iwywgPIlgw
NSC7ZbpXvFY8rWRDkugOe63V3z2fcv9TP8baEM3+w6kEFu2MIivDys5sNcYL5CNM9IoIhcOU8xCE
ZUSVTAglALUMbWzrXqu2ZaWYSQdOTIz9Rqzn4H2XkkP0bwsbAq/MWsMIN4u1KFbKaEZiIqdyR2Be
XOzYq+O4fX/RpK7ldYoqdmZuwP84HveIVfpbmvDx8ZO/pg2VTgcmplaNeE8yQ5A7/ivyWTt+PVDI
GPAlJQRkPK/SkLImmJAk5LqpDrQtpEbpmkGsF2Q9GEjkDhw7H2sEXQcNuzDqrvSuJv5NZJTlBJDL
h8Xkz4ffZ3s/+euYo+UGAN/Y/7Trzzdp6P72v8X1jec7tjLS2s/350NuOcCa6HKxzAW7BGWrwENr
ehW1/dHbPmchOh3VhqLdLcnB08tVtJNJBdLL60TIOk+8BpwtOikZ6+4y84OkG0shZxxVj3YvPhNi
969qK8EtGjDOSw3fI580rQ0ZU8LXCYcEa9MLP0Hyap1bcffd3wx/+1k7agqe0XXjgjK/60NDXy/9
9IuocuJVeH13xUMHBRPscT3w6FVsi2mpxkmaKD5MaoP7aq8pv+N+BWIiFHeDSZ8FVs6MVTZZF5eT
NBWIWjhheC6BmCpQ2mVT9DJnIxGU3chIkgtyZVIdJjbevhgYaSVx3rjZMkOw+FCgHJuGLTgU1Zg7
xC/YZGk9cEjL00W0Z4e0ad0DLYpVXklzYZ1rP6L48t8R9VT0UiLhse/Vw9ZeNJnL2GXs3Ge1tkjx
s13iSKf8evdzsdfayR7dXvnCOzGnBlBXn3HNLAOOaWJIXIqShcAH+4+HasIzwpTxM3inoHDgA1DD
wYtuhBiivjKiXFOjE9WgbEAOoE+uz7nYMGvN1eEjWBPMiG+aF04RkdCGpxsblu8HLizwO13uwKvt
gIbEddUQBhRH0eRTRumEWrJmLRPW3cxJr3oXgWZ/imH+q8veiuPeVX57uPqq/IWK06ky7I6B0ce7
y0yqHeSd4xCqcF4reD3yPEkqruny5hXOCMf2KMopSBgqKAx9KqlIIZ8Uj2cTX6BrZWU74kme7XXf
j48kAVtVDomkE8L6FIx7trCxtESc+rbU9viStX80pV595wH0Em0qmtW/eGqeZU+V3OImNkHYPgTl
4I8TLJ2Kzx+FNhxl7QMplgB2zydpa/eW36K1DMP24/6OCxdptslvuLY7Fa+ZXCmf0w32VsuutRdw
HT6f18CW5zc1a1xxmKBeAVchRKgDiOTYRPnw/5G1XQPf/vzdkCJEH+ikRi/LFus8aIXB/8kldckd
JAks2PB0S2Vnx6KV3tHLmzMl9JP0YNddBKVbZSdfx2XjlUIF8AQ2nIyICVF0+rj8kLxIWGUyqReK
g2A3YyO+AqWbDsVMyGIJaxeXWIDcrN5n9e7XJEXmERqt6oOiW6/ZQwITnptd7EVUDsLd8sHjt/Wd
P+FPeoqRIybthxvOl36cKX1J/SQVBpFKpMA630C/uzSr3B9Hda1E+M7m2iL/2rJAePTf7ipe7m1j
hHxYkbG8Vs2zmXoIaElV4Q7ZIDC/5KOab14nTEob/0blCkOL7Jrb863XQMrcin76LHX0iWtQb+yo
1eTGL6ZojBsT2Uf00+iN/MdY8T7sV+xJH0mD1chvnxyqgcr2AevbFm2UyZoIW86QBSrgEmfLNnaj
ouHczEf2MtX233qgukSfsUxFG2M8dJgfoVsM87xPkWfnrBAeayca6azAk7VznlRosLmZl6tL2UJV
jEWg7hujrn/5vKa8TZ382Nw3AzL/Xd6umut7T46aBBBXMIPIVOAeDnZAAmmHsiffpuUy9ukkVsyu
yW/gmQLr8bEHuAPLCMxbiNEckKvdkq940JYwajzl5MYwyfdInVBo7uwuALZrEYvhph7/kTVEfxLy
K5D0abB7JqmtZjFrmR70CxgUaB1boiHs+G0oQUETL8I31RDGMJnvmVhmtaxPUEt8hmmq/7koqhty
He/QufIaYzqwW/tL5hk7/OeMY5Ky/KbqSPqVUvEuCm8jkC1m+uIQ2HByfZ07nEOpxIlzNJSvRGTb
LlH9z18DTZ9B1WYsMjLYJ917HNMN0qYZ4Ha3qhSk5yXtQ+ygANzwfC+iBiEYbrWaKvrEHeH15G0+
LK3TF7+mt8uvpyZFFEm/3Lwj+KqVGgI1nzv4f97qDqCBgcCNI2Pm8lHvibPqG9R3328Vn84mJ9E1
dZegAT/jPRSTNA3fBW+1xD5HpZmph+5ZLk5PybBk3uWzkCgM0YQDsmDKUL5Qie/6FOxJ8hlcwLEi
JIOUvo751UWs2j7JoO/4tOiquWT2P2BVSd9iL52J7R++BNiqc3ng1nclpbC6s8Ldn+23HK2TF8lm
KxZ53pTV8VypoHjM5FMtdtMkFDrYJknrvUP8Ush9VWw/ObKewp6iY+WyuoyNlNjph1cFi3b06Yd1
F9YuSORvnuvQZ9RuaErWf5npL1XIXTRN4zeyepjfLB5/651JRIImIPNnMfIwEstjv6Sjaz+wwaCX
9RbZaJ5USFWf4mHQO1vzlUUnSdtTRFIDCPC9H6j6yf+WQtIoYWcz2GQnFjKZUSCl2YsQHMSm8+Kd
AaqlMxdqsca+temhM3jOQPwoLNnC48Gn1HEqaT/CGMZuxto81N3tpvAEdO7DGesfOL6sDk/DxABS
n2IaYxqW24gHoYTozjHh+eHzcFz27MoNBp0rJtipyzNsjfDkaRzSRsiUFDmQ1nenw2PmksZ3VKy7
J9y+ISJS3tviKaNUcGE4QPneqG/A39x13iPh7zC5nVsW6g5CEW9jca8oMBMHo9FRsXtqn5I5O8oB
hgxZXcpFaDivNL/ykl3AeTyiGjzoKnL/b3LGj9IJmeAMwahn31R+Aufp6VF1JFMPXdI/5/pKUKbq
QUbZgC264NLrtEC4KHR5yP7NcJ0KcqxCyADYEaqWnQrmWZxDj6gAJHyMrePmZej1gZWfR3Cslnhr
yVGvpRRM2LwpIEn2QqXr3rd5Ev5HXRgiGc4cG+RF118kpvwemmLjXIcOOlCykny0Vd0SCk2/9H/g
a5NUAK1SxdPNOhFLLTc/UJYZgdmYfFObJN+dy5bPXHnyzqLg8YVFJyhwp47+1zXlQAGFhr/yUO1b
by2rVqrwFvDhL5GnUQ+z0ORcWVGzDFyEVcid1GmzpWvmPmOT539splmAjZs0w0/5ATEuxZXPOc7k
h1PNilZ+6U9P+QPro60rc7ZDqFAGT3axVH34QFtSKJviZWaYVH1kTWNXZhWffRFdBgUX/hth+u7B
TrXk3mVtbM75kA1T5CPLqzgrKsqCFN8CzqjnuQxgj2xOyoQdPbG0Hu4V4DoiQ9ptUKUWVzAxdE64
HjUuiea38m3vrrYdXLwZxPJ3XkVs0kRrXOOI8TSVdRSatHsBZBvluJLBSGSvEgcOFBLUX9m/cNfu
IXAvhrku/YWiMrS6rKoF3Ocqxbkq/HSYZ3Vvcny5V+O3sF14r1d0ceLR5rrUtEX1uZEDon5uIL78
EjjzfJMxcYodoAht1SZqrYkdkuZ1t5uJwUxQeQUfZr1EhlnpmBkzG7mEuUVFfBZcEcGYhlE1R3Ou
Q92mc0dPJTswscYMrjR3xksVCwXqpj52VlFYLasnjJlywsZYyDJDw0lNFIodfPNMQ0gbBu4ODrWh
4gS332dv4ErV3kr2GtB10Hp/mc93q8HGzuanmW76wmRekzSojwFLyyZ8CyZVT8OF8UsQ66Ea3eT8
QKh82kv3cVbDzbi1J+nCvLe8tNvKOeNq6TQNSIKTNHEpnCbHgO3h5Y7TFLrF46V4rZNxU71ggLML
kAz4dakfx9uV7E0gPL+ta1c7yDLB4m2MegA35g2Xt9tjTeSWKoNEyzCPL7LKFJhShc62spZxP40b
oOiUCWrWdMM2iyt7ds5Fle7i9oEbMbC8ZZ4mNhv/wm7ICifUvT59DTwbuUppoIImsAJ0pUuYFDOM
lZ8btJUkTa2p8gyrB0Cxl+ZaY3e+FsZGsxozKDaOvBZD/zHAz+NFwQZ6SmnyUpo0zm7yHCCNA2Jw
Aqy8D3CAQanCyKPO1T+BFkF/WV/rKbeP+JoWrCZLh5lHqjIEo+Ks+aLjGsEN7UagNAITl6qKYRgr
5mmi+w4sj87RgezJe4Fqw1YONJpkjlSUh0D5VLQfADCk+XgIo4G68akMqrYbioJvAgjmE6wcLmku
71S94s/t0EchfqQm0oKZ7gdoqDBMsP+uJ3SKLi4bCCsk2w3FqU81VRGM4UzaF4OdAT2s6v+h2gN8
2fd/7NeRG1xdfTEAYBJnOXo8Yeg3YbAY9pmzTgwMilVhyv+QVx53zbAp8LidBMlLuS/CIifgj6RI
MYTa84TgqegyRhsv5pSXNnKGUa3pFP5lacyOT93dO5ATVDPE1Fxf5OBM4SC1+C4PwQqRTaKo8TJ8
1l65/pgwIzKQGMN258KEQfo0B34oVqXd3p9kfZqoWPEbI7zDCjWxnvhATWkbAJxY/CEABM7w3smx
0/SaHoUXmlWciGQ171TA6UPDjYeV17nxdp6IFDwE/6e9dDO8sSW8nNfOWE+gbYyBBul/8Y9Meflo
ChFu2SSygTNgihtQ/qExnzP5Hva0rGVKu59oeovxTH0b+xYiVP/IzAnvbMVy3tYuuYikKR3AouvP
DF18KSZOt+Bou9TBmuHUMFF7r5+AMHIgM3faXR9jCc9H7ODjcYaNZMiSJf54S+RfqXVA4/L1R6Nw
NG4hvw9VOHo66kIhv64Z6ljF69xPs50XpKDhn1RS5VTzNvdyYT77c9u22qaem6a26GGuaJ7ocklp
dvy2S3r7ZFo5ztapVBMsZSeqON7Hm+EFBDIdRQrJMb6jfj04shuEGoza8q47o0WMOK15achKyFyd
/1aZFcSDhY6NH8wgvDJ/I7l0/fJpfFHXiNNkbtLM7t2LiHtE/JnUs8LASHsl43SB1/tz9dZDx+6C
XgjURvyqzkFJZHQHAWYhh28nhJ+Inzh4VPdKCyYupBMKgPsFTziQUfQsxSjGQ9iDbk7em0ghDuTo
OzSscbzw9yLd0JeE6FUT20J8kvDRsUBI/83gS+zP4CxBwNuYZmKMN5AyAXvJiANM5Zpvi/OyNKjS
hTt12Dc+R6GgS44i59umZRlzPRtF1yFI7pf386GOI3LOsps57DIi8Q7Oycl3KzUNjWHl9J3gOvLB
v3zfV4WwQ7H9zfIXZozllvU3pzgnUcPiSUDZvKLXG8JkBkzS96PgjKk3NTBfB/G7qa2qTpNzkMGA
7ulTnuDJPZJJGvOYQvn+xFEHlJnYKAkbWaDaKLh4v5p3wUClNSKokd5D1S7D17PIrS3lUx6VlCj/
Or9695n5qVqCramiYXQz8RQvKcWZK3GKdRu0YmJkwaixABVlZZ9EocbLVFJ0VyXlLibZwhku6JGU
0JHZ1RQTvWa/WXMt8h514S57hNM5Mh+/SYNG0XKUBtL6PTj8YJ0meykyBHV7mhN7G7qZc8+xqCXC
ZRaAJFM8Vb4p60GiFcRR/+qMEucqAbDevA9JF2icvaGDNR+OHd8bk5HfNAb4IMFHbEmwpfmEas0K
eRMZfH2DT+Mjf4anAK7T8wFcYXVAMpbbJHxWzXBlBukUwjSEBkKcOm25KPDxARPEGKjJSFcYNRx+
gN6tdV//iR/Rdt2BQycgZas/8awJ9VOiH/q+z1z8jHjBErfoL/DrXcwaI/xZHiUxKb+ZyJF5x53v
XMAgy3v1KXl5civVpNiUWq2HKzVLtsc4vIakjKQ4Ze5B3MGMSb4giuygZZ8+Disbs9I44CvbCkpg
F0L3CPbYLYhHQsv/tRpKv3qCpIjbli4DnU2wVaZ9WFEzHsr60kYCHqlS5wKr8CfJLdC8Y7dhv40a
/E4KzugzPjtGxhVI9RZCTk21T5edeVhTiY1zVOaX+5wdI4CWgOtikACyy5u586NkS3XSSjsObd+D
9JYPBrMHu8tYCF+NmoICLwdO6FTaQFgvvoOC6TQTEyZimZtUJqY0WR7GRKTOKMopJrIVbGa6w5+G
h16KMVfW8eznoU+U+d4Ltwtiy7v5P8P8J0vH0MqWYUH1v6dDv1N7LQzw4cu1G1iqvAzDJNjh8qp1
fT+Q3SH78MIBM8Sk2SMaI66f+4N57VYwtp8n8Rwv2ZejU0MGje0QWU1znhAprXUWD1sWk1NU4s2g
RmPb7CPctqRT2LzfRpulTEgVReFuCnS4jIzTIfKe3ZP7kLepiW/XiECJbaLXO16gtl/VF2u3Mj17
zaUUfPfyomEDlL43A7mUe7ViSNYL4SX+H6KFhMuwgh0lnEom0SC4z1Ue/9ZAOq5X0UjKm6HD0fqu
TXv2qbg3TbTHPZtPZfRkcyJw0f3Mf7hBIug/LZ5Qi6RuWGt+odBU33fOTtWT2wtHMP21jfp9nbi0
o5+TpuCUHQo3MNdhyvDVDtZEBrOznUXCvvU5hR6Zxmmm4I8z7xGMbqacsUb2JYrKK4kVx0sb0Sz8
HRkP+9KT+n5Txvxhnulh7DnRpzvrFSdVzL+sy9dJzSKfP+MhFnw9WoaREHYjH52il/n3MCEfsPkd
kRs14BxFRNlLgMwai5U55jQXaTevYnXw7o4c/07+dxh94UCQh/fLulv3WXqc2I89znZKuaFdr3XW
Qikq5ohuOZOxSSDF7BNGmzmMdt66PdZQizWOtK96KnIYdGwSj3k29m4Gu3MxSJzmCRULxLa4Xykd
Oj+KshfEU1sKL+r48PLBQF4/KzRiagt0w4pleU/FSwrm0tFfiC8SC4VJOo3aPRwQNcCra5wd6pHD
spcfc4O1ceQsGq8dSiHtzutoXvsaVjcY/dvOjAROyK9Cmpjlaf6PNp2rpUr52OlFn4vSy/i0oDna
IbdvngAUueXk2+kSWRv2bIc2L5DuVQYeDXYTMyMjkL2jiJda2I0YpkVdvlUo1MQBERXimEzF2PAn
GY6Y3gYnAAeZjNSIRerW6nA+fYnl/1Wr4RiLAEpJkDqRPMwalpWkpesmwoC34q9pxthDUnrOzf0F
cSKabkfTqQvjsZUGlEfCC/us2xgy+/ZxImbWGIb/pNPU6iVSLuZ3hP8V0acLxj5KK+2KhrDR4b48
Dely0PCActFcXV1hH9gvsoENe+DlA2NFoJgv4V7HC7siPKegCfTD3u2ZRbVaM13DlZeQwy6EuB+t
TzPE1/neDVHBqu3J/SBMCW5aOykpxP53gfrYJOQnKDYu5XhZ6O6vJwfgTX0cEdezCBwjJ1OMFdQZ
KawUQ/1YMpwjgoANh+im7KPyq9lpr6En+n0T4iWKVQTCa/Qt2UJsAMPIywt2ZK3Qi9bUqRUP3ZQc
zdNe+7glb0VUtAe2v1PEQM8PDleQlrRQ0vJfqfssicd9+kg4bSP1choUE7bnsHcOmqZEbhjjyGS/
xyV114J52gEZX2OguDML+70eLOZnpAVPW0VFR7+I9GP2hV7MAsZwTE2B5kZP6w1EsrLxs9WeDdI8
v3EfBwyPLxzVW4mvUNeYyldo9xZ0VuM7i7qZbBfqwloWIgtEWC5zorXW1j4cRmsUGI/Pj7lIB/LG
7rjHoa7hQxS3FpUlumpBFFQByhYspzHEiF9s1s/I9rhF1fjo6O5izh3/TjAcxd/2SwG9iubVk8ME
1N5I3ctxsgkH00Ss9iGZ6onIqpky6zja7xr4jeNhtIfjMG2Nb6FNcWaQwlVm6Qi9gTJ6NeFAUR9Z
RxkO54i0nyC9o76fjMtKtk2rce3rnHuwacMdNQNtGgQnBpzk5QiZvr1HMUotRxjDl6efWY5T3BEe
hGncwLaWQ2gbigdr6GQMzJgnkT6hmdAjwaT/KIiO527aJ+X1v3rtOsyqQYq7jFa0BPK7uIAy/y0a
+ZsXxgb2azk1JJba3XKmom4CdE+J9qCSOyw30r8YsDNLr+kqzPqdOjHcK6eLmXwbkJj9tc+ix4Ko
oxI/XeU5Sc8doks2+mv0wFFk8R/fSwRt8mU0GUDy6pp/mPIHlSOVHk7DW3CIo3ZyBXGrf+Kg1L2e
WfleDoVxOEL9tavKKXiD37OP2sntWdN1c4TjGddgTKnnmx8AkITOOsdhv4qcwoyMZQdcOEtXrnlT
dTieZv1/aHXL9zkCYEiGr9f1Vfuf1YF02g3flxjrlKyJt1WWL3Wj5zVYT98fqiQLi5FtY5ky0Lzy
NH0Bb/iiBGRAFlqiJEPiMv/yvO+zA+f6hcgHWKT6dDHISSML6PCaN7hd6bz2ygZ7lqSMOsCxQLVt
f7k9BSe52P0wtUKqEC9/lZ+HQ0qSqBuK9+lrSywhk2t85AZ/W0g67DI3UmqlsM4KWGgAifsDACYE
9jv3NZa4545Oz58QXYfz6n5L4TaV+xe1GUQGqEgLFDFccOe8SKugOs3K3ObTrqMZOGmirjQ6givm
aSvC7pi/hsdtU6FHDGlfKZWdkmqeWGgHTWACadn6xQqcZvNt+AGs6l6O29/UpH9qSU7MQiNktbPB
qaERXc3jpSXPSvqIpH9Pj8heWmfEcxokg7kShAlNmbMsuw6XF5GuBbBdB4Ve2PmL6+0hzzhq48Wz
jkN2YrOX3pElWy+oiSlGLu7nAFDXev9/xOzL/s7tLgis/SMen07lnKucgcctiyQGtoIMJCDNgcGd
SFPbakxLvlXvzWPdUG/5vPTk6Fv/tBw8MXvvjNgxW2thmpP99CkdZ0BVDgFGal9Wg3TAjhthRuZQ
xO4fILMXPmlqQJbr7tFuXqT+f6JAiR9/GxGWdwCUoi31G0nwnNpNfTQiwD9MxnJAeKaa1nLsbsuO
Fr71Asg3nmf9QhYnTNgbfgETYvbzZSxuKdcBrNMXwDrPfw6yZsr2iJzY5+NTjhP1ULFdeMlQNZnE
fAym4/Wh/QirwVqIMy64JNbaL0IPY12Np/qBw4519vevpUZoPQIJLcNlmUSNlt3ZnwqizLzbWC23
hDOprL3VnrVnW7rHzebpJBgKcZrRzG4WzuXqzEqjGBAoo4sJ1NFnJkPhemQKlZa0Xc7YEXeNbPBB
Tb1fihAGYCeKEsOUvFnXrTQVa9bgpIXVFbN1gujKtet9ZLFASfIWp6cXLhE5NnOygWxUymM0OcEY
9RoaapwCqQLS6NLGYzbX4UYBKKlXCBQ/ZoO6o84XCexz0+NJ6LRjqilJLaxjbt44X1RLSqOZrzfH
iSMZEGbVVOcnSTU4exZdfEtpx5oGCRrElPyM1tnpi7HdvbIz6xkhLgp5inkKE6zg92lKEHbNWpIg
Xvil7luoZsslwdnDihrqDFzhZ2v7d6WQKU2eLn22WFIfrXs/ypTSdwVRrrfIhgv5AomSrcrJaS/t
PNYzHV5daoJL6M0V37p7VcMCBriytUvHLsNG1IrQojSEmc0nAuibRhmgUrYOF7xkYgWXXQopPgMH
R6UyNFjh4937YY2Qqlgf2HbUqSYGmDJQL8WIVBFJDMFgpGKNR2bBvmAngYyMsk2ng8oh3aNpbxvA
RPc7K+W6m4ZHjVjIO1hGSgEwb1WcdmwaT1eujecij4GaUEpBYQ2cpPPaWlIp4BWzIanbCJs7i2P5
36VU689frb9hNtN09DPRQ0PdB1NzRbodfFB9jN9jjTzcKBDTc87lgUxYD18opzAQveh0u/xIxYkI
dHXuKQB65Tjz6Wqw2dmy997Q5qqECDg+DbxWdxTyl5YD45ev0sjJl04H78EbmY3rvanjESHP5BSY
5EBStE+qjHJRsXwvIppB/SftBIXyyDK5qGsT3AkaOhbsjMMekhkjtrJ8k9TP57zFLA91lMW35V1O
yLWkhhw/onv2rVSPfhvDNc2U066KDe35Ro5P9fC2zCCPL5AGsbmkiiF5o3Pt7HAvOzCCCdmU8Zli
cuKc0GrkUIfZUUkC1maA+GyxAAoJMNiklOU9xfLZb8Vkfycd5V71xdGbDBgrWCAq1xhKvnfqG2GY
2uBWRSZREerdiynJSrnr6PbcoIJ2N+W9q6r8eBmVuPg4lGRA6DD0oCXz5JkfQMZuI80RCN8cLsUc
DKbE34KQfZZkXrn6rXw0kYd0E4Ovt01u73h1v2od8KLPCZcvlaRku4uzk1m0W+mEog7wuITWhwBk
xXYWsswatiS/Siezof38TTv41ERX1/ilSEHkk/0ozPADwaI34ZTb9tYQigBhl7+ytPmnvUAUhkkt
e0w7SB7hatimaeHe7REcn/2BK+PP8qcArxWI47/77RHbXRywO29LTG1XqL+YpMQ3K2Lels+v0260
5i2TB7D4eh4rRxu7k+0JetsdO5GZK6aK//2fsSqU+zkPSZkK9WQAVznbzI3gpGcxT23VC4fS//fA
Xv1bIplAThbAoZvEhg2pYS9oU3Kp2kKMYEBAwkJnWjREKnJ49IreMIuNtcdhdghaGbKbIgusMTxV
O/OZpjxu/gQlDHjP8DaUWqTTddCARi/EAKx/qX+tRYxqGP8dKM/Kp1atFJpenvpPlKQ0OwOEgAEJ
UloUy9IJrrxCCgm9ickGB+9czuvMkJhcHxGppVHKkrWngyWO7xIvXK7IXBOphDuJKwatAZxqH7Ar
HRPq5BFO3N8QKTlF70Aask0Knf9Q7ctzQ2BLT8m3u/grkW1vzjpf/qb8fNG18XuFkSxpvfglg/AA
hK/gH7x6ZCWlD5+tIO/k5cMu118lHc4MoaT47jtGBUkmpkmo4B3do+sRzXD2K2032//cPkyeblj+
7MiLxTGZTkfY2ABWrwcCCRwra5tyRbICHPZgc7IrZYX4dGUfqI3REfE/aVa1pIHpWrRpRLIjl69h
rAQfOWcpTC4ynlyJgxou88t9aFW7/qrYGcQLl5doTRuIXviFIvdsAnatD9SDVb57Blx5DIkFT3rz
BFmYfRAr4TVBkIUEpSfvOxC7xaS8eU63hqnmiGsOJQRNjglLfIwGSq+NaICErvNGKVyfsJJn3scq
TuVAMauRsFtvSiVkAtbMvpKhvyTB73pT1GJsbTs3yH4C26RoizzGzttWPKn1h1b6RUpxpbbVhLG+
suY3miq+/0KBmMKp16O12/nfBf5zuSGWI2XA2ZKE+XA4H9MZAZ/PRJGBvH+v6/+T0HZu0z7xKzv7
MLaAPa4J35hwtRBGroUMzCm6MEO1gfrlpJWhterk1MIyc+VfKPfvTSyDHt+eVkKlfEjDHCHmKbxI
uSJNxgLZ4Etw/1MWqMfHG66YVnuovi/JiYFFqMSSfpVFSxxfy3Lu1yrHZZsKCAal1mDsCbj3nHdK
34mXrvEIUzd+pI4CRbq6h6S3XOQ2V1cB1LZW1xN1iHenILaNrDjJQsWHjq8ONrXY/u5y/xYZR/ET
0PReFlVnYBIb+pWVkYrOIB72aprl018SfGrXcEfAzu7Q+Vj0pgjGqyjRzIjpJYuaXIR9B0Bw7zI6
FiXu97p+si/na1K6LKEJO+D2Cbba+bIS8sAY1uEV+z+zxzO0MWhbQQkM1rrVvxtRJ6eD5gsfsO1E
LAk56VrftMdn74fUq83ksGZwD4MFTyalm4QRpWStGzFk0B507BwkqkWnnN6yE0+I3PUEigJBjQK1
8BZdKYKjkusWXCoBl9RMKiHx06i/8eEMVoFn7rDLUWx3auHrCGIWvco/0qaoPMUpBZiEYDjKccji
hiY3QDhYY3gCP4X2HKtmK0L648BuJK1t249f8t1ZxfQt/IOQ5oHLI54p9u+rVepd5yj7CAXhdpEc
/VbgTUUT5VXNlG4gB1E4gB7YKsRchHTTQpRuHbeoi1aDLt1TgmqL0sCsk3AaZiGY1FSkNl3pbUx+
JLhyT8xCjU/2F6cB191T5pzbBpa7rb7wJIqNu/oAnCiVAyBne9ZA+6sD2DAAWMMffn+OPB9ph7ms
mAQ9Awk1sRER06NNXWFbNtG/n+4PcPsICtv6/P3Bxuon6xWTHJW7AIXR2s6FPMz0R2rFCFFfOoWx
YLjKLOn6C0WP60iEn8KJl8w8K80l5UtY2e6yRUIvy7TFE2xdaMxiUGVUpDKLzyhyaMPXB+WhFr4x
M6g3EqJNxqzregueNvhE1GnhrsIIV16bAVphOh2kmSHRUzREWINsBDgQj5Sw0j+m4EAYiz2nRVI3
hYZvCDQkbBfFoIoX6jpYcDJxLSP0FYkBhD5OzeE0CmY66ehDp5DPunr2KfdfC9EvVh7Glera3hkp
zLUJ6wKRxm+7M1ONuq7V5E3jSBMwr8Zt6r7tMJH8qCyVF/G3yDxt1UWtIi5lCwdGYT2oruoMYenV
6U0uof/xPLXSO6dVSj37Q78uLYU3hgeIbizH4stevcndjQqMyYv+ChGTY055tdieyQp+PZvDVGgq
P1qoJikQu3l1estmPhN5xkEkj2V6Z59qnGCy4sGiKgtcSIERKva+9Sx9JWY08ORvyDLgS3yU1Bxd
VnTVleI/e4NSxUj3liXha+udMXVUx3ZGLwjzeyy3iX+NpCHT54yl+svXzXxk8mDh+5pnzxJBUQT8
rGwWznQROWCzmAUy3dhDKKH5dUdcsY21pT2MCdpioyx6UgY/vM6sFhWx49PtfSoKFsAIhgpy1w7C
FaZWX3z/Cc6xx2z8WPTk24t6VnwDwf1yoHBve9b6mCKKazSXEwuVa7a93+lNuaG1bqbPu+tqUs+o
JMP4aSy7/lqkhB5MackXVLBnXyK1lXLv5z8Uz0k6EsQ0z9GqDV4LXcbhjguldejzg6BGxv60CavY
3N9tPnRTAU6YhBD0fYQXRF9+BnPUQD/Hq9Wou3D+eKG+RMQyvElSFI9OlS3LPfHRe+FjaC585gfv
TbisyKfTKJvLEuaomn1ZyU4zhOgiU85YNHoqSHoW/Cn1INdPOEI0qjkU28p0LbROXZedKxNXpZA8
bkemnP+HZ6eUqoQrPXzlRlAkZsFlaDd+o3thtTCv36oIFSKbJzhh57DYy5Yk8rjpWbhicSoULhy2
krc7Fqy44DXotYlAD+B/NQdc89sSXYcxhzCe70xNp2SI0wLkvRlnoHegyhZH5gHWk38X9O2PMWxi
bEJXRd3012d9aw1VliL9niAlvvyaScCA3ThuoYwx6NysP9JgwoxpIlK8e6Er2a8lVLCFcf/5DJp/
B5Ly/Hk3ijS7p4iREDfVv9Zp4Zey2TuDctKs0UZIJ1LrfAqSqBpdCRxk8cshDooxS/qUXsE6ff4U
w9FeE8y6gR6oT/djDqyScz2ICnCJfeP6/QshGUAMEAzj36pqE79f0G8QFDESlWan1xTTsg6n+ghb
YKljfP91wMsME0S4dsHJIZvkiZQqb550bfNvrqdYaGS7AXoTcTAvb+B4BfKVaJ1pWsYKWCAlWadF
9LKe3mdmloluzBKioqHQltqYQ/hkMXc5xf7uEZUi2NowhLfhu4MkSLe+HFWPoK80P9FkkGp1PJft
jV1ffyAn7195j3XuI9PMY6Qp8r5gYYAVRaVCH5QNOFL4CwLDE/M7PUCmc8yps/srWzQyPt+qXGBv
oS+4F3S0fJZse4JBMGX1YOqmllx7Vf5CnH4XJoPelobr+PEGCkyO88uIi1ilWv69few0vN1KO7ae
zcYlAEBSoRRjxw62ABk4Ro8uLTyx4WK41+NhcOdmUhkuQx01Oe6/+J+v48ZXUXBZ4StIwiJD5IZp
gVrmgg+NmC5F+p5AllGbA7+sQXBUOhWbGCUtfR8SpXtnv5EiCgx9jTS4IIM6cjJvBf+5wXqVBEVW
v44Dxk6icwMFTE17LpMasaQ1mDgG8UJ/9SAf41wEFOneZaiuqZf/q2PNryftUgvdt/ONaJHJt8ur
Rr9D72bgvHuuBG0TUuXkG+3SwPCnxTsN7GJw51WUYS+Lxz1ta/PR6EOnGCQTsjHu07yrh8YWKu57
tAr33IUoP9hcOl9oO+CJoDb03nl+lJOcZHwXqsTH651O3mQfbW0p4NeRSUqMDJ99R2wcSZhqwuxF
dfZkk+llsNGSdXqJnNaZvkUPUaHeo8Jjf2aCJsCdUMksswvYv4EVuaReBkbwmIAAMzKspKRKgWcj
SDoeSawLY0PdY6SWwoPsCA1nJs/Tcrki5BjmLhXGF/8EXMpaz2hizHowvOnuq12g1PB6tZ/1kk7t
/YlvvnXb68zweUtWSq+n0xRU556mrVnDn61kdIQeymKmBAqhItPgLjL0eFafGDnqYWOI57IiJLG7
nK6OUEycLXBsOpKy0OImsyWkr6MKlffuBmTT3Zz5xr/wW8ycfKA1VvPpI6UqpMjxM8a0FSCrSIZI
XBQOA9q/CVXpfKZ9peWEUjoCdM7OrAADQAlMEGlvHWZJoGGrS+gssarBtxx/5jkoGEs5sHx/MFwl
NyrzrBKFqlqT7n/foA8XcS/QEU01Iotq6tbgswBe3UEOZcyQ0CNGmZ24V9H6QoR9epq9zsuWLGsT
z2tzjiWqQNcU3GdCSlPwSfh1dB48Tzl28tXe6noMOVudpwPLIuoFcHJJngDuvCbxHLpGPcXM6rpk
avNCpBQa6Wh/5jiHaOro1Ivaq+viCP5SzcAMjp4NBWIGw1bfZXDGn+ErDg2bkY7nhXiituQfiYeG
+WCrmQuB2QuwIeDJqYYVcX4GnO5OKgZxgUFWgvLZdgvZB7xYp5zQe8tH0DwLtF08d60DIAdmqX7z
IHUJWE3xWX5Dzuc+oBbZTQdkzehRSX1vfFx2/vgTEfp1J8S/VxXvecfmellG2J1eTcGh75JEGlP/
IRywl9SRxmJXf0SVeaPnwDGY/4ERneQWQjv7zAwUbVSHn+0DoBMeuI12UOiV57fIJ7VZA8+XPC46
EFLraTUqaD1FNdo6PP7pPvKmkG9jRQ110V16CudlllynnXLCOF7wPTGcK2C8f7V5CbEinSLIQLDL
Eu0SbCFrplG5XFWQpxsva6qH9zDKNWdZ5RZfOcWxjQvqMVY8trnAnX4jI0k51bbDNsgfTD2V+gJD
ykPxxJQkCMs9LJFc2ZvJY1TvTN2HoBDAqQpdezNb0i3UCW7DRat4aSFRcJvNwtbOUvkGZaUZDI7r
KV4cDILPZlbjIHAwUMauldIg6mxVamlz3hsOOqIqLuon1dWMLUnC4R8H6kdTLOlCdXfNYGovQ+kZ
4G+HKdL2KvOZjQNy9cLJBrlosZvp982yr6ev3HYLiluFEX21TAaBvhnu6dEXUdxh34J4nOgHBtvC
ECsaCAYmPy/toxPSbvxvxyI7PQJH7Yd76B5MPS8DraUJRBatG3MdWXdfaNbij3BmynpLD5abzoz4
Blyy3bC9wpnMm6GvrUGZhEDkz5FZ3UNk2nqcr8yvsHnerkFUj23iT+sLXXlyyk955OKapzxsDeMD
7ET2u3BsPf1C4rYIMSB0Hcslcy9GNDLk3t/7kiCXOm8G/vjkYK0JX5G/OYdku+lnUoeWZqWTBcFM
m4S9+j46y3smemZ32UfLZeXAUtEP5yxtProPxggakWuxz8AFhXa3DD2+gSvG5ddboxp7er9agyXk
eVApX89Bb25VxlrRs+zOdA+2srMAV2dBvNJk+VS8hPAa1itXo2crJiRRdC0YConp9casC+RKM/Qa
V9zNiUb2Rpo3Lx2JnVHdmITuuuwOyuKMqVCnihraeyIzGh9scJbukRliZWJtPqrq1DQtwvxiGJUY
giSK6BEeqrJSVX3NUUMzIV1d/o9O2tPoYVM6rQPtuuwPF7+q4WByN4b9NQC58imnI+5ovEASiO5S
WI7eunG3CAHIrtXsmcyDI2CWvxkX3FDfqaVPUIx7u5foPV+sv0LFYJlQ+IEP7hUV0Gb/3IQeO6g+
Nd0HLXiGKHKqHawajZNE9rvVxy7YvNRCygSabstSJIulnEyaCKq6EakauDv7KQ7bMkNoisIplo/1
b/6u92RZuBBn/XGsu/8xICxwOQUkgGI96kSyRLOjtY9Ca/XKtzxhytj3TYE/PeaZosjGnsaBCDzP
cjKjkOBHdSDoEmoX0wUpV/wqGRTRitjxvzmLIOsr08mks7mbb1gfIgYzFZx2mWfhIbUZZUvjE/0n
pcpxGMCTEgqEHzwQ7f61zpSsc7yiberO6xf86wDd1Kak6kcyfYGqe6Z20ZO7//uH4ExDZdgLQDJX
eTl/kMfXFujdlf+jl7j0HUsvCAy4jjPm3yjLFqx/6m80rKaIXzj9XVqiiIxvQ7v45RHt/PTCjsbP
RbjQs1We2/Vsom3vOk8/EfcoLA4Ue2a0w0+s+hQ7vJo+CW6/kexLd0S4h5PVranMYujneWyQSjxQ
WmUhzC5GDzwNKVfAi1Dkk3SNbSjFkFthnO3TAglkn3+0cfyplCsLus4NbQJcwgxrmBM1IqpgFWeh
l63tgfFvt9UbAlEGiQysLcwBPaFhB9UYeN6Zp3ahAyADhYpJpRPO43Y1PbVzcu1b4c7VSqUT1LH+
zxWQkzBPNqBLKe/8KMgVwSxJq8Z3hTGjTXS2vRriviJs6yhPVywp2MQXD2I/7vRsy7WqSWnKAgSJ
yhViZYkY9X8lGKvOcerl9orjkRY3s2GsJq3E4LH6RRgAf7pSAKtrQ9d4W67Y5oc4Zk97PpufgpM4
+XeHC1T4x2eGsh26D1uGYG5h3m7kjFd0FFSLg+QzOyLoEVmfSGHRas8z7lGBhC5Mvjinjkcr8r30
fxLpO7sHnkTKUNkKHYCXKu+qSGU0FqIjfBiKXuTP2DM4v4sro7SdEzdE3SLpmyHON7423nMHJIbT
kc5MTN1T4AxHUjABGiDpjnqu94B6abMui80yf0CVKgbroLlyK/Z8yOvD2PktroOxrhVj2euZPtdP
YD6xsBdBL91WQ83lWmWzd6utqmixnziaMHUysEs4yWSjFeJRitKHtkLAjHF8NU1jjUOwQW9WFPC+
CS0moVtBRXuEI15bbGifeW12bL3+a/Lk2l9HPOY59VLNqP96QL5Vf+xH9WxT/zXSvDHmlpYTOiac
naouq30vrf2s/SvLHRaUjuRG6ETljD6md00sghgk8JQB+DB0r6CYac5yWfdJA7Pk9Oo8EL0gH0RA
pnYicMd/j8ng/sMSyiXqrKzGi7kGzLOOvEGbGhhprHJM50TVw6nlIHqE1Dlv95gy1jVbEJBPk4B4
nT8F5PA8ZsNz+UId6ijh1YnfQ/2DtkObLXx3lu4PMVDVR7TBjwjDZEny8aPUR/olBOBo2rrpJ9UJ
xn8LgQwaEk0zCfaqAxMctHX7ckp45hCOoEbiYSZZc01bcJmwSxdLeh9l1WAg2RVNsvgnnF5TFUq9
OJUXTOVj8bJ8Y7U3WnxV+2jd+DzL/AlLs1+WS5kxMeScTUZO7eBsOGWUKdF0IsyvgXky5d6Fj3WL
K+WI+0d+J2A9r1vjLucNg90yG9GusAiFoeYUZFYCQsC1m2Fb+9cs4JXWhyNX26xvkp4W1cYlo851
f7Ry6l90FZ2Pm6rpWX6qxBjxKenGLWrwcL6W8x+U82yl+YgUvIl6lQ0WGWf2eg8bgztR3l8Y8lc8
3OU1iuxc/gVt8sgo6WYAJBMV06UtkbTnqQ1xeGl3q/HoxegURiSXtUieLkGhWhWRbsgo6aTOsBPs
6taMtujklsuZPUW8+AucfjbdlHhr0bbdaLTJj0ThqitdKe3rrWvVdD8kOE91jBl+Kv+YbsxHN7Cb
WHt5SmbQ/vLkd/tei2WEUTJSnCJheSvISSoVU0XrbXJGOtGQsbkmINixB3Gbh7aKkGs8aDNXhNwb
fRuM4FOT5ZR1OD+xtvYQa5/WydCIv2rKrD3+KgXZqt5rHMeeV9wauwCzdWJHxSO0RMSGP0imDUPH
BCcE+QhJLCtcolA9FU7KGuHeM1jlgNPuiNy7xU3+L8xfStYJFG1P3Pg2xw7GMnX6tjjDsT1kQAuw
gPMzNdV+p0j+wLX89utc1HjpEmiYk66R9JYbyf4kX/z25vR+ulm3lWJ9HJtX75gYJmiys3nTKwSm
iPJoXWs9DHIYeW0j9qoNdtI2DEPaW5aoxLk21iqP1bnWWxbMhQNwkG3DnGZO9GLI+WPUZMbyCvqX
9cSJfmyidqwgNueiZZK5UGU6bTM/msfyUJfyKC/i74zjTy8qLSKMw39AGBFEBqu5fBVtnVW1ELwn
upL5qK7CbkAq9YnI2e+viUNiX1bguEmZ87yNQmprLBN3C4xyPwkiwo+C74pOi0ot1MZU9Wr4E5+A
7EnGrMzIyvN41HyavNbKP5mlMKZiJxPBbv49KKtRCeGofjZFfwOTsy5ng8eh0bDl8HVbZbnOHHT1
h/LWrtfuCKQR7DylB2+Eyhsm2ib9SQFZkxgx7GOYrrkoHjImv0t3BT1EZO++sKDay6VhWZQCIwce
naPlq67t/0vkBTyJaGgvcfK6DaukyUEpnAxPvi9xi+J60qyoYO34xfvXC4p2425L8eKNZ6sX+DbC
xFSCwyMjeHl0Bk9WMqsmQtnU7/L2tMmQ/oUXALbG2KDToXFT6GOBckgOHJ+rWC2iXTlEXfj4zd3U
qXSuIe7xiAO2H8t8B4mbxQpRA5UeCWjfULNCxL47LLxi6TtQFrbvg0lhp68adMTaiw1q2WbI5fRm
fMr/8zcslw3ChTuMDpknLhCyOE2DiWLhVYE6TwFVIcfkolVFIcc30LLxMOT1umlREP5Bf1yTFDzs
3l3UgenUnCQDbbziCEJkl42ibXf2qN0GbuaeAxxLeY5kuXyanSIJufTcRNirerdokogeQIq8AycH
+g6oravtwzGlbkHs5OPPBwCsRtj7SKRROYjVlT/uxgQ9VT9aQniOpyxxXIq3/YC06IpZhXbjCTI3
hUdHDgSa176PseVXDvTJ5mz5Q4z3B2sCnILqHqdx05GLrrl1HzSXumo15z4d0s+kyZi1oy92ltAf
elWCaBcwvCig67Hz9K7JQgyAmHYWgueHsmCihQK2Il7CwwmAuYj67dxvlTbKFYppI536FSizdwjS
EiNMKD+lW0SC5GGiih1vEiGpSfE2yVkLPruo3SPlRtKem0hMEaA6PaG4LpVZpbwi3Okv25WNDyhd
hWoPMeqcRZfZjOA7tOJpNFw3bElzT2QCaPZRnY8Dwu32UvzISih/kX4YYetNARvmy6Onao9UMkZx
a8D7PIUhc7gXJTxlGnuRlIc5KQoDmVL7UnsFXLAwgk4HLKKh8UAxroHZR+S66xPStAuQ7HhH1SrJ
nwGWH3St27JY//RRAg3BlEQ5SXobg18xneAyf8ifx7ZZLKDWX2VdLLi+VDz1Hk62Xy0Tukwh8XCT
blR2S4wKP2ff1+4rM+QSOUQYqYgDmZYP3bNnmA5eF4ivcM+zHKQv7t7hHKpZ6hseR7RfZva9GH7L
LooRyIXXE8tJ6XmloeuRsc7dXfUVdiOMGT/R1NHn+xGRxAIUKEaOjZZNAO79ec3+6+BL9wjtjUel
71+jrh7Si11uKeHn0jhKO3rw/e4K31DXXt3ho7UDgERuozMALbPHQBLH+cKPT4OY5jhXFayVN/9W
NddJvpo6fISsopbFJoKxsiZcfqTwnq2qyGMyh3MTacKkGNTK1pRrE9J8U+CWIywQbwy3enaNHq4M
sEySPsI4GdO55htoXferrqbo2mj9hbrd5arg40roUgzqzpPWI5Yoz1L7qAkVWPFpZkedqzMQPZDS
BAQCDgPEwv1iQRC7tLtQn8oHUQfluQ5H2I6nJ3Sx7v1BDflT2iAfifP6kU+CsORB7ixuD6T67XVW
y0IWW4shD97nGpQajVZK9XdXQwjxhcMyEgZQHSpSTs5L/PEKmN4tFUfjP+QsfxcoiDGcawbDUFNK
GyThQ0ykwxydyJicdrGHUUYAMK0jwXVuFe5apNae3GlRwWy+gI/q3DyXplvXgrdpRzejUNkk/cT8
TaI52HlkY1jG+IDO3PCiClhwoDv+3wSFCE9RhXA2UY6fie4TvHjIO868kr1Tfg+wTFbqchWrlyuZ
MJLGcJLyMXtQyacaxM+oOgoSC57SwATjADZuo+bOZb3SyjtXg+1eewvIZ6A135O7eFu/jNJLvX/6
hgBVVP9rdy4jN8z5xQo3WmORzEFO0DTu3Sz/g+G+OsXYkE4Hbdk3t+rauUKrh9vGEYO8ZilLH+Nk
T0qx7BdfodBRAzyQeGK81CsfmNBrJMNnn63RL/rwR5E2IlmKcnURHFN69kmwMg2jzBcl3p++8XQ4
nvbL1Q3Bmh0rxuDMMmR9e8nuA28PoIqHL5lgbUpT2AxPNMEsJm1uHesaaLMv6o7Wr6v3klEJh+yT
D4yvSIBqoOyHFUOpP8/8iGim2RI5r+gTEB9Rv53n8z/0cOHtaN4KaUvMs29ZwIFVj1UN8oJuyYEW
hWqAWz+VrZJ+xg1WuZHJ6d5xxxo6J7a3Ea8S5TFqe57jMjEhHost/K1TI8BkqkVV4Kva4zycpxl9
fRtg3G0dA0ikfTTbnJb/9GuyqO8n6H4gAVOVfWcAYl95WTa9o2ksiJxWlyMDlC0+IeGCfNhDwccV
TS+5xk6YOk7ptJguQWb3bjk1ezMELtb1fxsz4/nB1lbcX/XjV6CQXlw3MLpw101sfDu3wvgbaArP
Y67EcXJEfr/tnZ3CnwsBdJ7pJfSa0K3q88T4mp+JBwqQGRj94k3J6jKhoVX76aFM+ASHGhprz+V1
H/GB38uT1TvciUUajoMVBuhRu+D9RjDijPPSfXVW1+z0hzL3c61qK2QMrlf6KQ1Sp0rczSBiT3Wb
wKgioGqpmqCW/VrnDj/GW7Yt+uQLc4aL81mZDXbltmpR3j+w7hJSykGqrX0N89X0YEMNXmoZHt6e
Wjqw1EFBiT+BA4KvbfsoZtB4X60LuB40stXMYl8FKtk7BCbTICMywjOMcGgL4Nc9bPRD8VluZbmB
8Bxi8oS98qo3fF71ebFc1Bp355DDjBF6EYkgb9onTXiwdocfPDS1EdmN95YIWbdWJGpWILijCPwk
XGiqp/FdvY7nW6fEv/bRvlhpEx0D9OqrEiN4jsBAS5e9fDsynh19TxbzHOMABnsDNZQaWV0IS7En
guZK50ROxZhgbT5uG4vBI52uJhfrH0xsNaCHoLZ4clD8ne+W+eo77sjdg3/fYlsbD0FaL2mMVEEd
J2XlMP9B3oja8lwB2Ctn957HGE4cL0lT575FENh29htfp7pPjM5RyVHXW9m7KbRSRZrlJolEfBeH
HM4Q8vpBbz34O62anc6Od18GkI6nojLqbHGQsGi81OgQmpW9vMi9uNP/GusJmMoqcTDvPSpWm7rQ
NdFAq7YhEzesZ2xVonxHnvpm5mGdWckDUfdWJpzyqkZjqoLkKUqUPEUSkHD6z6edL+oDFZUdSCuu
l2k6uuR8XRib120E/QkhyzCdO6gWOA3EWv4ChbCa7PJUzgucYMz4fG9DwQCACa+Fse4oqnhMjbZm
Vy6agBjuXqsisqecpND02ottWeBToWyRiWGA2C80LlIxPKqLsZ6gAQ3MAnWqxHATsrCOohC9HY+f
T1neX+80Nh/zh5+WYHs5gbH57NXoNHmF2aYNkTSTFeMLH0iUikYjkoZd3zZDG9U9zz70JUHp+kSn
1FUcxpkLq3nvD6ue0JPwIaeuv3S0vuaTVSQYg3dTkZZq1ai2HB1HxNPBuqDpV0yoeOpJZlJV45Ot
gFZJbPLTLVD5kDajcIc2DNfsLnJUCX4WJkx3dXwD4PhgY03UD3ian0Jin31QQin5ljmFSbq3G4rR
sgxZ3Fq/++mlgzTHZ7bLAh1JWvJPl8vApDt6YB48EzlxJIgVGeIcxAMfARpKYhOhSHXnnPJua7wW
CDXVs3McIdRtEw8UPGRC4V6rOViLzp3/XW4xDpQLpATpWY5p1t1vAyhKayYb3snQJDduGQB+EEbm
mEm1+zmoKu6PQte3xe+8ok/fsAeVmLkGIMGVm4vm0egB+1hxVyiQXRi8e920VsM/ToTOeUuOeDty
FqhK7F/GgpoUewaRL5YPZK8k+rKQ1qJvL/nOWFY+37u2PRcGKICAxEOc5baotHzoNcO4jzsuaN1j
mvJdkPB8aHBN50dGoHHUbZTf5xze7vSGT8IEgFcDtUqs252Te25uLxiag7Sd2vzo5zM4D1R01yAT
BAv5WlpOxof3vZ4WRp449CddbfOZuGkFyTucVDKHB9/SJmDZ9yNjDOq4As/L+3rGvLv8jOSqqy2a
HylgyweQDZ2n9rOzksMSvjL/iXzxr8sKD+wevcRk6NYA8qzirvpwarEfYxD1cKCJQC+pcg7Lec8x
ikUNzZ9/qPnHkK0Ono4LQRuL8DxWtiRpYyYRWZgzLIqKyILR2mTLTiIecge0CVz4DfirOW26+m8f
4wOBm+BY76ixHYtUe98+maVdFrLP8RfyR7DSN7t9sPv/czkjqz787tRsDs7PHYQVist1i+x2xG2W
nH8gFZfj3blC3pfvC40KCpQQB/OXjOy3L1+r8/qmnVObN5nnYDKTOEfbA5iQZRX1uVEDTJkmjdVm
xptkb35fTh+eQ+2/Yk6uleGWHH3dCSUIOw26W3NCqxtuNKDoFQqgtAI7deoscyEjFhuwQ5JTQg1N
6lPu1hxo0zH1XLLuSpAHUtpHw/Jahfz/H1j8t3kve2VdvGNpernmOu9W+bj8p4YmP3ZHT2InW3Gm
tz46VkHKY1ROeLoRryNdf63AyqYvdgvQYxP5nQmtZmdytb7HYf/d8+v/VeLbVUdTr/rN/oJQGlZc
UQ5rwXhZrbdea9U36GRmcYWbv1sNKLvioa+ViPnjeOfxm9JgJbO2fxZp9M3yhwpF+g12lGR3q2T6
Qqdc20vZzGBCWw7/v+C1x0/A1d3g0BOFneicX3huSkrEzjXe9vWNzoHN27id2SYwv+PRXGirGOrC
qahrAiYn76FV85uxpPjIkXGXzYoHp0MliG1C+FE8xpMY4fnHtUxKTqKBSu5McqScjNxbx3WX588H
uWpmta580libIP7MVhMsCtPo4dkjj1BptHFsnF1kTBgtOjNdjt4EwCXCTmsuMruwb+OyXHnCbDN4
MOfw7EjL0+dYRQscfr0NP8rXmmr50yCumRZ5U2Ry0uo2Ba+4jZ0RQAbF1YN8EIZ+I/je0yaXFHcQ
tYh6QodIZ2+yVGrnTg8U35Q1X7CXwwCXRpxUXpEWnuAm5jJcDNHZJC24Hl8ysi4O7Upoa2JGz9a4
cMfpkEfJjz2sakzISNY3Vq8OBrSz5PyHKWOrnEK5axuzYJtyF1b3r08qKivR++/zr4e1cjmUFiRb
PXG6T21b2OFH9BiWEeA+Es/fbR+XZXiLjAtM/0X2k1sHgchA8bYfRnvflRGj1F6cEBWAmjFuHwMY
Uw0okpc9IEZ3AbSEEhvgMMGO/zZPTEGoKL3DeMCPPcPWqIYPu3GO5MlKA4kDr9zq0Jt2SM0xhaoj
kn3cgOrJJkFCZjWZZOHfw+dbSnmBPKfTaOMO19FCFo9ZhC0Bz+M378+DttDwzCwtbyeBCvXXrGHv
CT6ukiaxJg251IH3vAAfYO8Y6Lpo6oHmaXv9k8wI0b7Rh8D3vPJg2c9CoAJ6hu8I3FgmTvYiJvjL
9uNoiAPH+0DEHyz2gfYBVTffdixpdf1GWIAPFn2dOOZdxFHJ7U3V71sY3s1XQREJUXN++0YS6vgx
SKPbMx9xGNYDHM8IqonzDr6aHphr2i3yET+QVDyL326sSMN8wC6gujbtFbbLNeDDsAEB19WHay04
OalPuW2ANTB24e4ACQoBKyabE2wZra2CywklJzDvojkB7S8Il5fXKvbeDzOlTQe4Cl2/eVaJazYl
nG8buk5BVPIeeTfTI7Dy745wYvkpmCbQ9qJadw5kQkJclTq68wxcd1ni9MhMMtMV5tXqsrPxu3Rx
m8oocw1y6uL+uxci1kZM9MXY9Wyhy5jtSLoLnxZRQxxlCo0S2EeGxCAZWpZ2L6TmwUivMwUV5AQX
eA+57JQ8Idx6xwK7ZagpI1szMMgUUt16GE+Z62QwPNWdn96nfwPUIUlezSeTdsdEmiiNjPbi0W4I
MEhpXvYEBBoPoUpbn5mwp3IWSLoZGbuA67t9Jo0pZbQA4hbI4tqC9PtMOrbhU2aK173YzRWaG0+z
QPQwHB9BFh6V0/XI/ouebu2/InL0qjxhR2ouYBJbSVxvQPWxd8QLddFdKIyTojIXlE9fzexLcIIa
UwHCcEZtcRdANoi3WXKeunLdoM8o9G2pa1uaquZBO0y2mhhvRQWzxSSo18IWMA2QjGfv256Ptz5u
i1GAEAZtZvyUXDjYUkGPFYS2CtRWKjZdCKGNr/3EpB8Y9AudJhdAP15gXSePyJRq6RUdubCHI2Jv
nOWxGVNARM1Ygo7E/MFyFIOIU8+aYPbpr4fO0GddM0qdLAPhC5rWASuf7KP47Ocv6EQJZIHKvCps
B1oLlCc1gu9x+J+SF2ArelhlnjH94QemAS3G4A3MBOsZW/e8Z2XWrV7S9XUb4tSWS062A92Eo31n
ANGz+VjwJk+hGArXjnS8OTjkcg/orrvAqLQW4x/PqyfINKEyzi4q4Ovit2LAOrNVZozNXfGoL8fr
e4djTRsMDrhsLt52Lfa4klSSvvRbDR2Zy2S3Iim+UhG4/7dQA+iTpVv8gT3hocXy9Hvperrm4cTi
ZqeSNlA/Xoi5voTji6QoqNILTB1a3qGmcfrOgYIS88xhmo3BI/tjMZGVqjDpdiGW6ckyqEmmCCoh
IohWDVOxr8Pi6pN2+PbSMCdqPZc8rNM2zdBkqQ5nijWj5umF3mmaZg42DQJc0a70F14PwunJDVKM
vSRuWlWn5sM6jbRksH4S5J8cBw2+xHPfTId6lrMYHwSllWV45cd9c0H0kXXBmlA/+q0mxDwYpTfv
r6dUWYo9i+QnEhNNsB+adHPQjdey4vKsN4mNNJsafb1Lc9MBdcbDNVq8FFQaLgZFbNZOjlDclUei
o0lc6IHXJ2thnTolCswt+42ogPtwFdZTe/0vPnbS8jtt4+ltbxWQfM/IljdG9H82+21pjG5NOlYE
gbm+8WHOum1yaVr06iis/000JeC80RlcZ5JUiYUSzU7FAOizlBJbKyKPhhamYaauoegiD7MCs/ru
c8U6KdmXnDzkrmbCfvESPL3vmVbvzKX8mBien7UQ0iuI1n4OBJa7oZXH6geblXzbERt8pzeQW3he
kL1XymC8Gp/LnjkSZHooLh8UQEu1JXYVjTZGtNYJRwdkD6lj64HtvtFSguxsEgrxCvjvUPPs7MoY
p+vjIGqkMpjiFoW0WfYK0TmmW3Z+y6VVXl1NNfsS0X1dL5Jbb/R9AfBQIeJ4wVbRMP5+gEz5URze
0OOjQ86oi31cuGY0zhu6bKAJnDEH1f9nL1fhG1a/GWTNhaRlA/65+zlVr1NMpMtr5e0anQGkrviI
nqj3uOp7LT7l2UcfZfeANTYVc3lOvrGu6V/6oFEmf6NRMRZHOkGI/HJZx0OI5ZU4LLMv9lGWs1kk
JrS24wS5C4Muipr4e0m9QDQZaoLnKNsq9XlkpPTNp+8ARFvdy8pnk1/sAacflXNyAwvprSwFBX/j
xROiLR+vQIUJLUisttiQYs5tTEZ/5KUM0SJNoewaWK5loDS8IT88dW/zO8bdDI7Cy5f8DBd6Wc1u
kREIfaH1PQL0DYRYUEZcnfJyyfKsgNE0PaCb12HU1xSeWWPEjFH/a1lDuEZd64yxoR8p/77EEZsY
6s7W0Sg2q9GB5Eh47wjxl3H1txzIG7N11XQWlc7b0D2TwU/qVMpNtFYjI8/VCVTMks/j3/ij5ChA
19jSY5978aZI6iNzFMgme+C+t/uPyvr3DKGUMK8IRH2MHTdDkwxXdTA4696d01kkckNT1RRkpVXx
ebdBldrcPH3s47VfWMOCDY1ZEOMT4pcrniCiw+PCor0xP63qBu6Th5mUwU2U8g5QgDpqU721qb7H
ESn12LnuDNPw83EGlDdRl2knBuZHpoo4eXbaVeQG4DRdjdJrbCiCNirQF2tA1oVMKzcvR4nX2AL4
A6opMx46Z3gOMCubn1NZY87TOrgiEg09QB/AYP0p5JpadRdcHN1Y02FOnMBJddS0LGxHDY7I395Y
46Seefk/IibBWytntzenaPKJlKouKcuYPnQ4X/O8rGXEKyFn7WIjYQ/xKDemFVd8xTqzlA3Toif9
WcaKZYrOGN+OIqVwDQaX4nMk3Jdkmbl2pJ42NyPQQ5ZfebKR9LjsbSrle9g3uvESE8boNqcYvymn
NTAyJph7Hwi0Vqnqm0H8VXtZFlB3+EGj7CMMzmRZHVK0vvOarTeVr1PrMAR75mEm+Lk959Dl2HKa
8eDmzLkw4unapgZ9He4IMiECqwvq2Xvdz44JSznOEf4UoYmRQKyZEeKpvseCO6D1upd+UYLXv7g3
N8X6RaGh2v8XIglv6lGYnFtuhTh8ZRZdverY0qUA6dT8WTb7qLvCPenoR53ifgGlMA/LaEzyMWBp
MZsvDY/dbJWknIhLeZ9To+PAERU7huu3FXRj/9QsQ7KaYkF3uwP93pSPbYN2UyRNQnzbMXnlXKdK
3hnbx5jkCTu8VjusIVzP3SviyvDOijZS8SE9jkAMDOKW0OSqZmCLKGzjQbAXkYNNrt9C4T9D+bUV
zKz3vQUAAtfGg8FHRgRujHHEqifA7IrjdrKBaJH44ryCBMjJgcmdo0JHywvQpQLJ7EJzUQ7aOE/x
7XiOxqlNYzkOObt89pzTIeRhPRRddLU6DR2+bQFus9aSaKDsDVdj/HA4+3ujsSk1aBOPxaqsDWbS
ZKQQ4p1CJVoBwnrIOd3St6wX2TGqOYwKuB7ho5HuYc4zRAN7FAWBY/Kmr3FDx4iStYaTWpb8inXA
kHKfy1TqUJUVuLaOisi5k30ISyU4DrHemIxQtNJuR6Hz3TvNRut1m0UuMIyWMoYJrVUMwyXSxcMm
PlVuEalWtyv/bhFFHApuMPjzhCdpbyxKZeO9j8BY50gO127uQNqO2CAWrrG7P8QUYLh7Kx1dTVQ2
k96K7CuxAJjhE3MCZdglXxDdBVFRfyPDVYnz4ByN9AwKpwMqYNwzB2pq6ghdHCvVFtEMcMQv6rth
U2DvbZL9ePCb1xCLowqDMJt2QZUhSQI2ZRoyt2feH24X2Bbglht7e7oYL2UMOdwPXDkhS00T3SOm
R0RLROEaxpUxFeQ2hKdOYIbapGrtsWlm0Z18FtYk458bja3zTtd1k0nBOl0puI3L/0OoJBtrZj75
480gl47IHWkgOdAbMuxR/77Q+youwQXoi4Y9YGejkjcux72ieIC2nYHr2vHboX8EfLf+HTUtOAhY
gYRk/rt6F04lPDatCsh/Dn0fqpECv5bqHZ0MpmyTSYXtn5JcRm7QFWInC5S7fTCPCf7CzBoPPm/0
VbBGaZXQl8bjODfbWxrDkZ+wbjgGJrLI71PPrpLeg8w0XPsu4rk0o0CZ+PnPppE6WWK+gb5uzwIx
wjZyC4+BLqdMDFCYbT5kjOqcSjZu8oWWz0TKdA9v2fwk2AZDvqlSFEO13/FkeHhWy2xfJBYSIEMC
HofPHOJxcgXtKztN20+SB7wRC277X8JJIigZjthfoPxFhKcefIKexLk2s+6JlHRlZWFA7trp++9z
i/9LABI41PebpM0yoEDhn9uyBDw2OzcdRGcRp4Bh9fsnyJgFXcTx1yZr6pjHEK29nq9514Rcd563
M7RKvvyZHtoFPcLSaXfsDXwIPv546ngFqvCx0aOFhEgYZMxrH1pfcujU83pC8Ks9Zfp7kRX5GVsT
J8edWaCWzIrcU/p2ByC0mcVwbsb/3QplKVWyguUv7OD7ZbgsFMc+bSW+Q0kJdrWg+AuZ9YRn6zLk
AFgILYSCIObXKbYP/mCgje47hObRqQSeXf6JaDUXNVBoLBrSDQSmABxp5dJk/gwd2txX8r4tkCaR
nSWKOQs4brSU2QQkPqtQfqUJNV2l+U+kpVj0Nu2vIwc2H/IAGEYbV8asK6JyPZchjjG+b/O1fEBs
vaFjtLc3r1xGlYsIAprhiytr2hKogOxuIRts+hmd5Efr1HnJeZfkdGGQR1qeMv+9FK2t1lcs4BAk
nW6COCKwaA2/zvBT2kkCSgoNnyqM3m8tGeCEJDF+DeTzm7yZ2jJgT5+7SLcjEJD8fuqFEIADkmm6
9oAv99hy+RmCnM0Rn/7N/Jkd1MMzcIBUx7x3Dn1Ndk0w2EX0GPnL2lm+6C88G3mdfObIo9EyFsT7
Yym0fH/lPiA6aKn4veHciTyy7UQBuaEm/h9mVl2IF2dcpCmPw+slVvgAeicSbeyqhlj6nd/zOJJV
n4tlsZ+moaUMftaW4HjJVfgCru80TAvxb/YVsMcMXJRX5xfzs1BvP+PMGA4VTomWYt+NiuubMSF5
kPXVN5PRWZUciR42jVFLB3YXxye00leyX0AfmfYf0U/tUP3ocMNz9k/z0XDOlbnMfm+q64yglBun
5oSu/I+S6DX9pxLIfev6mGgVPFcEnt/uW5xKTEC+nYPEEBkcCw0RqQvCxN5/bFmCL8mLNbEMEAhU
9E7QLJBtHI8T/VB4GlUR2i5DJ8rUPLHS93fsg0HZoHSRtlo9YDQJr89Bq3kAMobm9gNNC83rGhkf
Zl37e5eRuMfa246oL4ikwfumkwPYLCQTGTibrZ8HG8669phELFGJPBfgJx01tJilVAH/mQGzGCfs
qMQ0U26uzZuHn8GJHU9qJArfJ266B5lDgXm3LE6MAfs84+JNn1+9QAeGOKB1wFMXufb3mjS5P/Eh
7egPCZs8KPfTyR3N8HI2Qa8jZRT4fKpVDlBa0N6dP2fuExF8ZdMgD1HPQUvedBsVktL2qOxETAQW
min9FR7xpf87EWXfufaJs9K2ZLHGZqr0qjkkRzueYQUg2iz2dW8tJHZ6sFj1RrGP3ABzxipgIQVD
QMIjj140qQTOWHcC1sBcteBR+WaRWRZWIaLT5RoXM992dc1gRIT/lZc3SPee51bVnK1B4k69OHEr
REz/5rGDLvkDituNLcGXTmPZfK0JjgpJw7VL+DdN1FHtRdtN3T4OgAA4sR2mJVFPErCyowQQ8R1G
mZkf0Kk9rymsRaNtlQFvCR8U/oYvrqIZ354JXBJjZWhkkBvTbxvm80Kb1vit8R0aOqdr1NNYiHQh
LrToWXfIufTDjnPu388BvuK4nHfT7Es0LCfsgiZtspgxe9wL7pg6aYrvAE+3rr4yvtLEj6t3ApAN
oD9L/EsVElygmfntpvf9hngzt+yJIpMVPwMWYARVD1CNxFERNJnILaNQj563Ek7KR6XD8yb93xOE
KXmvAz1Yqb/MBgb4P8q8hunibpnFzAbp8dvDZlEamRiaSdq8x47KvXkHD7q+4PPZy3S5D4g1uyMa
93Rl+hb9Npg4vKFJNcnrJTQXcpft1GiAMXOreImNosYbA9z6lsZYaX5EIo+TVJJPMsu/dZqFOb18
wQh/jtroY5ktOt3BCOC5cvg6vbxICqe68wPZ5sftAEtnAx30xwWaO4mzpXp6ApGQWpH6DHpnaJDB
HwqaGMQBdwszOsFO6XNo1FCAJ5uvKF7Q/9+WNSxTc3bZHwKUkQIqOtUczqwiTJuxR5TdlRhxu5dV
hl8NCvtgPYjynUcdJm6K8hIxF2xXR79eLy8h3rVftXay95EFMS9AOjFp8GOGYCdVAZAqd++0ozsl
S12HrMt/lL2xtSQbc2BKvktdheYaPOOj41AMCOVU9vHzM1Co+ls/cD1vEaF1lXfXEYJ5ofUI5jd6
z9lpHg+T3QUEGI3UEWhV0ekUQtZKEQbxMMTcowcVUIghXy+jr1j5lGmvJF36v1kLcjOfCxh0VHb1
aUqvBKUmSWsgBuvp36YPqNM4KGSXlSZNvy6NjsHdKRtLD1xcGPNzJI9I/aD8jeYRkEiTfEDGuAgW
4SrAk11+Io0LLW+/BvEJkDAjhYbepKrUmsrOkRbczsDdqfCMak3Xm+jhydmNRaisyemaH2vBfyyE
N4tg2+/5Tf2vWtNbdhNF/poDeHtyh7J0/i9ebu4KopuFe95eowksZV1XQqQbDrHBW+qQcTZOeF/b
XbDlGXqdOHVwj1klNBuApQXIRjDISk6Ojr9EX1sAky7Ac7wCCuWn1RhSS9Gcf4kmXZdMg1Oop/mm
RfFuSYqrulUOoRtumDKy9jbJel8hogDuhTKUatxwwT4ZIKPS/CpMIaSVj1jHEJouF5TcBekxVqZV
1pMXz+B6Rz1le3DTO9Rg/bBVd6cvq8s7x1Yp7RKu02EjhvMOJ0t56/bNBBEdhv/unXHcOMaYZzGo
1yqvRsTltYJ/Qlozk2Doq6fjZMKEF7hcplphNZRlbvExRAG+s6b5RJ6p7QMAyB0IkqqXIg3Odn33
jeasbt9lF8DDeAfm1WAh5mNxGw8m7tVq+vULzUPcDjFZkHQaeHGwJuC9CHMyIB6yWeqVsvJ3Dnw7
oIbOtoNueiUMly6YntemI/sdKQRP8o28p/vx5tVCXJ1OvNgeCzvZg5dX7OFsVJ6KqI6FQJB0QGMN
2i3MHwZM9WPwMZMcxxigSqEUJsOcc0On4AScYlm8a1r3qqU8UUeiZ5r1wHz3IjOeBMKrT0ZHbx8S
epH6rSJOJ5tABRQAM/wgLp6zzkKKNtVB+n0v5QRCu7Zui9HfOBQNWCVv4W/u+hatLdZoDJ10pg/6
IJ7mi7rgBY7fdAbAbTm0fVg0ELn6T/qxUz50p0H03YrkS4nIoNt7pAh2RS9EvAXC4FX3/iXXLomo
3/PrNl6KoYQ5SgrVMlAKt2Zgv/lb0+TxTVvHrUsxbvGm9Ug+KdsI9IGbZZ0iJHc/IAbqHNpV/2z2
e9ya7WwdJ+CBswtzisPxl+QLwGxebi0vNNRywpqevrWiN5EnayhR074koFKCyoZfzdsFNyVhi5JA
k+iGYTFtvZxwUp0yzCC5iD1Xu7za1hOr8TthoCNree7jvPHlwmahXYdJxS64MCQaGh1Jj0ailSHs
zRkET9sUi/vyD8zRrCnk7fIYf0qKDikymskxkriLt/E73D+KQl0AG/WQ1nTn2oTPH8tatmtVCIwc
cn0iaLWTEmYraNc6m+M+SugnLJcDjD4runpLyCYPPd7X7hE+e9cWbIOR+W52qStUpEygpiVAHhDa
6mbLSc171K+WKYMAIK7piGMSKV1cGSK5bytnn9dzhc1DALcfwcbFbdQC3q9hUvp0YPLc0JLvt0yp
nrbudAlWaeqkfwjhUvpQW7oFMzOACGmZpkvjg2Nltbwtj0++VDEeROiHjnjoGNwxx/E+EYMOseKE
c6w9PKa5ZnvhhMUvPMZFS5ig4ZAIbDCqnrvlF6/M/Oytx4KV8dY77mxDxs6rM6okVRB3GUYZcdSH
HTagVrKFB/a5iantCtJZi+DSzB2iSVlHk00srMqFVWi9CAsvTmqYFB7hLHb0Ex8W7l/C3rsloxE/
QROPtbJNpLB2KKWP2Acq8yY9StrbB5oaTXTyjugRr5rcyEqk1syqNBedyLuTn8d7tQFWTADw3z3K
PRXIj/IDY7UV+RNpUcL2d706uQCYDLVMc+b0Zc9FarP7fq9MevFGwKSpT3ig0Vvp48QcF58S/iBt
woETJJ+yn1Vyn84h2ANOnHbyvoJ2g/uKxsa+d1DKr5uWntrh6DOVkgFXxtezvoH2B6+lykDVmWlh
yL43tL0OREhTjfy8jd4F+nw5p1ciIws5NXrPzIDK+WN1LhJgiTTjUh6YYtv4mJcs3D5SkhFSMDyE
pIGEsfCc2OFsDWzscoRPazhbCzBYudosq75c4FcjNh5rM+5+qVCMIA6jgScJiVlO7Pr32oMjjFiv
lhC+mC6sf7jkuHuiOXFC4Iq9zDXiym3aiuIiRY67x/o4BF43IYjKY2kwAWWldspNvceX4Z5XtUW0
eSlUZiBR8l6g6oqm+SJIkC01naVSU24BjEQe7xE5HYBLqiBCsLb2IU8MIonOP/f86lpGhrd08QJD
hhNSwt3ND+yuuDi4ULnZMbzpEFqb1KBbw3+9rtKQD8vo71W9y0bVV9NIc7FqI4gU/KpEYEWyPCwh
+d2gLT62Yo5U2O+PWqB+pWDAohhbnbyo1kCGQooHJ0B/YW9K17xFnVA+qZKlctQaR07EJAwJNjLE
z4jfmF7kyQItRO9msFc1xfJxzFMsvGZbryzrgAM1ycoBE/xauhixNkS6KNoGCty8E9VqKU68HmQE
/c3Cow3ZOcs1kB3Y65XN9t45zRC6i7Owp+Xb+uhuMEf0fj93Ml4nz1n8lXAn7fHwYZ+AQ7O/MJxZ
kVSdy5UyZylPUoZBl6/5uyDqd9UXcV8F0cw3XlNCNGM984H81B70Bxbss4sHsI4frajg0L+TkIBV
gHuTFDz0dLorkE4IMbTW5DTXVgLGnJs9CzEC5WYI4hyx7KNYFjFaf1SU5u9MtuNnQn5UVLZ5AYeS
F4JTJBOlNU1sRpT4NsZ5lagJlalo4Ct36monRAgt5yU2SfsZWKkLXIZgjwLWBs9k3RzMGEumcCb9
lj1rUgPMVoNIXZY5LSj446JlwZEsJz00nQvU7/xoIJP3gERImf7vL/stDJY7lD7xU3W6bprTn2P0
WBfa2YKKiUflNhRLQbWmKFenL3NKqg5byT/pZ7ewesYzG+ey5HmC6fU/7cE12OQWQqFi1VeZ8kr/
VqfT8K9NpWdWmrpw0CCNpz+sDrZJFS5dy8+oLODBQRv19EbgjUyUHpca+sULvhv42w3NXXeM6NmC
PlcG+jK6dupkAeMR+b+LqU8hClXkhrjT9DChUyK7QMylH8b4AnGympum7Tj+/wiwUo6tnLqbmXyV
eP/C72UGm3xmA6mNyX9xZNzzUQDcRrHBy6rqeUfBrT6f1K3mGbxEr+EzYb5/McMQjTXM5hMSSojc
Vl7plNDZNeRdxuZp4pxS5alLefRbZMgcAOZ7EX3tSMvSadJA4lkKHnFst0/BxAL5MGLh5odqxeUw
Jfd4XRMxJdarzFEQDxQTUhOXd/ABMVaybqwo0K70zdZ0ZS3VrJxEQI6RSybjxsF23nm0XPFNQqEy
yz1d159FcsjLsr5S3MTRazx2l15VJcUlT3X0BFPx551fEnGgLWALCHZTUpk/6zOMx8HkGEwKw492
DT6Mbp+kJqdGhDO/R6GwMV5zog9xQ3vDRrSYYQPkDzDQK7t+HH1ldexw3BIgR8pmZH65hnOK88vq
1/CjlQKNZahwOQ+FmpOsak9sN7U4TJjOSG15ZTUiQRdTtbskiZrA4w2dirLDdd5ufF6/GITNXaAJ
baDvNro+oUALPldj9GpFnhmEQ8/oat/LXFjlqNpQ5pFfa8A0Ck4zd2xWgkJJfCG3MjI+050MBRTY
fHhpRPgqG9UvSJyED+D6GbMKPM9ORkLolOF2YYILmsIKhjcFEDg5Fm5j2yehU80IAu/j67poImkx
h+UenYdmGfJdO0hGjsOiO1KYnLl337y138wm+oztV81E3WlLCMbls6cGzleG1RMX1bGspW0AJ5NP
8tm347iAwat6tW7vJ77K7GeBt7FR8UeTx5DbJitl9SexbtZT9QM1I/9D39iTw301llOc95LUPf7a
xI+Y7FHXaMUiuhMF7brdVparTj02z5FBhJhsDu6s5oaMzY7yi8V4u08EJemLn0yA+klzs9AIMd//
SFZU5c8cAWz76agIYuCDvDugZZ5aZNiin/Am17E+bEAosEnsVNi6Se6YfS6tRRgx3VU1O/kolFf9
LwICk6Dx7A3mTFA6sGLmIkxehHGH70c0bWiQeqMeo6YziPzPRAwCG6gU+tcZ7iyHGzOHEfpGXDqP
0oL6fqoOKXELdwV/cvhkPBROO3Gn79yJ6+GBptFB9Vf80OyBP+Klm3pH/4DFYklWY4Bskz9907sp
RFnlSlukjPIQDu3Kc7LXo2kExiOGgu54UkvoML3zDjUWh2bzNXy0HtOAQFMHJ1hbbGPv8e57lejH
MmUYuDyGQv9AcoZRgC6PeK/vuLQQJO84Wl099jQVEEQAXnatakqWJ5s7AXsbHuoLi+eHonc0qrUV
dAEW11zwWbXHHURvzt3M/NxFQAKYOtVKHc+5bF0niYOMjaRmt0UDQoO4hc+96JTkPL21S5P06Eeo
U26gIM9tNqmVXouLUuFSNVIINd0FvPQwO5cv5kDnmJB3ODAF2FlfxVwfCn/iNir2yS70h62gP7+w
46fMYwvr+FhXltK7NEeWZcRtkVp5r7upQ2AEPsBkiGRTemnlCTwDWpC0uqtGkd6sNqLEpV3gRhFr
LVB0g31brGbb+eOV/tgIhSmpP0dYF5TEazXI0BEo2rx0I4o6awqlzFHcXMlgA864Q/FIJLIfSey3
aUViwUQD1gXhfa34eTbusYewqQIwX/3DTieqbaKpaLHTaPyKk/z1C+NJpPYqsT9Mhj2DO2wGSY4H
CRVctrAgXIP634ne6AgiU2KXt0zKUWf/zMYC70V+m79U4iYXUs2jXlZBZAHEoTZ7yQ87jHxV5Fde
NcP5/gTDZ+i1FqYdM1TmwQ8JQf4U4XiPmHDQb9ti8w+pDiadvAeOUpUeHJPmUYUMDiHB72kaPN7J
Bd0QlCWdqc/OCMIz8ARLDDr0iLM8yz5qh6P47S0vUCTEHns1/3GcgGspMe5kuPw6Lm7akZko9fJc
zG8o2vdwE3xNucw39mRY4ajym5km3G48g0qhYIy76C3b6FzTNrRXCReV/ZU3gM7g1MUVgvvUPBrA
Yyc7KvunTeyGCqjjWYKCS7zn7XZB480rhaEjZ7wh1tDNuYMDCkcuyQnfQ/1BDO3y5ejA7JvxpHnU
QdOkdbdgn9J8IgqwYsgs8ZIU33g9fxR/I5Zw4Pmdd/Bx1XoYt4T4s0OgadRDVFr5g2W6mwbTmtjP
CO+h0y3jq9ap7PXWRYX3KaZfatDOVbF5vyAATNIpDC1oTkN8Or6M1sEuMd7on3kZKQ4qlsCZk+8v
sL+ncXL1XffZrHaxpgUcB0ZLL9vcfS/xoGaimQyAWwZMVY1YiXYMOLGpS8+6eThhN2SrjxqGfsu0
1Ln03wPkN4sWrzG2s3HeXD0/AA/FDRHgHgiZP3eMUOBzU3DjvOoAwqRBCasbusYbZUCQMZPeNWpp
EgAWIsGnF/ffpjRyRjYjpudk17jNrss3FLux1bN5w0cB2g/t5/TQ9GzbtQwawrhEC4mxu4PVKJes
c2g5ozBAtFQwvtMrQkfznKJO+cOgOh0xu5NRODmyPkmwAxpxzyCm/iXzWlVEmtgwml9Fz3Iae5Ku
W+mHiwWzikvqbEl3vcOxAmeXjhKN2mg/b0o56SkZLyRQzpOBFkOP3rZwjPJJAY+uT0GioRWBvOaj
LlaaoQD0jYaP+Fp6A/acrcqVtn/CoaeJMvGnQtIYn0G9vuig9qSrO3+OrpjLqeLyivpQpbJxZ9X7
ONjSeR913PVsXHSqQbEzwlyQVCUFWDU+YPltTV75jjKaJxUM4VLPTqzF6devxW6ZKC2kwM5Obh6K
wq1EJY5TAUGaPPYA0F9UoatNjfJUzyqAyiuZB8oT8Ta8tkofbj/yImwi8fHytTdI0IkF5MhReHYV
c2KUi714OzcgPp/SzkQQffqKm5vHlmXrULTLgiq/ZEU5oCHodFiASQ7gXqioKzKZyLYuHsZD/BuU
Aasx8ZJyJkgMfHg+181jqxZgMj3y6JUu4tcb3U74QSaCru96o8nHxU2EN1o9wgTYis/K8Qer9YBQ
/1eBy1Pxy7SETbOu8FYPM8+HvbBvUwVsqNb3osKsy1WbJLV1Ulb8rnUmQ6n21Tk/E8aey7EMnpZ0
T25Ts4PgrpGVZsC+TFvITrpz7gQjlaBvSzM+JybkdCASnjJIJmAYvFpHnWnQB91dx8TZLgk5shaG
xh71XQvBLsWibLOpJsuTcOo9opO0EvdPN6mDQQWjrGAvsCoHNTBD5xdHc8NuicpD8ml0TXBYFPQs
b2GbEXYqIJrtQRElONsvx3LRFX30OQ3hmrFyHeeaa3HOYYlnXI8AYAAuNBfaoOhwKgE4gi1nf/Ca
Iylc6xjpjXl/QzEEGoTjQBBrm/nXysKzjGlbmWXEAVp2aoHkJ4VK9hCMhfjY718TEwasY8gT58ds
pAsUoJYj/vMj/f+JbnutO0oV86a1FBGh1jrTDI580j573q95MhjcK9i/h3xxMN4P07QAWl6wp3uM
hCBTdthx/n8XSb9vZjVHy2b35H93YbeqQ32bFbLQ2nydmtFdCjZZDtVnTD7bRI2ebFK4CL0XJYes
vDDmLX+4ASuuxESBu3z6Uckim1+KaFvAAyRLeH1mqe71KCA66NKI1LWyfkF+dvajjEppHnajrdGu
HohKvsDtn/dz9rAZe+9Zs2NCzcHoVHFoDZH4uSMUvLsI+69XRRho2Q5cpHlpJvxPbmXSrw6D8LHC
oLuYNvbbxKgqnlxdZKypDG/Yn8AHEq62cTELDDkOSi/0di/+fFshvts+ae5hDIvDz4SpA3jS07Zq
/ZWdvdo7UDLIHhodXFxN8JpOLuU7A07zyQ+HwTODVWUYlndY8MSUPE1i/gBFV3BKVainWMER4duz
Z2/lDG1nsEHzk0ZEgtBOnaN/VpbmqBmReqVjNfhFBqwdrfaPDcW8A261i1ZCCb0HAS7T/RnETHi3
C2WhZ8LmTlYJdAbUEI2/l45F3KL90O0IZoIXvxVyu9/XOzhyL10xAVWkc+LvlYPOj84XjqUSHRFP
HmcwApFECiRo7ZWDdSrzuxKsxGV/OkTrrv36Cp605wUhd/f01yfPB6W60uHKLdK76t/Jckt+XtPg
M3zw3ohfwshjS6N3SFLTnoA03sKbJ/4J1Js6o+QB1y/qk5qxn9nUNZSJS6MFP5iapLPct8qAiI8k
eZHgyu+GBn2BDghSGguvdfEPH3z4KV6nylfN17ITHno6XDl4cUTfdbMsRnZ1JpkFZdhtUTXXRCW4
49/hG0FiZwcwa//RUPBE8hgSv/Wogik+wE6ZDTAFtUi39w5DWhmhSaJ4olMSYV58QjoQUpm0hXEj
F8ze6btX3hx9qzjHXCS4a66XZFUPog7aKk/Z882O1zPfaMmpJ4nP4nhSApqVjxsI3KZxyWBdiJEk
EShPZySXLWCFT9ZLdUYj/vaKRVAj7hkWoBwPojBnWY21N2DoKSX/YYxyj/zLOiFeP24TLPGAlg+3
Adnp3emttpwpIrsI7KAYVIPvxexhQwaVUNVq/nbXrhHo4esEXL60XrDx9CQD0gLIU24VlnxKGD+w
c7mJifMUZnWRodi53R5Ai5C+SfHjLhye9FW1I7rIA3WCyLke/zwFmOH1zmWSB0+J/0V85F8l6TDZ
oF8+SA5Gr5vKsJVYIYKeEe6BRImUV3akaos/j9ZRaBj5XSmkB4x53GbgS/M+hB8/tj+ifv7lXITW
+Z6CB05QekiNc6Kkqp4nhXeGAGQ3jte3gvXtlPJRi9TJ7D12aAbhIcRc4Ck4sJ5moOji/laUxlOI
mozymExku2OkIaml6Gt1v9tUNNAT5xiMVRmB0OO2Mr7esx2eGS3O1ZRsD0LeTfd4Te0GF1hN2hXn
TB9Bk7u79Rug5vsldKwVqXxrlh454J181a46cBUmL9Dw6+iSlPEeU2dE25RB7XG1laUhfiE8yg2m
Vou2X5KyKSnuIqJDaJllzEE01ep5RBMbjs16xfpv14EnA3fHQhfIziObSFfQnBrAENT13vIrbsGp
uynVpGIJzDoIhZnb5l8If9Zym4+D+i9EpLmp4yOltDB61CsL2TStbgu36thvdlc7E4q8ENhoS4MP
hiGSpEAXbknE6wI3brOzwXjCSY5/ELf8bUoAQVLQi0yK9kp/tfhJC3dDqrUKOGSdmVml4GJ/KJ9Y
07Vn0PvB3RssKutFzuVi2U5CQz3smWKoChlIstWRuvHYfc23zTdZFlPpPDV1MbUmqkmbvTm7Q1zv
0QWH6xLQkjvaKtNytR0NeQ/fJqL1fVh05HIyPW60D+xlFe9rJLzyX9VaIGIP1SsCTg7ZAHp/MjZY
4DmNrIu/wCgV/5eoCTmd9fb0tUZgOIp/kyBB7XYF22Ml/eQ7Gks7xTHHn/9CkFpd6vjm6HX95DH8
rkEK0h7kV1cyzDlEcIhvU2zS3+OEK5TEt041A7KybZJH6I/3cgMt7MqPv9pUrOgFvxqUcfD2piLa
5e+Ph6OwemF4YuyLXRJxFkJ9TV+wFNJP3yV00UlK3TCqKI96PqGu+M/0k6R02a2mtEgIu/DuXbyw
i/kZ7Z9co9iEFlj5add2xabb9cmB7qX506R4Gg2ilfh5JVZSkcSIPV6P8FA4vYUqe7asvLucuZqE
wnYZduatqvj0hm9VOoU1nlKGO7UUiEbTU/mRkEyP6mhubSF4qP+RMkSbY873Lga+Sl2St+5RZtbw
dqT0oQIQrK81TbZzuU0JTak48UHcYutWeb3JVo0Pe1R1U26QCMJK9Lo9Avjn9TP7Pgva6VSpDW3h
yCdSiIm1mGi+lZi+SXBtd4A0w0yO3EdD1n1lcOkySXdJIgx3msGUifgcSg7vblrFyNkT4XNfvTGf
And2CSfuqDlQv4ZJ808nW0DfEY/0mata/7RsPWxYqrUEOXlVa/V5fG9Vw1JGlpbzqAS45NEUEMzy
n3HvgFYF5J1oDMnBUL+OD5uP0Y/VcJIL6OfPq1zDK+WA358IqPo0xrg5hb2FhCw0EgEHkXzul8GW
aVurIDb/4l27rJrlaAfHrTRzJAGH7QBnbJlIM1S9xbzjejaGZg4pA/wW9sQsdF6QQShKssMguGxD
9TzBfufj6Y11l9gZBess7K/mSd/OgDonygookbVbaef14+ihMTATILfIeC5Ah3w5/BbNPP9qNH3I
8dGE9oE6hNCqQaPazjExhVmsT8NVUmFot0Bb5LknlHQ73WOy4ERGGan2iIH8lYQbfSLMJcnikqnG
G+DpALN4VZshlZIvORlpp+9zIF+n5HXayuTvWSy0v9SH66MqPrKPTAejLzokwvKdd+F+x3zrsIyy
ilRVVuW3qdkggRJeogn3PFdTC+uv0n65klzQmxUVs3ezZj6THiRq1GAF79/9Dgd4Y600H5gx/OCp
iJc12L+mf0l9z000P+Hicy0Rnbc93sUKiPuORAEv3mztLrmmjRyomwZhV+o+123b91u8pLVw+4zH
tA6vfiAVNvd5nj1r48tHQKzk9vxWe7ms+lzCFlQF+1KIE+ZPBHrLIwbv137u1klrKk2B3V2ecMA0
GFFqbesntbnppD6XEWQ04F6oXckScjDg+py/9SgYwI7p96tDmHv70/hzz7TnulceSDIkgO8fvLLj
2DKkdSrD+J5TD/6xWvZMyiRkxowbU8PK9UPgAwNVBGPshQh47ImH3RN6s8SDhYCl2zl1zhkheYtq
6yC7fiuqeN8nucup/NgblFBRQF1ilfTl+o7HUm5+WtTV1tLGJ8jpMCBXrp+sie6ck3GMLX7Qb1UL
hzfy1aDaWLOhLDUauYjiLE0LqFzQ43iesfO59axMBn0v694+e8iCUcrH+4d+7f3GkvrHlFwHSphf
uDP7h6Az3riZt+1JKBHEuCrd1p+0Ee9i98OvuEO/Ji3prGTithKDPQ+/RBfrbWIz1+BMcRM5lVmb
cO8ACGLOt0S1FWZ6Rj21WLapAl0xFtos0TYsto27Xuw10JT4qf0A7xKmOjtgAcHsA81oC9mFY7C5
p6AlNplBs926eC9c2JhPwQPieXYVcAvWEgR673jNujclMaxVbh27c56NZ6OzC9RcS429Zv8VA8oL
4JLSYaSURZSdbOqwJYfwi0ERj/TOLt/XwK7UCmlYxYfRpwRie2Ao1y/tmKH0EGD8Adfe+Lz7RmUB
5T+9JYNUiCMXd/askc5HY9wNyriy82QHFYpJy8PdWxMG99dtNQTrZyDdyGQVSNNNHScnancyoy8j
MEiJCcySAlPE8dggGsfYODoA32L9wgObOl5vEaWJf1OopMlesW8qMRHa9zbqV/Aa8hRzqkMerQHn
2eBFSQTp4gHZHYed9cAFlm4aiXvFZ65E3e+99QomkIjf2c6MMHl5n9lPNWs9651/ZsJ92/4X3Ljo
g0MvdIHuqg4Rnep/K930a2xyC6iOarRketsYK/I0NooBEAd9JSXeVGvoISZsloKRiheKk8COpeU7
DXbO4ka0/NjX8yJL3keWKgLEEXAsj/DDgZsKOn3ITCpQ9U7YptACYEwTbL7fjBuUUJhkD6MynfjT
i7lABIGwM/ULqCB7N/mxOPZsu9m0a+T0132JNARxoVlPCht0wq8BGffy7VEimd6qY1nlOJdmYi6O
GAClDQYcZHIdOuB7V8bRrF5wcu0goPHWoiP0uyz72p9rhRWv7ZBdmue3UCwxjUAZlKYDR5/egfsn
mO6tr//v2tClt7vGGf92L3esfoO1ONnCfTllSWUL9tSucVmfflyW7H5G9OBGVPyGJt64FiHocMR/
P2mhPXqC0Oz80BAvV1pc3GXJwybVtE8PA6vjv0biJEmgwpXaxHyMlr3BK/MDTP1Rgh+uhLdMO3rW
BZ8Isdbqq8TnEqumhpQ0KZKRozYPFQOH7o5xNuG8pYgTi+auPhdRWT1oEftEhtMfmfGVEaJgKYzV
TYW9LIuXV3lWM51wacVK2D0RxqbMrgIhBQMkAoe8py1/IGVmGs/TFylpKEJiDWgYY0CamEbxD7kq
/Q6BXa8PsRuBzFOvSkA3rgtDLeflJn6rXsQbVlBM5oNQoR3mN0UddylHNkDzOuccMjGkgLtFmAyC
/FPLr08SvoHpPFxlS/1dAqx9jNu8iEbCAQ+u5X+NmoNVNvK4lq6gkzKHc9tbuH5HB5ORglvzFlat
GHpsqUWpJaWhH0gBcqoxAD1XGLUwNG9aotMCpqMLYdAXO7tA/FaQzHu5RnikGDUryOuizOXJtFob
+vD3kRCuktUXA48tWMnFcYFOmvQpvmc/kEYVPx+0+qetRW4PEOfaBqJGDY33tUgWYnD1drrsQ9Up
chHi31UF8JnvcXtbtl2BEBKDfSgiwsfDDPYu91y9pWzD7pCBPSZXUpu69bRNtP1aJ4Rkif/v+19O
D71kGn1Kv17QCyu+SXXnmau9BVgaw8IY6R46MDt+ZXtyLsHPZ5MuLYdNWtmZNHQ5zv2lqergNGtS
WYH8x0lAmEXkDvg/4JjkBk0WiSAkRupc0q0uzlzsP4bDRYeP4zNGmZieu4Up/UVAfqEPjiarqQaA
bqvgZadQ1laaqqCxjypXbQcn3OriJfdHhT9jGX1aS8bqTdbR4OvuWeIk3+Wyk46RRMrtTD/TQOEb
J3pkDdShcHHYk5yy65hLwmLL/hSaNzNORXxbnKf8RilCSa+Ie86nD/XQCLrAmZ/gvPnXb+N4T0Vm
hFL3y2dBNtRorZ4IEaXH0C68T0WcNykLiFYfSErR4lFMf2PbPSMwEUy13EqzWI+QoA+JotVchOkk
RJ1QKDr/9E2RsbxJFdN9IUSVH5d0P8EJjaKdZ4BAf/+D4rRi4/BqfcG4zHQDYZI2vpJtEStOli4S
/NgYDiQqsQpMJ1z5XTgVCwZu/n+BvQYMfFmCwsgSSAZQ7462pKf96Jnax4U4nlgIa+y7VEDiz+dx
YdklzwIUWwdQsBVSgUNI7bnTIIBfxSS2DFiGtBeJs+eaTHgDmwJXXO0gHsa6jGDyL341ret2MTR/
qXvSxmP1UvmMIVUzt/MIX5VIAVXK7cx/o/mOKT3ytcvAtD+UOcyrnq7zxhLFKs0lae7ZjIrsEFiN
OK6lIV/rUzcUsSJaqcEzbq/YU5kKyYWrZd75zQJF7FhRwy3DX3YT2P2jKf9rp3cPrwNzqBhKsdTV
OA0s6CUIErdklHBgDcrG/Ez/fn2VPq6elvQeJ0nkf/JS/ScPnqhFupfnhmX17q42eMXB6RXhqXq+
L1vHujcnPtu39ISGbkrb0Xo9rZ2YLEBylVgjvUKCpqqSipWauNjbuSvFepo3IF+KxzourqzU5CXV
+3MSzrzpiy1a9drJDVb587h5YqqwwZr6FIHRd9zfytEgwAVrpSwtORowAHKyVO//MBdhVCSqWHkY
dDesMzUEczSyJKMFAFwRcrmFef7BsdDkUlwKbQ2BfbIxTTVmJjvhWQ9uPiGc+tDkGtcB+BftMsoh
Y5xT7rVAu22lYJml3pf1pwbHXRp8DAHi5Yvfa56bQ4QrKP82un0U36j//2PZ26jf2bKH59Yhpu0Z
tAqYMKEBD2ZoqPbVxEISDW0w9xBfv+GTQKHNlxxLLqBXiVe0Jbm0NYgvbWJD6yhHUDgPb5lHMEdb
WERl5q2a4paHU6yGYwtNnAfyFwiQwUfu2iheG41nHLQELbzDyE5l32YNbRCScQtuoaT3JfXyehki
gASZKVagJmKRvPTfdmGaIerPsWuoUi0phi+yPvVJKqgw5yJ0X6nDqUeoPagknQ12s4LmhAwzvXNn
zH1grwqzNecAbvKOf99U/ehjgrSKQ8Pp31FbgvkYTe0Gkon43qRjmOdQHYEh6mHvy9VLjpvN0iVi
2ojTMdi8JzSgTHonp34LU8yMd1cF5+G+8p8BPj3pJJqwd5Kel7n+L+Z0L874fe1qVwwevZoOYHGV
YYAAQU+ylqnFegxYoVtgWS8fplfsbbodMevHwqH9Nk9NRGXjxzzM9Afkf8BmuX3EKJsTXPIonyGl
DYOOpXWpngNiDY3NPmEg6B7Kkn450agXOYMgPZuD89NQzDtskWkaD9kcGKYDxedG7AYLJI8z0m4A
Q3GrFam/s20HEnbYqvH0kPRRtNwHZ+yKFdcPt9U4IBvR8FtE5viKcYj2umU2Ndibl6oRKsccDxTb
7JVwtpcH/RmoD8ApvB4W0NYaIxw1ChH9wIihQXPhTHL66SI3S/r2EhpHN5pDWvAJ29k1+NcOas8j
3HdMug4eSKO4W2jDriCP5I/el+NhXKlp5n/u7+Octxhreq7ft17dQ0UmorXUrKulg8bjXb+Py952
1JKzMSTWIG4ffcXzfVf5V5KRPAfrgKp+Etl2yxwUdxLsv50Ci78Fk9pBQsaEo2O7KWyiF93vaIN0
qWuL6uFdlKKVzKjl+3bHHpyssBiCHznPnScSEkPjZnTSnZef5ZVM/UGp/I6jsQqt8bYFGr9EZzqM
/JI1KVr/OAz24THs9nLkPuGnArg5T5No4Fbk2KLPb/aas0IRe8Ql5vWRBVX5wRyEj0Z5MjkkaN5q
NRg5zsyS9oEgydHw9fEvpUKgGEDDVHYLWt2SHiZMKM8zK/dbgWUGb452Ki0rybdto3q6zfyDNCm+
Wuqdr87i8B5qf6GeyFQ+6M0StNFBGKr+XtDQrm7T4z8qMSv//P2OeeiYDS6qrCxQM2243bdRHLlr
+pz1k4GMyKoXyCvSyydeNkCQ7TFgmpx3PJpJjzJjxHEq2RIjII2Gvr2D0wMw7pzq+aKpK/pgCCDV
KfE9zJgTbWAeLwqpgF6tFyp4wTt8AOhZG7m/y1Nf3y/kPaLO4mar8sFqGENSlSl/HARvd+srzJi2
kGGaYArASsPmlJrHduymE/VFLTZFgiHC8ICwxOH7qBbV+8cRLFxtB/iXbpDXuEg5fHSf7S5rFsG4
/Jvvk+IXlgX2ciFlDQlQJaaRWIoQIDP7WRFKcTgW16Uq52nY6zVKPaykHG5uNqbz7C7ZQauM3/Ig
MiqbB/1HcIkUUUCtm+AObZ+xmUJ/ZBaUaDbx1Mhz3S8VLNkDgX8eJQRyBy1wHoncrTTnBfRWJv4T
Ir+wd+N05c0xB2tNQq33RKWyM/dKLFp40v3RoWPPU848rC520DMwaB7w5wt7I3iuXEZ2r7g5jlNC
KjcQBOW9JfWlLGZL4xyxBM7O0wwWulO769FCAm+ojBbH5+OdZn7HOOkGq+mJqrvLShoCr0ms8mFP
t4jVzJUWlANEC3nTWIl3pCfc3o25HkKgbmCHb6yzHJG03Q9yLKEmCRcHgy7JPmek7aaG+j3BqXA0
jm7g+oWTTZFspqwSN9QxcB5NeCtLR3qyv/lAYVIVQhU7hRfORzsxwgnuIx9lAtxE50Ouf1XZ8TA0
DWNC80n8H7Vl9/JeQEM/Gdh6izHoq4mHMRfHVEHA3GuTyJbVIDwVREF0f131f67c5hTb1vjDr2vI
LH7NFSgIUz7Bg7sir9zXbCT+LmiR+0FnK3LLqBk/sTWFWUQjzpS/odDxa4NznN2J2+KlXjyrdUGt
SJbPlhQBlv9hZ3vJXwPebHu5pfGzb4ym/TdMMDtXTfPDt9Bv5104kvMVteavhCO+W/osqpizs3Dq
p0Ufr9UDRL5lu+P8NO6MCibLgmZpVPMHtTjsO8cyAdHhBCrpOMx0TqchhBsCjyHqI4ixZFuKrz9M
qeOUOG4Zhasd+xMQFHuqzn7tQRqgiJhxNtT9y4muihLgBXJWEUGIMLjcVuBqaVVrkHi3bUd9PaeH
pzdZlDQEkoNNIABcShBwHO3SMJEYHZqK4TTNd938xrtZ2gNvCOUONHofrXiz0C1D5RuLhZuEmoUI
yClPB/+j6MAdRVeq/EZeQMPx71/JKQ7bQw98ya1ti4D3XIPi2VMZYzr0IvKtzHqDyr8G7/mYyKqg
Xy1OQc2X77ZDwhbPVYjSj4SUT8Mhc+PQ+KVdLEMeacLs3v8ZXHU3pk0vfnEZT6qqKwMi+qRh8KJy
zt6MbyKjQLqCe30l3VMdyxugCOBc4YzGSsf06g0eC1tQDur74Ng4QMf/GjVNkJjerSA0ZaTuJz/v
YUnN8eWQ4E5rlmeQ/UYwb5yjD5urGDYGl5eDL6C2f2AKQFC0auM0LLUs+zVS670XkZZjbNmFt3hr
j5q5tu9/Lu4MX9XPiockLs+sH25veYzlEsA6n2EjtfzGkl5xCJeHkeWWreA/0g7Ymb8GEUB/Ktv4
V/oijMQg3U4rxKNIrfHjrjsxv9g9+wjg/ekJumiQiZkQ6eQttZXeEbtfocE6cTOk66/g4Q3BObZB
wg8uEj1h4Q7YGf/g5dgk7BzpKYZm6mRBnvntG+xoj8Ct61FOYUoZjnTR7pxsN+K5J3cICvwQZOh+
8IrHci5LjU4KWqks/VqiRla2665uu4mx/geLfufZVJDKAFxV1w4FW8y5AQZuTLQR3l0uPvshpvsH
jZyipGC1IpriEfGuzeT3vzvoQUysA37LJu9jJ1W2wNB+dxYk8k6EJkiqPX0JZZPPCD5/LSNC+YY4
XXPY5MP4lspVOWTaTPcgygFp3sJBwnQPjq8MefSoM4xkSw1DoOUmT8uTrerhvLzqlHTr/C60+GI2
xd5GUcp2YH6SyO/31xLVl4IgUTpdE1JIaMvyIY0rUazxQo3AKmJKJrnbYnF8LSM2Gz5faOEO0RLw
2XUF/xKIdYR1fzeEFIYEBdgSelLEk6gsHE2Rt3yAKYACIswczgSt4jT6ogAV5CvOuTXehJ/W66Cz
8ANZsL72ciHOWwuo8YBcLEv0kK4bOcLSmblScok6IBP44qExNcYEHvgYvoQKfA2i1GCSWjygFxAZ
NNZ4dZ/Ar4JT+EH1H6aCgSZX3A6f8PumWgl7LaLTbTDf4gBD5ZxXRdp8CLj6Xv7j+/mz9WSkt/fq
38/qDztbzM5sUrPwhTUiL/sWRgkaZzLaOZcU7inOBQKZvU7zerxFDCWpBnxBZZawZFqgwaU5XkiM
LwZw90uj5h48Ykkz7Y76aLEWdwILWRcqTXVXXCIPiTbsMn/ju5oPjySSl50Yjh2zu9JAOcTA1qkl
stmJYwImk8hOoK1vgforDBi5lFvcIG9fASmdUPk7KNkWRGIb8xf4lqzLTGG03iscjkGgzBfvr60L
JfiK+NrD8AdCgUCWXtmeqU5cut+U5smS3kG+9euEYbxe3q7OxoZabzYYHHLBdur6fL43ZBADi3pB
TdSah705t349w2I656JmeJtDiu4nF+s/nUCJ+XEP3oA22s8x2z8tGJZbmdy3LY6rh1J5kAhXjGur
/0lmqpPKr/1di8MGmhgMAq6VEtmfbvfqStwvx0ZmSNlaZA1cw9dlvpqLWRsrNfIvcLM/WBlkLB9y
L9Pku1K6V17BVijyYVfU8lEl5hWQYENaW0eMHv7dVMKBrSUix8IiB4tuYfdW174WQpc+tPPgqtUa
rERlg02/Jc5uklFEa12M2K7uf/DW6kxuN7ppyoeiP+Kdq72/CtgcQ7VwEQVCOTyASe56VeQRTGHG
62iOx+HHLFU560HoIwXYCu9JRZVkVPpw5RJmsBvjLaVGRDdCdFNvWkpJ7CJ0m75Ag8keoKkvoM/8
Bn6xSJ92vWllQ2Sth1iyt0jPRz3SPRzzWd1VVkqU/U8f8H1JWu6+j0kKWW7kyquRybwdKDuD/pQU
y9sckFVziHHCWRIh5P6ODxn98uqrCOEZ15qGfcfPLzhieeIst1lKJbSnjXUPJZkOD95BtCMWPeKe
YyfzF/D5qWxyBaMzTdRxBmBkFhHslzRFztG8Zfyyt+AyWyjcDn3bksAqBEEPwWDcHgNC7rWGXPwX
Tl1Lbz399ZniTCOLYHEkQKf1ecE0kxsWbZQJEJyVnfLHLks2aFRwzkosMUbvsaSu3X80XlfRB2Fk
bSi/GEzGLLf830feVMD2AgN/LRnk8l9SHFPKbwD1CA4v2/D34/XotAS1r8T+VhbTvv0DEpki+IyB
yrSmrpfrOdZ6OVpmi5ZBC7VGMkZLtJG/r2MjAouBJO/Uvd/Ab6rt1TVrytfpVhSj+msKOiQxorfh
Ubd1sHp8lRtrUBwo4SXb4IctS1Td2C8f6DxnencgfUHYcRTKXTYau6d3eMP1DXjUZ1Y8VBfvNX0Y
8sSzEp/HwoI5NftCaqHLjy4Cyu879XY3ISI63TtsZsUVUQdxT4QDcx1xAdhq+GL/2Tkda+GY2WfG
CDWF4xnhBuBW+C2row0sZSnGYoUrofCMc0aGOO68/dhFELL1BaVjnLXoOxtX4KT7AQt7aTQEXBhF
0q3JUwBGdrTwzvNmRIiVqoSscpdWFDQNWHXml9EQpR9Y1G4PzXblUx9QU+18oq9BpWfljQREIXvJ
o4n71hS24/tHhnH+qlgeotvzN+/5Wdd8sHcgXW4v6Pkc2ddz5gdNWdVSmvKP4qUgGGgKq4VaurNk
wsJNgFsdcXYGVdiqRcEWjHGW98mkwh75/cWWNd7hUEHP23o4/58/XE0gvq1kF4WFmBgNP6mxoQL8
kut0FCtCSpeiZ9sCPIPC2YTYFV1DcrggiT5hnWN6n5nm3ivpG4DwPwQ01g0rttLwP6vWrLOd+tGa
nEzs/EmFyXcn3fXgbVN5iMFuBM4v9slpK9xwYgLSC6+Ez5kCDcNsj0Dn20z8NQJw8SRkcZa2Ynh+
2kb6XOGDo2zcDnUqh25eUh3PT2G5NuD/25lDY7oeB/vb0ceEOwhpk9iVxZFbB/JoMwvedZ4iBMpx
oAI+QHos7k0ERSTnVuFkz1rkgsfaz+nhBynUkkM/zQbs9okOfJm9HshzIpd7xRlwvbJgrKY49cYA
sgjNloiPoKqNiypc4+C9bJc1xXHeBRzHnwcPFnP8mfMEYe4sGNrkUyMTpedyWMd3DI8SwO/y/JRB
Jgrbx1DUpIzDiT35sfVDrCiTAcFOYEuYWuyWJT/EHTCOp3p6lG84LQAPoSEVRYRMuGXEK9NQu4sN
8/cBkIBklo1SMFCrl1z++s5bY4zPuLSzz9RQHMM78Ups+ErE17KP+7VJcfix9ViQ9Y9mhFxQYFCg
g6rOKWlyAwm9ar4YnVz2tPfOkJ2lNOv5bz5DzC1iqJ6MjUU1fTwmapAVm5Xf9ctsN0DPX+gGf2zN
UV+U4I/z+nD+x3qgbRH/LMQ8DOIBtUYEc8hpGgX7hRaSTD8p81QACGjf7Ins4LqNWC4i5bitYOaY
pOjkXwtMd9uj2JjYKC74zqMFXfQkSYcy9LtkFPHaj77nMZCQng8wcxgbCZl/Pu5axVaez0dGSTpA
r1koNAB3a54S3FmmezU5VIg4fEQSB0dKJ1hAnp4jSjatE7Wh/sEmevQTxRoXzHSfboq8X1SWYQAH
D8dhgDX4TOYMaxgkCRTbaw2NODTWCRPrPQyJfzsA0NrShy3r7V8X0lwlwN/RWLP7RT83Kywa6hdd
fZuyiWisUJaznmFADWRc1bxcY+3lCns8GUSTOwnaK3zPqUAqYouiSox7F/UcVDGGoStnuuArRzUV
CWijk3fwgi1MZ/wzes5JtENkIWrcYNnsUZuNFuZAZ3IT6S8MEqm+zWmx7+gEeJXuhlSY7pbSMHdr
0uRyBKRQe8Dh1yupRGxTAWyDf9wNs95278Vq/65B0RwhZEr4ksjsmKyorrvQY1byjDyinvEbzpXL
JqHguM2+tcXjx0v/pEz4g7Q5rmWljJTOnZ4LJ6G5JoEzA13k8+/K1fSUY15cCfaJjXSfupSvQLTo
xuN3kItMgzsq0DXZdyQiAVhrxDc/7Lga8UQUa9JtjRmVgoX6iv7YzrgbPz9gPTi5NRKAdrZEhXov
J9siMMw0uevDI6PtE3dJiNXKW52Iy9sN68lXqA+9T1Wn8Te53FJJX/hLdO5gQ0wHGnTRr9EOfQEV
JCzODMLsHOOSLhllXYUESi8nHSGqd2P36FKbjq3WIEcbN2ft7U1bPEUKRSxz/cajyOaKDtK6j90x
gPDzfRongH+py39q6/uKrIe+RKzn0S6kCNuZfVo7aCGpM8SdNfR0ESvYFR5UuNQpRzk/qB/b/SWN
w41yG+wOemYVbBaJa/LuiGXX8n3kQhj6sJaoq9EGJHNR0W+n6qmGQ2aU0mY3/qC2Xrzpol30RjRC
TuRkW0Grt5fccfpSYHRZD0L2+OuvinqtuKjmjyL1snMNmW0cfQmGmLrUpAv2ohqwO5D0FHCNNDLX
Tdf75HqCnr0O1bfoO8sE0d8VC7UszW6ptFKtuoXHyvWPYH78WCYlmn+Rn8sLNBqbcsjkWpT+f0Br
PbB7nzFcbQEjlATPnFhH/G6Elvv0Sv3ATmSTmEm7Jl736F0QxYOxsFqf+fSjPZJr//lQglDG6/Y1
KW+7PV4dv1RDmtHXnSkBmvNC+e14CAvgw9ktUvCmN8izXp0hX7spxrJYGy1z0xJdwdpCqm+mDxql
dCaGzyWAxon3Z4tYs0oVV8Tyxt5CS4PDwgadYmE+t4ZtPXbCfCHqetXs3oB+nQRtM5/HFO2iUsNV
B2qKnPqwHbYRP4NsPeGf5HiUzjbOb/F5R4aP2icqjKQ2ebMJzZ+aceOi3bj3X7Z7MkUJfg3PoxjU
gmdHeAfKvWlOl4fEzKFbqYVA3a7cKGzVufy6r2NLEhdmSGuhRtVuT6aRBBzX1Go4VBjqufhv6l9f
NnDtyaO0u776CrNgignOIWFUKJfbmBJDcNATYax9fx/hv2C3oNJCojlrhnrdILb0RJwVYryfbJg6
jA3mkDh4feQvBfTZFz/0/yp7fL5pxj5tiuIM5PlwgchytZsmIEtf4bMqw9COZUfcsCovVsBqR1GV
3dBQEzKDDHWXnMJYTUPP1Tg1jjTfm4z+MS1OonArxccElZuwX4v+7e/b51lrA37k7YB5qD//iIUS
uHSVnbAYVuRBKFuBH5D2maA7VU8pZoeNfUlpPC4vmgn6u3VX8Dxk004Uxn3cDpvojSl9BZXPQFLG
1GIVKAWaBjWFX77woJfHi5HKHlYfvbW/XiVdEGqrEJnfuets69gYOWXvm9ytp8sKZuYxodnKdM7z
G6dJW7mq5krVnx2ESGaiyIneRq8kpn4WOpe0TPoiKE6aCtBZZxvv+mklf3bgmxvBVIWh2ofwOeh5
UkBcCrCBdFpKVnZu8E91Sjfd8FKXL67lRuGnJNwfulHzsQrwp3vJzJGYTQzGHcrhvcfvkmVA6NP5
tgOuHHntr9b4zfgFLf5CegbW2RHyur17B6IISjxpztysW58B9Ze3g18YSmlcLJXNx44w3g6ymZBG
m677lAWlArs9Q6RFpK3zr1mP9/9DnX1S+CITwf2IOsDlOhLIWGS6YyuHTu2JlXIW/Y/meuYiMwZd
e8X4fOku+M8InDQpKs/V6c6tnyjseSGi+ezj2zi54oSbMtAOe4JJKZLXjJtyFDpISK/4Y7JWKhjU
BL+mA7jQpo9o1zu2hTcl4glt9OSZpaHwWrbPeVihzvSlJRq9ALWKpFcVlroA18yRESawz77q4Bdi
00J5/pEr9pkBrFWI9ESg76KIEc90pg6CCOcBgy/7REGFO5H21s4IhOG1Z1nkH/Db5KkweAz+1ZLU
Xiq6jOFDz4yn+okl/pN3lRmfzHh/vmlKlsjmJpeq9Q3x3sb/jmb8rJeKG5+/AivqlnOCtvw73e81
77iz1flTiLkXAWbjhb6BPeDAo1LJuS3vt2tiyRVtbRmtzbtM6xRuoI2Amwo4BqLglpLbgqGQdCuC
FdK8WidSlX9alOrVd5oPM+oRYn0aOn8nvWRN1UKYYWs0iCA1sv8BQNoD11HTG4hHUCGKwfGmFt/h
cYrnNNwuyqesqzqDncLbRtbnPRA05ZJhYuChWWuQ8eEJXNBo6tRvIrIrOqh5NR27aKWhrHGxQrfA
8osDSTxFXp0zsY0KSQxq195O1iMKTGWJWjuJojwLiLqJ8uBbrS0+QfKNtBLd8LhcNAQ4S6+bPnTq
Vad8Qm6kPLdcfPWH1og/yPMNmc7ziha+UzpccDfHoAAFt96uKb5vzVLWRgNbAM4EMCQJW8FpuUSU
A8DzG41KQlmj1owM76z8DWYa5srzFFJj971UnKXiUIzYIoL+1knE2hP4AGmdkXuUhOUbE8IL5r0E
PL1pZIotIFA5E09uBDruDQyp8ErRJepbqzI+qEVR5Xotv9fsqIhV40Zu3LGlAOoIoNLNUPOzq0Cz
S61PanwAhUxOu4YtBeB4qPlbmAeFBl7cVPv6TzQg+qbMSaYE7uJzdRz9n8oOB7ui3uqFZlAh0r38
hUyNJFLWBaH+GEfhStpTThT+/De3KOtCSLV14CqgfexmoWmj82OvA39rEHXvw3F98gB9+55L9hpS
fldQiqGvy9YsQGuSttyn8YrlOexUY+/SOdxtPPSZIZG9EhwNANKIBY5SDK9EEnueG72R4FTmkQVl
Isv21mEVvNJS+B4MqJKsUyUTIDpLjyX/Nkmqq92GTrsbbTADvTgjdNx4Jq/rULUuap2w/RzRBdTk
vyywAbmxm7KtdVmdazPxVw6egXPI4vVCFWt+D+KedXKdBJz4xi1WR9AwZCyUX7sjZOmVkV4ynLQl
99hVWsM4vKVdjPCvj0oSBJvvGSOVDa7BLlV2idSs+GhIFiV4Kzf/7mfK2HQJoq12IDBoWQ1EhMex
OUlfJDi6yOpnFkoD19XVYvpXs6i0/X4RPSM64DCBYKv4bbU6P17rph7EUXS25jeoGwszyaEuk3m/
az0tdjt8PbscqunkWGyJht/djfZ5lQ/K9FmQ4KMwQ02zdlmg+mSbr5W70Y+J23cbd+HOYUDPhI+S
1Sln2ekIEFyTJofnvisYw0KQgSaeKgHQGtGzT2/scmgP1PtfD2lgB3vPY9k9Ek2Zo72+4wWZCD7U
YfgL9lvN0L1DHKPiA708lZVhegduGc1ch705AJHr7E4CoGhUuon854xIdJq0NPiMIda6oEBV4S2T
kJFzuoOcUASaJuonHn492Q0TENiCROQGbS0GpqLU9EJaEbVts9t6IW5L+fb5XjdDzyPsh3f1swkI
Gq1WreW5a6jfJ/CfZp1s8IUGM+gHZR7Lkr5UKePMw01lizALDIHgGwzYoLKTNlxZGh5oH9XOPReU
Pc6yi0y1wUVE4l8N8fnu17B8HWkbwM+JwPt/bmUE209gxXzaBHGALijCzl7xl1It6TmBsY9VZrmU
9ctNyXNEo/L3No4B//Jxi/s+iNHZoYQVxKLwrHl9LBsdHQZitb0EkdRXdKZF+N6EGjbeYWv4J05l
Yv+sd3UPLgIyELYrciyOLNRKxxDCkzNXbN3nwlHsYsji17l9lpjEG3/TvxqTdTW/hZJ4bD20nA6D
7G87BTbde40nmymZyYwTP1v14NSG5LcG8PWPXHlrsuLz/ULcQPBtC214etdz+XWz1vH7Xw0CX4aM
YlHGo7B76O3v3S5bu169G2MUxd/NdwJoqvqxtpEHnc1pIwXk0k5COtq8kjAxlBEgyZlXDL9nOnq6
73h4mxaPtf0Agi1CulVEmC9S2WnCl+A7ejnST56aAgna9fQV+ytLgHh8Ckq8MczTVLWUNcUWbgyY
pukPazS0GmQ8fBAkI01qYnQObeYNGPRy95RsxEbHpCe+iPGf1E6VrNp8E6K+LfursWcUYgU2XN5h
dc/K3Crcdp+u/PTishWVBbWokCAgJD9VE7NU7CCKuT1+0GfLZQrLkXtKe0sPH5mfxaJBXdou8lpF
tAnlf2PEyAqhscJ4Ig2KfrfpqCas70gw8gyU1AFnsDaIpyBwkqUHvXoLPzZD1LonwhVhuZA5uf9B
iFUMRixSB5oMb3tDIL2qsrM1DHYsvDFffb7h4Z9DkS25dw0WFDvr39E3oHdV01IVAouvZhUwAbHS
PM9D9XclW8aI2ZBm1d2Q4gnUb0MCbsUf7vEh6uxLRXV8W2v0Lxdz0RiGAYFjmAi1hVv0IiE7tqpW
kMR92pb5PzBTVZsaHChS0cR5muDJyVfR7oUqDZhqpydMWegFoAC354hKis8Z9ipQfbm7KSwWffnv
T8EFKa4/2iSYGn1iXkQyFLoLvqa/7Kk4zJeFzWvSDvepGvtID/T4ds9BJXavyKTj2Q2sbvrQjzuz
UDUjAfQ8o1cLqqg98Sr2hLsRfBG5PHZkGnD+LpSYZd3tNYKFR4IA80P58jytOtqsO+V2u9PTioCM
0X7eos+V/hbl5ogmruvvIOEUfHqjB9F617/3GsGKDdDwwu4aGsSi3oJbsoljE9+C0l3KTmzQiYiL
frExkEf4oQFKnP2nXX4JKJCJqzehkXLaXXi9nw8TK2Ch/BTn7iNnHyZpaZ9YNPTNwBfTHGVmgkPS
Xyh1CYjm+IDCfhB0uDJOhGjJasWXtYF1CXh+qWG+tOM8kWKZNM+5sOBXqIP6oom+Ws+iYbju+QD1
7T4wTknqse+dLoiWI5vG5yZnxduz96qL6TRVZIE+MqnQrUR1owwVKVJBtya7WhIjP7BUqfm8STmy
D09/BORWEXV1MlST65MjCj/NpxGv0MFt0rp5n2nvYYioEVBh9BLC0u0FbMANj4uZbH0Pc3Rym+Ga
aXCDsqtCWGKQsa+44/60nxwM4mIZoUYYJ6ElKka7Mblz9EQJM0NBpdk0KxHgPhheBeTk00am206P
tz4GThTAdnKIQv2tyWc5R8CCHlYYY5R+n6QiCqptD8eciDyjS5ICDltf47azC+EttIYeFDUCFGY4
rhoJcZ/oXW1xMdOkXn3ICPxaWrHHNn8CdUYpb3jGm74sYqyIyPYR6PZ1hdiB3iJY34Zw0uEpvEnq
pFWn2Ex+NiCA7yprIPDsjpZbyEfmq/FAVK5Q4V2oCNivSS2OU7WnEOUKkcl1ZqFpDFyyHTU/WLfn
fwQIbD/SQVXPaHdZmtfEXxToGd2KtrQwYRO9lL9gg0DDAdoimN9x33wTh0r83fKDGX5EO08bBaA+
igfBh5Y/3HUe2lNEyafZN045doCIapD4ZbCb8Z92//IQqLCY1ob9FRs8SpsjV0oBL7SPKMwK2T7p
GEcTyOsRQFo7BhKc5sWdU5VBOuLeoACVlp9w6MPuN4KjalYDPNIukJTKBInoRp476CVKFKrDFm0f
fvTztWsdxcCjZddEgBBeHk3ObssgJRtsKBUzjRBcTDmuhzMLE51O1xCYXibVLS1vFyuBFmssC+8z
UtHDYZxK940Og5wSU6OrO5swz/8d7sqQ/r9e4pvQZlXWYQr03IeE2kynzUvzM1ZL4PCMZdYl9eaB
80uArS/i5neB4jsyzUk38JY+rerctlLAwTMbkcPdAMSN35ll/stlhL4Qy/HClZWnb/Fpg7yYSaP5
wAO3kaRBTYjI/XMWZN5ghN5/S4jnJMJGaKCgS8aZvHZupzPihuFr+rEpExjv3RpXk0aMLuLQBbbA
pQw6EtqT2tKSNe+oWCV6SSs++JbqWZmDymIsDIz1k4+iP9IKOQDbNLyJu/ineELWFgOJqx7bpRo3
F2+h9imQwWRFmlsbaZUhGNIf0cg0/JtrA7N3ezgLU9aVuOOP3KdcNEPZy/ODRlBvOfJ4uExOLm+0
5CxYANLWgBvPNMXGK9gdwt0aZlS+ApSNFZlA3sLMiVKE0OPBaLDkbobgI1lGK9ooM7z9t1WCTIyT
vn+rxRIkFciUiVAOxALdeenTM9kBprC+PrwEMJsVO/96+c/H6kxRd+TfLyTp1Q2HfMrUHtvB7Z3K
Yuh4M1xfX/8wJh7ln4vVHVOf/nUfpmPD71MIr5cloYLcJnhwnGt4MyWd+sJrOuI5G/bU9R2yFnvV
fxaxdpoCw69ozP9pxZKHtMjWOo/7/2Qgiz7LmPQMWYwIka8T+r2pn8pIlYZSMdAYp1+iGAE5nw8W
Npi66gQvZOg2qtmV9pehjfFerSMqFgiJCOFlfCmA7ruZVsKbGEdcf0aFURq+Grj67YY2KxNIfkm9
co4M+fs4DSGaCy6YcRNFlHx1RZWHVcD4c+M1bUUTKXEoZqdL4sd2tAawyOrb+t26yat0zvpOYjv9
OcnRJUK/GLhedkLDohiYD7D/UjLnPWDCdlpCdIxN0cnXP8mWnTcMtX8sYA6QFJiTKmuPjMELYgWo
QsrDDDaUnl1fAL5PYHXJGSGafLPUZ68RH151EHTMz4ExemMbLxSxVmUL2jpdgQmveLX7uRSQRVGo
d5ZeQ2Up9+UQmEaj+ULHr6bAksXu5L3nWAy/54L3yMLSGlx3a7YheorRWSXsI1LIVi/yUNFThYTu
S/8h/LKJsWUQeC5J5G8dL361OscYaMebGR9czvg9GE84bASvP2e4dWhnSYBpi6NzjlNPdnYFlaHY
WUHUVct1xE85gvuQ2k6BW0MsjdBu7A0lX7THLANagBO5L0jq21n2CK6zybJxBHnteceFqOvTZX1R
ToAyzOjTjdRBC5W6YDD27YagrrD3k3hmtGGbwrExbWpuB0jFN4ANfpaPmQYBzezD5XKIqvzZlklo
TH55kuQ9d3UnbzUQ+pPbGUb//ZaTz3siy7b111Z7wjvFwlEB9HsxG7F14tmm7Pmx953EBZuoRWa8
Xu+y1IBFsqnZByw+FieF9JLP+M/S6Cegn5BXn3sqOLRbb42RJ4S9IMxASanuxy41AV1ANsxXWfbJ
8EQzTQAxnQEuMUKvrV4QnVofsGrgjqRrEHWNI1YXhQT0Df1o2wv3ro3THUM3ql2jCO19XZkxC4J/
PsrdHGDZZN+2CboqNm9l/FXfLexJhmTBUbZiT+nyRBo3vR3Z8Qotg8JFIAKCSfj6cmjdo8z3iV7J
d3nJL2IRylmG5IQDQSaKN4sQQi+abwVuaCGHCIuab9ChgW262qDOQbBAp5/LGz390xAq4AbmKlT6
OJEa+5Z4nAlMwuzEAjXR4UeE5a8+DVVN+YkoIbTHaA1XwHua6NXsXl3wd9f5PRFhPYegN+67vQwj
XkydcwCRVOrb8sn2Qm2iKBGmdJcxgFUhyuVZdGouqeJMyopWC35zRnvxnYMuuycQIZhYEtp2UFho
GXmldShTbTIT6z+wLcOJg/cO8GkfC2nGpJJ4s1pYIeCmAr5sNpl6ejlgB9TCRXoDmLD1lVgPJBvW
ywtUssbuO7alEVyPZTaxjQ5JV57G4de6I3dvssUcsOd3cei9hdSqmGoxL+AuVP3chNPiWscB6AA0
fTBK10GJFFqQ+jPed0c6v85t9TERU60qw7i4TjPsvoE5fX1Lz0igb3+hK7EKh9tZt5oF0AYG5d6f
Ld6iSbh0b5nJo0ZeTEEqR8fpiqMNZDyi1K6s8vZBXqqr3/XtSK8SeZ/1jvfej63wqmcimrBWQHEN
54SrnYCcVOa+4XAQS8ATFmRnQIUUlG4hZK1yKhOGslJG41djgYDHtHoyU0Uvybim/mCwXykwNHH7
pzevwr9bTLBF/qSj3rnrKGiflwILegFt441ntaxCkmELV57PofnTWvk55PpZbkorngYvdOM1Kfgt
kSrdJ84yIaQI7ReBmXqxrOt1j/2EkPasl9UaOWIUB5E79U081fAN8cCCF+TVGyb29iSV/uQcp2d2
HhDlm4grXBw6dKRgeVnUhOng25+OwBwifNQHJw/mMCBZn59xCYmzVDR+fyrD9ARe1t6jvmPr/QRR
kRp2bV+vWIfBAgTztgNmN0pst0llxekO33B+1hAFJXfNiB1JKHqLI7ic2954BCPRzVo5nS7mHfMY
0GftJadBSbOUqkf7R96cAQSLBUBpBzLf/L4Ms6d75v0c9KBHGOXPoHqv+AiS0fR3/P/QsyCxHW/I
Q54vyS0NepdYebV/hS3E4v/TKbo99tGmUTdsBHoQpV4+UmodKcnRJxR/cfg1PLQNoyK/vo6UHf6M
ne51nheErxfLerVTEKqQMrq/ZYZKxBGr/4FUAICCmgrAO6sBHRBi6skX0JGl3IYmaiXMRVwdbhKE
izLpJTeEZwhfhveiWvXjyzy/iDScynXWbOrH1n1ZN0oTHmImcEZmsgknJa+4Oxm1DML2AZQr9wOh
HwUr0Y/EmYqymLwgWa7IPfeRg9YrNfshhfOmmK0WVlpxkOqc8D4yO0SgrItSNpQImsiAhvqhv/f4
c33/WlALTRGlRJgsHZtlI2ILN3agXAH1a0uH3e2pwPbGQVour4J/26UVaxkdkJMOfXUj9sD2AWuh
cuP1Z6Jc3P1xrfY+rMGSEl18zD91rj51jc7zjobChWSUIJysTT2esMir33Ehe1j0mpQqdGags5C6
V6ZfdPCvQ/vMqC1HfGw+7YQm0x2k2kGKOm2l/GmYcLHexq7rZdNZ0LwzwBhgv48PSPpef/8Y0HGb
N1HWJah3Jp+bhAB7Lif3uuJjJ6vCB0JtuLBXyDu1n0sIbGoNYHvrog02AZLrw9JmBHjyP+DQNxVA
SBNpmLY7NeXBX9NASIxpEpy3k0TAZzmg0yC3V4W37lakARdf0GNl/BTEXocaOJ7gSZXIbVsXXXIA
q0liLGBNaz14Qhlk+jMpxA4OE4GvutlIrdeYZiGya59Axe2SGepmW767tjXRnPdnBdmcnKRLN3Iv
9Uds7f/ip5KD7a3NGe4jwKOznRpIWAFFXMVTgCMoMPNxKHQlvOsuf5/dgfEZkvBtKyp6L5eH8oje
0EUJx/f/GZdAd5YT08hZ+BTo4d3q3rrlm8AGiAvi5elOr0hqWPb6/lu1CzAl3sI5y1d/iqhaCfYB
inE4DVnmjL4vEGN2bVED16uS2M4N2uDHPfBO6d/pUml+Jlat0DFLYAvNSaejeN82oZSEYank2nD2
o8lEX1s956XKtlsUqsRBPtMjzlcarvVG3oJZT7QWHZ7ldv+xWMMUvQkW916DJP8sp+4JZCuyIrtL
7YUOgJgBaETnNUdsZE+lqSMcwNumLV+GCwxwibKeceR6SSgZqbtQ5lLqDoGQnMRfS0eYWZ5bMHXe
fm9W9Xjhh3hj8gYgdwHQXVf/BVSlC8yKm4VD+emBO0L/xxuFyYDosAS3ScWiPqbrXfsWQvQVprPd
3oA+xkA7gWsLDR7OjGRruBB+Ozu3PC2GHk4NiuAwYo/xk0jxWTW9QHFb4lV0PU6gzkdr9htJaKKt
pr9/DLvLuup8cpvA8wHH81tjroekLzsQGoZKmVok2pNcz9eoXIr6REJ2kFGzVn/Se6PO5B/qLi8e
RbJuprzCUivhttA7UA7n0vtiLIlcN5o4YrMi8hL+TCgLwUZMe5JyZXpVoLSGp9Z5Zc9TuIsxIGdZ
uHHXKd9AaKVyiOGvnr8tzsngit2YVwl6yDg1gKYcuIcSCOvfu6WmdE0ZyqKVltOj32TEB8FjbmqO
nK2d58B3YW1LhLnKyw9DdL57f8EteYlSL5TNuR5sqTV6fo5OTCpAY8HERYc7Gr9Iq0GQFsHdFIwU
topeAVVlXz1jg6iH/wWdDyU6QyDqERnMKE+tLDiZejDmWQlPUVwm+5lRtGzxYEmO3pAn1lOpv12N
Pcc6dM2DqFW5ttm6epedeGFN7fnKzIWTHtZvxosw2QkMOATEh0JRt0zOYVmfsoaTr5MvuIxX8VfX
YoKbt6QqinpT0HUj6QXZJnhrnyH3IDUX4XxFjossqE0auM2rBlI1I2croYZK/pEWBByDmmHMzDcD
xZNftwfsC1vfNFN0NCo7QN2hvZKlLqqgtP1c8ulK30ws1KyIPDM2wK6AwCF1w+m4qaYGM7uQVqQu
TniwdiAXsAmVq0gFin8SOXOFSSUK7GBQGEq5puRYtf1K0pfmd8Zcb5D6SD7x5TqFayveYbY2sW2D
62UOcyAR/Dghkzx4rg6QVR8nft5znrWzdAugWu2Z05DWZSrz8wGFXEj4mk2hm0TANzp/dIKESKM0
xOwzuOYT2owgGRg3l3dY/qTw2oiXqfSXQh5FZWAF8nQbYH+aCEwMac6tzjoPEg3xJDQuJ01subTz
HsWmgm2jot9Ysl3TkUYGNAVhY2CPRa2Wl84BCTwAXPzjQWZp0lamu5RJdx3/Yts0BNSS8knH/iSW
8BYhtRP8DwRCJlYkENZ6e1VslU3VOoIrG6BN/WayHfc5IXjV3POnSPT4hFPTieGvFzcl5SaN6u3h
H2qzQ6KGe8E7lMC0pFSRh/8DpRbAcDVsbN1am0V2rELSNluKE/8NJn2usBtW4gtIqu9gkf1zKdUT
g9yi4o8U4ythb20KBYjSNhqjapcPsLIl7eYK3Ra5bFJyf/IBmQtjNkHxXySGWYh+/O/7r71EjyEn
e4J2ceFBxkYalSimW1GWt/193ZN+N8208zxX7Hw6fucNwtP2RdjfrE1cSIUSOfcyDrIhS35ttZvR
jpqSKl6XM/o3+puPQkdnzYulsifcy9ATto6CKc1RRpMcs9H09i5lQr+sjbVzD9SXAownHkTo7uEb
MpXWpTdfibEsONNIUjGFZPKWhPhjebh6nZfyiWY/m7vjv0NTghKBjQgY+9tAR/9eX22b00upvPCO
y7N+RebfbN+NF1qdX/Y/Y6KY/4RpOyv3Op0zjHkMRScCSUInMfAogipBG/sHVMPgrHMtX00Bg/a6
mi6AISWrhS1hpjhtI3r1/CF3S0qgFTfo3heboMWl2lqpHZ7pd6zL+YxrDob66g3SqcbHOHW2SGhS
4xK/WDhk6p1wUQ+0jbadYjKLRaGlRoQYMUo4RdP71rUpQ7UgxZE2mPGvk87AsNDkIIUaqdIBUmoJ
wCEhqp5/TAhYIGgoQ/akjB6n+fjHn4Q/VlRJqStQf+u6hUiXJYxFBAYNQV2qlKNrzDK8rvIksnmd
Q32xw/LJMniQ2bpbvCEAZd1+OM9yDlANfzb1JKSdeIYEGxley3Wt59Wy6BD1qm1IRMcJdE9H2gRU
a6cGQ0/inIOqbfDfgMOfIMAGvS4+FQTKfhLiGJhsxIe1+uHz+9Xs9bu4dyyW+7HbZ0xIXa8nvnAb
Jb17Bu5TNB/CJa0fU5VyY1KE9lnKtPZEvNGlUYSfbon7Yc6DM8blTclIq1NBfy8u3GiJ5m5/pfPo
IU4wwx1WjCr8fps03yBBQIDQg/awaQsW3C+IpiQfuMS+hYj5X5hj5j6iQ1wJRxsoQGMUGG659VPM
bUOQ4/obfjw/4IjLL/EL04r4716RyRoR5olkENPXcnmOQhcEGAMPq3DBVvj4LKxHmK8FWjiOfDYd
MSF2MihfePpWaPEa+Esm3qmrodPrtnUuwauYx59T7i/chA5f5Ss7vmDCoEwomjlRPRLS8WY6XrSr
F/BJKv+Cpxc7+L8209l5+xqdvLMjv2lwJHAhN3c5zPzvGmMbpOWdCz6WIG0M/6lgDJqG8OCh6fEI
g1kzrUCyLbAdEj2gvDlCmO6HbYNr+Wq3FR48pWfw1TBo45W4p5QXIAjFYcRzsiGw7DovTzUwGppU
OBKcQUy0hey2YuNOCsX70ceKDnZvlqYryTVVLiM1jXoUlsdXJWheb5CQEuRRcIiAfaoziUVIcVzo
+6PwHt3VTnpPZRerGvvKeLG2h99afFaI/72L7KhIsk0y2ZhcX+JXW0pnpjWF7/kWhX8wVAH2oOa7
bpJD4IpI6QUG+uo6ujrzn3f38P83PmpOwm11LmcA98O3xILIPWiGWrar9hxChPaZCGUTgVvugdFZ
BndxkZaKrYOpuAzHbWIeWLAhENr8WA+PJgQc2YgWjEt4PyyUq8akzszTmU9PpzqsHoi5MFDFUjpq
odASfnwRG2HaxUgkdBHc531ssiwM1EFbEE4ry76QoYGBk6MUvPFIP5npDzvyjkWqMZ9d3oIT1mHi
09caGnTDrCj61DDsKFU2jXcB9m0F52zLFGMv2UWnYRlJ1LW5KhlQLWPUVssbopWz1HrgkRCWbglg
CqSQchH0aOpsitrfKxAzu3FycEUCH9RSp2rVaOfA9O+HzRwnWEuKB5bVFdT79AbxRspRD392qUVY
XKc9amvQ/aDLUjan1bZ8nkAwFGB13pu1vaJlGcUVdiOow8gJQJqU4+S/OHtCKP0Ne6zeS9NmSGO9
84G0MpdQhdHotvt4BKoWHidfn/8eKJ8Tbjf0cmsSa/yxRCWZn/YQIiiB9q0omGG3psQADebjN9zv
QNXTClIFWvMBY5lNsdAqQTFQhdEhvc0JbU8LZQxwLbkkX75XVSwQtXQPOhTCp9YFGiDHIJi9iigF
Xua039S07dZTczcKuFGqv4odIg4k6CADYKwTzCMzmNz6iZ4JUm2syK2NWwKMvYsfobrTEwT2YUtK
QKodiWb3tYKxfdBbv9akfhhWNrz69UpmDki92pKvM9cGDD7Z0aG+qWmje7ZlYqsVoXFAJe0O7zLj
Xt4nEFwEo/QKHFwV/od6i9ad4D97wk09bh88IIC3VZbL/FJqBVMqeTWnAeDqlC4wwSsmGY07qhOC
e35Gib/fdHep4AuD7w9wUhCPdX/fqDGoozBxJ893xSbDtCTw5uD3JxadiLLyo0FZzSOyXGMvOJrh
mp3hF4cWL5sRozMmPesT3lODmoLCiYswoMi3QXRIi0ol8whgkw6O61LBcNx9L1viL3uVfdQ4inVQ
IwQiWIBuVYjuI6r/5I+lj2X0LmCXhliHh4qIQYOF3bu42IfkK9hcqLkJ9pS6DWVIodcBaUrGiXLf
ZJ8eiJNdbAXFtMLVYHP3vGPRKLNLfsKAsDbeNjifwBNr6iXliorrvcG09r7gLjgvB/iyjlTYK59i
BsbAJ33sEFU4FxmAOhNGlhDOtqghPU0N/x9VK4oGgCqTZQAqtxuYkItp6MlH/ghPiJgimpIJDmlZ
ueQ0kZ9rRbhYXIGM8hGPBNzPSkYX7WNW3v2uD0RC9RSBlUvtpw7tN7lR8L2jDe9ujLnJhvEHM8fX
DK/ibUdtgGMeWTm7UbVUfI7hZ9UMVmEQiMDopMOSH/hML7uEL1iQ7K5piARM+IyNdDxSmjZI+lzo
0rMjWfaLPuxVmJmjSHlK5SCqYqSylb0d03GSsU2UZkQ/BKUh9wxRJMe5H1hL51ERd4g8PimFNYJj
g2dXRH2OgHWA1PGUdJdZv9UysVKHmzs9+6SRfFz/YlLeio6l+Rw35H4zBxtGnbJBYnudVf1/1r/A
VwyMNZlrPcxrpCXjL5lVbPoGWOqpx4o9G81emosL6M4JrwCGGQcT+CcTtu+xcEKt5aHSTdqjNz8u
pcQU6Th5sSyNAlj5krCEM57uizE1OrI5qJCT4/Q9Rrc5atVJiLoEExrZRYr2hVO44y7k7BeBq4iH
GVxJ9uDsV92/0838xurR7wRzJ6HnxpebDx/+4tBnJkkIz4ffU4XS484/qZKGlRGrhJdyKhD+ouB7
bYUIrX4dlJHsVBYArMJf1wG6rVt8tnG3mTungDSFbiFPdd1zDKSeHasAbVwzNGYm88Ii8WgOupYf
ucybLgXW/4mIASEZM2SrAvjOZ8SSMYjtNV4ZS3DxLwmUGtqXHllIsS7J0Z4zg+8zVlepCvX0VtM+
A46BdViQ83ctv/T+va6Da38orUoIboK2rRB70+GgQNO2jg3Grh0d+h8nO+xLyt1zXm3/oWyq7NSz
aFIGduB4OYIPbEDMUmDs9i0ER/JmVoVzdXHOLe9oQV8QfKBTmiFrzgLLJ29T7ZhNC8COsAYxK3b2
acxVvauIIzNH4p+Zcd9LS47bYpl9j85MeJcCcj1gfGp6TmilJopJFnOTJnsAytoubDe7RNte8vnk
s27wLcfwdprqLnYTbLjcMzOZZjoCEsMJpxtMKNxqlsFDGFJRJNUTAaBhTeiTuJixvBgyuH6UVGFn
wqKMuS/cLatDlKnX7iZ7BPemizf0OFWQsOsRls36VIWjrC75DOOj0Xmk7F3inhQP3LE9xG0BVvNn
KjoNFO7fC4y7syb3NjWanFldK4mlPimS7Y0bvuzQeuKdFALSQ5MlWTCdI5pRxFw/FExYTAETPfxJ
j/i9d+vRg/y+sHZYO4PPY9B/dg/vIs/5O7s1RynsLQ9IAypKM5co/n49CzAOCub5VN3UaWH8/vc6
1C6MgO8Rq/4iOwFD8Hj/giMiQY40V3kG/HU3MZK1iUJgb9xyPYPyergYY38jXiiiWukkwify3+vR
S4qQ/NRsQOnIzorMxGEKD3HMjvSaq2deoydbkf9LVZcVcB/TjIV+V2e/DlPIOi+IL4gheeyAh+k7
yvJbmDOXUtu/pYuE5dW5806U0/PUom/s6pgf3+piTYetP4wzAgd5vC+dii3mMplITlcBqmLfF8FW
kaQfrqxwTRbHruX741Vhynqa9KwawpSqNO31Lb9XhAa7SKhhToDO5ED9oQQahk4/xMA24zNpxOhp
uBOK9dbrzzTMFWerzgeUoJu6ilUXUrQxSwY1joVGUeL26WKhkA9UKuXb1XK/x/IcZ/uf5q7QX41x
ardv3qJ/3Kf1nPx6muMNjXPFw2VhenOinzrJth6/xoyme9+paPniwl1LgOfY2BF9XxcdfeVWuZJX
04YVMBj6UYvqCJiZ0Rr5be9F1Yvolynhfx4DLXNIgR4PqhHCyOtL2ZN/3YKjYuCSGTGKiClUpgSl
HY/X7uZrWpROunTyBwuVk82uaI22Xw2s97iwFKOmvBpV9SKcd9n6TPf/yWmoxpuTXO+GEqUbuuBq
Omkt1D35NV8lN/wz7nS84ALTHOK/L5+iiDFR71pHp6RcmuF24d9nrKffVVHV9xLJ6Txr3VDHVRWA
vT6J+iGuWMB1H1j1nPl6LRex2Pj8G2sLSbt5+9CV4QR8JwNMf0xrzs2a/Nw2iBpf0xWYQBzxw8Rj
mFyzeQSv3YQb6XvNHceDGFV9AQsNjsKcTWzYlnqrrQbIc7owPQcWHtEcmLiBFnF+MccXMtID3Sqi
P5t5cF9ERX6vca8XQ3+KJ3/8QyXqLRR9vlNShEa6nFJdWoaJ98PTVKihaFB8dyd+NJG25tAGkYAh
e3mhgz2e91UNF/q3AmLfBkHSLfyJ3ot9EEYvwVCo/FGrgpIbDJTumhKQrfzvzJmlW2qnni8pKhSR
4x+P5ssyGpkjNtjQtFX2Kr7m8OiOKgdLxYCTKKj06znEP0OfQaG6+HusLApXuzxqVK8E/iGLauFK
zFHIvFffpKlhoYQoCyYznGv/fpZoXWJuiphMH9a63ftSoBiKKe1ZrqT738fwbhpXbWXSW9Mwpw7f
emXetJ5M+hwGiVamJJb6lOi45gtr58ykhynHMYWBZ51Yw6JGHLfeEyEqtXffOHLKLZjpWCN34ffB
D3Cero2rVyVvv/NAzd8XBvDxvsQ+yaw9e+wGGUTdFrpaV8tCna3S6yAI+yfqWQKnYfXNy10UWeoT
FwcxeHt2BbTGLNlm9H9kJ1jtUB/XOV9p/hPSFarSai47xBW7B+Z82u7ujv1qT9NzEu4FXTaIPpSb
ZLhAfRHaVVg863sREyRD/q/8kGZ+Gsj0jd07B4u476EOxYR1oLx4RzwNjdmc7OQLI81sj0RfsBqa
q1zKU37g8nIIh0bcmLdxxtmvnUoEM58sTDsjnEOv+vAZ9MGLJZmE+5G/M7XuI/duD+IktsTqzCRB
Fn8WurlZCslj08Ei8Bx1IW3LiBsZ289oZNYXuA3663ynfNcZ5mrXvUvknMuaHbwz3NigDwNKHapS
Gncqg0jE+1UUwmAsekUxb0bHug4DoW6eGx4eMEjp73ajZZSD4bPBUu9DOhaT0/DqCwKbAdk5zLxI
98VQ5zftU+VB0VB+AScw0sMFYe9F4p705oUV0PFZdmDryn5h4l2Qrs99zymMLAggvFkRPBGzhU+1
s/CM0kzN99mAX0juZTP3XfN4JA7JYCENWLqrb9LPU8xOMq0YVkeZidW4zbr6HQsIgFSSU8I9Qnxg
XX70QPGULssW1rTkdFEU9TU+Zkq+57BLqr3NSw892GKb0MOwLUKnpsZw/0Ic0CnmsgwnVo+5qjqB
CL6RN561aPJEuRURZFRD8aCby8LyqdUT+6/e1FKUbWYGKwmK8IdV3DYqxp/4WzR2yevanRy67MrH
yLudy6OOiq8zKJRZMqDgZqpxS+OrvcgfgDB5JfTrHHYW0ErqibWXC9S0fX+tv7cganQNbkIyRg+7
nx9FAoOMvnpY3Npww4B6WuzpTrbbp3EO2BOfTfJ6AYLD0OBoMxTjm4BjnCMUuUtzvF10QyW9awY7
JZlauLXyS37QE6bfmUWeHeZe2JNbdls2cBcPqsRSEM/INWuSSf2YJMIyMGcPxCaBHRarZqAzexWr
leuZC9M2UNifvQIe9xKDxmZbsDSa5ROdYcTCMf9I2arq6cESlbvSL8nqItWaoRu0nKOgZ73wEdAY
qGww16qO9mjHjcxQ05LkEx1MuU0IUvcbO9ZvX8i9+03cbVKGKcCGpkWdtfweWfCyDQZZr/q08xd6
AxZPscfYsvq92CZShY0/cNS/yI9Z6Pz1zBf7x7iv/1S7vN9TdjmyQp46EWBa6VYWNwa11dB64V4x
HHrlRv7hmDPmG8M2zfsaO5rYMUm9J413ZzeUiHrEW1m2J2wRom3NbMRWd3tJ4DiQlIIvxfQsV8Mh
4XxS0+7e4VOaAucsxQqmcqbIWindrAM/tb1qbEj3Cguvi7+VQ/BuLvsC5IRVmK7hqD+FDdtVxtrY
hDZlqeVdSrIqMdSH4duvAR4zGe+fgN1jFKYlRxXxRdolnDLz9yByly4gNk64sWJPhFokreZrryfl
XH145gUpRTZ/66qRSUpqDNykhecD5+GQpsGm9H0NETgpljWlMgEkHAElaIl2VsoWBWnAvFQjrFgN
YUZj5/SH9imTvK706g8H4qee6lA4nfEFTsw49xPgcj6DzeN02tj7aE8S7zosG3+A+uxNxV6rVHEa
4+2IwsUbjM1ZovekzhWJCwwhNdlQoWBTKg0BZEt5AvYCMEDGCPjDKMrxNiu8WBgv1pHZbW+y7VZ7
Rph4CGEQIPX9fVJQH9/FdCMJ00Zr97DR2LfyoovhmVhzyQ2WZQoZ9FI7FPWy4UKYsOh1OW9cbotP
NecxRvEv7Om2B2Bm2vZ91UMclhEFyUJ3XQG0Gs/dfkjKSGze8MB5qJSdnAR405vVrQa4xCGwMSWZ
qkZT7/WGfMSHlodYxu3t6QZJRVySZEgHj5St+M8oNUQr5lP/qgAUFGYyCbkxXDPGU0oq7ilD9pM7
J/P8wiyncYHE4fQ0Tp/n8a2jpujjiO5ixcfqnlwwlc4IWUWN2ncczGa0qv79iFn8gWAMpPh+mo34
WwVEuw+UHjAu5Pk2+7PqQmG2YCL3No3g1HNlcqoW1sTJ+szPZCunPJVk92SAjlFM8UxeHNgPtNAC
tZdqq2Oerr+EXA5ZA8sW+ddWzpk4bVC/N4dK/hVW9flQmonOgjTNpN+TuQKykNBdyYKACPV/Lx4E
qkJiSzqzICj8VAlfj+m3bDHsYgKuKe9UUPRwkLqY8bIlKEie6yWNbUh+ywrtFHWUiUOiAwaY8GUb
j/SqFodUVxIcKxEo558r1DvjHi0N6SFab+fGkm+UIpQYW1MnJZUb1QWnlL58cqU5z7NqKNYSfSK7
OhzTr4kdi6+HROV7TZu2eH+EVwWa9Zvc0G2rxGpPamFNLataBZsx+voLHUGR7kXy9Na+B4liZsaa
+M+Xs5QHActk7WXf3WQ19DeqHeNqHnKewDKRFSwCDAPPTgaNsFmayGSA+D4tETIEsXwmd7upWfgb
NhRPWYIIj1ey4iK6mv6Up9Aj8ykYqXygzxQ3g/z3jfpumSJo57i5pmRbOwQ4QeD7fQFblnFtT0Js
nMm05kyxRW0T5iEQ6NHDkaRVIwzTya5xLDyJ3ilG+/ByiZgCeaNL01aJUtDb2Vzp2Dctd+LZOG5w
948C60iwKicOQKEwPwwxoDCZ7H1f5ekUFTyGkQiZ4Tbib6ZErG92v7U9mjpLH1ZmcYnMu/t4VoZG
hjLNkTUaXxP4KJkdh0+HLI+rXlY29fand7U6M/UQyT+y929j2su177DlL1VV25Es3nZ/HEx5NluS
kgupzy28Wg7ijXUd8sI/H+ge7HROwmO0hmBZ0Dizi/OgdHsHPUT9xo9fFknnJEHLQbn23uXge1Gt
wMK5lJz+VwgHeuY+o6wFNtsvRRjBsUOO6yqh8/nLsYmOn9spWlzJO6gRyTb8DYvv8CWtO0vhAmxz
un3dmQmvZGOAIgfhXy0ko+2wDWWarrdh2914lgLdHn2BoF8nsjDO8DXCSCxHb1kpvo7JOKSdJiR/
lJTNLjgojCKwOadVIGTTbYjfyZ5ioLdegee2C7HDGXVdKU5l9uNOziGfCdDbcRdML48kyCh/5PC4
OMHydTMlP86WYufQr56KVL2AdvaugCBTBa/7xVsVOBjGfhbHF+j45NZ77XCCm59X2UA5hSf/hmfG
/iZMGNF0ggjkuNhwKY1bSThROCsbP8OrWwHTaBlp8J9vUstZhWypFFX/ZTVEiVCIGRDqVFqkfm9E
cmzGTMMNXx/DhNh4Ti806J1JgloighchQlNB908BvvcdsQzVB70ldR7nVHqg4CVbfgo7KQpj9i1T
Z2vkwQx0LLF8qxenKSjWTTGgt9JRoqqJarFzFiQTiJpDdHYrhLKE49yOo/nUpOlLgO4d58PXtbyk
MoMae4tmmzZ0LtloR9SFtuPNw9CCjVr1ATsx72znjja1mPwhCjDVlYSaMoJNmSW9mFmrjp4qTXhr
Oau3Bzka3E2iCHESk0X2QTItYeRbh/4JP4xQLK8gK61YqHllp8PQxkGiyxXTVUjygxZEIfUcl6Gl
O0h/tx1ZTRM6oBp7sV9prgzThUb1MR4LdGRqUdtHhrEcKjOcXuLGTeoGiarGKfpja9NdtXqUc626
6Wn5JLoTJcDpVaDF0ClryEEJIToCZHC/p6Djld5XnAmHWoaLxD1D73dcaEyzQVYS65rUehOq2iUt
ApxGiDCDsNN5T5wDCYTE7YER1ADymv7xMEsJ3KCMxLCMHqSiJpgBsKXp1sFAMlV55je0z2JImWFu
uRa5A6H71F+6N21ES+podpcVhpFH6GfWNg+BXlUDpEtsWe5gz/cObLGHG4nFAetxDhCB7/c51RUL
0qrIl7c16oATldkNBKnnnnTQsMKoAHEgpgF5Qp2jK6rDBFVTLUuL7MJNjTOvbH6/qERVybv0zzV1
UkaGKiNwFELaBIjy//YOqsDwBsbX/IC2Ur3S7TQ1kX0UOt1L8WXREiwPv8Urk8M37U90UVUmlJlZ
bNsTsf6sIpfSEd/07GilCnjfvaCyEvgQNRe3VwIBg4ZCpiW0x3ongwh/UKT5mFwrbVPV3ZySXxtU
iLjSQM4A0ABWYauUvlbkDGotjP6x57R9EeP3SppyQV1Nv1B8bGhpyrwjoHZkw7kU6iFt1NnHXqBF
aScUCxykXuVIrkiIIRNxjOocV3dvMKDgsLh1hSyTMLYdGghDmyAXG40rnABON72tsLrg9HZ0LiCX
rA5DeQiQKbVWi8m8JfERSvBaaCyRudVWOW3fzXuxd29E0Uww4Y7Y/bi/WQ2nPCPmDUPunxo6nAh3
UYCASRMdqpIpCKVIjgsO4tyN8dmIbLOIoC+cby1OIbcgeRGMgY1IxewAX2meLyHde0NgkAIHVMX+
wN2uxdiD4jVUuEJS0Nfxz8v6ViVyvkSLrt/CMAlCvNreQeVxoEtKvMGAblR43aCOq2DLOXzEQtvN
BfVJyGzO5E8ZCrduqlUbyntP700Ogd6xPOuU6R9ymwKHwxs1okyi+dZSdPUF0HMRHv/fwjIG3L4J
BYAeUxdMNWOabRt+2e2oD7NHXsim88zt10zVOtWKkhFHzSYvexMjz5D4qE2uNjOsWsAtAIYb6sff
jBC0ka+ysME2LAG61QM9zq4XfPJHg5yQSOFYCzCU4vJGKmZXgFhRj5VwA29gKYfnuq+VIXkHZIgo
bS8WQpYR3TGu0LC/e/V8VRLF+LsacXQI0PCcYdtzzQ3t2Y7O92Udw2k4IxmHkOFdehlRxaAzWdeQ
z5faoVQwMH7sopsjQgbiW1JZyD8aSXxUp3GDx0JekNmITRQtiop5yQu0QKOYaGZdymGBTri/VKE5
K6686al3ismM+4XqyWg9F3zR8cweinYUppNwxlwP3cuw5YBe6FKolA3SfR7t6VHM0mrdW0TABU4V
gC/dBtOxugPDRA50YJ7GbRHN7/OUqxWJ5LIspfT19mK/g+ns/lFuxa2lmkOKFGzRGYSFTakdFPrs
NvuoNCy/HI4AI6elNwcVx8pgyMoP2Ut24GYfn87EQrRvzcTDvXTOxWYM/othRP1Tv425F2v6w9TU
G9JVSiVzzwHQ2DVeYJ99HR00yUESZxH/RjKUuOZFy3sOcBjSUBvB6vlNCyWUix5GuiA6yjpha9lg
e8wTAb0LomGe6PLydWjojmRCw41k0JOVmfFVzgGZg13mVOow2auZ4dNNCFPdm2IfTENDIgrEdx41
KHooM2B67Wi+tnSo2AZjolz07PFDZx8Cbm+yG7I7q7Rckwq+M72R9+dy7JTnUHWiJIxHqSREEF6p
wnwCzJ/0UJf2/+AXP/L7/Weua1cD9wR/w4rJJ+SgBU2VW1deTM/Euj+/ouMH0wIk9sE49uG92YYk
sRvFP9i9vJeBMYBfgsIE98UXmYWMeApBo8rHCSTVMB+E0vhm1aGnZWeIxaWHxJUfuv6HKuLV7RjJ
kWEh/cM3Y928iulEQNwfh3oK7x5k124WVF8L/PjtU9MDd5QftUkX+o6aUUpaeiP8JEt3U1hP8Cxn
IigWyXRyyrR0eDKbCXCZ4gXbc6K0QB2nGxriWHGQRhOgoDORhphOjAPRUPGtpJ+FhAJSjAh4PYzv
R7gagQXzzUh0gTtoCzq3tifcc63ASDe8WtQQalOuq8NyV8UgMqNpeyj3t23FOpy5wWTvlAFTMhm5
4bym0pvl/NlCZWAYpKt82aj/h/UifO4FTv7Cffj8n/fSXp21zxy4CBJ5twwvaBCuWIFNvuK/GNli
iWZpk6TTWTp3/5nFdIPB6IelGTWh/sHeo02b9cggYM1zMz6y1HCcla0tUlirWpQOVXGO/3gcAosd
nM1UjzKzdb5Vrm3UYdBLwitYTaI7F1wTG/xYioD5Km01cnJgtbr7ch92wTvOAInXnfPsSGn7Leog
I047GQB3m6ZTgOzpZKsGywrqErC+/3j4pbQsX9zxV81OnoD4piLw2Ja78rI/5+0D3JH/ZLSgYckG
SA9cchy4U8b06h8yYiNDi36LVpc4Hi1/2VW5Gd2tv9BnNYC5MxnmKPRUpUbi8EhNEktkbqyUvpPL
KN/yOJE/MABNqH/fu3GOOIYH499i2SuGZWWVL5SvCc6lZGEkv6DuKz8ny6AMzhp+h6kGKjMjJNyG
JWEV1HfGKPcsDRLnjbq0PiOtuKCy36P/kVy75Pf/4sTcsM7ydw8hN47CkJyBtzntW4QHrq4d2I86
/S70HqTH1kQxyFWq9wuEZFvjWaOFW8d7V8E+6bpXdHSEquIIj6cM0CaeOFWNsyLEXAyMcKQaIFDO
GPTJgZc3RN70gpZNklOkA+Sq8U3CXEfFIsoo+WgAKvp8U9tyOYbiZYHF+Gk3lFQfeY7mqnNBpmMp
QjE28eisWVDLY5WiyyK4TXhhntY8RY65V3mS5v4vTH8jcAqY1huaa5fP2Mm1JRpl0ffdX86odbUo
7jNvlBZ0UVqVUGJ9oBwdokkg0yeI/uMv/CwZFvPtI8wzK1+OD9og6UcU+ALpBuTUxQyHnE1aq5kj
ZlcKBBrWe6qDYVRjpzWRdtiPC5RgAYleodCAX/nJB+ULOXgHQ8S8CHOlCnOjfu/MM7L9MmQdiTUE
clh/o1ND+hTEip13gj7s2JdNCXCRnlID04SsxeV6loWbwG5fp5nyYKUbcbi5qEfeK3wPEajLbSwH
lfw5PqH+517bAcLmAuU8JEduc5wMploZHxc/Eiv3Z0XFwoSOJmif4jonRtiXHT1wYFa5OD52/tTt
Og8Nc+7+arpIZxTkFmsDQqyALGInZEGuwm4oZF8kwW3bfD3gdD6jhCWpoGWhMZmw+GjWAoveldTf
Fw9kuaui+LP34nZEq+dut4sLgM1yAQt7yyZ8cPWRF0jnAtE2mN87YWASt+VSbm+o66eE2BJ/2VbA
Rj5xM330dVurQ/rUqVo3ar65sZ5uym2L7iAtGkVAlScXNe4h9Mi88SpXwC3Vx1b7pVuipsYnxzaf
AH5h0B228I2BARWPfI4xBRb9RtO9Lc9jKBmQtblv6KuE7vRqBPWaHwbK8V4g7H+j7zKgJce8aSxh
r1YEjJ0qjPstiT5fmw3oHCxNmQX2zvUed398wxLy76+PfMGfOSikrUsHCh3VcH1lu5M2DaxSbGqE
ilS/CtRKuu4eTUXmXMSpzX2wUkhug0qyho8o6s8zcSQSW2yadM4D2DswSsLEIMH/OMTxpQlGbXet
GolReFrbMePO6IRmaTcTDisy3EvdfCbHdBNlgLQckDBpirtFOSy+yWIdI1ejMPD6yT7Sz9MZfsoU
9r1vt/1sKW9vga1tIg/2ZBf4BZeTt01An7RcvIworhvpS2UhbyUa6+abq6dBwXNyben0PFh6OFQp
FoaufVYU20XS0lQ1Go7Hl7b6Nte1ncqEHygEtg7OqSdcXpCSg+c0lCIIwqyK1zqb1yvTdoBJQFUL
rrFaFhSsqTV2huIchPMSGYRO+UqVOp5tYl7pziOfuR5ymx2lNW+60v4V8NfHdUvZe5aTp8QTdivG
/7Y9/mIwqkmzZ8kAr/eQ65iIrO+hhxqnCyYdJK4qpR/AmT2RvvWiyPKfgpmJ1pACqh9yYkrVYUkr
Ph+Bz/l/3ZsWpgPsOY2m9tRhmNQjlx39Qd0eEsVs5GbGMG0uNMGFKU/tAbtblx17XUEQvdV3GpLJ
xE+n8yZ00gG/03cy2QqGmPJG3qZpf4FPrbH0A2itrDioUKlaeYCFJP8zkQek5h39RAwonjpsdB+k
tcvfLIM+1oqS8FkdwuTBBnD+roypVoHSQ4BSzz2cvWE0/bd6lFeIjEEuft+5pYjKcMOXfNa+IgDR
FDaPyZnlwVumNG6F6vp0RORSc38ild+5/57KSuoEd/qgpHiqo5P4trs0Ug57xKEYGGWCGBcJucJ4
+LPyqGkt75pDfl3DwXDf6Z3zF7VtEbmdVeMgM69DVFs4fkUBwXFUQKckT5zch4qq2eerRM1DKMT4
a5QrwlxO/irV5GIUtAQQXJHGkLQ/X/0x7AaJFCzUwDB4Ihn5W3THlwMYZWhaAsHbqx3UA8s2KBbU
o0oUbdITRnxnV1tCX0I677MpSkxF+Ria3ghnjvu5YljpFWQlsL5QjFXUuD/CNlDZpeCI4Xk6Di6w
2teNyBecg07wDsJhUiyZdV/qYNdXO/xVxXh84dvqD+ErJ9LmxicGKJd7LfLH6xHE/nt229upae2M
v/VpSzswRb16yQnpn3MokFY6RzsXj8edDEQApkfc7Dbzcjig+uBFOVG8OclKvRUAtx97Y7Ob6f7l
dDja7IXT/tV1TkPSIL7kHEWmHd71CvLSBnw9/Vm8/7RkufRmUV0PIkNkU5td7+rLIxFP1x8qe8kb
N/vpWB3/Yn3C+lmN616l7h3oXh10DcROQRfL+bDeCpec7lsFVRP2+ar1ISxRNDM1mHASSBkmY1fN
vh0xX2m575Lep6loqrPJ8tpA8qQBcAPke6HiCye94PhBHamjrG12PJ0PMewR4c3eCiRKDcY4OIsp
I0gHoe/sKt34JdklElRBJCqwFgQKXSwrFyC7tUDa31z2326C46osityCK+V4OK1VNqH52Wj1Oi9L
mPdOw6p6gvSskqRMXhq7xnGyLiiNVC5qoqvxoNil3FnEDKSL8f9mVFPZ8KQlBjpTyMhCDm4j4yKT
GP02Iwn59+mjchMGVhEpjzsEEPaZCjW09Gi4JyXMDZD4U0ZJp4qYtGQqC0ohVWQNk53tHfsE6l2i
fbNIFoqh+nZWpdlayV67zKBXKeJSsYnUoy4l+YZwHLOrpWe8lqr4g2196LX+iezN5hL3M3/N2ELc
V8OvUlD/MdilS2xOXH2laA/fx78YoCUrGxiEQI03sbf+K3pg/VMRn+yg/XYYoRRSP+8w9EeKLkhT
0puenRgzjA/gdAqXWenZXWlEDXs9zbD2T7DYB34rcs+5BsSbDgRnhNysKQ7Lo0rdP1YeipiPBABJ
SOKWC/GE8ZtecvSfVkYnFe9sNpJwKNlcNaLqwszFbe+7ZpAuGf0YHOvn3Iz15bYaLohDW6DCW5rS
OTHhlc72EB9TCaJ3mckW4GHCmmSAmTG4QPaU164XcfmL76Os8VEs35CoL1jVXmyC92XpEuB8Rirn
SsIrURYSZc79xmLYSjqADekh4DgMOaJevnya6TWAjVk5sW8Eck88xefnMT/ke1VlONs/c7/bDHWu
gDwQJF77H/58lL8+vdysmawTkNUjiU1DnnaOuL11V4G+BPreXaD/V7+eqP02+DlZ3xHEJOhdAJs2
7Z7h9rNSzW/HwX/ZlBiY/F5nm58oUT2LhiW84O3Yu5tBp/GPregyDvOwwb7CxPH2HB0IqPHJJ1TV
tV/cbwQXivmpmB7/Qla5XDhC1G6f66+n8ZQk+Z+Gl79My56HTbhl9qK6rsXvnYdN61aTKPwJ06S1
t6AqHqd1AuO9ZdnA+Ti57JMJtq0EDpvfL0ppvzlDBYYiwV4DI2xbnBsw3VV3svbCoPtrVlj6Neq1
LoB1Q2V1KKfy2J62kHQrQFxV15iZBoxH9FBuwUdq6vZpZB//Nq25iSqtnfgscVfpiodFuU6i0VIP
qg8pVioeSIpfcDAm1K2QzGu+TXjOJJEid8oJZHiFs4fuogC15WMWkwvWDLKkrR941ukXq1n5lMby
IcsWb979f7H9h0LZaJG1iD81JNaYyEe7WY3n2LKY8A3RwScXkfF807PiAeY5I/S3ngXTo4XBEbbJ
z0QohEpQOvDFA8P1ejOXGtpDchz/7OdZKbfo0TA4KBn71AJ/qzT8qwNWgeOfNC5qDksiw+3IV0wt
KTfhMQfJuBexFvFpYXl9LBa2v3yckEbQA9EIhdfLI4P+g7P1Sm947iDl6Pm9DWZPxlmWMe3SRLUf
54R6VcEiRP/5dsbWJR+/2hwmxwmSKzgck+NWtGo8RymqO9G7X7wgwQI6FCr29gsRMRbAvrEKCC7y
RYOM9Bs6XhY4liaH/2Z4ELBH0I/Sqi4SSbUia5ZdyeN+4BXQ91i8w7HNv12Oa99ZryvdVXfXxA3D
Q6+citacIsvyrcdASXY5pTE2nm1WLeAn3y8N5RbaviFb2CqjFJbOvqGIa44WDRIOvaZ6KJ331K5L
VHt8tsgpY7ATyAseJBJgmK5jSAVMQw4BIL9SHnfUSKHO0A71sLkCzVLSoE5sMfeN4CzEqwvG4X/J
JbM7pxJYWapHNGehRWpy3h7CTfgmwTJt5Ilm5FlG7PHIXYb2iGjm+HG3dT3wc/9vJSomX/tAWqlT
EcuPUCaMsZv+aiCAmOOFL87RBmXhamyliv/xDdWlxbIuWQtTV7AENmTNAsI97suYSpL26r76mL71
3qMzs7V6PKeZl2QbYJsBJeSYSIrK1sq6izWEuonyL0tybiJkRnkuluz8yifqdayNdbWAP4Rgjb2F
x1/dsmQN6pDAvLRLHETXbXg0iOf2cDLcpmZK2YPTTphiYHVnjFcoTU8Ll6yTAHzpMTGcTd/zHQzh
xkuDXoHcbaDQViAuVBkcgGWjxqky70sfth1aknP+7Yx3K7lE3GFb0NmsmQ5AehIsKlzorF5KEuh6
lY2Wvo0mmxSNNfnDEmHbrD2kfTDxZakvaz+84+pdfJI7Y2hTvGWc0bHhpJpGNlLaPB5mU1rbYHrl
n6YAwQqgl0fnViXUTPu7+YPFODWYdUURjJoaPfRCUkq4C7kP+TqYK3ofnZhOG+Kn+P7JV7RCp3H8
TgnKGT98YGLnL0hiEjdUrl31AdlnkAYGMZwfMlhiE/TPI25VznUyxnGCJaYpZaUSE33PH+A8Ibqd
rGz8EYgx2L7VOe7wCcEQ5EOVHSU6V0wG4fIjH2N6n7cguLKpcxQLCTm1yQOY2FdppnFNSTcR1a1I
rOptRLrHNR16TWGJvCtN9xmv28UegekrKwkwldgJ+MNcwT5pJOg5xG7EznkSpqxc2PrI8gwYegJI
0i5BoFYHWsGT8upSex1HvYkvcCYIhu9ghvOwe1rwDRHKb6cWGjnmsbxO/BOZvGJHOLhJhARUxq/M
b5DmtIDk3yYpQjEvyLF8BZ36O7W3ObFTAQ/aW/95Xl6JTMtOZsmVtFHlM01z2nhx21rt4wlUgXdO
t52tG2/w8s0PXILFlo5PeQfJqEPSXM6IKZ4qg2wadZ80qZJyPccCNRDKO6sEJTpEH1gtJI/msYYN
T9UsvAm80/X2+XH10fElCBPaOQc8W6nCfsXHcKhWNclZGWrwUxOxLMnX37+nxit3KvtoIR2nQGD/
NxnoP95cwaEMjIXktgOSBgCX+Y1HvDqO7t1eilMbEGi3MskYSdYAmxHzIxWbF9iRe9bDSpBIAnJL
S5kRorSoyoSNUv7MgoRc8ybVJv2qJO1boYMKQBaReTclzKAE7+YuCjEQgRZz7kZsWiEK1rAFPtDf
lpQkE3XbL749JklUu1P2A2lM5jerUXq8UVmgV3kxb1TE3GsGUe+yIWB2PQez7ErfpSYgB4HvC1aH
AQDi8CIKF+2Nu3vaZXFmwikD9UvSXH/cDWKr+RDVg47VUvA2cuP5CN68EPYaRbtxBEA2FK0AVRYm
QEfyQhyRH0KIPC9HGga+Ie6l+9d/bqkLUbA9SkiwW9jqBgCTDoKMACQj4pPcZahJ1ZrqVvFHDP14
aIuMxeBPSLr7E2l5HzC+Uj/XsBJAXDwTjC5EdEXowQA1fKns6lqBH2YBNdkb//sMOsJWdW1Yy88A
U1NGwM+za6+mzY1XljWCcGZOw5M8kZbUC3QmbTXAuRD1E3jBYc2SqemXZb16Ndc73hUNiHFWt9NK
IZAL84bQ2hR8a0KRhTt2q8zcWNNEoLXNXlzsV8x41WDsspWYq/AFyiJ7ElTCeCBLzb8XyvgzsFSG
4z7PuOb8hAODEshTq1ba0JIxwVbRgdmvTvnWPZmUJoT4XJB9UNGobhuijvy7c10UIypTN7pEQa13
NpkTkOd0GntjJLi+C829bCpQpMyaeOejE0PUhDfA8GVGZ1lTahbdV7mfXKplmvufBEj2BKrnRKHH
kpeWHIkKJqi1ZotUrsGFT/F3Kdd1AbFsp+ylYSu3cTccZvc26JdPj1td2oByBQFn+h+ILE5eAOM7
h4GxanwhEXmxOVrSSKTqj9L1FWUPB77XxdmQjI3UO7RS1Z97fU2opQ+YAsXpSnhlyiTS63UIR8SI
w/eJJdR3TkxygTbqB4gBFa3QTz6DT0iD73kOrfdGqfQ0KflMprnGiUFmb1aPBMz9N0HHN5O6UD8E
J6jSYUkD/GUKBe0+Ut33nepgI5l0w1BrXprKNHUSI/M/s48vOHplsThuXFD/fNOS4quaJeH2J7dr
xqDn9l2lxm8I01zGTGKKU7qU0uJKQoT0sS2KnrIFQAWnStHMDENQHmUOy7XG4ydcSs0oGS8bWnyd
U5JkZXxq5wRIIMCFiguc6nP7JDmi+bic1hL6iirXtDoXrkLM7PT5EL89lr5i5GVwtlXYwgnaYzYe
gCpWBh7xylvk9BxXnXoCfsAkrptrW4wAF/JdyEiqZ/x4OLnN2aqIl+EoHOYw5MgVsriYSYqZ6jt8
jC0RRxd7NknBTBDaxNouD53HWh5GQtbXTFeF0bwDR53SNmamNd89W//LXNyH2RXaaKVfpXroUwnb
YJbka1AemKAe8TggMJEHFkMOtnAv8Al543nJsUMeD7nZZLtwwKIiu65lYQLkiBwrDIUg4yYS7wiG
jrbe/1EVn5SCRyBk4XAUfrUSkx9NFsxvADxFKOOi1ReAxbJMU8muz/24Oh8CVEbLTDQxzcy/KfMF
HJ2RFZe4SEfoKt4h6LNMZdJSk4PwEeZ4q6SY2Gtu3d6WgEDe2iMh+iM80uBDxw6w7/PwdG4XVuG8
SjKkaE6rjQZQb6I4gC3mNd1jgswkJGwagMReFkIGzV58sYnPJpLEjy0htnViP9vawUxAtFYlu/jx
/I+wtE80PqTXsuaDqb076xXSXV4PdRYOrmFm2Fzqk0Ofy7/MNm3M7JN9mz2Ntd9LxAFQPEZVxzW3
GMqQaiN08N7Q5C1weuKz2w9vbFidPDJM5KYQr4eiPYDpRU+Xxv3jrUq3laJaFNv7b55r3amecBR5
2mY9NJqb+llTT4/IPK6uFWQJYbJs436rsVQlebiyu1qpUJbVPE5kpaGHPD0YhZg7b7tUpJwj0U4J
gjJ67+otvdtnGu0S9/0XoeHZnqnRDXSYCnE3BbRil0wveifQ2KNhviSeAOlDX79Eucn22sfnFmFg
a3XG2S1m9kbwtB3mEdhSWDszvoOU6t2T5IxIEmVDm3GN7kOR1JhT9p98LqmFSGL3WjNHjewI/FtG
snhE8h3fdhMSVIDMaYAUGMr1zGI3WqbrA2TEOU3RBKx6GjgDVmVl/9dOiXN/kcGdpCpoF/GWl3E/
m9MyPpojrGPWvys4WE86EQLaJyN3gI/yE0D1KYuUmIUW2zmPc1DjwL1fuWxdrHJe5ZYYisTCgEVZ
if8GB5eYd/ywft1fmQuvKnRSXyLFcetqA3BY/OenQacHQmOis0X/6brQxIC0tqoXc64EPkX5NHLX
2XgwmlJ7hoEnIb0KLmq+SOY8naUDsRRzIL6J7PSOMEmJ3w+KBrGTKYxqi0ZTZnaUmOKDfJh6vOXh
Gqb5AehyG2qqOp1S45SkaGWShx1BTMJy68e3q+g4xrHbno5QsESSpP5YlRI7x+dLuem5trnSGIXU
+hdNweLkVowBpHbXpsON+BTsF51zQsQaWszhij86ps5jMh3My6KwFSfDr83XuLpNuaPx78wSD+m4
VZ1bUc5RcC/bxOIOh6pmKiz5U5KO3Wq3g5MsM4nJgqUq7SZ3oG49YjRVLPC9PNXV93uDq/SHnPaM
fdFD5E1Nncqr4Kh71ZrXufyQGIwoEQBjHX4GV18nLKencsXo7gBA0YCvfVJ8h5jSgehFZdp0sJuv
qEy/hWDoPh9135cj2Hq7NFJYKPwQp+FGPljo71ekczjliFEWGLPLUFxwMHY8CntWNCM+xUik4TMQ
qR/8lKT3IpgnqScv55n4XQPK1lTMf+N/+dqsRFSzBz5MhtRMCaeQ4RnBGGkfAAaxC9sUldKQont1
uYJFGgW+RUOFncdvI2cdZvv8kFdcBPQh7HH2ZnRD0mhxqLKUtr2F8v64R/1uH3anUhBYtbyln/eZ
d27Cz05SE2qipjpQIW+5FJC8TOxWszKxIDEWAKGhsFDMYJ5ezwVlmxIMgGUYF5qa8za7qMw5Na5A
rEG1MBESiuW1sqjHrNsgbtNIVqkTgO8z8HpVine6wLQcliUpsqYVTJXzbZ9Oly46FEmzE8J8tff6
AxQ4nkhtlOGJnZWKH7RPj67GfpgdzZ1DfZFYExPNv3QUNPQa3GyyouqHlt0FAolE46tsISfSdXzS
9odDXhpqN4JfRNZiE7sbaCHQsrG14K/ImfHg0I9XxdyuBCliQ0SyRf1Jpyk3qRdPtK/+X5hZFTUX
yL2RiqfY/+ZQBtDujE7lybMnlyKWcC/VU29ZBqkogTtIhtrZFuS6Z2HSxQ89WSdMDxMXyUAWj7ed
Byl1XfobG89Mj9AibHbdBU/bozWcbBKgZCkRpKxK3pOQiIgNcE8qLKwXRdnZR9g6/y/jX9wk36kd
oN5CjjUPz82nb+odF6QL0Tmg+/ZAAF6VvI6zcl1Zihdau2HVOhWsD9SFFoX7oN/Li+EDg/YkTEVi
ZjlnkWwkHV9GWkgkjkFWDs8UkvqtCt0OKPfrjWxVsYYKqztugHOO33QX52dPM8Vep1V+m/A0JvQc
st/frRkc8FPTlL+s0+vaMDAGKQ12Jfu7JiXhwwqF8ovOxwXyaPIC/Uf3QsgRP3fVsTcqQvL1XxcN
esFySxnROpgYQ72cBGklj1m1wFpRwkohS1UYDH+sQwlDAe4dko6KiKxwaUc/O3ouenjcVgpvAPBe
jD5hjVfKY4zdYGqO77etW1X8CCxslh1G3+WvdOSbZQL+oN7kavFdY9NYKWjEIETB4jJb7/iqoIMB
xvGJUPnpoX+nZm9E33qgSIER/JNFP3jgBBL1Z+/1wuaB7CiC6P57EZYglROUHxwxjQ3x58S/lE1P
UFPOEn+a96gG03ClBHQ6jUnJtegbqOCfix5fowh21nSVjjjh7RBHUfWhp89E+UoFp2KYdlI6jv8F
paecwBOEsUznTxrlbEOMm2TPxpY8wl8teIhDKNaKxmevnI32glRY8OjlYWr3rcyc0P5f2byftTL6
UpGQrPUCYbb29JCKkkj55pi24D8cTicqL9miEqRGZNTL9N4RveAkyq2fLebdJlEEeCGWUceQu4lI
Ya2Rnc8/T2zbjTGhLci0TjyvhRfpca/m+sDI4nGDVIRGDEvLBsg8iTdSOXXShVgYs5Oaenke57I/
CkfiQGwSX3EdcxnlKG6YzLTvYK9ZzO0OmbtPnLakVwcNa9zPZxpYzO+xyBP0ivafu+yw8TSeR+g1
3GGctDddfy+h+tUnuKvUYwvwunemYvdtfnty1V2O+F5z1GmKKW/sgMAzOOOT2nkZtD/pq55v1DkL
1q3RWFxxXaGzB6Lz1oYEAd8liIuesrYgs9w7PfbCFkCR2cg3QIbCPyCrvzF/7TK70KPns1vt/voz
Du3iTtTHSJQ08fhFr9yDUcHHbcARyA7HWtfjgEsXoRZbG6b7rIIj+6kP+ElTffBoiZRQYJKz7Mlb
Y7+LAoRXgvn3Wt7OzNmIK7b7xnwXhO2OdE7ZcCm7iARuwTzg7Wm6uBStlANZfrlAatxHpP+jcqGg
BWYa69FYA+h6fFuCX+aqKkVUbyay8t0DpoU5thhNBEUOJoJgb+YhRLxZHH5LKnTcygoBM2+exxQf
3SXPz7fdQwRxj88NWEwBMJtoDy4EhM6vxwKuiWcBPlOYozykgx3rBN5VuJbpL2AJHc4KPSRPJc0U
kR+g74yxSQz3acZlYPsoabL9+ftKjsnV4ygOnr+zdPGTQgooKej7GE78Z8q5Qnu+G84pJ+RAHzgt
NXMOEzzS4kMP+cQtE204wZE7Ctn0rS55sqaAjs1ZquikeASYiorNGvwQqDSGRIPUcDtaDdd8hX4X
9KnzSXu8hI1PMVJz4rR8hpfSEkjC7JK27PxL9YlsOoQBGVOTlQkMNb1vXbSNua/FCIFPgCPy+PcO
lYpcGBmY8LxQXr03S7hhFI4oh347cmDjmxvacKHNK98twtOyXyRNS//S8q4SyVthtkldCRTgoq96
HF12CiHdYM6/avvfStzxoHXdvGtVjat9R9B8vp7DF2PAT5fG37qYZad80PxnVLq20kBFEAHhHtKc
NhIk8ZUstUj1TFZPhqu9QV5H5Yq0D7sxQ7z9W377Y2tvA/uIkedaRnJP/00YNtpM86wIV/yOcr+s
GpBYIeGiX9xmKDNDgROITm+HMVzX9I0R6hIBrhHNb4TgXnTQEmge4m+34W7okMyv1j7WFPxcFLMe
zZxJyR6hGOP35Xsd9NtngYqquRsGXfS00GdG9y3YFR0/oBlSIsT9TzVRWXMLDdh8OtUkdUcEbURJ
cgnJ0pe9xBqmKzFj2/tPG9R0WW0FzHKzL2Rtjhe99WLZvxsV3F7PW30uPBd8mF/VC3D4ieVqdIm5
NByU+qN+FPmLyI7TtItpBPsQVLQIdGuzq7TSYWUF/8oLX+HZPfSYF+CpLtpP9RKZ8esNDNwzqXvA
o3K7TIdzqxEHMBuKprktX6iTqNGCD+BQE+TPJpIdFlyMQsAVEJta8G/HyysYJ6/BQEYogjOVLyxN
KUpJ6zqU0Ko6so1nWdhFPDKFKZipl6wWEyDTDUaDtxQQJSNFnQjBZTLFzS/vxfVXC2ZCD8T7dr7A
s48lhrdHP0NtEm51LDV3rRXkLSntU+DBkL4Kcr9kYxYO4D72TkNVK48dfc8nPChE0Bkr0I7EBtYx
py3h3Ll3BNKHj4vSnsH4YOWPb5TyZibBXYncWFLVocPiEelSqHErzXM0sz6aHZNHaB/BDfP81QS/
I4v4qqj+0qku/r3vI7YNHXwSuPFC7xpx4gDznODM99uCNn7DWaqp7Ylf6//Te6Hw1ftN2jUjmQ1c
LDJ9cr5MHo8pUkzV4owz4lKjhBkp0/xXqq7pkeC9wbqxTgSWfpS9k79XjI0Db40Yc5qMQKj0/QHm
rdfYxfbw44u/FIVEqhJG0LVSPxvKkH3+aPeY6hR4f4MLq7e80YMwdpsLZ0eyP82n1lpeoK3H4I6I
Ybs6CAmRI8YNkKUXqcMwKjBl7c6lqZJntrf9Pkmx3+UormkgUe8xSL6SFso7UGp+cO9bKLcCmdyn
KdlzqADxBZzWnvkXtDx64wyAqoD5DauMt/5zg6cWm/OHWcbG0ziKacL4gvXeVuwuE7OKwcJ2NOvk
mRgcQfDzUfFq5AQ3CWNlATqXga96w7PoH9d/hRDEqZOZb/Tp/dsYYP5ZQETANJ/P/3ITAVQhnrQq
1AjxBI5v8dFDLgDLMp6BQmKZlV44uLNteUtLIYpwujDlI/fcU3+dUq5DdnxSMebYncmvQlKuVveA
bdEm/EJhP6t2HsQ+mkRs+iQitzId1lve+cp1wkEmkFHZtQQEbzcaH6HYJMQA1hRMxyvz9hN+uNyX
Br/UVm+it4lj9PX3/YNz3SJPD/a96en71X406z2DzRFjj9UeQHKcJUfJncjibOeUjYj8a3BMo33I
V3GwyfA0/3g7Ld9C8E5FDQmTuUQECBeRGKzUwxq3L2CBUOGQM+3HaRLWUKLeZePDkmcjMvVf1AB0
QF+W3jkMF3eIoRMsLduBopTmzzLrShbCZ94MC9G3mQPH+saz/9dtcDU6LJ+ncE2nHHrQu749JULL
7f9OwxCUCgMwqJ7z3Onx+Hjh7YjZnDyBtRQEDnEmjl8rMMmRiKzJ/lCQ5pAPQeIVdTg45vxcId1a
Xr401OD7BO/80URlOr+1nnUlzh59Y3XtPXeLiuZ44qinogA/YzUBKM+fSjHThPETVhLNg8qEKLjY
bnjhRrrSQCDpVwdGM+Yntl0ptc8tZ/Tz8k3CVQJFAKE0UXmA464pryIk5RYkS+y0YvneOgDc8ecr
mpQUJaXn+T/kE1/PZB0tmzGnjTz1Px7a5yxSnxGVWuaokNY+QQsrDkI5uKhXiDJom39p6KVRqmdM
/OvUGBxI+/pNdQWlUvnQGmMWzyfhUfCAboCL78iyz16IVCP1O/gk4DIlLwbDzDJhvXkFkJ66n/AF
cNdE3dfOtXINu2GXvuXaJEb/D5XHLEDSOftxQzKERJ3giJXi8j4lbC6N6QZjbToZvfQe3sb2rBsM
Dlnl+kcaDkHOe9PrtBReKQwfEKO8mdKq6vJansShH4P+jJVQKIRXABx++7gd43zWoGSbi467zcYL
y19MxsEvtJIDhz4yvKsMGChrR/sVOcBOW0fYOfSPCTJNKaT+d4/Yw55YR0YUBKLYX6WDjDJIRdDr
c51IXsY7HIH0dXNCS7wC/sove9n/dJvd933GD5rXYDr5fu6CXCbZqPg5piApMPK0/nCFsRk14YX9
trhuViZ17AXT+kMyJgjcVf/Xciej4mdNPzjU8F+T6b6wM6NUeQHyXdu0Sp6E1rj7d+DXNEkZjxpD
4O3S5oDkk23wEAxREBMCyBl2OjbI3hAkIbuQtlVC+DFyT6UutnL/0nrNQNf25IBf3z9gn0cibHVh
ljrk/z1qRW4azANuerC6rGOXEaxmhm3EUeTvWfPzUklyvnvt/gzHQy4UTEu74/QmtsBzmU0gsKUr
CeHoO3DSl/nTCPeyscNUzrnh7YGTkCHvJxBiR78dAB/2uSZrgtOEujTEnxC0M3tYnkq4jmZDNXQc
vfC36DDrqFeCjQh2oG6NA2i4+r2Gl/jNkdUIsik2jiFUE2dIN++eCpOjHKHOndZ3scaGSiF/YOPu
7RygWVAnm160k4CShFgGZWpF5Lqeblmnz31lXixtgR5bSbSo02/CAU7Smk0yKJ4exj1qNtjjcgcZ
8x+O2aqc2Ozp5+GujCmrqB2SzastSYHjzFajyR33oM6GuyvY8+18VjzknaXHWeSMlic/IwyZgtuK
jankAGwSvAifU55lT6ckHVYv0Hd0BfnakHMTqSCEqHs+4CxsPz1vZ/NVYr4A5+yf4VrzgT13yXb5
G2vQ2kvV9YvrbQwHrbFo8+8mdbqDo96O4UmWpORAy5PM2EeX0hViZD2SIAZ3T7HP2F+2A7XjHFmU
P6uOoAXsPb8bcHzPWWJ0BEuTNvjBbqb3iOIyXM/Ssy5OGYSwspJTPkMXDkB9elnw/Zglqdhr4WJM
ofszE0MtMADYmyy+9Qh859SSJTG4HhBgdxErV3YBFJuYeI6o8VYzVXQ4W0uYWPeiPo8NSjW5pK+C
1qltWiL+6eoOw/p+i+N2Hv1CoinVVDK06uRQuWdCBEK9mSkH+g4+g3sMvfvWG3A5oho3OECDZ1Fo
Ox2UDFfhcNQY56MfxPh04J/fMS7u0Qstl/nPbYhM7cdi6Twky2BHgfWFOzscnkOXAj8SGk2o3w+z
LfGK/ypOm69R20o7imSYtbqk9Nw8jywpzxET59Y+CntPUFOBU6qjM00gKebJXf49cF2S/Nm2efC6
mdQzGkEZZ7ofoVC/TJ/UHNy6gZz017fBFNhcothA6qrXJ/B6lxFj8eMUegFFTp5onPwmznVxu0Zq
PRC2uGDGWC15zuHB7AJ/XkSUcFiJXvBPBqW/7Gv2xf3PIZGOchhQZ9HIORshkARXR2hXBRvCAGz4
Vorjgchfu0pgYk1oDRfRsKQblTjwgfQjHP553HY4PXveaUz1vXeYwCXMYSRGhfkWisxxW0pdZZpm
PrHghkGSqU/LtnAgNDwnZWJBGC6C+U5vpJ7Bkqg98c78qYi4VYdUXCAtERSQaiXcYPgqQYicM8qh
49JWRNUfQx71fbbUlqWrcYPi/U0QPpA8GYiyAdJWlth61+RMPW07yfT52QjwKRJ+HMAL47HI/DM8
sjRGusfkDK3v6Cdn1qirmdHxlubxW+XJLdsRMBYg4n4i0g8COL190TlEXF3UpOV6uH3+QSoJZWDg
k/nM74ONmJ1pd+wyHtSzxwgUWfwN+zP5V1fcJ6KUcDlwOFogOxQzFUDoHi8KHymNSKm08Z3uuC8X
B3TU3gpD9Lbl46LJjtc9NH20Nozg7aiOYpSjXZtScQM4bqkqz+JaIL+xpMzNcDh2fRNQb7gRgqVm
64ZHMJYYcVeHTi2p31cbizgXLSCKIJ4uJqg9i3N06oTT9FjWXAH5Oo0due0vlUWV9aMPLR/aYdsY
dSW3Ta38ow1Ypsx0tLoPveGtC4hb8Q4n9PsbF/HRBhHGvhWb2q68q/u6aK5tzLOmXy0MBSAr9nOb
69tIVMYHSil0cCCZ8M+4TS1OGyb1Qq+Jln0EYolzIxsoi9T4iwZUfoH44TntChP+j9hIIErODPaj
XQKz8+UefT/1OfasngwNX5VMhz5GagJOjC1RnLqbJOxkD3FV3GMKPAmZmkp22kmyBrT4Yl44gMnx
sD6TrP01UpeiovTD/106nzRSKL/V3ohxP1x9cnUUu60mUrdbaL+ovu/9nq6l9nOjuzGMQx+yuZtX
J2YmmTEQIGNAjx4OBuHO45uF/oTSUxRmINM22dDQpNZ1wpGbNpz1iqEP4gn6CvjYYmAyJg3cJIjq
eNpbPeEBtknINPBEgfPWL8mq9fimRbrryy4Y2QKiPMtQPwtj5gbrPKpF7GVFvrGLaAAchmI/vnPA
kjUbqFT/XQi2Y+xXlD+M1Xt9PI6tVA5o3v+oPO8M90KPdC9gSgtZ676p15NLwnIJZMJQtfnxC8Bd
Dbnggx1fcOv9GVLShAOxvElYHt+nkY0lBw966L39aFQ0qdxa9BxM3rYPteBym7Moij6cximdIsdJ
qE2OjReuKWfxLbTe+lX9om4RGyeqvaFZsVLG7CNibytyA4A86D0OEXdirrJ+Snk3fMesP34Lt3rJ
u3qZQy6O39NIAjMctJoTcTtFQNezX3UjL5O7dPiX8e1XRmC/oYYCN7ZtXiGuXbOhomARHhPT0WGO
lRjvOUgUqD88DkR0sqAelJxj+7WfHA+NPyTMaEzlcdBfSgAMlA0+8H6OLRJFt6znEJA+BufeBxWV
QaeMxPzFiTTRXPdbX1D9tzOYP8tCoa3Iepu7XT06OI36HpOeA2s6A5mJ8SD4jdvq+KBAGrHtt7Il
c5zsfh91GKNrgQYU7zb4iLJCsPXwvPcCpHvHn57bJwB6/JodpupegNzLnY7vBDeBpq3bVQsF+3HX
MFk/x1fRTp8caB8z8vQt0+AIoYY4+UkBk/Amq/rz3atK5rBL6D1l9i87PcDAySAf7hECrE6MXOld
Tn7pKYITj4zN9/SRR6o6MTXZiwVdlk7HLFDxBkVicBQYXhjSinursbSRMMF0emicK3r4nU+A71e2
aSb9um/KXKzxf9f01+b0SBhzry3A8DVhwOoSENqOZQ3ZduZKjDi6OJVr1iOMh0AbUMy5EvzdXmdA
rKmr8hCCGncJb0agmLWXfMwiR3autwCxcjAdl/Qn4RErxggq23D21W3nAetziJHE7Ox7yGS+BVei
3RduEKFGk7JCTNCE9QOCZwRVpwTRyPx6WZ2vb7CGr38jxylTeWqmiSfuN34NX6OR45EO7H/D6a1T
ybMc96HhKsSjJJIEUVnEZUV3BbyHN/z17djVI2kZgku1onlaGAs+KccRHMmvd8NcAMguVa7OakRN
AunyfuohcReEkk1yNtCLC4voIr+JnL9xJEhg242pHPCQMvmNlpPz/hYHhrUcMNo0Ug43jleUzhQK
ofjvovEGBJDitadD18ameoJr1LJeHky0NEGKRl1YbaTyvl/ZCmKz/u1F8utlNKW7N0UlS9SmgwCn
I3Q9s3aWEcHtLX0/F3oMlbAJbGHj0aBnUi727R0guvqTQ4M8siLOd9RwQRR6EauS9SWepu2DmcDY
/8G0K3m6+fzHujl9M2b0ZphMH7FW+axRSGljRGoyW0nHTv/4/0uiUmCPIskj4VecnBegKXpQXd+g
0S2oPsXny0ntjxYr9qdfwUlOggwUg0zdDevv5vmNDSedj42Q/3mIDrU8yUVswRQyAgllvHYyUH6P
nqBzdCJRmpbOlQyR99QHxrGZEDrYliIhuIBbzgMBIfWKFjzXA5A7ou4Jz3G/lThWjSiBAsVzDEtS
8hA4kT2JjtlCvGxogTRgXrz7XyYzvoUtJkxyDJxEaxPC+UI5m8+3P+9VAh7UMiFUPvN/Cjz1r6X1
0E2NtQo7wJCeW4xiMT8AoXoxvjKLDXCPM/YUypFTu5nk65ZBukZHo2ewAIseKEoNZ8hpb5qplYZm
9PSDLn8siek9+Y8fNRZwKlZsUrlU6yFchtBqyN8OVKdSD48+PrZdx8lGr0XxvwVva8vqILZsFezR
G48rWQokWMYe5Nx+12Hiy5tKb1Yfi4VVLwYsA+IXHQgm7IEoBEaVLReKl2ai0r+OSXiknR74/6Iq
gCl0QLhVJRPABNZlHne669OLqya3sFyvbwlQhXP6vR3gwkwc1m9hiq8oEaqlgW/HROFWmSE6dzQe
+Ux1wvUbhaT03PBOOFdgc/0uMcsVNdWoCox5rE+9IBSeiHNNAp2e5M62zgumod5W273UVkqmfoH3
o/niWGsXcaTcz+5Dq8eMHTPOhJzlHeqZ1xjif3c5IoraHT6uZB6rX4LWxxuOI3xR1/HioWl7fdIB
NBbtd9DPGOJbkVvbOOSJy3dh4RMUkcx71E+VylwlWu7XG3pg+BjCQBdigXZ2Kdu30dEPON3fzxX+
qEMBdMIddLGrqYwu0azBDlvIY1a4trMJhYurzN5gg1xQW37PzW8PgucQJoV6JeYHiWJLbiEP6U2s
pc3A6N0oiNJ1E+uLfVTjVu1OKa0xx4Kzei+9wVhI4UZ6gAeCvsD8rBh5D1SDbE90bRIUa5VXuSTR
BpCTbkskuzFpU79yKftKY9bV9XSm3anXlxiivJMiRRCU+tD8IdVIukAPQam7NGnuQEvnP0/iMck9
DYOzkJjVsgweSZfvAwwMtabAQah6uGstXMPZha6jCeEodBaQyO8OMFB4M1EhvR7Wao1Nu6JKRyW5
LT65oZxTZISg0ODSRXyo8nBwV3hghv1ar0wzl/cEKuLmR481zG5PgTwntKm6cEHjuoXWupbWNUaX
4zAUIbiL8mksEpen71qSmVpeszloocex/gTOFtu3Evd4fIUdXMQdxUWEKoCAfcAp+q8LDBT4xurh
AEUZ4qwH7apOPTi+zYd8HauPzcpnsSZ6drpxA3BjKL96XYpMi1NMEOCkQAPOnLN5E/2CuRFhZvc2
esk80X3wI1HAw4ASoZxe5od8t5+dOp/fgpofXU/aUkIepMNsNg+tl4362eIojLmOhSc9iYXc53pC
SR+Vku+bjmqm1MO9cZHV+wDIpcsJ45fSBFJKU+0Gz2JqyhHo5PGuZcXp0QGUIRU+Mo3vs3GzUsyv
mMnmQEypaLk0H0Ne67n6187T1GilliEC0fBZO5HWhq8mIAJCsiKv05EJB2gcfyg7rIiLwMGvvMOs
k1zSQsJs3RJQT4q7lFv+q7k4cerFIf4DAx8XknzHFQ9UkyhiZjX+lZpekyqknhpF0JNYZPBHcYjX
LySwXn48pi0FN3F0kMscGY8X4qwJ2N7TrTtVhvRej9enxQeFkaTN5gb6ArIVsIsGoA7xBlOzGSxT
4Avg27y6LYmCKNOdYL1xq4ZKGbd0FCMTPru/wa6439c1FChtVI3ZkzRHZAprayCbyYp0hQxMAByh
VUWwzkjTrhjOTMyo9IDKJP/llebQC5NS+5dc6LA33bxP1vT48eOwOOmN17/rCbUY3MRgkXZQWB+X
KNDKkKuV+gCy33uzP5V2eVUXk05/V3dphBf9tId7lYp0DFv/G3bZpvUM82Z+Vmh6iOmfbTkznGRr
R8TvbJydq8sEdZeu7vQ/O02vpOQFtZenAyzCmHPCGo2OdENhJPgKhB3tyc3Wtjp8liBfVcZgnKY6
BOMh1q+kH7bL/TLxiINT5d5Z11QtR2BM/wkkNqkDh4rxoKpYTcYB+rmAHzUr56Bj5J39HTRMUR97
7sL2COb9AHPNN9CHlhWDKOp1j75uygo3OY/+P96RBE3cUEwXHfQMo/85Fh5kIG1+vs0RkYu3YhD0
OBul1r7hPQISS1fMnT+UqcyTQS1KqR+7FkOYqgLxCfpb8PUJZQJuAH6MmcCiqpDl/sA+jT0MLwFB
FUQ7ctL9BSHnn19IH/a2michz7w7k+3Rh5AQdHNTGhcfhLlEgtSGl4xlizQSkGPwNGlnAWs4OHT6
uKLqHqmAaUSJFE6uM7D1EHmCDXTE78x4N+Ln/qNH1yvlKGEUTII/qP7yDLzLpQ7swoLo6Qz0hXfN
NtJey2/0p1JNjMeww5jxGOBoZSkT5wt7x/F58A599lHsbygJ4UyGanetQ4kJlFkwdMvMX6FrFlkx
FnrssQ0aFv8H8jPPD2ydd8rYDh7HL8ik+zrGWCtB5CrLOfUnpXBigItrObsg3rZ2XFR1PuO9gbMN
HI7GOl3EtX5lHanSI737lCMVr/vQy1ebZljoKfrVPNyJNkOpVAed8afUY9TmcjRoLhOeJ8S7UKY0
39EQeyKS9OVU8bs8Mdw8l54Vln6JatjsNn/O7YkbING+owDf7Ew4EZwLV72t0X7DBkN6GCtotYlM
IKUgmQYpNTxWGXAokAxWuEzJSGEcp29ahuSeaxjpSfyrQuRGMCCGWlkCGC548/tFuxnJLXJkqa83
9tt6uVkoRV2efmWfqJ1wViEcrozNhgO4elVSOe776qxjFNazXWVReTdNwuF3gwb1y2gVbMR+efJi
OcRgkQEEAUo6I3dG3k1f+T1eHGY8ijffxK6Z+oxAYc4o5ggf4h1M57vkkPsU3niYEbNPysBgGhkk
2icK11QEpbSyFxwDD0IIz3N+ZHOjepRGhvABaHu8fkjbFWjWVD0WpdKF9ZRV5ydYB/j5g6ssl2Tz
Lj7OEthh5qsXkCe6qMOfhhFQ48PV2oLtFjejjUIWXCuof0ZON9iY7ihWRVns/Tb7rNtuEI6wjeui
CkDWdkfahTt1ZNIs447n2taEaq9hDRbr4JAJa5Y9QmncCEi3ED/18x8EjH9uffVXazIkz1qWbDs4
z8duthD3WrBaCahz7tjTpyRSzQB6duYxXp8Y7/Y+70SkfyBrYMEPN99y7jpDuQb10GrgdjkA6WEm
p3LFRMB59d6t2uOqEQgs11C9VV2qFYOTP+RHlhO+rZUTJIkDn2A1xkebn9dvPR18vc1+lQDDHUwB
Dac4gPeggBnZgVMcXFKutIFbJL6xfR0IWnvDDWEWdVGppQw0x65CG2hZzUqBGUBiOW6+CwwQlyYT
caSQK4k3LdcKdXhIS3jQRxn65kJuhdSHJoeRrLxlJsGUk7qqbds5+UQwGkeseG6JqNy/QH9vxmkf
uphiAgq5R1toOxzp01PcSuj8SyqDky919KXBO6qXp8kZbIARdCFdDGkIL3cseQiXH09cKJGIUCTF
xEPFvN/WbM0mHL6gmFOC2gqI2qk7jjjycEzyysYPBygGzKGKgOZVvj9S8U0pEsgBgM8BT5NogP54
CraWQwUDyr2BWs+KD2ZJan1IB7ni+Qn9R0KW01Bzo1awwtqzpISYVFaSN2LbrQ/S6U/rACu3b+cu
JF+Hoj4LfoE2yMoemft++z3Y570Z+Piz7sjJsA2fxQGNZLlcNeQBVrgWF37DDGLGeGWPPES87FL7
4S1jiwU7SyFCZZyR9317ixisGQYARHxWYrzAMwQDGFjFi4YkOREuTOdvySw/S7NHYxbEaRX61LTA
whmx73NFgboOWPxafxoMa6XwaD1jhPOPp7AvVFfF8KBrpHWxGSAIWU1W7OSOFDYXepQRe63yS6Ul
G5RJZWTmwhLwJ0Gyt6xScMQ1wSSW4F51FOMd7JhsrpadAIHgqf5WQB1GTiXuuMkDbH/PVsUujFET
idmVvHWC6fvLVsrWrH4AegBXbMRsaT8MtTxW+GDtcjerCUs3BgK4iDjuduVBi1arn8AvFM11bjpY
NgNRUJ3/+Z+XfyJCUSyLdHX1M5MeiOvhgzNLU0j1r6iNXhKh3jsRPzBapC4k3PEDk68z0LSi4M3O
xIR2u+MpyvAdDTBioUaLi/tPu8EaislcddJw9/lkHoX/EHiFNB7Hiz6gt+HPHU5Sb+N0+CJ+wHPj
LWn8jRvKLmM+tELOHCKdFH3rozJZ41pCimrlS60KKfe8KkFTp82424XAEuvQ2Z6RHY/SbEKEHCnU
mimR/zXbC09LrGof+Tq3APBcXwfu40SsUGcK00IHM8NvTrd/ynBJ9J9391282oWchYgmuvc5GEu4
A+8T8gNH29s8+jDHHhKWAk3hVeGoP3vUlydDNwxjizbasAzDMIW/bSpahyoDCwjtaDGH69lNNCy6
ITld5B7wq5QF/Kzh+pxbuaFx1QH7B7/Gz7B7SoglReCPqeHhtp63EQU/45tyRCfMcjPoH+25B3B9
tLJo+dM6BWB2/XSznJDXgjQclRv9d7XgAaOA2xKum+vc4bbtqteEO7z4Y5dAMk/V/ljKW15ASKZa
n+9VHB1p3HPOoM3lg6P2MQRZtXLzJ8tidQyX5Ggn//8mYQlfp8Dr4YNeRGx+ccrxduRdjY0vPmy1
BCfHoL2Puj0og9YtrdD2SGXianUF4ICVR58/DDPSsuwxtUGzbw3jZQ92KlBj8En22cwtFLn+nkRX
uMEuuC+uM511t5ecgohOpNHJPxyOb18xooKWAoidniy4ty4XSKtoluxpZWqIH0jprx11Lrew99cy
ftBcYMGDpHfa675ucHY8lJ5cw4uZFunWy9UWvUQQFRT84msx0gfsaHHesf/8QiJGO2Kda5zSWlmR
l+9GvjmSlGbldiBVnepxV/JNqE8N2qvBUm7XVv8io7zX1mHAo2Qjl1JYTDkrlaKVFbYJ9pbka8jp
swAtYMcloecUJSpX/mN6BHBCV6UTQHraMjbBqcNVIB3cjY75CIEgaW1ZGGSpLpm//WPzwLQ/6Ym3
qKGXtH5Nasu1Ec4C3yaNFlMdmYWBtVH7xnJx+sVSsM84OcHnTrZB2OAyce/TsmIPgBu2qgePGt1Y
/D49KAxpwf+MW1fdfrMlBOtuIpMaVs9uA3F8Vx7DwIL8h65uc0NXquJqNfNgR3AIvNjTv/3Orntl
ufEXIT0vtUSS8fpOoBKSdJZIV0+ZkbArkK06VMSELKDzyAD/yhL4WqIL0/0/WXCVGybwXCgXV3OW
y/7QGcRWi1UVYvbZZ4UharzYGOlscjCbCWiXsRl/PVpa0KBm+ByHUeh84cglea5QuAyAMIx0AECr
8xHVp2fStYdtJkJ3z1kMj9Vxm9mh6mYYSImrD07mbBJb3C2tD34NwVX8andEF9tmx9Abfsm9uz9Q
8j3cmlYatqgRmhXx8FceOx19qvGoAr/ArXOtwpeEYveUfZZnmwBVtLx2t4VP3iUDa+38PoZV5/SL
kmjbgCsZekPlhhUrMGAMhahKn0g0oBU7XEepc4X9MKjckBScpKGkOhnBIy7qGyHpRzKEhBpcRBTj
iC9fTogvoOu7WbotPrE5ROZ4X6lJiiDmwQqQ5ivTj75G5SYmS2KUd/pxUy/FX4Lj5LIa98f2CrZT
hAMCYI+d9F0KeDc2gLUvZX2e5riMMeGzA/atIwMlysr2zIOdUGfs3g5bdIcwYupKPdT3F/OvegYx
LN1R5I9b2wMQSPWG8lf5UCZqZlh7jcD9OoIFSBsKMpNCGhCUrT+xdHnVfBULmzqhNigchJDTjjE1
i2FAXuUvPpzCxsORoTf0svO5dOyReE+qD+3kHKuMG7QM3VH5QsJ6vtNmCIBJq3hf5qRxalpIxr6S
gIsiOAJqmdL7/PT/47DUXoXwDVJaxpJ/TTIf/ehK0kNG2wGMyC+k6umsE+Uf2Dv4GZgNPO8Xh7Ie
oh6O7dNzYPWPf5uf2A/o/7WBmE9H6XE7p9ppapEDU2sa4Pyad5+/+Db/RtYhw+IZ816OAfJqcNLU
BNC/fOKzwDQMgRccajMlkDRsy/2bw9DhxG1U8zFNino7JHyEOUL9PUaWAZl/jGl8zsH2y63kBGs3
vV9ft3mmUzPKMl4eLXSFctnAE6oJckzJcgWrCgGpSJMYO8I0fPCK/4ys3RqTtwcczcLgE4s26Dex
rrtx+8/n9hZMG922k5jfzD/0yeLMEwao8PUOIqiE7v8YfrMw+AsKsE8Cj1Yv1qtAhe02Y1i8QPyY
Ij+EBm7660MNuDqpWmUqgOYlYvzVT+2uv1POyODdaTDcTaBSRrkB9fwMq2JrMe0ZIWSrw/TS4D2U
OkDbPucSUdOh7yaNHEII4aWMRqMAuczaldUqEa7TdLJ/hPXcg8Y4sKwso2JplZV2xcC1oAGZqk1R
QLvgcEcwebEzpUcXng3eNWs9pz/v2SU3meiPGiFgddnxvdrXFqK6S0FvWNAWGquM3Cfw036CHEa0
l9knYa8CrTtMv9v6PUncugbhX44uKdwokD299Abh4DHVeVgHCwY39M6FUDpDNvsjJu4DaJRj8AjS
wB0s5RxlizCc3O116/hZwQJUlx6IiqG73SkzS85WkkAoV5hrdR5jCJN7wpGqEdXB0Hgzgm1LbGd2
IbX/obmtKGC9pEit4BOoWa2dSP0cyYGgCg/9nlZWwsQ5xzFCVcesTD2zJW0571KIHhcsAQlShQR2
LDhGkBIqMEL+bdftLVOJgl/hfRRCJw0SdgElCarKeIq/XZK6lLs186KankQOwAlPza/tk84a6MMs
hfcKNlqdt7hVxF0q9bXdX2ZuBJ/hGFiNtfld+g+yd/nHrPPLWHiuo8GhOwiTn0ImUh1kN4d78VdI
+9qwAtvZPzakXZnT6CN49QpvOQkDxUTBrDhpH9jIfYLoeImzbqtgpDSTPglm4IlsrH6wlFrm0bDf
0ATy371a39GAAvDqioIBbWBGMfm3zel3HOPQGu+AEpYz6c9ZMlYqWfq9qbvUGnfQ/9WokokVB6qO
l+hCbpjUEmxQGGBUkgJjwfQL4qp86kTGAOhr/NlULB5f3C2SzLivzx+qQ92NqphXLY+D5mD/wYKc
J3/F4Yy0wBj2ptzpeTgeUy+NQCGe90DQUnNshWzeIX51Cx5BtjcV8A6ap6R4yZg6//vypQbOn2NM
Tz26y7cHFImc/Evf9FMw1vX6CCo4nXpB4R0ORpDvWAWzPuSLkTeOTkGT1gVg7ONfAwEFXT3Vbp/a
8gZOUkvt+VeA+TZgXjJIvP3lCUbR3TdBky/ki/XkTiKkDc6a0o5tvqE74gUg7hZm5OPTOG+/ZmrT
To6OropqLOQaF+134iq0zIM36DnDA1cLf1UFotk3wT0McOKxysSTrAzFEl+CkMTK839SUdekbRDE
LatfwWYumSW+nZXPLpbSqsMLL0qrpDayfCJT+ZqrIIxeiWuxMdaM5hpNQhbLm8fMgKUOmf5vNiOD
pnXv3AkTxsY28K2W9dnhLRl+LgkqaAV83dZl6z227gXB3NhQhHg/1L0XbS0hjIwGSsgUqObmKInP
oWs1tUvEHYotqhOrVczF+dmsfU+DAztOfzfMB9o87f8H9CiHwEKvmNkWl7eP3BQs4aMBvZbr09rX
e5YGsKAQJo4zsgtL9IOX+H9v3rmLZGuNJOntx/0dlM6++rM/ggrhDT3rnsVQewx9nXwkbOImBSUd
nWY390WowvPpAduINRvDNAhdm2iaLrQXbG2bFlEhhNUteH8AmNB62DYok4nqjyRarFVTLxQH5EYk
ugeU7sreYX/FBtTgDjrp6J1O1bi/thTiCxvdi0fCFAJhLJM3QufjmsyR8gaX7h0SMycBcbkBjhxY
lIi4FS3+72obLl2d7SCRuZ15RTVL7o/wN1ZY5rd2C2ilNRKqGSlqDXPwHeppTV8p26ZvBTMWYcjh
j7nt8kMvOX/lELzGo7aAohTtkC63pxQ/sw8m4YvYK9MYDuEw89Nt2RDbvUUHEu09Ow9HmXiAJyEO
/QHC60kflTyzzoWlr5rfdHIZHgvc6S5ykNQE0u/qAIg4D3NkA2y1yLs2X+nuoqQk8whn98bnwAnI
32Oh4jXPwnAkJwa24xiZeP9Hdr/VEhhvp0vwqwpkhrcQdMRt4KZ8U6+OvhyKHRd8pzlVDdlXr+Ce
6LE4qaP+FxwhW9bGmpC26jzq5PQlDriPHEEnBmnltqwqnuHKiyBu5zDnq3Go57UXC/s1j2h09AhY
14WAdwC+ZYgiG+rn0xPuQ6jCdIDLPWtSZuGbRNETSjnIkCUSUIIQfEr0pZWxEeFV/kTI0TDPL4uy
YSUEp9VTu1coNC5XLih+zRoTXmdMU05tuJLff5l+eYqb+wDhhmzmjyJ2V+p2oOGpfvNyq8seuyva
KMJR0bj1cyNBp23XcRFvcuhsOd2XcamgUkGckIMuxoi/r9gCMmqPywn66b5B7Dr59QPFrYNi10Zj
/WhzgeMJrt7VvrmcgjJvPfvajW/6oNLTVOUrVvsbJuPgIJSmVmLUr3pIjCvevq2anaOikCGHjh2D
xPKZSWtC9PlNJm9Mbbhb8pDe3zXSw7mCzlXQofkc5uRWpfuUi4RxnzH5jDeGSvWGk9E+ks0fx1xS
tqRRD6RAYxQuxzudUOImPnNPso6c+9WYJDp4S74XrpvBJsJ9ZlG6Ob/l0O+FjpHYnCRIXTP831Gm
zka+ezQAbGrohqGzZlTCUnWFVco/UqDWYIY9OCAKTepg25ztxDqJDHcbXP31vu5LTJcPd8Rd75yi
95+evDcz+ExjAdoKnI/gyYygG7uMsnAcuvSTf8kZNnpqVTcg7bWw6pA+PyAo6o0eAeaQP4F2xDOL
DMEuJfbdstd5JLSOyaUScc8FIW9xsyVoiRJgHVmswn9zXqjwjIsANx9YGzMZqfzAd0LvwF2jB1cB
H4FgL+S4ZhWHIb2z2kNdiBQJpboFDIYjVDJb7QKgnygKQPEHn0uPORqKDYjwGTaopZohE6/o+AJS
B/rERcn4bFctsYimKBcu/IMO8J4LCAFUCfPt4kvRAI1b6o5WztwO4ICmK9lV9XaGYC+ezvO2BJGU
XGeLvzKiF/3GzJ7f39FXAfoKi7k9AucvQlpqZWLhpAx8zJfxqV8UTFAkQWmMKZAORNgolVnsWB1Z
JmWdnjrDKPtpIOrAPaF8TceNBEey4KeEdRoiwIHmGYnT2YCUYmTHl8+hZ4RZQNxQOfdBM4hs8ZSt
tSKmw/aLCdkf8elQjMwH/t5QLgSsxWZeXBUJfhIUfcXPf/0M+zhNAMBtPXer3ajRYO4m8pgdljst
839ZqPO7T1opF41LtF7pJYNyIbbk3MNhU99FuorKQk9ioZmxpoqACHHyNeKsmFxM9GZH+hm1S6o1
NrU46wFEwmlCr+5zGfAjUWITy10KE21pS6JfWNxeQTsIGU+rEI7PFUv3P+8zBchcue2umJa5ipD1
WsSdhzyzxumSWgeI5ZDD2JhFeXhiKWcrU3M/UHffBITgEQ9jvaGzYHTHgiaUvXO7xdMIXtqgF+x6
ZsM83XelvuwhRk0vyCQny6YfpTunJJf2Zh5e4IuHLwI+zNKG3qpT9KFjVSl5KWEzFk7vT8mApmqk
7KcU2mac2WMQMBOBbL6QximSO6+U2Q//gJln3uPPaVQ9VUMmBAFnL5tOftcWiK1rnNQH3WyI2GkB
BN09DNrvuMSY9Hn50HxL6BUA1jDY0PgZlclsHK38BOG7biXu51bCOQkqD/nSD3HI12ZpgOHw8eSu
+KFPJ3s3R1LGSvvpM9OZmgWVuv11UZ9WWVkAZK3uS1QjEvALgqrCqwMRwJyBetMtRQQl8bwSt3c4
QlA+hUZ1uTFVtNfeoCwat2QIvFuvBxZRBrE1mYjsXIqFLrLxGUmuPvC8nbMqlFQcaJcrSBZkcJSM
IsVji0KF9qq2IlEmIEzrH7K+r1paGz8hQfd07xfd3dseQ5iV6rItnaG7Efn/6+Wv8JzG5LxW1eDV
nxlFG8ZoZab3/B+/mMh6pFB3m1fN0e29HIsTtyEBQnLffkPwp7tMA5PUATFFJtIIP6P2rI35nETs
qJ/S0XppTfLITW/CicUPfSjbRT+aO3DRytCvX2NjkCo4R2V/4QXs0lV4qKpsu8Tt/P23Wjwb3RBz
2Sf8DLjAKWjVI7mA9hR+zZA7QzGb4dVvjQ/uIuZcJbaXZIKKF6UJudo2jJSf8dd0q115D1dRDxv3
ZUQ1gWszqaWhKww9B/+jWSr6K1wclTVLjw1m061uvrypX7ari1+0vCaen99/4rapCN97ntrawhF+
eDc7/XX3XOc+EMYvOOyBxhmHfWEuYGOdHD5+Cfh9eMpNVYoKh6OUO96gcxKW+1ilcHMtSZQmXy8/
rsL7xzQrcCAuRfYwrUqAFsVlIJU/wRADff6uEnGnAV1I4sRpaBs1llQXxgfWp5Ra1bB/CsFgYNYr
QkSi1jll/beTq5k1cQOour/H4W+27sYVZR/B0MmPyvvto4T44YoPXdNGPys3+9Rs2r2oe262lSd+
cXEfxLVBre3OVTHpXtpCpZpy4b3acABYGoqLlTZVXBFw+HPiF1n+x/9dA0YvOm/xv/80lzrboGOv
rlrXkcV43+TPtR3fiJYikIPCdre7Gs0DxI7zdoB7pDcyLVLHM1gk/7U3pZlTwGxbI4E8tmkscXY2
rLxCA530zrxSLgNysNDjP63RdfsnnUao2iYMEuB4QHaHFvNIvcAmt76J2v2YUsyf7Twqh46i9UL/
Rh5lJQtaOJZ/RLTa383QVJkPgOH1yOYCxUQ6FFC9qfrgOCsY3Nev93fexEd5DVQ/xyu1cbkr5yWZ
Y0k7VDAIn4UXrqCSxatWLqEoKSf0oFP+Zw90yl3wxxi9x8tZtI6x2mqcsON503ThOLcSK6Gpy6rc
GT7N9DWjttmjQcDTXWGkft5+Zky0rbgHOpLzk5p8wKwfHUKXY+l9klAW63nBuXqh6YYL4wFXUrPO
FXSgjo1b/9AHn9HyOkxGzVe4mrE6pLWFlHpZYTZ5F5y83+hB5wmPlzO8vNHrVlLFdrSjp0RwVlYI
2jgakmR0AOAnkLii1tR3mqX/qUcY85BtNeoAXQBYXPQX2XthfoJdcViPRB4QOxb5JL1ka+f4xtYI
fHw5dbYMhRg4C2pL1bH3AFLeLbS86+Uv7EKEb8QMzUPzzcWvBdFrYyi0uUu0yN52GK9O1CyZ6QHy
Po5Z1X6TvhKDtTlZSW2Hpd8HjK0ojyh+/HqqW695dW84cKkvP663v0NDOiP5hd23aBOmbW2ICsY3
Xgxu76zLfZI3Lx3BnTmfODz1BjSfQIT0peP3anZcm25uoOyv/sHScF60x7PihJcZLWJBCkT9jLvS
R1gug4vI8CvTOvmsrbUaSiL/6ICxxKkf//IrE1FSI3EU+1M9At5jKBsL5OalZPuyJVz8r0Yk+Iuw
fcXcpmxFn9br2sNT4b4ZuY2VSTbFnaIKNSGvasUkg68i8LSolKgZylIHmp7xjta4sRbF+RAmzEta
dqcOSCgUbqKl3IIRqmrjmFXbDEL3CSo9HeKGEMe8i7J3KGCon7xVBkzRxxLmrtcJ8wP6Mwg7S7ye
ZWw3NKWCX+DD6mKq679ymX7CxK/2Nj0WiRYROH1iAvTkmVfeI2xq3RVb9yLR0OswkRah1k8cTylG
gPVRddcKOLXiBXZoOz6tiXctaF4kL3Rs8TXx7Dylcpt+cyaydE12XUaaleZYf+iVvEFwInWnY+UH
wrSX/jQpKaVcCuctSONDW2dALvYsqQ9MNnjg0ZuHAC7YPYzr4DsKYAUM5YQHq4QLLnsywD6Zq/9V
boYisDgMFP67lKHbU8GUiR1R4MS9VCSrq95Qzs3zmQ+JHEOF/9VFvDUW4WM2M4nrnMWRbX4+zeQ3
oXWSNiTokAucuCYd67C9wJCyev74cwkD3ioY2036QmfwcBCURJ83QTZrfXgczw7j6Mfu9sfGTVX3
DXkOsyZB33Ah8JqKkUfIcm+/nAhVhiNtxV3yy5f9qt3RmYEJcae1UQMFtvPmExEX3rKQtWUis8ip
7hnOcurO0Li0OD7iMTxgoOpRikVRZqaQSorKp/DAbQUmQ1C3ZbGrkuDqUqSQmDD1qngd6/WcD2a8
NHwVW9U2OqE8l3gL7J0XHT70wt5Yea1ZmcbHC+zTJZ1p3FgGRJM67wNEJNeawh7TUCAilpEhAP36
7Xaxyl2Gd6sj8uoSt+UwpoX7zktjmFMR1WIC46/ig66FyzspffSxi+jSif8MY44LNjiFQ5qkz8GT
fV0Sdm9eLqev4XhoaI+T/2XFQT3LQpgGGWtymM/zHr3detfYCMcBFRkgq69ZKbl/dWxpN0fC3gGe
OrFzuRPzulkwFwZ8EwcpqvrxbV3wMN+C8yikEDxP5XNE8krA0MD3jlvQzQfh/T5dDmtlBwGOZXmS
a0f/VQA98XMhozVjep6uKPsND7YCR/qJRXkR5x2fXXcfw2C0U9/2JDTOfu4SQPqOmaOkWLB1T1NQ
RhBhcgszde9WqKvJTJraLeXFd+X/j+3uF+v5lkbk/uzIhUjwhcwhyitGtaHVLKbWY85l17xbVpAY
u8cdHIvee90UirpYDMYG/qS1DeFQYVbMnLzhzy0iYBrMdQqkxVaeylCG23jpYLBZ+pjAX7pmMtL7
gNkAe5tQ67gxKgpoOxki8fEQUFjjzwWSFBpWUjGXlu9hGmWTQI5oJKxwSP8Qoys6xM/xWrng5npe
7cj4p0M7QjIZl9NJMCvuWResxWx1xprNEeuTmhPFc/YKz6irZuiHdUaT/pozvuXIHUm7MHIqr9Y+
DUhkY0zoel3YrNP86J8qkXAKGopbbo4aNNgxelEER+UFpTdnW3GFqeMLa+4w+7tXHxITmy/UBE0L
P2lCnwGB7E+58/K4XOU0NNe7X/RYgjypdbLyRF3hLpqJw+z3x5z/3nDWUXwldVNkmZbrI+mhQKyv
DeoOFFSn+4r4Clnfa7rSep9gdFRexUO9/2QHQxmPm19Nrs5HZflUBXI1oKoMM4gY/Zmr/qde9KgW
UoeGeTaW+Vda07ciudNA73BiNmw2aVp4/vjjHTCIJW+pklUrBpok+/E4YRfb4wRuGUWNI1fu5Vjz
prrJW+ovIygythrnD3bLhipaM5nxACMWBbw08f7f73lm8WBNsLmPDHw2s41dmNEbV4ZMsNB+k3cy
RxIRbJkuxgkHsoomJT5Ah6Bh7LkoCIgTwcbPOGnbcz7dB9av0M95uKa5uBzMmfxPf/+bzmgW+s2b
v0IiMmaiPGT+Jvrp8PqrExNzOhssuJs4cdrz9bsap0EK6UHcSKVh9s4iyRCTJJKajkVHRUReiow1
xd+1u6ziFaMS7Ig9reIQBB5OvTl69M0AELf/pj0KefoadHvWLEzGOgI6gZKXRQjs/eb+99qGbyxQ
iYCz8wH+9xftqpqr95BEgz/VSrR6gTzml0N+CctemVeeMtFr8myrgJPr6uOErghQH74CH3YVo8Si
jHc5pf/9U1ZPVNFLkv0UFnGuvlxY44/s3s1ubj3nlg8NqOuTqHkazmInOB4WPvj3BQV7EIzdZBv3
v91LcbgTdrBHQriIXY49OFqBof0+ntKIePIWT96Kgb0KuPBTFs7nOtN+c1HHUh4LgJXYu15C1xYf
aGEI5hh1AafL66xO2JB7E+hz4Zt0I1TmRwR3/2zfWBVQiJu1S1MrDyT/Ee5WBfg8MDYjwe0Ra6bW
IJ/4UU3V2ZiajIIRmOJf/JQKNjy55t7Jhn+IFv5Ua1ORTAWi+5GUjlyOHwHCLqp3aiBb+PmUTMc5
5Kg9yW3PIfwFusmkZ3ISgvXMtUZo9IgXJAtzaUHG/Jt6KoFOnMfITiMieyx+VIJ6sV1Jw2ua6exm
X8mj4wrcto9QxaMUKkLJr/Gl6yvI6A3iJ4tszZBNVQM3KMc7OLr06ryDwh71psdTbwsVEsWgJBXd
sMaWU4xoHkuoumSg1U40WIXifyMmzlAgUGfFA9UQhnuEOOWK7uPDVnQ0yvaXT6abewPfSIQ263bY
h6F9Y/PnOC2Gl9oE2LgArZP7eFydi0ztOO06LRklKU+bPIOvDlVOKb/0JC403dT1pHOAKNMnIh6M
g7Y8kQ8as/cg2pLEiAwgcshqxC+ozAXZo69eB9dsZqAL2kp1QXchp2+berbr1CdELF/zq2xgjkDq
iebU2y7YWz1I0GuRb3rT6PhQX4V5I60/RNrflsRcRak3/3YY1CvT3QBPWLH67w/fX6w5Z4NUVilb
qbcCHbA196lybx5XpEiu+QqIt7sIw+00MvYvkJfHmxBCCER1l/zYtwVFwyxItP42r+Cs3Yd+D8Fz
iOei/DYoEuzyx8QtdL7G+FqpbKXzgLSdjmjSHrw25/1dPgrS2oeTyLsoayepj0m20lhW/m0stGcN
A2lTkYn/7l1UYtddRZk9eNnlATz9l9xoJFMib4lBAKP3RAPBqjIfWjcS5rbQwwCX8s2yoV8Jtzs0
odKsofFbWcCtW5+d6gBEH9ihscTrA+L4uHD/vyvnEYXfywOnfmJ8Ho8JvN47F4k9N+BxmmeAXGNn
hk9CdpX/ak+l2JWEEytVe0t49a2h8IErkob3MbNH/Nb07M2mnMzZ1xPfVCAiiimvIFVV681vqu2E
WoFMDo+M6lyQhpir4WpHnEqkJhOnr+MF+95S9BbRyD6f6xlgK83OoaPd/vEEX5+7SdgCNg/wrUtk
gdjw2IprcwKUxxIsrrxXwqfscOIAeIJrs/dU2/sibngTpJdzU7kprvoJScedmOZl5oMJSpb4ly8l
oXypif0RMBI4d25Q6S4pPeRu3VTBm5oQIR4uS4Q71xoMPYG5mYQrcRaizzHRIgg5xlZ1lhFX1nAh
Kb5dgPdsrdNaRYq8BRg4P/vXJZMxSwxIn4+oL9DGnahKhe3MERCIaTAySCf4e20wfxFY4CNlYavl
LGJD80Zt2GHNXHsYd+oenoEs9yqcUTHd+ULHBKfShHn+UKLgglR2VuC1lfU2rMNYl7X3rOJWbhWL
a65b84FrzcAym6qciLnb9ndLsngKn80ynu8bVdvMS0IrlMbsr9qcdDoaK60/TQykCrqpd/lplxwu
ULt+pvZRyxBJUZOh+gZhZYO2lMlF6T3h3dxVw0vavBHfQXCab7VOl8Ybvm4UmfVdslyUkGzZzx0q
P0XiC2y4y7chF0yQ4SEcIxcQqw+cyXxdteeb+dO9l+rw67O2i3yVAr0IQYWVYFT2eyxcF5gqUl00
ansVW2JOTzEQ1MCg1mMky9Zf8kY7ya+eo6vBBCS6+SjkPKqJCLxt2UPykRIwC6CrgK2IakA838Bw
AtXyopEnej+VgmsgcWwIM2h6lFeyMVohhB6TMnvxQYbUIgOSiQxUYFzj2SxOS02l74GAfYUfgY2P
nWft06d5uQMjr080cVLSJoneXblEta913yA3E4p2zCMzg5uCmw3LZg51DQ0FWvw+8TdQsTVLdUEX
G8VZkuGZFTNZaNeVIteFZMoLYs9gjB2dFCiiR7WhvZGTR5N2556YyALCCoUFwEjAojfVVYAM1sbE
xVGxQgl79N2HuHP4qXbtKFxbGilB4a1zz3wa+0n20KhVHC9zBQTcxtTs7HDOCVq9y3JYZUNhLszy
j0xHId0zFI6Ngrx7yeaTa6AWSYsyP1Bspf82V+roVIbT3UT/233Lue+9lhP4ksltKMQEHdwtvOM/
NnWWKBiS3MO1KCo2uFYkoUJMHcYQsVm7gfaZC2HL6nUDJ73XevI2/Ghz7xowICO/yl/SG8h4h1Ih
Z6839i3NgKf9+pIaErkfD4rj1QMHClEW9W4s4bIUx7nFGJhWgoVgL6Lj70lU/0b5NmZo4CujdzBk
1kAefXsUOZxeX5rxcLjCn5uCMFRyCYW3QY277qldSLXf8igTpkuvSd/lCetO8u+R+0FV6eOzyynw
iB1rYsyKHdYKeV8q8ugxcPJ9JwIp9MbGYF6Eoqng9tquZxuU5kA51T51e7MbfBAxjGxViHNz6tzB
1QXjf+LwEO8Tfuxz+tEEzIogeeS1pBtxfugtSH0607tz2wVIHXKYdNU+1amPxxaUrfxk+ih6v3uJ
5fP/mqUe0AePrbF9111csLLtzVJA54libQIg2cdFpxM++3A5fBBoCAbAvz9PDDkkfMuz02xTB2+B
kywUAVpm7i65kIdrixfztth6dP+NQcQGWGEs1aLrt7lj8t67x14GCXm5SKaxEg2m3Qg2z+7b5G47
IR7va/8SMNXQqWgeLYYPUnjcfcz7G5BBec1M57XTc3uJkPz7fffea9DaJBOhSGF0XEcIo0wTGZRi
syYyNcbjoWPT36O/4poJMhpV6WKWRDvJ0oiHLblEYj2qykoQN4QX/PRcVmxX4zqXcv8QDT14EJP/
8yhEO0iT/lJjjWrDsWSWBRrtdHoVPzogzJtRFIxnra7xyFCBFmw6sxue+gI/GYYzvXRmw37gKQFJ
3OwSFrJ4V3a37lGf/BXNpdcuaRg/cuqPZI1qaV4aiYxAThBrg5DdLjigI4DMVK+KMTLsAggj7gJv
yfIBMc2fgSVO6Y6sdQs82irnyIagkbHoIfTFZ0BHqcaBZWcKMj56noBpFv/qe5IdCvgnJ2XLCVsz
sjprxY+2fAndoon35hbhatDpFTVxec890M2Pc8jfaBWcicqODrgc+LmHNp5khqHGbzMp9z97Gv8n
FQM/LiOuYRtWJdYn2OoZ/hVzSXtmSgOv638ch/SzZX8AifyP8ul1R4+OATGOLNLNVLL3ilDQlA7o
OKwej3zg1PNUWMVV5bjXvVbPCPZ+JSof2e6kh+siKBtBnpt4nZPp4bHvDc8OpHyYJX9YJbfckWJi
FxRqspT67q40yxBsTPypNuvNpVQB32YcmH1R/d/0J/VgCntlaFh+rRILtACHCF1z2gbxkdkWq5Uk
vgyOW9YC9udCgCHfUiNbDwujsJ8qH6pHGKdYXHi4FhFvg4DkOAlEfLVZgbJLfqi9+hYZ92s7zu0L
7pKthwB0d1sic8yDxCn323/KLLmdDv1b6TE5mIaEiC/RUZgFeruqs/eaRdfqQ8gLKAhhLkJoeD0P
6CtJb6J7oF3NSLuB8hot7W7PSqWT64KPb1gCUY4K+xyO8gkb6RhU/+5fcKq7VEeN4l5k/+FPG/gb
oGKcLPulssKGmJ99QEkjUDuQrt+TJLAnK/bKUijj+wovsqg70/bR6SSNr94iu9iftCHUT2W+FgU0
6uMzfcdGxhJ9BlFrL0pkHsEzmZNHX9jZM6BJ956Wz6zGKfBHCTxGZf8bbdED7fVg1PrFn7LjupBa
Xb2JmhvcZuH1VomPtL2f7HZeo5/Q5V/TKyGxth/4o/py8X9bEqJTW/LIK3o9FTmELOQdGvS6LGM7
uAEZcop8ZMMsFVCe9Mi1eO2mB1ITPg+2PuOBXXii/vSQ5ZrZjhdTBhb6XI5TkCj6ucqGoUwznZXd
SY99mRv/xLN28cZyjE/P3UJWb6aYPyV0yffvIBc+OIDmPGZetueUSTHGGnxR8lKImi05LA0MU/Qf
DQAmvGxa2ftdgcKwiiHL3S++hIL34mZeAAyWaLgTqDMuvjEjR3i7krT0w7UrG5dw2A7G8R0yiYH2
1i9nAQvncf4U+/duc5bqCGEl0SKAJ+3Zb1uJL+VHjMuotNndFpHvsvbCLfKggdRWtRENQoKz4UY+
L90FPiOjEIdXMWQglQYcc6iaTk9i2lyOQzTtDy8g48K5rM1tVxDznPEAlntLZgCex2WTH673x/H/
m9sseqiMqbgiYAIWiKkNVBRiuof+q8Y9HMPFuH/UsLyDSFEVtaHXYJ13K+b5vNiX1iu/bAC19QHU
yrac4WDOEY0K6AjKIkeD3ArFSi/VKboRoQkD81qzTlEm5mJIbwWUWNeWbmFzQ+ytSp9Wgf8is0bb
Y9GtsYOdusQdD0cRasiYIcxqR1HlkeVIeQWaWJbGyo2Zy9pTvxGffGx/2Z0Gke0tZGkHeVlavKl+
R94nzOOEoPRR2KZsnADSKR25T6kAInIK4i3U5NBPLOLGiRk6E2jILy5OGCzFWYQYkNo06a3pl5NH
3YOzLBOdKkQZ22ap+yS8elb/nl1X9MnJbqZgjZL8HFlmcNyREA6mpgr94c06Mm02dnjPBuumXniG
TTo8EXsz4t+R/IYtQstAePUclKxp3rhfk+cVlBLwlKG0zqNrxE63qLXkr3nXpRzi2KejyRlOb9eB
Y2yQYhFN2kgU4npCs60NrMxg9C83Oz3VCp8DSJ2XrSeb3L+S8mrzR7IsoEFXeZzH6COekq+Ipvwk
dKOTsfYryh/XHCpxv/7eNL+htC5z+DaxKTfw/JX0yrlNvZYPQYva2J++C1sfe3db7UWGvdEGzU23
DJvJocVOOPjpDIof/a8kDPd3BSlzIMCxMVaSnOEng+qLBGSiSQfpgJnUhpm01gxKOxi9DMdbDDjl
nlpE0lHi9DZBzrJAZiJG8K3OjUPIlkFu0eQCa6dm1DTNU567Ojx7DUEE6uP+2PvhgJw54QvTA/WL
TLcRJ7eX4lZSpaDkxnE2XH6GmNyS1uY2i0FOkzFQ/rA+6T1StslhZ1kOl/K6JREGpI69NOfLvtXF
UnkYuwo5fy5hia15SrcgLSZS13NouAF/Q6DIHH8pzalYY2j2NqnrfT+wYwYLTeg0f8FkCPJpzChF
jwfhehpy24mkTTG2UIgfXL3jHlz2n0mpjfLWAq5YJzplxsz4GzUhfVHZ9xZLbCJTVNCfJ3aZHJbW
t1clfe+Y62s1CSFpwgi8zwpGU6jj5CC2owsjtFSkE2lG0RrVy4RAI4dhDHSvDUh/l2t/pYptFN7V
xa395Yfrl0S7PR+y+Xr1h4UQXf2HY0ibVJ3RQvXZ3iCIhmbu84DXFQR+z+jbZ68RQEaA0N2JDwfV
FhNXbvHMEHjZTSgWOCvEHftMyFh2XqZWmGGYeJniJmxIm3EhU9s3Up3oAdjvKipDKFav9DYxHCHH
idVTzvqiE0NAXbWzwj2fJL2c1O5YtOnjlYUZ65xBUxTubfayFjpVYWaycPp0mjV4gHIAe8ORJNov
G8/o7ewvfzX4T9Wu+qD6LcC4f3ckYBU8zJK6hgW+oafYf+z+mGsVF52usCEOUb1YBOfO82OStHb6
z0RMrb4eTq0J0TFPErbQh1fUa1cKIxe8wQLUOY5gHdHlztMzLdV9Qe4CZFj6IrUCPrZZOaUuEMFZ
pJTRhYxCMLppm7qAWVojzq/vDgGxTHrpnHHt162NjjiegKEyW+7Rk/D7rXsMEPwnhL9tqR3vDAf6
74p2NSGFiBIIsdzsoBmH4Iz715Pi88Idyxv/QDDEGLWBRW4BEjQd7+Iorl9P+yUdpVZpXwTP+uSt
TpBJqUw2svefhJjDZj6sMG1/VOuTLK+0NlCiodKbg9coUyHFj4KegfZysme1Ld7FInSBujYiVA6t
rQp9lxQAhd0nr/rnv76NUzNw+Kc9I3Oc2uIdStecBSKR7hXYu3u9R6rKIQz0wQyM7OPb/VSN0THg
HlDo5XiXCltfs/WGRAW/a5kJOjQMo40OVIj6tExycopiMNakNEtDzsD19n8BdAp9i8eLiECsw7cQ
TcqlPrTIrsWJQcI6fYoYep1wCWpmTtJXTu2nbsmG6yhBKrLDHS+alUDMuiDL66Byf3EHmNaJcBfc
RZDSSc8JDj4rlMaoKVWLrKA2v5uwbT3Yuk8nsiZpBi/QEIK3nJn/TqbBi4nLOKvE+NQgylh+F//b
sTwtBGfzXkzh6a0aCMOuUl2Z5A5+IoESQ6arl1UbMLAiGTK1wYvkzU8PCZ8U6m5x4uCWL9sfYPO/
4ON/b4dnek9W78edzoZ3mY4T9vuxIakc6ccUsz0CgXEB4Tlqg8gn7IiTrHmpVYqGf6fNd2gd5sOK
gSO9vSFlcP000nprvCP2qKrYufh5BJzIFXFa47CfgvqirBYcTbFmSiJDKNmVhr5UbR4M0MHMutPh
RblSUT4VOwz3QHfGJBfOvGDe7PNmclHgoVoQKGaTLaraMSA5qL5Jv/iCgsRo2Vyw4h7g8NqZUQ6x
QWF1Z7YuGi4dcYmgzs76qIKlRtBaXqwrnusOAbFk2rV21k5XeRzEpXjqAg9od1r6tEXEBApIfw0P
xTRvOiMtEIbVqC4bDD/naX7a5pdkNwH31gOmcY3ouxF6ybucNHB/c46UsZzk/dEruoV2FgzDYko2
UqnJtDshS9cM5DD+mcWMTmBFmKI2LDrPT2emM8B26DTz/hjRH+HXUVoTs6dFKWJfW5w3iygSjVoW
WORod58Gdb9uwrkvrSOZl6HfHr2QlGzleaaEosxWkkE22/+ydAo9rF1hDR0ypsssELybo2vUeZRf
NLId+71EFOsZxHKM6eDFBLpxEXz2TBEwPLWk24m/5xqcHAHES5cDEGAK6j7p86ixjzvrIb9agNq+
ToLpk1hLxRutlSC5RK+ZoX2Br0TjMpZOmQC88PKpeu2z668wwPLEmygTFqTmusJpDiHmmKlHcXM+
nnIrrRAhQtMINxLAX/bYbta0UURGnOOLYDkkC77z/CSnh/MmlaBISC5Dct+YE9Y5rR6xn1ZJZ6tK
HRhakEsXhh1QAk5U4blIDDHki9ZsUdgA7vKMkKmIMXPEGC5kcfxWLpADkXkOf0ixMQb10pDjYUpL
9QKT2QVaSnnbAiNOJQf3Qf2svBv3OMAB17sYi3LtrwI+79zSIuK9KrRMrGeQarn1yHVgGyDymWc/
W1U5LK5QjkZclI8VIgxvVOB1pj+CAEy7pysCIEv4GDw90BmRpiLAG4fKoz33WrN6pRTM3GiDOngJ
IJ2wDD2eglrW7EEvYV39Pyn3CFFNLd8ilYHIpFSUMGGGhHcPjXOrqrMTtIsutwVrg13u/YYw6vUk
n0da46FfMsAp6sJ4YjlHW+X1hRBxUEpXUqWjAgOHvkShMjpsZgpkDgQlNEu1rBuZfbyxGW9a5/2t
dkf71W//0ed9tih3CvUZO7e8VbCJie51Q0XcTB0+FkYVL/tN68qXKbkSlTY08W0P14nb95qhrvs5
b94CtXnR3KOHS2IOJDzB9LQawshFnnkEeo2ZI8aMSNtB690Ku2Yht8dSYhd4XoL2djoQvASASmKu
HIg+68HRah6x6Mwy/N8337ZBhvzGISIHYtf8qWvYXacov+cmzUcnCyAXUoeveLJduufWymP7FOCY
1uWgefTsi/s6gj4f7S+bQI+GNuutng1vgwWSxyBl/WvrWg6xJLjjTMykK1ZAJT7JxATIvoj7oqb1
f5ANWu26vU8w/wJBwlSNyRcH+UxxelOJKswYczMEvh78W0Mle12N6FNcEbRnPUJ+TSV+sb7UbcXk
0QB+tuP93zjOUKGoKZh5vPWnr82S1UPrpIoguILELG/gJtX4TtP2yXR1HuppoorRjJIxzkDCEgI+
U964vgV4Jn3MrlouUfVO+cFdGrcWwzP8DGZx6l1JRq7HBrFLAFB9sfd+wr37S77voBt+rFSMdGMI
Ww5E9x9mPqkWG6dtknioCfuwFmiyd+MUP72qybRpJrCn1Cs8Sc86cP/HIR9+40dAQZlHvuvQ8/2M
Lf22xXiiw8xQR6UUoV52oAsDStr2zldom+v2iGIxBEG0TciqEHBTK2kqQL0Taphv74tjJiKqkepo
zRCEyyZ2OQBqQ1IRF8Md8//Wj65IOnWZRC3FVqOzF/i50AI1MJEwZRo9sD30/CfmH9JQM0M3U8I9
JcXEUhXQSZNtslFAJiSSboavuGROm3WPt5+HCOF6nlMp42IQUqsfVK3sxWdnFJG3DAM7VlqiBHuv
wqf1Ej5P6M/9WuWiHcjLU2TmOs5TPdA7fQmr9DvhNaaJ7yfF/vX7IHwMJmZ8YOpjXZzWklJEYEoj
+Me3ckaJAx6RYteh77Ux9eyY7yg8G8xpN+5W3Q7LrxvMffsGikhlbj7DRVHesd8GKjoNmCfYtHLs
DuYCi7ZugW+pg4F8+au0FA13Qkw5O/XIe6D6RWJBUbNMYYq5jDN/9D/8PwQVTCFf9ZOe0I3Mn4fx
CrcGY2gHgSLqqnGwreJJI54H7eGH0Tp5nqd0WVVPIoe4G50lzFDGo7usmQ8Ts+/VeZ2zq/LgnVfs
z1I/Oki6auudrrZRYN7OCzawC+A9xdZKzHuNFkN/G/692uH8/7BDHppYKFzduCapQy68OA8yxFxu
oVLMP7I/d0urFHKeMyMDUMT7SqBBoa0pGXeoU+m309TZ4/DaeBALrcTDvNJ9AXcXWoTEHHhXk+LE
U0Ar4njqdzKJZkaoiIj+u7KlgKjt+HxM/f6lJEm877JckgxXHuYqnsMGb23eK6QeTaAZU/qAXEW/
t/6zTA6UZbAzi952h1BgPj6pbg8eYfPrmq4B16EpQpVxXxN09vr/8xBQ4Ox6w3bswkRA9AMX+YIq
BktkabPhE/6HH+1qWDldcPvc6/oEfCmqCm1Yx4m4/HJJ/HaQBZu2RMS46onc/9+8GqQbQxlIFL7g
/JJmZX6X4PWYkEGVoXhlJ9wRO4Ar1rDppM3tvBHmzj6CzFdLqRfj8avzxfexXwhdOVbdoBpvQIjB
z9gGzWSV5m4HGRESVo+/tz12zGrWSOHj5PYCxFlc4yzBa14F7Aga8RM1Mk5L4rFyECuksDb3taHe
qalE4bZwXNF4sxLHjYVxLg6du19sMeW1SLm+GAloPWHDxuEpaSagGvQlbN8gAmTp6MDjkSEVsBab
Tteqy/6Y347BpYip6BQKwbpOO8RNOfzvAPQaMjBlPAH23ltPOevEoImpBLeqCDj/PFiliBYi4wy7
iMp/EUWZ5W9sQyyp0l/w0W1Q2Hlyf6kAtj2HhDljNwaTV88QvRTRi4Jkk74I1PJF640WWCu9NITI
NQ7kQIvfudIV2i3MSM4gm1/d9oHI964rlTW8lj6wSvFK/q0Zmum4GyXGY6GrfxjdKP+j7iiJTc4F
SQmZXV8TT7SnJIN3XhUR2eJcXlK1FDrBrSEax3x5qjNLttYTX7sQYqriq8UFmEwwE4GILJCbgZtV
AmLoQkuriKHkA87VL97jCcc8+Ap/m1l49xn47gPlCOGr/YeBkZ+jHu+MKWexPZh353VdLGxD2b2a
dOnxIUY5WG2lovHqGsHhDHzNUqm/U2pesUlIdC15GD464pyUgLl6/J494dYXTQcGSdNWn50vt7VK
B3Oa4B077nMTB3F//PWzngUxa14Fa1+5NwSTnvdfZV70OiJcNGtXwzCHEFpup5LB0YIhYVf3/ZTS
g7E0PLjCAIWGWWKkYt8Q50ls6Yxo6x0Ebx62QCtRuFV+HdJR7ibiN6IDPKcPb++qCLBGngdwDAkE
/Wy2PPxsMUz0rE95KWX3VUk47vKB8sn0bZdqflRhrr4LPJGuM3+wCFNEafpBKAqt07EPFtlL3Dv7
Q5diBCxcNTG9RX70ON+YdT/nB2mMLnxjcZX+E+IhC4gfESZgbFVdrOIkNyFOn9P2D9x2YG/3JhEX
A2iNYUwzjCQ+xreLcYYMY4AYmjiXSfo2OEKE6ZAoFFpLYoKzQgB8IxSiBtFrl56QhhNhuIUdBYZx
qBz207zPbECFe3DYKoJPe1emRAJjol1mzJICn51iUiG8YrBUE/6KEHpYU9ism3pVThB74S+pPK2t
m/BwbkqbWizb62+ymuNMDwImDkwv2DqzkvbySIwJRlvjqCXpPVrYs4xHY6kEzDJUpRffQTEhizer
qbBHPgifuKSKdSProrNljMA0Ti4C0jKeP0xgUVOoVwmA902KkCl4VUpFtcQ7W9CMwUJiR0TCuch8
AxwQkx1BRWxSwo2BPAZcbYu0HVhRCS8v5iigWOcDKYJhG73pQdvbrQD3lYFfZi6a/dlvPAIjCFnu
dnfTwa14ZWrFEEu3Guqdk0L2YlYy4FwcAQAJVkDAwDBLS6yJiFnDbbWWAYHn02PMQ5B1Mkpc5PcZ
wGnBDTV1cFDjMrOSkdW0HyTW2TekiVqSZKwCWUxmdK9vdizCfsAhMJdYpE0xAwAwwZstA5/b+L6U
J+Ty7JlUpFvVy2SwpXwuIQ7cqYdY7oV8myUkbEUmqWUD+rzPoIVFAVY2E2ZJ69+KLHisPRhei/Dk
4hV2Zml4SFi1tqcgVWdNZSzNbsfGfP5sp9u3zW9Miq+ZKI6KyTg6+U44S1EPlX6kEECu1iFPPgLw
U4wRCNDU2VvQe+7n9zL7p0anM6c1ePudC3fgeGAQFOhxpCJR+VgJC2G8XG+BJekwIA4X43XXg6g2
JXlO+/dcjKrdy1CepXmtPAQLGNfxBp0aj45pD03oFzgiBbZQ/tz3rTY4z3ieo4k3yHF4GEp3aHYg
t6mnV4uoRHUp4vCElIJy199DodMaKeYHSDKcMdaaJ5k7jUN1MwVDHDDJC7I5hJ4OfSGmx39PIfFg
p4FDMLAdkRIp3cnRVfrW7d6RUem0b0fpe1GKUEc6AISkMqShsXDwPsXcKWoi97HeFF1PrhJueB7Y
Oa2Ar8smV/d/4YAZNcxkeFcdfYIWu3EYLQIYWfhpr6sTGIY0OGyVPz3A5aPHGnN7wdcmXRLfw1gu
oiFWVNgBKQViWmhECN8+XqcHXcjpfYD8KL0F9C3QgPfIaxDTmp1Uqy78mSJVx+q4ff5H5Hk2HnrU
8CREi/Ddp+BYqAjOp5kh+653WB+fw5haasl1kQoEV0cujIy1/QdyWJDValvyaHEDa5cf2mTNcy1B
X96RCpubKt0dhZsofyiHKejFYI/i/mW+aC/8K2rwl1iKV66UyqFZ4YurXGUYEQ83pQ+hL9rwmPOI
M++YV9wOx4i1Dkhhc0GYVuCmswc+09myReD9p1Yp3Uq9IKak7m+EzIXzvrmo+YSuB1srQfSNEkfG
sQ/fDuBjsdCQZQ2SR9lpnNLrAxz8I8ALjIIOWj+EpxVFKAqd1ls2kw5+M79s3KqKEeSnGxdl+yVS
R8uvmu3Gt8XmqbN/PBs3hQ8VEYvC87+33UYbSiroBJhR1BAJQ21lU56txWM/1qoJkDFbYDCKLeOv
SdCk0fjyw+GrEm4Mx9QOagAygiSvxb/wvc+3O9Dj2xPw2NEM+Tt2NkxZzvH7shP3k4rHHF57ZH+Y
lHHu+d6dpC2l/DtNVa0EADLFtpuzPrWjdb0Lv69FhJGQRYe6ItDdRNqdnH1+UmNac057orpaNWDQ
XITkWjcMwg62Mfnn2h0DhXxGWqCnSkuhdbJNsShFR/NCx0YIs/zq43eWw+2SYOtojVpqvQ9UXqKi
+VMO7rnrmRGIB3wWCqTtBlpA6JWOQGramK/6mtj9S3LcUbg8C5sXovtkwWGlQ1ThQHeSylcU2Nu1
oCc5O/XpYnYId7gjG8Gud94BGnx9mzjIfkJCdfaqFxgwSwaPCXGVGMlvWjRnmyNV3H8nLOoxkIWd
JkUiXjtKtXmzKLjz4gre25H08GjwQT3gLhB4cLcjgR4X9JAQ+Q3pNC+gZKMeKdFmX/u5Ylinif+D
NLVwjaZvjyx2RSNEVxjFUrI9vsHxs6E99Kg1W8fnOuKLKpIlJt0PFBZyu+v8h5XnfFXUdKBw0kSH
WBDKA6YBbYfUKqKRN/TlATTuG4spXlitZmhdJQHTSeJrcMAjX43YrQUkPz3+IixCC2lf+EpCfYmq
c14gKC5vmSVRVpt8mg5E7g6/HVW1nwNgBJcGlNPkBqRvIkYIVXzxhnKXZTAlEG/kV77hdlCqLBMi
VDq2vwnWcWblifjGImtdKhaoLPMwGT4Lo1h+kk2+wN8NSwwX5gCrgSmWHdcWOF2GvY6pPCQyB2RN
owsGJxfQAFrUSTy2ibyTUGbgf9rmOs8mDL+A7wal62+Na96gFioBpkXAIEbNmZVBvBgrDroFZNfR
kHaFUSR1YUNqi+Ed8Nf4a10yF9nGp4XGUEYJbZWmsre9TffawDxrRTEXW29kIFJK75rXdGulbQOg
dDl0pCba3nSs9aMvqRVa7NnOE942d+W4MMv84W3D8x1tWt3hSLMbPOzCftlUjrkQLDvoaGmfWKSW
jT8PIpRKlFEoFZHxpPebuRrekudTbrsr7aW+9NZdAzVWne+J05f1SrGpT7EkSDvbCYeDvss/nUIs
pN2sORVSszPdbDw4kuKeK/zJYf4SsLuaUai3pWlSZAjbw22HCS7D2mW9+aGAFtea/lKJIKTmOH+h
E0xdFnvjWphTeQKXvhkVouUDveHcOS3PF1awfPjQmZwUWLSDx7KrJU3dt5hSlRemAvHChzrnTfaM
CLW4o8NXC1b5XN+KDZgXDNzE6i7nc0R/og4Ebq6Pqjd9jMI9Ls7GLfu3rBnSOyT1HO04RrdqWUYs
MmBPOfcpGfX9q6uowLBBr1YbvdyKxecpaK4AiQnDoZ+NPP0OOw3IJipfQmiEdrh0KqiwuvHxfrsQ
NzH23LlaDuwLZe961eEXpeUvEA3h7mi+uSGDknBWHYUN7iEVGFhJT32Q0FmBQG9ED8ySbSbIzJny
9j2p5k8mcMOCoY2MOlr2u+9fjiHr+nF7+uaKqS9P1hvdW2D6t6d6mWbcQxzjOco585xasKF3Cdlh
KFIQBr0QMVWtdYi/OlO+gbboLvqB98EAwKs5lZJwosd5jPvN6ZbkARYr4n+obKEii7Exla/ERppV
jbGcdZrRfc2itXx4LYi/uo6zIEs6bJ7k4BPXgAJyB7WFRgwlk9ZQUVCei1Yqr6LIQxQJnaSVtsG8
mPyEPDDeg32qQzLhJ8/BCzilbkNP57FU5xO8YG2jN5D6BhE9YRav2tYqLx2Jln0vdxFp/iLl2KBf
U7sAjnssLXBrgMDYy5gFgBJTxpFXYMuDtiRX9HOEUksvjV6TIh4x8/M/9oun4iRL+WyubUduey11
4/W2XO92tI2cFLIBEiEmzJAXiKRWT8c65rD95fxmCHnShUT+0d+UMJUDppUjUA7hOBBqsfMPTqCf
2C8ROCezDFsizvHmGjEEbqFVJSIJLa0tC9Ib5DzdMPlX1hn6aXjlTiM1y9/LoHRzsDe7WuIYsWOo
0I6fyr/vRRDTPEzgEEqzeCn0hBwxqbIelIoRyM+yfa4XyIzSj/b1JU8iFFqmJQz1jpLxf6RjUvDQ
J3pc7XP9R6MD5HZP8gUT3ls+myE0qnmV7xoGpPlHDKbJw/GjDvSbTpd56zpkvN2MTsgnO5TBKKgc
qhH8YDRKhdxaSrouxSu8vJjKRfnWlFnslT+N3VvUsbpsKd4rX2T6yzePPjBSnyPzDCWpjwcFXKh0
2+LBiBZZdkVpz4BLEgnpNIDbPppnhupKT0t9bdHfdrUqjVNk7r0KmVskohCWRt1AxpIwleBYVgcN
irDgCa+IqYSn9FGH7GE8Igu0S4rItOzhTlRivJ0NheNURXI0WRPKImKNn78MK5G1UA3hi2MUqEss
ULYuz5jc/J96U2hN90Mb8yIB16X6vDy+dW8KBZbaNXAFY1q+KGuBqzkj8VXHRn3UP4R9TUTi0hdy
eGVHNho+xuS4bYO43j7aM1DuCP9MvAjRpY/tQdlEIUfpuyLOU058U69z9iB2FBzSn9ZnvlCzI03N
NsK2k69ui/3zdKx7jD5xwaRCjPykDlLm8gmDu1hBAXpBvM4bTHZAv5s2yfGwQKVENflt+uP0Q1gQ
CHRPWrQt+RUBXREz/AZUF7DhgfJ5TxSeDW82RyqYnOrBKfnvdZBKC/zB/P8vVSsO21L+GwwnHTCO
HOXlXiEI9Js69q5rSJxTC7tAVpAr8ByFh1n1PVuWT5cEaDRIMk3o0ghZHy24ghDZT+BmybC9Mbk7
qVitqoSNZvER2E9CSHv7B2L9vwlprd+Eh5Yb6ZJlyL7GwlMz8gqcPoGWP20+QlegnQetvorhldj6
Sh9oS05sgNAEtSXFn1VkmjAzfnxhLyiTXZ8z5wbYlX9An77SiTaxeO87QpxMnSEO9DF4WQ+MwDe0
jRZbr3TGn8DpJc8KH8liwqHQ70vb/lhS8LtEFqA8VF3isUKLzM1df1VsxlTSad8guWEsz6JiEuDw
lULlhzFosnOlaDA6VuN4GduULbDGXdv0JHG0thvVXVX30FJCf8XULOXQBisrFQefkoTTb6oTZdjR
3a0jIHqTMoMqYlSH8GYd68qi+SFRzVQzqMiNtQcVzDR0FNrzLgLV0Lz1avAkgI+FOOGXPSIvYYmi
pB7EuFUHgXleD94YC7gQbmVDFSjx+yknms50TW/bFz4PhS0ZxXUIzuQe8med5PVd5zhELHeH579p
dfwtuZ4I9MLCvQ0XXXRhvcNjehr8MkwBdpA3W+UUe3J41YaRVOhX/2sRXHzuvz/olhoX2D3NV6Ak
zMABWiCs9OLmN8djltbUvlwL4ByfT7n5WFhLVqRcOCVncKfdVq6F29KvO7bk2HGTqHaxLCnlNmPO
yPerKZZeLHlQH+W80nAOedrH+mVR2Yp0zcGnfMmiwXg2Mk5UujKEhmmVQnsffL590es2kga0rHUP
LtnTmwGBbcXZpRzf4qNV/fo0yEllK7jEg9DK8+qvDSfrsqt6xJ+hXT/ZD0y+zmXQczJ9bEg55V4N
ctNjta9p4RkTnwZ5by0lATVdY+c8Lrs1rFlPqVX4g+viyvF8kF9/3LtOm+RohSDY3tZnmFsa+qt9
//BqAJzOtqld9wzFj8JmhaxsMWlbQvrr99x7OIjDnc5DKeuCW8YhihtsR0aAdeos6gbAkypekM9g
b+Cuzld/Lc5Otq/AZ7dSfeJHeHnVK1Hh/Lfl4g5vm9gYrMXwRhvN6rjApemHWWmqoAixDOd6w6HI
sJSQeF9deSyFyVdFjJvsCARDML48EPxK38YLX5FIVtKxDbCoOa/zXKsxF+b9FSGxfBOT8SXOOADn
Mb5EieYDvRmS+xG2SXcM1kX1yPjceYhY+7ypHcE1aO9oikSUdCNnWcMG793+vzsc85O35gFQd94p
V4LU7BSOu/IETbEUnIGOtgcJKCL/uETgwvslAKxEufWxUKyS9DchttYrU1w/zeSywE8jmwGzLTB4
y4XF+g8nLfVwl/zLMCKxSGV8YR355W2RA+VV7+p/F3OsO9QvHbr/Z9RMTwQP5mcZOTlbGFI0cQDm
JbGEic4ZrQpQGjArWaMl2puaSYva5OK6CTn62n2C9KwiIvCelN5b3RUt5zxHxzn+M20myaALKbIp
AUPY5hSNXzs0slTeaSconuvRahDObxz8IRY4rJ7ZujIYEZMs/qHXLSLlZbwa0GO6bQcsZtL9I+g2
Ik4kaKLp2I7+NqQRoDopDSSPcXVozj4QZ1Kno2NI1up6uPa8t63JU8PiiVxhtK0zZldbiNK31ka5
dHfsWdJx9svS6BgPi6ziyspnIJNfJfjIpnTw0RjsGGbq+p4AKnJ01QwTjhXyU24oRPSkha7XasaH
cbZzvIPM2O2Xne0bVigSOd6kZyE8MmTbKfRJF8+QvqpbgA2uMYH/Nff5HEIWXAw1edePELX3fsDf
pnRDdf36qpHmcmT8l28p8oOjUh+ZZxlKQfanFs3b4WExSnvkV960MugljdDallJI7w0TJdQrZURH
ZnAq0m/XObrvEC4ZsL7QyyGTh1UA1VJGz3qG0MRnoUMnpNurp0wuQwh+j17AUyW2YZMQMgNKPTX/
0esxtPxuKLEt+pQFicyS97OquCo/+hNnKHz+0vcpLdPMXHE0Vb8JtgURgXJs0lgByYpihlk4R0Sk
3lRkT/oiMIZIkwJHeCwpTwlBx7Hr/dRqEhTepwBkO1Y6oxMdNiiK6qk4BcB34r5vDMCwImA5xnqV
6zY0DkyhKPFk2jMPjuven+iihZDv5WtQPbL6Zct+nuJu+xyCzAs67B7fboJ4UyTd/cR3nZXNZO4a
5jyFxTlxwzDCUt4RpQZ7Qd4cooMj5htXj0xEjbZXGfIlNspSkU7Jcw+6nk56i3/rc32QTnFRsEyF
JEBUqDW4UEO1OBlyZNCVm1XM99qusizupt87dzW+NcE9qoBHvb5q5meuwFWZC1MCnHQR3oL1ib54
dCzK/B0nQXwUaH7fmShf4zg/+etPrHKajXAsAGOhx0VvY3FeHu4InzBw2tE2XvV0taFRiqcdbdTp
5c2uyvsz690HWR70czO0gsXoTn5J8yRbtLc8VxBr5Gq7GujynIxEZ1Aa7pT4lzMLpKObsbSkiC91
nDBQp6+8ezkr+n/FwT0Qt8N7PnGS8Cvpu9oE/GzPIzGx7hXAmSrY7mEpqDEalXTqEshrr/QZe6u7
/qHUgi5PH14pdCns3sDfiA/oRwHC/PpBsIp/ZODvif8t19tx2lXlZstoGOSCA/GTonctnXUwn830
9AFRY0Se5yqPjdD0kh0iDG7BMK6w8VYEbkCu6XF5zRtVPve36cW6e3MTjW5LiOmyt4rbszrwk8Zn
JQtat8Ngd2zYBxgOD7ArTM8nCYwfkFOqjACoanKqzv845HjnpMnmhLmZLwpB2mnQmZ0zgYEhpiFx
40NhNq8Lo9WfS8JiW130YHdJJu253PKb4/LBvRvyTZ6vU7odcpHuzcMoZkvCHGecfzAFoTGc38AU
fnmD/8vGY7Rs5Ej2bYPo5E1ppkBW7uTLbBJOU6nr15MsnepGcOar0zKgnH7RZc4o3ICwJ/27ZZSx
ZznLQnXsnoPY1mlblD9OIaCQ9byw1EgpCiMrU+ITqx7Zdk4roJxrGmttGZa43vkneTsha79JXN6k
t3YUXlfl2K//qYbKnSSrIvceeFBicCcu0q46S8SjROVvgPDhX7AKEH1zZFjo4xU7uLw9VCvjfBQD
KbTVePPHveLloZ+vpXVJJco1gGgrQGeRJEpaXocbU2D1yQbJrv0n3N4XokGrHq077DxKbaXFELB7
WaYQc/lDIGQa87gKvDe2Q1wZagy332G4JAI6E++YjDsZzvfDkZZWr12V9VHe/JzbKbADXNNGfcz9
5K7AM7+KXs+5nqqBeuM/mq2vGGwqfkZTuGjIsqBhIelJZAjofkNRzcEGdJtS5Bfn8+9BPJLOCQZp
NVCw7y3qBLZJIw5DyjBDNczJ37ZCLrXxSHlV0Ge96Bn9tmTwRdK6f6r5YRDCpdfSi17dpQlucpQN
x2zr/MvEHXP7qla54+Y+IkinZRwnyxmhn0R6IbalIzTZdOaE9mRwELcoKsQfF06dVvspcNDd8l5t
OqJ+t3OWh3/6sy7XJJC4ejTOG1z6wxLOCIWUZc5C49AHfyIdv6D6Mguo0c35dV9GObORy/snRdj+
/3cuy/8+TougklBSd/4Lo7SgW11+8il23qQOO4Lb6p2zO2e2urvFU3hADXcflYsdAts2Ra0GXC1x
zpxEqtxueg8Vf5LsDUME0uF75b7K9pwN8cMwiC31aDNDH98C5kaARLxa2JmirjRxE1SGWtYaZWsu
ph01Nsabug+PYnPMDczfX8Ak3xxSqsPSiCMwmMWNnIxCU6M6590Yoqec2LqAOVCxDFxWDrKaG3Ot
4owfqIHnovjHlM7V/LBE7TRDq2yBTBJQUwUm6CFxHvUmRkb52ikb3RNjT0dALxqq4z1d9a25h4V4
FL27vQKMwyJ9tKCI+RUR2+fcWiKe7v9vnqN4Sn+tJ8oYUgDTUiKT3WAbN6bH/HKuywoUlQrAYG7L
yW8hE0YCAFmrviw98s1CjC63ag5AQS6fkHf1Nu3O/KpuVwCIQ+Yp8l3uKpkEYPOy5jyPUIrXBOeC
xkZo+MjcbQfnyUf7p8/Jajn0aK6P6a4usOrs5BvrxlzubGyw0cfdwLOnapGc3sQJAC0fqTKM2gNX
culWpk1qSt6owJV3Qpl/YtBb83Jod+8i9yG9R4XMZrcEca1ysodsfcByDydgxdVovwrDVsq0IQ9w
nLN+54XQD745Nv6wNZYpWM9Tt3A5zl6sO6lqoB9HZZ7f6Yk9NAJBI6TiPdFNOf1O7pnUi7hrYFv8
rTTt6fAv/2DV4ZEGmgjTjy6SejqmnSOEy5icBg6I5hrHs6XEShN99G1g12hjR2Iui8rtQG2aQayb
QfK9p0ydqfIeneru6Cd7THY6kqSDFyL6t6g/pvIyKdgeZZT/QajpWuopPXeLQPR39oc/pIQbLv7Y
bUpfV4NZ7dOBMCX2CBLAlPM8JkxrSPGklRyu+WzUDBen0OvVF7KY6j0Ba4D+ypTqgjxQ2p24Nth7
QHVTMQWYSefnhGmgL43TdpNL8t+EzjfU5mwnflmIz67hJNI5K5JoIhjYceqESvwudbzyz1MvcU6U
qBwbLq07MKcKRiLaNcH0+ug9WI4NymDdM0PhtsjvaHqA9SRDbdZVoGSFQJPiDifuPiCMtMjcLnMM
WcBlOKT3wg8Qn6HyeKnrJyY68tkArxEaakRzHBZZT5RwKlNM6R7xLTaJUmKL9Ho7wRoJ2Z13Zi+a
B7uX9SoQ+JdAbqV1U7T508S5sa66NTv1unzTlTj9ruOiqfGnY2guAt3oIH7Zwr4WPThFCCqiQ0bb
YbcRSv/k7e5o/ThHPf3n3Dp7k+q+RMDGUTO6lHRZidut49F9ze3ohF+sPM5edvfVzUcy0R0n6Y4y
8NTvTcmSQHE9TbK0V2lIsl79V/dzSsu8y1SNX0rfZN+BLFFvDscL0dNj2qFEALJIYcAOEAtyhTal
sq/i/98De9KV2l12MApgw1iKq+EdwoNNkUDldhltJAVQvTC8aXXcZb6RWUfXDgepU2awWccwxyTX
5j7ZNxMjB05WFJUNqbwkFZ016g8pkUSRlGGd0VLSoJPxTBglTJeYb5TC3UOIBJmmH0AH12mgglc7
v0b1d4oroSisIkdBR6GC7pw9/fpLzdcksVCF1QyZpW1JG4f4ltD66B5fgbPkY3MQf6LFkGtwHMQu
4KrNmkKe0wId+8zEoSx5VVoO4bjy+nrdty5SlvT9lD8VJvp26Z8jaTkeM3Gxmqzv8ZlJP9QijGvI
3PwCCzhHZmC2SR9hQV9kAHgKLOHr6eqK0KhPXaqcOurUfCr25XadaHktnhl9t5ovXhzwPCw8r0sG
QTDKU3FL1zZQI+3ar4VPL73wSrdwZiPy2y/NEPNu8hLhv8Xap0WCcGDM4IxI1fPLoZz3+UInXTzz
4m0gB9iid/p9nsq5KuOwoybkn2xA2B4s1SDYMveciUffQa+AhpdHTrE/+3tH6ABDqprdE7K4NXHg
PKeiI9162ICNN1ppkmxLbY+K9qL9P9kK0pdf+Ipj8+W8RSzDi6ryZTWDP68ubzRGRAH2I3VRA0zz
oTv6eyz9p4ogTw3IBqCzPOCEVZjtFqLcFNbFVZ20V4qyQUJsvegKBKu/fqBbzaUFKMk+Fy9BKb+y
VoFXeXTU7Csp4fQTVEoDBmJjagbCULUmtBgZMVhZl9arLQop7S8lUKUTlplD31u12Ta4rMo3VtFL
9t7q4DeEG4DRo9uBVOgqvj5XnCZA7JVgPhZnE3fHeL2dik7VqqSss1zzJiXplkCDQB8Ph4Usgwjn
Q67BSJP2pcxpo1oLzKMP3w6iZkwXyjkwL+ht2EJc703pPGuHVZcz8RKPERaZDGQhQHA/s1+ruq6h
hGcxSYGZkY9Gk4BlygKnCtL4eXmgGXNRB9dTeVa4FinKYzrLvAyBHWyHv8nYaCjzQLlrKEKVecrO
p2aGvg23MzEJs9u4/kiCE9a+vb2Yx3j4P7JCoccsTI5eKsk5yovlu09qS/vri1fpPNTW4UzYZQBW
GDwKOH83PU3AIDGelHeYtJWmf1JQxXJGsncPOU30zkGd9rRkJk8POPsbKi4Nsie5B6crX1SCnUgs
ZVZhr9ewp6nnT41VKUchETxtJuMofSyy1bLEyi+kAwTg/RWT48T+W/x5gj9UQhCCz+P6iFJgoN0q
AvHd8jErTwVKHZC3iugSx4SMkPhQQfw8+6r/NOY7lGDEz9RB7U+lx4pTpCQVMFa6sScoSrIydSi1
OnRvdbQW063WIf+kojYN+mXJtUl7+FFK4KOVPb+zzLKGlJyv3IFlRt1tF+1dkJW13smU3SAiruHF
VhIJp5Yr5CowhheBSNebSAZ3Kbx9OfSzHsC7su0KFQclpJJ9MjbLxtRmOXuvZrjgt/R73CAPzBgD
JY+xC0bvS4QctdxDrcYHTJAdTGa2t0bPAXraBAcSnZhQSIbyxpSsPPaJSIfcCiJisGiquuV9L5mo
bGlRaLJH6dZZRhI3EADLXFptWoVHGZxJ8kOhxxpW6FpJj9EEXiGR1N5n5A8dLQI+PFq1QkQVuBaM
jBmlgW+L8JNrDb+cbHjzJLknuOThwhnaxRWaYUynN+7RKDroPffQN6Zm8IzOhNZDHVad4F0uH6m0
4Q5ChrgFg55G4WyUd4S0qziB8Tfr7qCbsnocI3fHm945tOugKUeylj1s9PnJp+73GB4ai7pWX9KP
11ikunf9w1iZ2ZGgrKiH8pymmcJwxrEPqDDibxkE47jZwrT1FhRF6D1D7Gi4ANXlHCBcEJ20mlx5
1Fs8dRf85gFoqsOAaBtZ0TM4x1MgMQCQ3ZEbpw2O6AYoXSuQU7BUbGQ8v1T0PYlec90ATWtOwL43
BzccR14ltPdRgrnGoYZGlJ65JXBJ41Pg4t+jI+PPXWOLYGoFRGm3uklslqzeVMJceJ2XRE6LVKZk
q3NN/0aUNIwp8Ea3jrick1lyHomJB9Fo85OE7kmuP3/1ykmaAkrjsskHq/PcAhS8Rr/vU28j4IXS
qYQWR2tVIQ9kPLnCU13wmnLlIaKHZMhCOQiMlXV5cx2n4Z9uwLTWrbeYbxpHdV0AGk/zw1iRtqHC
zvUDmVaGhkdvYuyCJSCGd87q+lhz4uw6vtzT0Ow0cj7PUqudsaalqcUqyXBY6Jo8ypek5o6FyMp6
O6sjbAUHI3x3dFbWe8mU2buLrR8+kf8SmIW/ddyqKAN+YgcIJ09OMpW7+1cEtNoi5E4RpOUeKT+r
nQH1X3vQBRulEFxmHjrvOWZresavrzoIIgkQL1J0xPZouJ7aoKbD0f0k0IGfA/MmLMKoSYrRYiiN
HmlFbuXdGddxd1G4kQOljNwuVwBK/wtqEVomHTYR71CkA+lrjYf0t3wNSsXSHFf1bijKkJCwyqUp
aSV2VGGzcPmAxq0q8QIvg9XtWlxUN4pdRn4Ab7OHdRMdRCS1hBnfCjbd3IekSOc8Gk78IqLFhfIC
Bo1LeKOxmSA/Vx6AClktXcKPvrjyhEoIWW/TgGMTZZ7bMmF5xPa4rrTmKDkX7TDyEPHreFdgQ0Np
NtY/NN+NiNMFvI9D4BkB7NkOrcb4tN1bA7Af1xItHwQWdSow+Lja8ta9k683//uE8PIAHDK5D20K
tZVwE9tz0/kTr8v73Ut9ywakVYOVZ4mZNDoK3R9gJcK9Rw+02do+2CsVyPBwZDZe8jnw/cp7YdM8
Ks+lC2hFkZ17DcbX6I85b5iu9AzmuhHe1i5WNwv9nljJyA3EQMtnyzFefniSWWI+ObUWCMM2z+RF
1u7IIEq7jRWbU6oEpQvH0yxV1fyM3Ak0lG2nCxDwy8/glCbynU1v7RXaqUJwwzgW5/SgHilV6hWK
rh+PWrU7VO7z7Z+CP0HmnAbad+SoEs/BFUIwAHnO3lJ2ic2Nc+7XjzMMCwMwf6dfcoO+5F8+xuUh
XoINsBnRT0jHP0xgz/30GrAWv/sQD8E5wf4ULupaShWFX0Wr0xsRyJAqwOgdsoYmtr2fiEoBtdCO
juXVM2UJFN4jlNtflZ7tLS5qcwQqrEziG0b9pjo5s0IjGd/T310dwr6q/KbLtFoEX72/xfzldHnZ
HDYbXKR/A74wABaLx654VbY56YIMf84GMZWYngAUBxXnyaiiQjqh1bCtqSaYvYxxG1CVikIxcAbo
ySxOZ72wHsF7ks2Bau6ATGTtNAYv0zL4y2deQMNoFRl/m5cgSeRIxWxNyUjAi2ASYtdWxJrYQxW3
ZF3BNU76NnSq/x3bjqKIYGa6+0tDfqLJDWzreX+U/ttR/TsbXvPaHFjb5GgIgwBH7miK1MOJLZFY
Xgpb1L5u/FFCXiyq0ifuz64feooFQJqJlxRxKpZSDKSzQQ9NFUewzuAF7xPybupcBK/JIrMetd7E
kfWWbHTsB+LCPrBvh5zZ09Vkc9NvJViBMOxliUIc3KvVEwZPkkXCWH/4+C56jsitiLCpW9iJjbka
+7foRfi9N4eE85TyIr/XapmCTyqbZsC2KNtnMZjvJRQRNqz7B65tNtaNptbafhePoVBii4RugaCz
hSR1E7AoQUwAAGgBNgqlCEv8usD4vUmV5DIdWsXiBnoYwpRv2Wmg2V8F0hNThmwhm7fL1/GzsEuw
IM9g9ZvQpZiyLF4f8+t20bwGD08Y5xAU4nvoSWGu16kprK6VIDtEd9DvVI2Rc7Hr3HC+qeAqTXLT
K0IWLsd4yKYASPYMfmkg0WhcxqC4BZhEi/6FOeOE3qa7HtrRylF7PnelTGkprEXFWDhszaDs8L7b
XQBSsb4e5EGkc/2IMa5S5b+rrLN3uv/n0o7VjLJk+tiFzneWZjewPdgzn2r/x5LpVRY/aaMkoTuw
4b6n2g8HX36b4e+QF/nMw8MkMvl991h65U4dC3pU+0eV8X7kiMrEonix+emn1oLpF3CDiCuVpFsn
uz1rLny771XkUCwqq7l2PySiv+Lg20oM9ObpD98tR3r0dMq18+2C/ngsIahYbkSd5opQWxxle/L8
zoM0gLZ2LArLo4Dc9h0rxVj5Ke6Zz+ktvdN0566vcTAt8lgb6xmdtfAAQBZGgybPZ28Ix3ka2iS6
f5RvwglelN7Ec6E0Z3X0TnuBtPD1pYJ9xGyBAYURbXmrvinybVimY/38UzzLJjLuQpSZpt0cBip+
oMMTpTZl5ix/Exxdz/y2pE6RQtDT1hClMIf/rSwCfI0CQ729JHcQJBvtnPt+ak1TCPlUrBmrE+9W
97xtIxnPxDfESJXkdiUtxSUmi5UjPV6z2ZIOB3rWk1dQwiZKe5r1C2V4hECFUI1ugP+738hsEJH6
vVY2S2wVQ7LkVHAj8K4Zb4/ns4dWGa3SYcRwBpFnRi8mrG6wggeTeVkKkIxNLmrBsnMUYYjXQcIS
LsjYGmxfNzC3ZyIWbfX9ZqNOvgT9ayWi3Jva1RADAtwCLffRVbXCAJkx/jOuN/+OzpP09iUsM4sI
JbFucYS+S0++oe/5Zdp31/gYxeKR8sardYnkz6HYYY274mUoUzVlRYWIzUTxplTWfZttAgI0aNWj
yNLdBZrZ57XPKQ5WcTWHz3ZXie0TRMKlH6dbPPm8AJzELU5CHi6DxPJQWDGhP2L8FaGh9cyDcHWA
hSSlpAGdrwbKRDJIPj7LU3rdgdzg7C66p27te+DGO0uy7Q8hwdZHCyuxtH0szUjYNJQHYqTlzdLL
zfQ1xB58zOqStBKwK/Bf4BJtwTC5WGVEM8Es/7Q8AxpYUu5Ek5HJhuhS9y892VCV7JcVcCjCdMbn
8T7u13YK7kbsevQvfnW5DecfmgmFP9qhygpl8fofAcELk0+FmpR2fK8d3qsyKBaboqb8isFYFeE4
7t1eFCcsRjddL2vGzuq08rPl/jijU95igSxfI4v7sAdCySIhd8g6RoFPje+mDDk8BpZZ4TmpBKyk
juT15aLy9RGPVllz42ZVaK/RP9j3ngRwSQD4ER4n1bSHIOeGsSOXpbVHxcbfEV82bZMxuf6vPZR9
hpZYjgE6BHlc9KVT1JUym/NEyLWMuqnV1M8G+muL4B7R5HFsRRWyOmNxxkl6LxADObkJ9mhcA30n
Jj3efu1bqrwrceKJMZnKjUDPNRNkGg+mu9qeGqHtxWNfUzoh2hTwsyusJUT2Y0F5B/kjeXTL/CQ6
IN3T5mtPXwxagafL1CD8a5AvaOZh+OfK25lCseyDZTzbJf8X1gf5gKQCYFc2JR6fdRq6QMRktSC8
cxheY60J9QlWghbTWMmuK/x3Whog4y9WauA0+4LucOddkKhezhM0TbDr0uQiMLA6WHDHLdM4ymWh
HA4dTUNX1L0mS2RpGA+rNpor8PxqvzWOQqZcVqc8vScRHEadpwWmgdPOvHuFXoAhNPExqNiW2RH8
tl7CseDExsa3HBUqmEOyBBfZBOtwbu84gT+C06Iz6NU/AxYhbnYJLOtk5KB5r7jRmzggfQUInRDk
u8ldWO+f7sToFHm/EwaCNL4j0luLZ+8ysM7WxYiskZTD5Km0ngLwL3/5XgGpEsunFEidzuRQqiKx
sy144rSdnAcK0yhBKh+wyprGfwmjG5zO/1Qq/BGRxTec23KJ8IfzImwzble79FbPKvif1/7w1XwZ
arBa5nIPAtrjL0Nul0cpeLoW0khEvYuIvoKd0O61FSRCaUvChO9UPk2ouwS70jR8GTvVKb8j2YG9
wpaHjOkE75pwdNNFBSfrRoGgR74JL1J1Dn0IoocNv7Ix9Z8VfsW0AAYcle5zJ8BYMpxIv5y7m64Q
QcNqx/GJQ+W9yVaGkGp7Vy7BUEyTewN6RH5Ux7OrY3dfCvUYPSRNx7ugDpk+hNhJqmDG82a8vlEp
4gqtzaFHssuFM4GLAFh7RVNQdj9IvZ0e+5kR7J6v0DY7MeQs7/T+7d4M+0skOu56CJde9pdZnUst
QcPAj+6FGWw5tkwK6Ybx6eTmA9tJDDEXRD9iB2Ae52D32SIapstQ7CWr6FuIfSfC4U0t8B4BE1bX
slnFmjPDBfbspBlmeSOBIC/kda5+PECuNP4xNSKFVXa+2CD4sxHcan9nkfYRDQQTaLyPJQfL0tKb
W8X/ayfHayT8w/s8q6lDh/Ul4U4SoAyIbNSRx0ZBU6wVv2vW2uPmhHRif536YGFMSGrmoVQMSwrA
al9IKt2OIA5/JMd5dK7t3AuXuI8RDi754CVqG41LfMdsut3h8AOVnbvV28YLKWORLsIxo2Q614n9
sd6t1Px2w8ZSa37i0/31e+JjpNtxNxEVNY5f4iFnDUVcuJpHx8XEa6wEl8FmZIojzrGhJBWmJosk
QyM8UzcMSsOH744nk8zsYRriCEU7mu/I9Ri4b+uwzSibVTtcMuYS1owtOTqFIVAdjryiZQEFYlnX
N3PDrE1XBmssIsbWzQ80msfIuCy2Y/qJe0ywG5lFGklAlhl6zjwzl45r6PfnhCXFDLXtizSTy83J
EYl1P6XA8z3oBVIX/912acGx0TTo9JApaCkzDrzzX+oHLolsXmLJu+sBhi+G+2QpdC+mfyeLB6J7
tsFDhpBClwRTchEjJaInN9FRu7Yqkfs8cwfoBSTj6G/939p4Zqtgds3wVOX7QV6MwGne+KSLcS0j
Y/RrQojg7xDTyIxkd4sRfkkvlLiWbVIUgZ2wDkJqzheqh5TYxwzmaPsSOpx1xWFKbBwv+ES+Gha7
vdjsaGX+b19EOlPxDflOzCTbOeDwUjuBdw7HY5TrLyQx6mF8GbB9JZ4tkkyysvIwbgvpLYV2rXsQ
mEXHIypx1v2W0Xe12L3pvkI/7wqP+nMfTsmoUWPC84pyaEDYZrbhUEExWgvQavukXVJisBj8BZLW
feVlN0C1ugKHM2+Orx/ne1EZSDfy176UoDAb1ZGIOSC2y2OSXh+Pe7EOJRqaDZPs/xp2lWho6xA1
0u+7D4kFytKbEZebbe6z+gPSrJvFrYgOCDK39/CEB+mJxlwk67t9KG6Hh1JC6PM8ZO5N/PVERLuO
Gk+asCcQo1H1tGn9CCHLyV6HAn2p88OF60Re5DXOyCaV4rLO/tWqI8Q1Gr8sSbjyZr+OhJZgO5mh
q1I8p8NtEpoaNEogx4xJEWvuiFd+2zo9fAm70MBoZcuefyRphJqiuGNdyDlkbnsmZ8swUc8+1PiI
UX4UdlHMUxOeykKnBnCOA1QsE0vMt9LLva5wcqIGQpUNKVAoF8gF61ja9bcppmQrDbkyrjfziQ4D
hnwjtIuUlFWIeifKw98lk3Gqwq+b17YgugL1m5SrWunAX0LEacqQmBirR1JJ460i+8s0UZ+feKvU
iUzr/ZE+aEaniuFu0NvjpaYvswNiPGWzxTbveHwN7niwDKAt7S7hhSVQpYwUoAd9LgOjlAdtu9J7
MVPKlNNQi9yVqKzrLxSEWFwyvrKlUolpBJ0bLIi4TRiuiboXlb3R+RqizifqyWNR2SgZeQtnk9z4
gilWBUQXGhN7rcgr1/Njv1SobZ1Wd+jwd5dQyhvGua7koFOUOlhGcaF+FLqeSRt0Pn32py1iMqZm
GIP3Jbdj5vvdW0QfhbiU4QBaBdSu9GgEPSvsVdbncENUja2ceUo6rJcWECbbOqqiduYR90AW/L8W
o+APnQcLcFQYcsmyd6ZrmWlQUKErXzcKNw6vjOKRy7fDxe8w0zMtfjd8YxCNbdh+qGN+gesoIoTj
dPLYasPhhkeyHaRCq//RlZ/Oqa6u8ekguQEdjjqRNnizN7NEGOjGtkEOK+fLLKt+sZ6EV6aMNqvO
dlTbqXCOt9YYM5fsi1j/0aCSBdq+734xEuk9gCNd/Cs323Dj3yGq+YF2zKH/Q2pN5HG3GQ5m0lVB
8iA/A+/43etLerZkLUyyCb53yyC/zl9FoCKjLJNqaV9XBggb+5kbBvwlhFEMZUh/uCfd0N/ne2eW
Y6cPCUMRJwdSXBgUPHIeGjVn8P1lP620INI1ojZBoPjLwy5Y8iqnTOjOZ7Z/eo8Y6i7t9EqFtbn6
g4OYZ2YEPP/wkH+il/3leq/oALWnafoPDFq+ssruJL/L0q4AoG6B9cgaNi7y6XHQzo4fGCrcURd/
6N8gtd1bEBy0RtKw2mrdGlwK9FSBIQ/ItBWV1s3U3o/1ob1bVxo6eGvy7Y/U3yCt2BsWFjaa4wEh
pS4cJdLzinSbDa/MRN5YVRS6wGFbUiEv4nA1pSpxHAXv6v3UEuXxUF7O+4lgDi3jts/S9f2NDEGk
Ik+h0o+p/6r56PXkKt0yGaeOY97/8zoRBUU4PRB3ZOTFko5iRxAAh1m/vF5F34jrfaYIg3ouHdRr
TwJaJG/So6xGNGUdFawF4rZoC6AlDaTHBmOx08n/dqu+uGacV/0mjT3ZHixpzk6ZRjNIj/nL1Rjh
sh1io+VP0j1+qBYRe1vFS7qUnddWUXCEQWEWEUU1nDNEhN0WpaDT+Gtk0kR5INGFX9hVTf2toOqK
U9W/KKWiYpBo/LAtkoXYP1FFDZSzxmoYo/hSGtAxPSQKKOX18gTImiwr9Q+ycxMb1QpkeBnVN05B
eZNI5HJMOcI17jNE24Xv8obgRO8SwHx0r0wlrJLHLmiv5fzUtuTIwSFPYO4lxoXY/Em0LAjgiUWG
gm4hG9pRfHvbq28OzSpw9cCV+iU7PX8W0+VXbXoZ7D/0+Nd5IoJl1gwrT7QFA48yVgL9zxXe/Ezt
M5RtZ8PrtkdumeeMHXTB+lo38hxXlYDmEIKMbtaC6DFsB/Ev7vUxdBa2Wjw3TwehTNjPUua3/+Qv
0LJCCEsgvxEhgl0FxBkycmy6WGOxif8OgQQdh0RJ6eIGKy7KaAQngn2ttnBYHvL6Ys+OTu61cIWJ
uTXfIowpVgeHOrJPQhtrbTUr1lyHEhQcaDUZ/b3sRFtUIWG/FmVhHHNbtSoXI3deHIUij2ZYV5Ht
8EKXpfSXFzbMJUHumDEQ+myroUVymFwCC5uAJ5g+k9TKUVT+U/Rz28ysuqDRPsZYN24gwXnFoP9k
jxe7Svcpv7+agoqz9bSrklUdZBJM5bqtCKHgGPPNKPsHb7+sMq8qxtIypak0dj9HpNMlQkoSOC8y
S9hZkauVEM1WvoUjCYhDBogkLxkGa8g0vueymCB17akXrXdpj8sDVYAvpVHweAZJWgATWxFlkEG9
cSZvkuLlahoCPu8/YufPM6jT7byu6wmu9wmxDkPJk8PQndZL6F2XqyoW46WEw6NTHWC0AlDxhhgu
m7o5D38ke+yR/dEup2RfmFGLX7d31IG3gzTtvIjsSkG/YMs/8HdQ3IcNPFr7EZeM7/MC6Htj75vR
b3ecoR3czPMkUyvcd4JG1ANMTdY9IP4YLvjJd8Ixl500eueGFNVuj2LuAv5cdu+s4ogdwwo4ymCb
DlYQ77sR1VHmhb68XQw+PxTOLGefsIoc9rlRHnAR0wLKXOKxRIvafGhbAjvDVaYo1KRapICGOPkX
sMWjJA/HGNtY3VK0NgWvyFCjXHtn+37e6YszfHyKFvcbi3Ftm2PNP+53KOKUvuQUy3DUnmeOS+3x
MGxkiDq6lJHt31o7p3wJiUqrxh2C0nwq62cSE6kkyOhzZJQYgzHxkNju7qBPYy/qHy1eY2HruuST
m3qCW9mebpjInVEVZOQTiONg7sd+6j930REU4e7QlNGd9HI/OYi21+N5uVTDsViY724WnnzFEqk1
d92AhM3Ev5FPOV2xkqpYtWl/NSgYTJmxmsWNQw0elvF73eE6LXu51vwxMzeS3Gjj6snPjHy1USFL
Y680lhYIVFzTJIfHvR4ckDa+TeXMym9PScJtWcuoZnyoo8WSKvOTI5ZAJB6uO+R6TOrH01kUDrBZ
PrD7aBT8oxVAneYhI6u5J01gPj+uJiMjUhpvOPFolMreBX0LrQFV2CEHxUKyB9p+PzIGedw4WyRF
XehZ61O7HI4lirB0ivxR+aVC/Zo5F07ei7b7knYAAJ+c5vEv8GJEZzgIkKWVp2zE8qi85o73F+Pk
1242hs9sQak8N5WA4annSynalQ+CG6bswhl1H6HdlK45fYKkupPZvy3Sd7XJuqQLUyRDH/QbMvjM
op8d7aBI46IE95hjapxOfx/s6C6xpj01jSQVpRF08HbFGqjbyZdcgtbAO+eGcKppoCbJi3PLyHky
FYk1laKpdchBCTcW5qHUOAjceEEMnFtGs+oRwdIUlpx47yEeWrYMUr8c4LlAyppodoS1RPIOVhE1
VS4o1NUKqbaUMiBnTZzkwjUyX/Mo5ZdFfRYFPNEjiip6dQ71AkAbPD50AAsMWcE5d2bcP6HELt5h
Xhc1az8w9DXVAtrPDqOcadv8qQpdJHXNr2VHuRtTB07mO1ywfllH3kLpMKFnIH+GTsw99Mi5HSi9
kreN55kX1cT+GGLCE6K/yb1s3Erjmq1gAch+Ji4fR6qUEimkYergAzCLBR5K0jO2X+OLwd27MMIj
Q/ht9ykj5G3SD4VWiwuvzHfkDG2Izr0gn62jQG+Ww9oAjSdcSz82cpEghlCn2oIZ1ajy01flyZw7
KXPgw2b/DjoO4IGRTmIDzZj4nzSWMrVlIRxixYY035O7uukFblcodLs2dpaNVBSpe1Z1vTPvreS1
gL7TRImTFkPEoGZpPkPJUuzDr5sJm6RDe/OuHjlOFksb3U4lImTF4m5PGVdXOyDRmfwUHlexOO27
lAs9qlPXeiWeKU4E6UkthmEYBmUK8b01qpr7kDEmJpxMGrmx5x4bmkNcmQVuM65efMT+fV05LbWy
rWJB2RAV7KRME1ymj/2NTCCU3wK6OzRXiDsF0OFLwA8iuP1i4ja3XwvDE8d6p9tDzVZ0BeoFiJ21
sM4HJo9U2dDiGaM2Es7r9pAw8paHHmNOlKh47UXhMcNRdnwLJnxriqNts9aGXEvImR3+HkbBoaCy
4ok8GbHHZ1lvbPmTNzEgBFam2wgrEEVSiF6EGrNGW5Mfn1zCVNPc3355Td3qyPsMUD3kSz+7Ivj3
LrBLA7CJofwS59QyBKXQjifzHYQ1RMBXxM7N34VeVvjXGJU2e/Qr/y2X131NVxyBpc4pBjUBIRos
PO8TO87k43+dWVFKThWwOdJYrsaZdxrju3v3NIasa5MI5e8BB7TMJ8MlGwXhLIdo8ijRwJUS64K0
gx58ybCagNakv+bNv8+8wXn8xRZQx0TbWEMfWrb424ZUM/f15gMb5nPwKrPD2MUKgKtII8li66i1
5/WIRDupoVaYBQLCnsJ7tt0ELT7qtXQ3ifwqP5As+6tsOxeXO6r+7UE98gHmesu8Sh+wjyCU0IcH
pJftPI1FeBpKGLE8bhv/7/O4BGRMtZES+DFFrgFczXKSHqFaWXsSVwEN6l5QL5Enl04DOnLsxS7c
v37dySZRXiZoshGkf+1AxCHQ25oRTzu3gzwUH8tWQwdk4z/j+ktc6v63W9EAGck6mtLepXp7SI4r
chMI1wnAzMoXtDXAJFm6kooPWwhfRy+vuooIALfa0t6uj0Si9lMSMTgiEqOXkEusPqGjv/aCahzv
K4ylk/5OfAQQo0f21p7usHjs7ev0vhOwXW5C7q0Lryga8zVrAFJ5RN9DrJD5XYbGsShPoGW5LPFE
NVsi+5QEGByO6ucOZePO0eoM2iICnmq+0taZlEPVdK0fInW1q4twEI7clG4s3Mm07vgO+PdBopRi
8emKi6InRHUvLJw33M4IiFjH+Oc2ZXZFxJKE6vY/XB4/EiwkcZ0U0ZOTDQmHqQafus5/eSoXa/1M
LwK20z+BloAIesICdMCtERhlHlMjy+Crrn8FycqwZZKkNIGeukqNGjUKxMFTL+4IZlliGYyNXzxT
OVNN1OzlgavK5DCweogon12Qfpt3R7FGbbmrjG9NYmewC06kIc/aO42CRvYdG8XTdQqBuI/7dY7Q
TYeYj4CqjzbxmAwp27HJO359h7RwuIQnsv/zeBkLdfwbsQr3yKQWLp9ZdwXAxWbuzfdBxarsdtpX
AX8IB83apu24Uwpe4iTN+WthZOpHQ1/iHLBlrF80V+4OIBuloSjfDrVUVEbs2FfvJ3D5aYcjl6eo
bng8kPhcBCDDM+RguSQ8mrfnC4FirdmE282jkSub9QKTFPY60Q7tH9QjB4u9j4Uzz+Q/psdKEZcb
A6EG+uJYW/24g9iNXb+1VNseQnHpA6EMGU7wMsaMIkk4VA9v8gHUpdrOn9K3zsPwhEyITRO9L/Ld
vU02tpXCw7XD56vXmxKmr4GsLGs4/XVav2J0nAYohXk0hh3L150NCdD69HuCeZhEnRka+okg7Qzm
eRrZn6Ly76lpxUptgggMeOdtFlNUaHDpMzI+07RGL+tIaG3gx0+0H/37Y5zdMGRWnIbGyr3a3vRE
LU2BtFlU8aO7cz0yBYY41Zdc/EublvhWCRfUfOj3V3EozEjQP5FeCeDTgF2HTIrmKEM0wmCjw8k7
1YMhU2fb8Yg3WYEAWsJQxv63scFW67ftrErBIkzEvOZmL8/H1qTNu+dmxr+IcyjtpNfBoT//+PfU
CP13gxjm7rBs8CUZ5xNkHUd+KlWA3QHtK4k9i1YPj2bdpzdUFneOp8uMQk5ggRCbtx8euga0yp8b
7E0TpSFa+J+PjO1MRPyxH+yAk97OmoVBm639KUmYOn2p2UWwXYYRy21TNhnePo4rflI5SFLs9tWm
Qsb4Sdq5g3uC7CUpn5KP7vqicOLtuF86rhucYwLLz0wsniaRdxlWhT4UAc4UaVQTylaiwimbvymj
/CPsH8xr2mAE0L3Gc2UhsjQBLzYWjcFjvpv2iXHeJI4adql/lllwPdSZxoB2SaDw9CGXeJMukKkX
8hg+TMWf+/zkPrscd5aUZXzZ7pPHzmkaBjRVObs77jhAN2BoAnySD8OZ3H/4EprvR/LsnSfOfy2G
Ab8SYbc7vJrYe9vb8Tm/0rC30h443ZzSZVx/6nagiukm4vjYHI3FJq0Y7YI2yq9eyexc0yH8bLyq
3syLLGzHCCcoZaSYOk9wUYjObR5SQdQQnUTcbxiXZUkV4ASUYNmF6hrPkTZubb1pDejfHjfY6EXo
pYlkWw6a0P3l3b5vNh5VLlWL8SDN7q8i3cnAvLAWLAEgm+/8WXTP+pU93m8YlGC5j0GzPqrHoMpb
3O55iYKIq4ifHKmNOzsNHVZsyppfZkaICKX8sS3lCtSahhEAjRoTM+YWPs18S020OpDUsLs78A2i
NWZo0Ap1+Svese4RV8ox2vWN38Hft38xkcI70iA1esBlPhmYCiSq/Bb12TovEqCGbOJ565U10YYJ
P+tojmth/FtzAx6Slf+qDnjHPg29yywl2iXJ8yJ4e2nl7rdgkkahJDUPNwiIKMRwtCWLgETcXmmC
UuaVm/jds0CbUf25ws0toJRNh89yA+fhry1gDe14p2DflNj1+AwlxgBAKO5F5tQODZdPO7VxOj3t
8Eqm70SrmJsKKPdwfWl1Bdh2VhlfdRjGQWX1O4nrf/+uhWizzw3OSfjzhVVM0BcGbfAyYM+dpm84
6VpZTKssuIDuQFjUewpZKk1sh5mlGVnSSfYIHNDQgDLxG1CNy9ZF4cGOQLZwTxEuc5gcF6vBEMeE
KqAD+1LZZN7fsqrnxzuUS+8IWnYzw3Ozwv5MlefK+cAQCN92dakQGlKnPglsqv+tn5f/OofrhEd9
xQw83RsuDvMknY+9EaRLjLWdAmUE5dNzbt16oInkwkORJnFY7TJdR93GV6eToQqrFb8Is5ZF0V6q
17n7I7wUYUgYH12GX9+17cWaAhIp5gsQ2y0gTStgyryDiPlsEU4EI8UdR3Vc0NusIlWExs221eLJ
5xYn2oGXf3JfcQDPgu24NhXq9wfL03H/g0Jt4cfJoqyAMCcw0S2akGJWZt2ChEO0GL+K1gwOcms/
I8Q9QaYaxIJAzTdidw6JpjXIduK9MNY+IcdtlfpT/yOzxp7nWdJoljVfL5zifj0mbncCepgB0pwb
DNKcyJvz60GRUBzh1kKR3sKbxG8oiOdCMv+qzkKu2OIAIxO595n3623WBr5MSZRMIbSOtD9c2wDt
aiX9Zk3XtlrU0Vy9bdZhkta637RLxI3n6z5YZYtfsoIPwxJB3gXJjd60bwzfx1WVupwIhlnCyrmv
mNg6iIvQ9dcKSOWJV5cvk5FbNHyPQsL3NiCLic0q9pHRf5P5CGK7JtEg0k+0Wso0fulcQBXCPBrR
8gJG3ssFwx/ga4d926AjVfKBEYGnGU/kmSCzq3ASzqOhDGyccRuDiD0Bbe4PakHBiSo5R6O2KrZO
NDQdr+SkVtT7vLRx//ACJoCaoCFbLmhdhAgLQjAiloHstDHwelEM+PDYdG/0XREz1oS7XaXfXGgL
ZuKX8RLA30pa7iGdiQ+iX7oFR5MfSmPsA79y0JrRK4u31bNnMJARXXRswg+v0OmaTXY8Jr679ohy
9KOxGqhXAMa2O+zimlg2w1EGLimGYaTOpGfO0U87Qn0iYogs+K9VGDjJdRbwXY3FKX0woPq0ZKOP
my/uWAPcn9r8h1np+4DbW0V+N1Q0xg+dyf1uj3rhmz7ZsZv5g22E1p+D8wkZAPwMMJA+DvaU8WTO
IeE5sBziZSl+1U9Pb8DZNxXU2twZt8uvwWwVk2aWcTYfNUfV0k0XeGvmlWg2ncWinxJpwtfd401s
nbvi+0579nCdg1VyoPImyg2l+Z9nrx1Q9RL04CQHmtiMzHJrRcItJ2Fs9+yt6mRnxbDDMkYJj6NL
x7f/JaijbZ1btCbmRWY3O8ezR1uy8b/yr727PeHy7Ti2zmNjeabZSwioHvlnlDSrAMcEwhRTDJi0
pyyKG3omfC+o6J6QQH+MIUU2j/hIoOthNGCKsmdV1tCef8YBi8Tq+a1t7vcrfe/+FqRg/+g8V4GQ
qR8wFiUFkrA3c50820x8byEjqydhwgc2f3PbZNIZOdcbToqRnjgzuwnqIpPfAEXZent0ZQEKyz8S
Gjmrj+q/4TyCwyC51sWKsniS2JC/MjQh4Ic1knvp8nGAPu5rNjtP2T1DUZcqIowDyityxs5j2MiR
lba2L79JCOy2L2fiBEdr8Fhjs8+Y2EQoN8rK6LBQVOjyTyG1eWlE4rdVoyjN13MRDcrO3xB40trX
HzDMylF2xnYNiRD5NvT9Uwe8sQwZAzAvdWhgUwBbrPeM0peDJFlUA9nrzpwnLAZuiiz2E7FWYEo7
uycCzu+ZZGPAWFOL36wk98CmtHyimMOhX6tR502hpcVCwuegu5sxjEu++YnDxGCFrNP220zoCxkT
rF+CcAtS46gBS7yCvH/730BYWh/x6CGxpnKConCMxzzdBzDtzQSxljK970UsbYpmqII4NvEHfPHN
XLyzTRfrlgOwkznNPiMKnecng/1SkRw5ZsLBSwTI+DXPbo4U4Kb0uzPDFbJZlWiDw00WlPp1iB/0
Sgpds5v9WNtTifgPt5Ot2Rb77XpWAzfxnQOZM2+9Ha3IW0RqEWhmQigKcAPIsYIJ9kllUfMRPfJb
KnQbO9zd5JezaJxDUnKRw8pg616x1cTE4EglpDIPamzZPIOPNNHCADlhP1h/Y/alMEZdmAppUwIV
ArTqPjl6x7xpUZhHUBGjXhOdCxrlX2fojKQq6kI8ichMZ9lS4/czKF2i9pSQv+5VEcwq1LwFxFQf
ISa7sf7outoFiwLM3cN+vWF1RGW47CWAsK2mgGgjKXrr1RE4KRqyp8G+wG8K4iMAi+6z1Y9OOsiA
j3MR2DBiCIo0KNxKAM4J6sTAquCa5PFFMEyycxQzswIJxvKJ3UuGpHRI13P0nrnZPeYkza/Xr4gd
m4D2S6dc457uAN2kVdmD4X3ZKtjocs+6shAX6Fbo/PNxRpJMFkK8IxFyUMIBBCRCAmAga4Wddy+h
LQDmSf6VJWgz501xu3iddpX/ej596sF/AF5yKm5nd8gR04m2AmldWVHN0oSfp/8WvWDweP6+VgB4
KS8ZplB4bdwVeQFFcDFazVrzwyJ8y9azmHeg8e9u6eI86i1bxRbtf3vhM3Ed1MA1AndonaBaBPhK
pri4H1ZJqkKUONaFxR5P+69R4DEWdTpLGEG051QazwR/oHFEf2kuyiMAXez77X0owqtXjLQ8iYxr
nNvIxLnxxaYzmKxosQdyp5Aevc+G97XOazGVkKooeByiNqJfojAfR5g0mNac/XOTzSbfAtMAG8OV
hzNYDGFRWFtRC1Lrdy+5fPbOs/fiC2og4M5YOoQx9LbQ5JeGqKb554YGO5Y9HKnM4ff3f4KprCAp
BRYRXBf2ATxkWhxZnAXC76TbMz9Z9dO+vfcHNTSR8vJq8npfjyhkjxxYFdpGTj80Cf9a7iRQdeq5
OwoERDpIbi8qv+VCF6yaDooUenH+OEZQAX1pnRWCjzzOPKbXv8Sb8gdKSXvqjTUhqB1aT/IlwW2K
FcTSMewmSdnQIqeH2JNUba5tuOt6upeCvVk92bmiMeiTAk2CvnpPYWQJyp27ylXMkBXb01kIWhcW
gJXkDOJTt7yLdIIENzH+XbI7wqTlrnzBB4tiOUUszwmKnhsJeHLb3zXpp0Utawc3G0OyuzI0XkQ8
LTnRZ0M6u3WK3mMmuNRgf6bZpF/gquAWlLJ0ZEs1M6LtSs2OY9NZQEuglENr97pmuaRDzAt/655r
tT2ZTo4uEbonGUhfFAkMQGIx/AZ7EXoSIw7vn5roVCj4uVH6tdEanRNaxJLc9TkWsxnhpwlt5KWb
L23DVqKHK6AYTc6t00Z7kQURYDr2DRzX5ZfY/OkAuM8J4RNeBwE0VhtuK4lLhnqQ++fkT2hLesB3
Xu2wJpIEab9AUazFgpblUNyk4TXHilEedQQPqumq+5+cJGV4PHMn4hNd20ia7Jrkz7FmtKcl5tfl
f134GzCMeYhw9mmzKSFWUfkLQfT3j8LTsNo2xPEv4AUPaf8h4/8JHcNFzOYjoWd5YQXD8Z9wg8G+
BtszS31H3KVOpja7BBgKA6maFAUeeiLzE+2okAosaIN6+2GsGXAqu4b3rwlXN8TtPFH6UFv2iRCv
+uA78WKDZEXhNxw8Ao5ACyO7XlQkGXy4xbN6ERQqe7zbeqlULDtibL0frD3WzEQqoZ6xALb4cEuc
uIJMLY8NAda9Zl5DwebW3EU5Zonx5nlRFb8ib5aMI72uZoM+yAAG9m4IXUABqhqiDHMPEquUP5ON
yNIRflihzk2jUQIA6LDvDQ6ba7kpi52kkl/CzWHeuV11FX5gBAzi/EauquHDbdHWxUbI1UTiXUiq
J9UQAICtxGw9G0wOLZeoUDpfDi5o7WXdhEBj30WjrX8ZbHa3rmQ03BszDBQprSuhaa23e2t+MNdZ
gQ1ituJ9pfAQmd5oV6T03LjEXhx6wmgfO/wiiEppgAQ+UCxQ1YqsSbo41i+I3hv4RgloyxZ0poEY
tueiL0EhYklpxf6/91525t2xBkMe1XQpsu1gyqkAgwHRT+oHisxmDVJvu8RUHgOlGk2zTC9kIIwd
M3WT+03piT4nwNhRKdDdhfBQVUw1zXeV15r2LxvOA6TNL7i06+vKdqZShKKnAaqb9ZRHI9ci80GE
sglxy8LtCLHOsSq5kUaZSUph6xHA4wwqm/AbYxuGehPpwdVFdBQI+4ZwIOjXAYDr/WVxBt3WK+hG
4PJ0/G5dZm483hNvti5ZPa5ds1jVHjIbGFGkNazo/j6EiS53m7TDz31W9V0heN0ADm8yQpQvGofH
UDvTvFROuqCc8vi7bEQDjPdrIiSm/rRP89spQthf3t/IFmapLy0kwiGyYL4m/flJgjl4S1nKflCd
djmt9eyKFXJiFkxqK5V0kGv4tEuknMbktbjggZYrx40Tce9kd1EKdT0Rk/5mkzEzf3NpRVwa/6KQ
O/IPh1bIQ2Z8xXW5KnlxSHpxmupsINaRus/v2J2PCxTjzo3Prjof+/pRuKZUGGoeagKw6bvmDFdG
vRBKC0zekx88dpyU82/5L4oqYC+rE/SyAmVBEnQO+j9cHHUfrkiGMwof4COZcOL/570UyLVDgX1Y
ZaitmKA4XR6SPFFz+88dXsQfUCfNGP0PykCD6K2CHytgAX1i/U+V+bLQTj5ac7QYnG8yKsZkR89D
3Oj3iGbGwAVj4EC11fe5BLWXlWuvG2SP9THcP8In8eAo2LzanfPz1IuA0ckvrh5Znz4Igsl5I2oP
t+pGLELWxVn3Auua45P/Q/L086IJcmGjmq5GVbv4RM/CchI6IZnUA4E/9lLrPuyQPBTRE3YyUwM5
MXAKduwPGIquR1nBT9Ggaxhdhb5RELS1cAZ886IaD8ykXjcV0LOqUtS4invnsHsQLURrc0O8wcf8
eWXTtDxUA2G7mVNPeG3xf628MBEzgK9fuuc5OweB7t04P3o/EcZq27cumpw/t3EeCDDlbylXiwHF
+PrL+lcXAIS0IVGH/iQrsq957rHgOBAbupMuyng6fOwKJIW7hkSSpv8papMi0qjtMz8GrHSXmZ5x
JlBEM+n/ifdKVuWwtHwqGavSHcpgepK1//9zG/8oB8HX4qzKDfkdtTN3JQgEooClnEZt7yQoP/mg
P8mtQKyzexBP2V4kt7lqNCmJAsRwLwho8eH4QttbSs4mWqqs2u7TyEKHeeAwH2OXGsRxnIt0aNr2
cFdvm6CnVrL79DwJeJcN3aqZ7TUgIbvJGi5OvA4jk1uwA4KewjtkgM2/enn2BqgPej4s5//rf//I
andiXDnrkI8t4xjCyUCmezZLO3fRANJ1idloqyZk5i3gM2xf+olRvTrMzH5q/s3Zjtj/CK5SuuQ2
WPJoUAHQA7PIDtTRk37zP9JJT5Dr+kOxV5rDPPB/GZJq9TGiMu0VwdEYVPtxFOodyEYNhQrzcLqz
ZGHzAtxkxDLka5CRwfCQ0KlNFsvQIgDLBJ4g5wYtSrsytiWFG0DDwc+ZARSqBzwPAeIAEPYJxvdA
M7IpYm1xg65vXXwzo5Br73xEb+vibEj9rtOAztwU5KUW165BTA8houo2nvKwumkoxerP7r+jlHkG
n6m1ophp+AlXWV/rrm7V2X+iLmEAPbFjUAtQpTc8pg32wK4uu9TEaB+nGoUzy38sTypMoH4QdUMZ
pQe564+ylpSVXKnpVVjqJbw55wKBKYrWsVy6SftCGgKtw3CIRlirpG/EFOarC4RJYzkAgYEwwTmp
ydbyc+21kwN83uBfaFBr3T9c9HGHPoKCvRPkOsaokJIIIQOF/nI+IKnsbslK+mwvVc/JKIcBUobY
+qKGYZ8ZkY+Sjkg8+viC+kxHBeGbaXHKzTcnt2wL1uyfOqwcBoODCMMvDRDWDcvoNb+4bTWwL01q
jctRbU1KNURokPZebBlU8M/WbLZnkknWrizWeuEZlG7OXlRZefTZMORH/7zra63VCqcywYYM74Wj
b3p9eP1IqI6Y5EUNnzRnCXEAxrrYoyweKax7s9tGz9Ej29WHNA8fHt1dpY7ECzTUVX0v/ljKGSNF
8FrlpQUY1H3IFJFjVnrFNCUEN7zCsEOCpLq/h72rIdBzgx86sbiq6IptdZJwpQKhmTwAOD741RER
I5jnjJLv0ktv4oKlZX5YPryaa6ZrqIWAMrZvhoFPPsBpbFOLDpMnfuJedpgvsJSxPfAxwQ339sGb
ml0tqf/FeIzC4Pk0ykfYWNAAIdXCguN0/8ln/LutPN7/bqO65C7z3MigqTaAoMGJchnKms0DYSZn
4rPpSyVPuZlmGnyRepT+ksBcDd7wmmHqpXuIShok8/BENKb6aQ2KOyxtYvtAMM6C+FNVh0ME49+h
oab5QSuammOKqsj42VcvQgQR/2A9E+2OZMRxeatyN11EbUNsrUfkvIPonNsNuA3w4d6oq5SNnBXf
YTz8z59muAoa/KQndj+7lXkpzZ0wgS534hDAZ1U+XzQi8ZjT8gPV+yke281JcXGF2YWvmpmlI1n1
Ho98HHNgpWf+LkURjtJxOVlSxoiL0p3MTXER8Q+ALk+W8NjRqpoRYYsixNHMgkzFYsVbCPjLF9IY
J6Znil7A2T3XmYkEDrw37rvyRQwnq4f/F89twgGZsstbFParB+fEdigRhpjcwI51aYBMWdzAvRoW
C0KncRiEy3gzsrvS5zQmrgKCLVGXLTQFVLTc+izKTcR2xXw+O1DoB9cjdzgySdLEwoBuZxXbkR1G
+pzMibmrNKp2Yh0EtLUbBZX0CKjD8HpN39Yq0R/YX05AKXugBRj/4tZaxwS39JJRolWbMLkeZN9a
I34SkbF7jCLLiyoHZcUX6v5ll2a2j5JIexGE16MgaVQKlWj7JfvgVRSj8t7xa4IbyTkGIYoBYyj1
pArhju0KLS1IAJkN5mVWIgwHngxhadzhmQ7tzImTXkIxQUUunSMDASDbUuXbOgS59RwW8oFTpV/7
qw+iFyycpSBE8A+hlRylylweWJIcZLbr2V3/tC0CSGRPtGkqZNzU5NEXvfxjSbdWmvaL+AGCnGZQ
GUr10wx7BD+j72/bjh5c+idQAwcvc5+8466ErDrGKV0hzCYDiLl0rdI4bhSktCN18OCxicOFBFIU
ZchELDpf1u6iPBwBXaSVjaXMt3AriG0+XlAEx9mkYzRZpUXrPf7fDrdXvClVmMhEo2dk0fAq2o8o
wYtpFCVsvOtrAuk99doYR4t/A0oIkx+BJ7vJJSVd7C1mJvqCqL5MOUKUm1vOPQtEv1a/iznpgjkR
5yWHHG7kI8/jpGyZiNZu8hGNDmoXmNmL31srL7bU0ly2mWvSSgAEbQLpbxLAdXETIpxvt4klhBTE
RNyASc4apsYoPE+JS15ZfS3u/NgQRl/bmoi/U4dcuBJ9Vnd70sRMMwvQm3EQ++3SVGeMpg+qgbaT
tw7Tb8d+vf2tuKA1VIbI+uYLmg8bFUFSacR10rzTi4udPAQVxPbq7oWreyERQog5okZL+yO8jPPq
BXiBVozwhYUyW0LDKSU903LGs5EOB+EkbhCP2uKngmB/2seFGjfnqSiZ1p63FhFzOq81DKn8zkUI
bXbi761xsIdr4Jww9kViD1r2HV0z+qDdKphHkZkvZpk4ttKjXw+Gs4y9pk/XnDjmSEpxkUyBkHUl
oZioyLMGKDzjM90nhwr/DpRjxqcL2xSexxhZsMs5KC6TLi/m+T5NlEZVTtTKOAFpmPKuKIqc16Vn
GV45tcl/ooEPWgJj0Wg+tBJwkJeHyM/imnA5TxFi8MSWBGCVlHR8f2iwhaYHDt9u2KkTdWS3oKW3
2G/m9TFvPT6E1tzXnl4TExqTSWTEGqTWFTP8n//jgr4T/a0/BOyIU6DVQ8WbcSuJtPrqrdQpRis9
RdLsVT+IRWlrwL2bZjbImLZru032ala0MfcjPyyLBeaeWqMhqLwPc0mB6MjZdljZRuR4Cd25B+71
msNRJPwyMnqTSYo0ZmdN6tF9/UiogkBo7oe26CDY7eHj/c/JFVT+DQ9YO0MfXJ9mDAyyQybLEkoT
wFzQixrg8vEU/JMNsGwYxbqjj9Nd9xru1mLW+216eLFgmgO6RPl17bYnhi4RrR2xNj0VMljllaZy
gAWAyst+xMpOU9pGQwJstw7c5aPVnGmpq/AofDDAPNm/y7gvKs4MLXoUOJJqgoMLkV0wFHT82n81
yiDbt59gjpJhWPBf2jy/Z4ofN6RZoyTgE0qCjDSWSpf/CSl4Stddn8H4zvgjrt1NTnTVpmY6+E6W
zdtu1yNMhGm9U0ylokDcZoQoRRpwAs03aCfm7Z+B1fwezJOaWHRbZkJ8CeUBDDRGxXAQCtjAE4tE
nNX+05R1srMxaRawSDyCfGBBYyrzN1fB44FFz5s3HHpLl1Ozfw48gLN5ai53EWE5nF04DeTRcLwd
uo0lEAbzf/nXB5/JmG0RBQN5brBxLC2Z3s4CYPgRmErdOWUOKlKFyxNoL1QGtyrCidRzospakQDK
BCIjbjLOLlDvngAMw3ODcLl2VcC5NtN+DY5hh1U6aSep/KjMTHMQ717D74ecVDs6L/ddoAxIIKd0
LkpnybZuRtt5566gc6on6lpS9xSeuAqwJci1FvDO2QOEFO+c6DNl7Q9ixFOwHf1eOwyXxEbVst1e
zC9M67J9JSV+Iga6y49JKD7JiZjglzSeYW854hrAxXv69znNj/mHANY2q/+wtkucE7/Wc6YMomuh
fph46Q5F/TlZgJy1s9zGGGwKDyurPycUei2ra5lW3bkPd/U1DZKZjXwMqlVhLW1g2RDEiz+VA9rN
3JLbWi9ZKcpY0Q2zQ4dhSxMjMR2kTfgE/sZI5qlgg+E59Q3ROWZyhiHb6bi91dWScvbFSbOGdw4k
IwFRLIZulOEuBvx2xN8mHtLHAAeyhzvcPjknUyuWhVLWziwFzRSMvgpbeapJ03z5lFaw79RG/T7V
BEILmzTLYfxDklNBBbpyk4TIftlKOnxCLJEsDMMuSqfFx/WDSP34a6vhT0KkmFSFh+BfLmM40xSE
y8Kj1HKmCEVf9Sf9ycIgiQCy30HhhJWPiGAdtoUeG9YMiXvrlMMW5g8URc3Pr2qTG6X4PXvitiBj
mJ/83Pw8uUfQnG0Tm3l80aduwPEwYBHkkgQM7aTYTHUOLyyU4A5asw9OF7y2sX9udDVS/z0lBERV
LfXYaDVHqYZMyReU8E96XWDe3oAlGMOaPHe56gOt92BG5qodGVcpjr1oXqDq6Fv0q/vRa1VgfIUp
SjFJn0BvBVrjNq5EJ8dJ92Lf+X1zoEi3yLnKB/8OAcHpds61YyO4GgtHnLy+YopY2meQgqKrgKHg
QHUqoHnIyo6jDYvq6F7G4ovtSRImAcL09/iuDV8lYT2JnfUvBLMmoqoRUo9FWiQBKt+IbkknfKBp
i0k7U2fMG4sGp0Is13rU0sFN7JmY13ntBgODmv7Hh1lK5WpZdBlPTcWBEzoJ2BO0vSkhOgXJSwCt
C+Id19en373LRvbTSuiYU7rL1tLSqdW76YhoGOFGUwNhQOibQRtgkKI/zoe4/dSCCFBzy0Ib+c5G
ZH+oNLQc+XhxMaWXrVRKq1M33ER1fSvYMsqUISBANuPaNqmbXhn5hdiKOoJ/tnL8PkG9n2rWHBNQ
QnVbljRQn9bubY0N5k/Rn0JLx4DBveqKRDYwy1heYNFLOfV5zGNvjhAcg+jLTcbq/CJM4OTVegUF
nw51S2qI2yQKr8WRECip/WRG8NI49mp3+KqqVYU8pL6y/cyp2lvkKjv0smXKY5+yTcQeHJiyk0Yx
lmAafFKqFYNp80QeDjh7simBo5DJiSpKiAsTyydWzyTKUvqUt2da5gxY5TjE1WrBiLk2Nq+tCE+J
hhziSu62k8AYhgREGNMuWFpLev3f7tGjb9iX4y0gEiDOVYb6r+idq9P3Noc5b+ge60FdPogUZdL3
Bkzxx0t79O1eRxls7lU+uIaxJKjdoNSMwob72drSGRSC7mA/TlWr/wEylole13az9SXqKEAO+x2L
eW1n+PwgPhkDYyHuZvmRJZQyG48rJ1puZ2swMwE56tgKNdD+OTZ8Gk/+wd7v+4Qi9xAUhK1pq1UB
rcZ4ZvvjP54TELZI0FGfcpZPq2M7lmWE9HR5Pl/Oyy+Sm5NN3oPSe/rJ0kas5Efa0MHZVEeDWGOZ
wKm32FNRTNrWRtDcpQnM8mFr3cpaEkQkalw8qSFjR27tvh2ISmApca7NjqlvZ4wRvmxTdO/NhixK
kVWv/7H8AiARXERXpQRfpixBco0P8TpDad88OeCd/Zt9sGEsMISpJbERHv4yp1IVcm+y0sxgF75n
fnpKmRTjlnCbc/1s9v/AmZv70OhYqh9bWpGeBFwfRyZcw2x2fKj/Uo1eNp83OfLOF93Jf/O38ZiC
0bITDBynlWp4GWNqU0QekUCRsWcFZm7+Ark4DnnSH7IpSzNBj7TEliMq26TSz/OrraFdTlL/XP++
fkVdSW0w4tFYdLuzeB0EGLvrE/j8Wfv+kwKnPJt27xKVZBaFrhwXyoE4mQ+8kmb6wM7T3rWY9rDy
1QC6zesEzanpx3imAi/H7A5vFXJS4k3jsXQ60yDb6EcpzpJ1pOeaEBRqC4HZq6jZecCQX/7BGYun
JcrZ0XOfbQJJeFmBjGBO8DBrkKqKf6Hr1nOuY8gZAy86vBgErC3bNw6zjjg+RV7Qsj6wNHTxMGSZ
LlEumb+YdsdPuK3GltkQCftuWFd1M5k+sGuS3UqGsizRv0hLuNPObyiRwPLjrdVzA10vjRi8Id6J
oxzPdR0oEp/9ceNsvg3xPieIEpx5OtxTZ+wqF3RzHNYOyIn+QJ0VVukeSuMQVS5nwCPxkLW0a6P1
j7ToIZb2tUO5DVyrNg6EIeDtvlUOzG8Vkzc24DshqNi3cwSLyM7EOhhDlid9EQSGputUN2NRMEI0
6Ctqv+deHBgKJW6dO0YvVd27/0eCEh2ISjZEkRR+nqZk2LJaEKgoS1vGV3H9iIFtJ/A+YLfu8X38
ExCz55AWYPQ3nwVPXuTcdwPuqgVl5GU0wzp5bmSWalUo2kEx2oeskOCxUGk3RYWiLb3QUjF2zPJO
HLtHd5tgnN85EPHieXN7ZOeMmICLpf588eqp3V0WWc2wLX4ksBMaqbvfESOLrkyWtxUXQltU5YfG
rkNK54TbJSrocpA4kk7g7hK8O6YBn24TDI5xwDZ/pqZshNRfddvXE3H3BnQhRRVr8abGQBXWYp22
1C47SKVJIcw4NYiK4P2EswIzl/V9eMTdQxGTCS6nNka1DpnoxMmzSuWrkh6YvVOa9FNYq8D0cX4P
fMUYsrb4jPrysYlRuA67xGu4KZowxUSB5KV9TNxnACUjb+F3AN9+xPOj6twMsVCjNn34swzXVqeF
QrfQfWZo4kAAeUPFsDNKs01Vqyna4iuhgSJp5+6xtNWiqWx9NCjOCc6l4AHS1rOk2dgBXOrgchAz
xPUKWzXS5nWEVnNQdxuym8niQi5GvTLnR9DBbk2rrk3O6We0ZiuBUufk8+zN4bfMXDcRshCy6mJt
V/+CoRCltL55zAciP9I74XgPEfyF+mYCKw7yWTpWpPNKX3zdeQ5MxNKeKS3Tj9SV8xe46fk4ne/6
XOMLTHTzAWkZ2PNuoYoUkfjP3EEFEWKY29S/Ilhp9NM68aCobo6LAvXRNC5IR5rHqQKekP+agT44
VJON+jUnbFzzLRrcbpQE0p7jEAXe2l8DVH2iQus0PT9mBCikgRCSW90q8cgc7iT0wDTey/gTGCdM
kNAAW9oTvNb0HBY6zZWZydQrbF9naGuyO13M3ustaUA1A1AyO37X0UM0n7OU5a7HyoDBp7LkPHkn
bZ4PXGb2H2luXlRvqc+TURaa0Yy1ieMi6AGwPBTAUpQqFBmtRJjn8V2TJoGAIIOPwUMX57+8ycbz
BeI2oH5O0PhcH3ZLX0/+fa21TpmF5NvrJH0PAtNvrjUpZPOl1RZtmtU0/quXkEJUoSUh/JuXTaqA
TpdOGGUBJjEAn8JhDTTGO+C5TEmCc/Eu+5UnOK42AuaEsyZEkBk9aBc+GlMY+XH7WmM0mGQvsycx
6VabJWF70fEkgBMw26oNGYmzhx/vOUeEdHMQEGWJ+ZcY+GDOLZvD3oZregyDwjJog5mRDRm5urs2
6vzuKqmhLCjpqHk1r3k5GI5v6XE5qjZJTXekG+E3vkSWJuWV7dz14wE04V0VA7ttY8x2FmOmZB1D
ugNDnff+t8JqxCCQsI/OYPZ1xhDdtbF3JjIo8HBIW67gz+gQFSsmZD+JyilQSbUk1RLT7FPmtNMH
mPTJak/tXkXKRQ0RKFVodpzbBSMb+FwwWvwK/vr/jdLuC/C+4dStpGUyCl2A7GtrL42u4ArYMmhK
krlGfdHBeqSBZZSwSFwPZBlhFc6kVmcz3oVF/KVV52S6zJ0kINU2b3iSbhWOZYzwRFrc3C4mUsf9
0N2Y5odRADHdgrYrwb/Cm9omxxEnLq/XFiswT1gvVTtM37os9OzjkgMWuTcXVIwDxrWCpxLtwOvI
+HTj/v6qhiqeaQRpviOnS4adMSoen94zm8tTsqs2RtLJgYiDQhSQ1E6NsyFm8WARCgiB01oZeEKK
Owkgh7ICyv9Jg7XCL1wo9CqlsSEK3LCpeTiOhROektXFKfho7lPF9JyRIpLfjb0AMjzB1PX5Fk9M
1ZQwOSnYoSiMZRaVyHlgTzrdmdLXWV6IJuNOr75zaOS7OPOvIjRl41K88sS7He25zIyV/qcETpwS
U/ufGk1dNFXcsD3oS6cw1azyuEhy1H6PVA3tSMNOAqLhOYW5ZbRhji0dXrcmlAMS21jfjEJf/klL
b06+YXacdD0WwFAzcSGlT7ByRdkwt/iPoR6lvvWKw8mz1MvGL9mTuDzbktv2jFKSQs4o1W/opqX6
6KBoWX8PPWxr76cPIn172lOIQrdzKnnAscM1TpfR3BkLQD1avnPAJ9PGuzMOwZDAR0zAQBqOJEW1
LMUF/A/4mRgWYQEbTq98SzMf76KKvX27npvqvtNt3mYvnOZOKqvybMu/zV/o50tAn/u4edQfdRso
OFhgwRFmcLmR1sSYvuZth/mDGCr2uyxYwB8lCN8IQfSSof/okPypdDA26hhdBdqjxH4M1UWlBSBh
gZLaN5J0x0WzBrAEAfq/ldYiBz1gyfgt411znZP5Vo+uGVaP/QtmNQU/PJ0ssPBsxLTVCJ0PlaNU
YsLvvJo1mKpKhmizeCInrrsCIbC3WQKMljtRakuKkXPUsB+x/ooChQq0Wb3KW0RH98VmYRF0Ue2q
vVHqoyI4Sl/wCI7qmYL71dnLLPkNSiWo4U1SeEBOGWMAXGv1xI2c8jrZ6OULr3t3F7Ci2tjTFhHw
ZN/TxZ6qTskfxn9phtHKBtjvQqriOt22lQBJWP/RCBdZW2ti/2d1HwHtps+uVVgxwhED/EDlfmh8
uoS5Vi87PSsuc559ulJBq9StwgmYzBahKsgryO46gxp9CKs5vGLMV9ReizYSIu21RkRIVj3/g/Hm
I5ztlChiaL3uwIcuiYcaOfuFcraQNKxlaJOkrC5NMGcFDlU0CZ2dMh+DHHmKcNOqH+dw1jqz0KY+
8rRg1ytBq11ARPsmjpIlZwgf2/W4F2GWfUFSJ7id95sNU0EuflwXdukmUmHcPXKP6twER64itJNt
V6CFWs93cM5U2s/OTRc5XMuXXqqnAMp1bk3qeiKvRdyaLpOaW1yMfcwBLFr27YJlbR2rLljStE6R
lj6+7rhS9ZMZrSkz0WFZ4G23kdfEo3we2dF03ZzQNGoz7bN5SYhJeXoT9UqiOdoHG1qga5yeOY52
z9RgwSU5PewqQgla6eUai+fvtLvXnOhjEFBXUdjKZ5DSLquEcXDi/EhHmhGz9RQiIbSEySLRMSHP
fM3eaIceXN+umdop71swshbM/7RHwety2an26GNCYE5lfBS+HmY184Qc8GilPSt4PuHYHKyJe83q
pTrKc9dIr6zL4SxdEkLyjjuiNO5iP91nNgtvz6gwQ/m0ncxFhQ9UHVMRPYZu/pPk7ljRTaDYH2J+
gd4BzFhcwj6FbFfsBETxTh0e6lEWUpvxAi0X826APYcoVSB1nEhLOUROa2o6FIbBrHg2Nw7Kheq5
hs89Skcp4Dv+1MyrovC8TeTxoAbGfM7udfwDQiqd2mnQbNjcdwsR4OZf14sGiDNXHrBe59QCRsUz
4bwZ4FRzg0uRxu2OrRiCNOBUlSlUYAtQ2mfjNjqPL61uNf5frH9NjM2tmNTCuX7BwPtehCjdehxO
NZvIA8MiYoP9IwhEQSXc05BcbQi9zBRxHslZNU1fjckvC/tTa+9Rt53WnF7pFyJWdTeCv/pVBItX
af2nVir33emCridlcL9Ony/r2ydYvHA3f886O67lcE3gP2Uiy9q3h1t7dPPJizSpNCtyryqc3ug9
eh5lFV3YVqd6JGu71QLlqSJvHRcB61nC2VZVVA/MEoqt0Rbplm2eyV32ePkAmUXUxVaYmVzQShXz
bbV1fmB4gRFWrj5G2J0Drg3dKDQ7MWw6hwTF1nl63WvKWu235buh7S+qiMNiNayIO2rrKM63oqg5
wE5GFn3vGf0skdEi1PRhelakbh2ttEBK0ejz57QzD1M3q5ivjVNjotNa/PZzrAZAXtbAfcwLJSGJ
HPvTjSV1Ptr/YgaHhV9ql7vGEeEqbrpYxbJG8AaCv9l16KAcVS/BCY3nfB0BUv4HfPZVFjvOd0R4
Mi961w1Zxg296BCcHBCGMyo4ClK2I0TfmT1zcXaY2ej/XgZJOyK0PqvbsoE/q13RBL2ORbxvFVvj
65onEOF7BWlqyJLsgZVI//IRW+bdSbADFVnwMIJzPfAATpHepUNMV8QkSl20VWtLHkQg54fwuGMl
fltqsEKu8N8KcGsjnDgbvgHTmfL1OciKAh4agr+euotIbLcMy59wHC2ap4smxlBnNgXNRX46fkKi
4HovFLIdmjQzesRfRNaL1MAfCc2DlPP+lUQa0IJDQS6vxIYcRpheXskK73UlR7rMgEai6G1An3wE
vlAyEUuTnExH4nEhmc1Hn0+FK50kkNbYdKDUJmHiI2/rC3gln24z2CApmETfkmWu+FXybqEtnXrp
pStLIYgL/8rtWu7qXYavuolqWT+mFyPjO0RPejk5GhAtQa13yax54zDJAqcAfHkI/d4EM6yhakJQ
h6O1w42WbuYRpj0eBP7+fxxCGzAL8sdj3BEAueNKVCohYMnvTvOROcSAFbgSkEDJ6BEqDs6+LuSO
FewvUFUFqKBrA09TSq2ONjoaBUZV8MGEnH5J0sv/5MWYTZnt6CYMb5pWDLvHhdgjNy8ezlTcIZyf
4x8RlaBNauF30nkq1R1VZe8RDd7p5mBpMoDoV50T6cOKUEbqaJ2sGxsqOu5OumAt3TfkvpAOjvuZ
ThDxUbUGZoOm9iQZUTkPDRs8PQFZLAVY4MBfjcZNGHB2/sbnHCUe+qw5lV/uUtYA4t66ll7E7O4j
Cs4zvytigfpsIdKZDq+RR1nglydUnszTEC0dvSQ8riPJ+AWXN7dZ3edhuIgr8Mv+T4VYeRXEyUSX
VSWUAyLybrRtK7NpzarNifZUWYqFIbpC9CZY1EbThIpPRBsIBTGh+dtC8LD4Mjed547L0gsVQ9kg
aNw+mwEsscyQpWdHfX+/vgbwvwlOx/Tfy1XXO3Wup+YgyzISPB92v0UlOwARcVGQ8ehq1hcdsJy+
jznHbP+SsFeDRowxu70um6iGV7I1EBshwYRkksl28oOJMhNdXfhV9lRCY8CZA+v1GzXUROBdHSBk
DF77ZgnrhXI4Ps6mKfhJmg1YyLoIiykXtM/NHH6A16pVDsK6OzwN+4NuffGvhgSxmxAqTypBc98L
Evat4kbAsk82ormnVQ7T8tJkDRb28URG/DNw9I+KSMp0qkUssWws/RdxukVTThW8VHK7tnk8Xd9D
hCob0Xduof9UCdllsQAv8bb/pcStt4Md/f+mY0yVSqVq0AeWI3tPt/wcEuthGmN7BwJ+klKvhcj1
7kmQFOfN4vK2/xTnPhjRTkRIzjB5uMyvO6iiJuAcXOSrRmguarwInnY4BaSfH/xoTRK/HMQhoXG3
ERGgGNjjZclb8PCJs/bGCU1EAUWIRACbv8ZDC5lyrSOFJcztvNo+Lq2OKgVbn+Iv8j5qY0z83aOv
ZFNajOK1HXLR3aALQiZSnGByfNZdxfA6Jz+Y0immcY9AMfGBTVafrHa2n4hQsNoPZx+U9j20YhQr
d5kOROXu05ScTa/5VBnRr0e6vVL9BnVCnzmRUlZbTmsPHPF6cUPu6cIlXtsPmw0OuTPBV0rqUzLe
OD4fAgzI1iIFmNgzXQVFHfEsm74+K0hBGI2czb7oXULJwzZyezflrcUTbyfBTtr/kUpDgMckQLqN
l0Yw0pjXBBt6NjSlQ9U6QsdJr9sN321eLHcMO9DdNcHwdnVbSgdpmev425cRIXQGSefuS/2fAXOK
Hg32uV2hnQXe7HSoaPvT8AU1TOLHA8P94NnNgPOtrvLHN9mWVDziepXB7JV6eFi0I66kvKEqvMiM
jmdPZWlz18iXiUcB1Kpa/thQpKy/wsYajXEgp3xy34lFeo+naaTDqWPyc8c2XPPew9ulDCJZWJYb
e/CItnNWVrBZIo2II98Sq6u1jOEKL2hjlK5J0SH+aLMmeo5tpuKiP/TYO7Gzeajrgq2VaY2b69wh
JVrBb8aBspAgGCvqqkdgranctl4icFbi4MIKt4uEKQNNaQq/R7rECxcAeGcT5jcIPshiUdzYPLYL
2DhDahVZtCuMfLQXghZY6p9rUDrKX0NzGEcxJ69ULMB+hLEcjeeWh+BsGJucni+Dqh+JGoCc7Ziz
STOO5jmc7MsK650hxYWCGA7pRic5oT6UEoXmSUOUJwC35e/j1FvycGUfBCIDja1w9/vLZXUZvBEj
UaTw3cT8cRAEWs71pgVCCs+6bZu+fCBpB5VXCdYbN4OpIYlt8L7PRbHaqH7EYkWivBdxMJZNZEvO
OZ6I/X9y4NchTlF+NAJjchloxvuZX0mLw6vGaaMm0DC20oD+Ob5DfBgw4kPURIVjxsXar3qSWhA5
prNF/vD5JpUCnIHAKQ7ePbFq9e/Lo17dRp164iP04X36nNg8FKBv20eWPeGX6PWL1PoVRkkt8OCD
r5WVRlcJE8umpjF8ezc7zzJ+UEmFAM9WOMVEjIIBLopj7sp8WBiu4s7dXObcUczTfRFOwvvpGnzv
pyv0n5bLkFaBjyKFjAQPJvVcwVVCpwlGt+bI8MQlhWhbc1wRtzmlZPgQo90yRmjgnHgRHWdu4e25
dWi5bwYx1AsTLNwPXTtjvsB5Gz0C/ztEztA4fng0PdyWw2zu2b0uDQLhnRzcGpAnwniw5OzSo5jb
pZVH2HMwp5bHs4eMabNjzer+0EPBQevsh2kduD06bRpDDljR7qH+9KqRrMc7M3J8TePjVAjWvVFW
uOCCZKD7zuJPBROWcf/QbLcHGbKfF2+qX9uOSKFHiyosnoHeqkVZxfo9OBNDzjAhwPDt0hH7EK5p
FNuM8hhJn72MOTeMZeCfOMAoJyz2PImqRq4u9cXx/ZVyMm3syfVFP+1Exhm02npvntT+hgCvk+gw
0trl4EsEzs6v/0lLHWNqBGBUw8valVu8YOKoOZhoDyl/xAJoO7C13XR8bgqMXK9r8dA1xf3kJT2u
Zy5ZomPadw0ItV4Mr8tN/PyVwC9akCKxbdnx/Vrz4Mnr6Zs+Z1RLtwsnbzFxme7vseZtHlBtt+eK
MkcLP8g297f4VanPbHKmAurvsE55n9dH7R9xUfOI7WdHGjsekhUI76gb9H1eq7XsmBgm8+ueBK27
zfK7Rx1FlSuKRheDfLCQZMwSsU58w+vXQ/GiX5LfisffM+8O/ETa0zGgnBI6VsfrzxKBIxwNYD6j
cP1elYbOz8PexAsyRUZ8rfrFSdrtO21DMknz5+7jNYD+5k2uRhKUcLUohDdLMniPHmbMgsTWQ8HR
qU8LSSRMIjHvitjKdG+jexVpQ0iOL5dTsNPyaZDn7/JGm+MRDUBUCazUAo0rpgjtPcOEwVHlAnTc
xYsMvPAcTiw9KDRXYn/y4EEKitCsP18zSOe6yjdd5/nDkSbR480SjH9cfbg39xTKajTlS/+0acQu
FAQJPOWbJvjE0elwGc/hFcHtvoRU2SmcJiVFgYWOL9oU++a4dE+HGPe2rscCgXFin1msgcm89IRO
Bs3O8U8gYaTHmkyiRikz2NJnLRjp24ecCCA/XuES9WS7J71UXC/InCzYwmXAJlXtrqY1AzjGLpgX
sljUYZLqd+X37Gbc3KJ9CdYvmCftAa4n2gME371Nn5LugJzeJc8nFDVxJApa90r8fbzDA11/F7B/
o0FRi1qzaeGch3nJJ38N5EqRJD4yXSJupH6EY2VKfBbJyxbkn3jSl/KG+LJtl1qFpEpksU5xf+01
9OYfPLpMjsL+JrZvgKHHPbSlCtFx0mPQsuiK2OWNI5JvU4S7x2mtH9IoAj8eMVj+qpSFXYPq2s2L
or9r2cdlVenl45tRVfBfZSy1zN+O9lhIX7RJhPUeyFkDO7zjJM1dN2SmcWrYtKBWpudHkP+KM3oT
awJlFbYX9M8gWQ/lkkYneCBkQiP4tko3fWhhtBI//j+cQ9JZXJs3U9paM8Mx6XanY3/cA8Cy8p3V
bReOW5xrvGgazmMg6Q6tv2vZH6yHkM5zfNTyU9F+Jcq6QhawohsuNxDvSd7oCVUgxyCzhTyTQIum
nX/dUK6HUaoI6G1Pqoj9L+0XLDVSHU8IS9LgMF+Cq9Q4NR9LKyXLiwUfj10zha7XuzIp/QIIw4W/
a+Xw2Z1q8cSeRBLOBYcveOpe+2W8+ovFpSzlQmGpUwdhU8JvT3nUttwO7bX8zAghkxeGRptSREW2
It547KN2ncEBz8whrHLXBoUTgp1HhGRIFnaU1SXR+X602oN5QobUXzCDZFDnxTMvzdwNsie77hJ+
ASSylWrUnYGl+iIAD5c9x0SQQknKRtCQd7KlBUsHw91wCYaY8WTFCFFODCDrm3aJcJxbcWxrk/Cf
g2hRQoM16CT6zmIe9dHK0umVw7YIMkJ2thwmOtplV23FMrBewPngUh/N4dRsAgT1LVCwj4mPE4fl
RgDBJl3tpFYCwalhJ5BIFvkvtXgNS9uPLK8S7W40pzshiGR3TN+bb16XtQpXUVaxXk3Gh8xuyvPD
M9MfHDP/5XoWVDVph/yCbam/nnS2cG10EJOPDAZUNbTDh+TZOL+A+4Qg2ScSbIcZw5TinzrPyFtT
4z4kH2UoGIqb4JFa/nAz8b8JwlLugg5JxrVr7r0F/ZABq9KcXUZ9j94yjS1ZFdR4pEq77lb0nTwl
l5vzMke7wOZzRRu29ZdEqDxjbu+gTIDNoQwewBKaeIIog+6TIszkP/719YodnASUL98naPhvlbtg
lz5/BtyPsn6hmjQejOxxT1bSVG4KAbNE+flDsTr5EkQObLEG/kspqL68gRjXBgYGFCAOwat5NLZB
Ya/6SvV1PhbunhRaS3Ng1LSSdOEUtQ8LWk9L08EodCrrVut20IuMTNyqeh7W9ItcJchLM9u+On6G
PgcveEIaigOF2vM5SueICOUM7m+Q8ehn7hZvE79mK1UVyocmNjqL7w6qULxZr6QoI2loMNPrJBof
EArVSKUMFzc0ZES3SueLtj+0pID+fah+6ryWDRMpcVQxn0hc3EKki+NdWQyW0nY1hn7Bgrs4rhMW
72SB+tfHRnrD+x4WjPh0H9skO2SS9COZnV5oknNXFCIP0IN127opi59WD6yu6IFBCCgNQOcDXVss
t8rUmrENBGSsYjsmgNPv57c2R/4J760/UOOjDQ9AMbJXcA7LwcQ7xid/KgywOghNuw8ZBwxYqmXg
oujn9itOXHebwQRGdc1XfJWAfek83jW2BomPJom7ehXfYcqoImEiwTxyJj7b1UsQekZHCSbNlbrL
OVYRAYdl0WrbHoDsHsZ99IZEF4CP4M2qxyxV6WtMy+QU6WEk6FTGRN6Y7GK3tK6U2E/FZky2exFW
9PIYkH9yG/LvgeoqTRWi4f0PatLK8zKnCLX5OZspJPqPuM+7THJRZTsTGT69/tnhIIk1Au04rz4H
7qs7PFKoWUCG0q6XxvbeEM5LK0wsHOjZ27UhVJPWYdZ9ZbYRYGE/zUTh1CFMGNWjaSXfJsXZkBWB
MwOyY/dhYlk8o33ZBNtnxMwl75VITrvttM2XoZFcGJG6vKMRgBRFD143+cVm5Jub8fj0fEcHWMot
S4PS/A8DVIVVobmBOWX76utS7Vi1Hitx/al9Snc7la0baNNmck9hR8QwAOx1XfBMyGsTirGWL24c
JApR6IXkVsLJRT/9aqs510ybuSatkrmds1wEKgVUVkKL4mqfs5UDjbpEuiBHMl4hjFW+4fVcrpj6
PC1zZTfwrmGS7+/GaQKDkzVUfC40cxZAXThph6mQTIcjRIwD7Rstnpokg1i0/hJpmc1tB+rxY0su
bG5+ti9pQwgdEiUjtrwnwwYbEfEI0+XApg+3zxRhmPRZUzc1e+h0qo+mA50rZ6ML8VZdJF9OpbQq
EspES3bHIY/jR/1CXdADlT7u8oWC4FtPc/x7lgOf8YcmiXvhEn4mgq7gypLbsjDtG4rk/Frsy12F
LuaFqFqxUCChNi7TBpoG31PhQ5VGUTu3Qv9tizispK0LMmjKNnyZRbnlAMkAo1XYS347xNmTcM8Z
Hd1NbF4XNTai9UuI200wvP477RMJ9yGTBEJ4Q1RkVck+TWDtSpGepyoanXYEBnJki8ToBTOKxq0V
Rm43uF2kP6Orl8c1ZxWaIOxmoqDwv20JUnrhwLBVTeusk2nmJpQLBdHWLSWT2lwHxOqDkFKl9XBo
UXaTTz2BZs3GozCdGSxwKAKZBgI6hmjcz0zfVddQyCr/Hyj1LadamPw4ib/TZXhUErM71tn87YDB
nkY4EoDYI9D4tv+7Crqkd8X+U7nk1mA6XCqhiTDMyFztwAttE50pa/J1N4KduVFapW7AqqVb1dH9
PwmWOTaph6ctGE6cqGx1Xah0/ceaUQw5WY/+PeY2Mj2SXDXtDb04pBrVTpC3sYdyVeIj8jNBVgEf
plYbjfeY2ifRRqQWCWNojXPnmBUJRuEQ4b0YY1ihsRk+uC3yn9vNBjzpMVT2bKAoo7+P0m4YWDpl
KWJtCDXho3mpNPhvIBpmAHi+YSlO8BOSOCR2vwf4XuQDtm0ACtL+h8cYvczeXMG8UXHOcIBcdLTJ
2YAOlj723mT7XypAkCFZT4rqcowwJBwiKdnozeeSt84xjryJqPmJaeFoh8m3Um0ntgAgRGvh9jzq
948k4d8NNZv5ohqighKpneGH84kwsYQgTH//q2ep2B5fEBWh4pVBgoihfSBlgrmy8htkysBreoxu
6wI2r/9JwZnyveblsA+qSHcs9QzFJgZr/730lrO2uWfMBfZtKhQazyNG8KiQjAnQsXQySyrl2Q4r
pQxU3I3TaQeWs2bthaIY8l0HqBXFf5L/RAbcZ6zKoMVu7qnfl111fdr8qySBb2//q89ifYaFzsbt
TDU1G7RPCutvoEN+GXVlOKwVetNkvyxVyd2ScuPjHt88+JHEWzl9iTiG3K7D7pDCDPjyITKciA01
nYriDt4DwC1KPPfNEMyzxmvM4O9c8a78p/eyhC5qoXaQyIAZ63lCYcngJ3RKcoEQb3z52DgtWr7b
Mrce2npDRB/ZOcJZLUaGxUfF8wQES2512z/C+4iUjnhsLLGKgGzercX4v4fQgqUEX2YBhQBg7bNH
iWITsNDZ/ouBRnyykQ/rzjm+fy7Bg014ovMPCrHcfiF4ffRL27ibINdIZUqHaTf7VzIQkG7yWHY4
o79RyR0pI0Hnx3TSv1m4m+2SITJijymREjAyC0Ap7Ike0YZmKl0SAUrp/QKBfq7XSGOXU6Jw34RZ
BrxGweoYQefxuEMX3xT89xxuSzTjv9/1okc94098W5su0JmNOU6Hofc+fR1WfS2uBUztqTL3VocW
JhOcWk96ooAvYcrbB39cJBYDffTC0uoYQib9mc1ZhXY7owNpc8RQf/2HDJStFC+SJwEkuvCutZFY
fXFysxV1zsKRMLpBLEB7ojaFod4J95aCe9k9BC6Ne4qrv+UZ7d0t7SGWYZ9s/0o8LXf/T3Sfqn93
aKUlmPHvikB4jKjAk+1SOFO/P/OzvzSqX4QQ4QsHD4717FLIBJxN7/qqAGXzTeqam/3PW4x4tMKi
5rv6nC6DLNAWRjk7rcR8JXaWPVKRhKZfyMMK7lO5xh4bZsFJUvFIZtmC5B84dI4pTaBtcwAEfLyB
bWCf47O+5zhupBprj7Yp38llWKeJsKTQhnjuAtQz4z9q03W9j8Hk0Xfp8YWiO0rHfGmpJnw3SWgU
byRTcK49P2SU+qFALuNpxykBewEpVNjCKsvCcRBNtSAT6MlE5mcG2r2qyfP1PyJHGHOGMpqOhLFX
Vp8hS1Lr960+IoZBZe718n4+PWKSILsv6Q+pbIPzovvJm2CaNPaoyQMPJ50rArLW0zeDYHNNwZV7
im1UJsUR89b7DUH5WTNr7x0SweFue6u8fqoblCwxDKL+pe34+hCJIlgt7G4RbFgT4oQLP7H/xLdL
RzqiYwN6uvHySRSGdt8FrFkp9ETEBIQvq9Rn2Fxv2FiFFLwzUm0V1+T0whlyi9hcB4hwzWIfBwCg
GI41+UI+3BbAVlhXKeBFGl2kyNU1uyem+r2JVRHGkP5JFaKV7ja6XgS8egBRX77bT+dbs7CcDUyG
MIPwo58IkqV6ay0J5wImNMExv3HZCcyplVpicy6HwH09vX4T7NE22bc8mzxANfH3MhKbef4cwJs5
2MCulnT7NWxvmFasFVJ+G5Gh+lblGrCThT/pGZ/o0dcGXSFuX10CpiRV9NkAe8YXS1jlqSve5pW/
65c1iUKaL8tL+DJz6BiZOML/vox5AcJBcNG4tka6W4BFJaeBGlWS6vpynhPp+UWU+6H2afa5B+HG
MGepTm8mVxr9KdoLb/Jvvhub9cxfsnSN2v+05uwggYkF742AHu83Da9QCJr+5sJhgPLEs65uZT3m
eElrPMatHAF9TK9d58p3Y5ybj1P/Iz7WSmf6wtQz1v7mcnhbhHpTB4NDmIv9ABcMg9xiuue7nYlW
cU2vxXG1pytHnHyKHOCDaLK3YTDpr+an1eCuPBgo3VOwxCFhvnMEu//kIpVyI5tb6a3O5n7Y0fNL
vAmgOpCqLFlZ15RavzhGMnibX08SJseDzQw0yZ+yDi/DaxFXENZqLpV1felYVrVGBZbxTjbMUblB
yjKfK7tRIrF+EwdpuQoP+GMPCTuK1iaYNj19tEhjTpE0qmj0OTv19eoEJObFEKGrHAEb5ovQKNVD
IYg/mt1lBUVWovdg5MvuXixozutJidja5BxaGXyvRohk57ZGlXuCvswB/3OtOcplU/6GcJgMD0G7
2JiF2JiN50f+nsD8nlSwBpJFjOMO9Oe6MGdQJAYRiCbcEjwmtfJuvyUUbeXY8p/jjS2vbKGBao0E
6r3k3KbRREubV9LUjmpAIqe3RH6lKGIKSEr7T6q37+/FTP3byqYvybDsG1sK5FKyn4zwG/TOmQdm
YQLBPCYeG2p7H+WBS1CG6VU0mJoXCYVALDeh/p8n6+YkAdAtBZdTLRoSURp2h9hzak+m517ZT9eg
vVt+6qhEgM6SyqKb1TAgvqU9VK+q+bW0dPTk32ZWLWCDZkRvhW/zdJfn56HHr+dTtdFhtVZSrK8y
h5UTXapxidNT7ybMeClQi15Qz9RDgAnky9eFAnLvbE5hHRk1PsSqm9iA3inmC/zA+cBNpo8r9MG0
kf9F223/8UdzioKQ5IF0qa0LUuoJ7fkPUBdmIkeDi677APN6izBoz49g0+KQJitG8B0AyB+o50iM
fLOVTLCI2TMHTE6EN9/xPO50qZSPmOp/MtqAvzVrRJ2kfx3lZN8PXXMxsQ76IlOW1asKL1ib88e3
tmm+49uWwJmuxFmvsymzwsJ/NTH/QiCnW4Kgqc4LDQgWFrk8rjt/SCEJR+ZOBnR4Pz7ZiMz2VXES
ffnKBS5VsVa9TBL9yMB9+aE7GWVGdtREiITHDB42J7h8XdJsZc7SiIpedmFyeLtIxjUDwfoe/j9W
U22ld7Pge26n+awmxm4MBjopJCClbHBMfzvJmBTvVcI94u6bT5xZc4j6021Lx//tv8gzkDEfAvPc
jWdF/CWmwKEJbLAsLn5/XcE01wPvthSkLyvfrteHaa5/kuzKOMyy1W4YoI8tVibQlKUY8f1KKjMK
PsDgls1gAtY9l0Z7yWmoqK5pdpsEPeHW8+6haOtklwQVyJsuDOUk03XL3cuQHmNVBpvjSAcMHBvV
g6/m/xWGj30iaMCiyCQOvC5Rwg8NNBcorFGJn9d+4WVI4XzS7vbdQW0lUcAiM3niymisR4JlZAwj
0nzVMaW9pAh9dijGoREcvk0d6Jq7e6p3AI2ZF6Epc4UQBkQ0vd/Wbd25IQRzGcqlKA9Ela0Bvsz5
vg9ANtf9vHbtNJ/PhN4LeeLUsC61ORgdmdz+2O0YsQV6q7JSfa2vkpmQmbLkw7GHlgtKnTIzCpYH
dH4zVbAg7Ve2+Grd6EgQ56Q/Lve13us4LBQp4L9vdJn/JUIACGoxM6JVmgDpcM9Je3BDJwm5Vb7w
9ax1Hfko3sXav0nKFwQfV7MiY4S0cZpqaZFMqxSI2kq6BFWRecHd/QYEe2HFXzuBOefonJD49Tm5
7UmbPZyDsgydRzG9pIn5XpPsQYiX2hN6erzOeynWOuJBFiU0RAMivJle3y7phZ3cMrPMVnHzyceO
lOaYki2rlegYnmFHt8PSoImUfrLucGs5qyb8+LQEpafxKAovE/n6PuYG8frRp/jLT2KELRKPZqN1
L7zuJZEaRfqKeMSk7al2V+6/vebu/Ng36vMe0o9X74andYKAfyEp4tOquOS63ziQz84dlyQmJZzm
7YnYIWKM2E+GSbUP8r5K3Ab8IfxcwcTE6Dz2nZxfY1nmP5Ug0+hkTzVjAIYf6XmlZ0PzItf6YX3n
tW5WhSJd9pWgCHEMFEOpsO2UKlKhEcGCtOfqdcWjgVJHzyIiSKW6owKyi0kzNkY7u0esR0lokk5z
C2Wm2bjDN1Xdl4Ci4IfK8lErDjUYLNSc1SdO+rO1ptzcAjlssGao0SyAr8HYe7i5/HFZKJNEG/Dt
6kWci7ELMjr8PgMQ7Zg1hFcf9Ut/9pUd1XQO9WkhDF2adSIw45umKkJUsg/XTpfpKgbsfm98JmrA
S6M8324lXbFOGmVmjRkj+/CmF/+7QWjjmqx5xT3OpY8kUC9e/Du2XYp/EtXbDr2kg8oFvNFpBLED
t59EeNXSFoIL2ys1qzmTIxIhC+YgMGpNAW25DaDb8y05ls1AxZpT1zbp5zNbZygJH98GSmiB3jnW
M9HP02DNlNKAovoP35+20v0M3pV2mfAjtfi6kEMjTf46t+bSJYbldlTaJT6+OFpA0QRMzG83jTlT
WHbc4593fjoSWowxZQGUvet3RJzFHLouSQkBWhQATti4dq08W91QA1Wg9101lNeH3ixGtWR9WPS1
GViPVTuQX3TMRicXvHXZZ5dvtHXKVhRhBDlehzMzd970Qr0giIUrXvVpE4UbTxuh17nfHy4YF0E4
bsRwc1aC+zYynsBy2xxSTzXCqJO8dwTQ0UsbzJNF0V0mHRD+M30q5ei7oNjfGYlBT/k0POcbptEz
ZJQa681uOG9dHKKprrz9vf32DZttkLI82xSm0icvINW62bgdrog0uGYumh2Akc0vYTOyPWH/wvvs
7M+Sfc35z72QSMNlxbdLbUIoH8i/Kb8+cr2hJw3Xidm2bPpLxA0mjLQwJM3fQXcbJDifaNtFlfLH
Zp59t3FnE06/fcQ0NhBbIYzNkjtSnR41+dcDcXdlohPVlnrI38LCKgnwi4AYhXRIc8GMRSnRLuQm
3dRODmLeJyiXkrNQEx0vukPLos1fjVoPC8i2teq7PpmV7K4cScQQgCtVd9p40Hm4DBI/QQzABIwe
ZwFykaCXgf3tjDUq4MYetEwrL28QXki3AX27KF5Fp4LWznE5NvvX7Rha4HJodn+sNIlFPNfNQmby
aHw0IfkQweeFpciVH+mg4sTW9D4/WKaxCoyfVGI8IpX5O8BNr3fdWYIG+OIFAUzo7HOj7MJeshKG
rzJ0Hvx8ij7YoIR0AXaMehGMgDGYeKGAB4x6JO+T2mhuGRZPi2RU3h6GggFGt/LZ/5EnVx3JIN5e
qEcoIXhInffI88F/TSGbIdF9HXTurLggWlDT4LST2iZIy3W83Rz5o+tYGDoBKS2Bu0XvIu+z+u7f
aimBTkz3AaQefAtJPF/cIcfyvRzq2L6uNGoMYBkYdxtOeGCmRinhdsHDVjMBV+r3QXYjVVkIGDId
N25Vt0wBApQXWpqXH2zKb6FDd/gv16a+ko5R5TkOLbRSjJZofsc6Z3c1t3/mxCKN4YOioBkjaVyb
XMYhcHqkumR6WmXo/dHLEsl+KMTkJvjJOTD2hcO6nQTXDIHYgd+KYRWZEBSbWFMEf33rYiLhRkRV
FpQp55XSAWwz2E1byGTxhJrc9+bJjUgLjcasxqSrePa2w6cJS7jEZyUm61Q29PSGQm0a7b565Zo0
HWip6/17YYahZ1aegV3s+8TdXL167fDEuPeT2pB+6oFzhernCELmVwTjuXGmdp8Ge4G83dT0JKnI
QxMoOv4L31vP9gDZx4f5B7Yl16T9Lq1a1u86cu106CjfHQE0V7qLJsTdcwZofNIW6FV0XOqsBjJl
NGrfQtvvXVNJpZhe4vmRTPGKy+44vvtFVw/3I7WO8qmP4aXTupqNMTjRB7Qnaiyir4wq9EjedwpO
eo/uF5nRQ1bhQhu3V2xn0fQ1M/zDvw8mYhEXBKGaPObRIGMhjejekzkdCpaQ8FA4jjkfYw0CeN/C
KWX3tf/5xm3bX6B3OoVAR2S+Sa9BJtFmYrJ8ds4ExWxkLS19CcmCyOWYKDojk7R1KElY8/ra5sYY
U9y4wt/skvfxgKiBrEETuQiNdGopZWitoKKLRKbk8UtgZHHzsT/oTNfbxFRRJGSL8s0GY+aDDWOU
4BFYFtTXINvFz25kqgUtf3emcxRI2kqK6hd45g4SMZxmgg4BIkZ+ywCuTOXzdic9cx90/I+3Bhls
YnDVAn6qptxvLzasgBaYMevOUd3a5KqCsmWGPkOTT2IYSDWypwW+wqJ6PvVH49+GGuVvQSzEy1hF
V/gCTct/z2q2Fbc5tMV2wmURkNr5frDJ25Gwh7NyLIuyWBQA181kEYIER9vQBti+JTMPY+r4ShEV
kTkBWI1jMdWZ8n1bRHtamam8XfI8cU//5lUfdBIuOUBqe/oNnpjhIGX5647S+7XXE5Eb8mg4X9vE
+jPbu566ZrSftESZtrqU23jpTj/DorP2qlZ9FzRdBvLPWuNJASK+8y7xB5FnjYNV6Z+WAnGuUJWM
Zjm0Z7kG8rL1dChAk++tSuMlAv2jEh9nFrmztL9/m2mMTUBJhG+yFSO5FQ5BBF1p+f7JBd7ePqDQ
baM3M3C14cIGUzaV8AZIKuwNniRstbXjSgbMPH69KigGt6Ik/bOW1Y4c26tDflzBsi9XxC6Yw8RY
FtDGbFk+Cu/277grmXqiblluo2lMjWuKGH88QVJl/H3S53YODGFt0g61P22T0Y+vT/YqLSNBoS6m
ta/YL/YnkuqNRVS0m3I6SlQf4hEd3sAv9JoB4tRo7JF/u0SPBCmH7bDO5f0BYRrdOuojfIGYWlBj
lFgmWwKKwP4vz3PfxBmWkm2vnAZxaOMaP9wz/r30/LLImkQ5bl2vem4kq3sQB8StsdTZZHMom1Wk
aQJ3ak1888yidiYlupfmClH38t0Stbco9+v7SqbVe4IVdHpfgnKm0wCbtVIQI8YnLIULvE6d7T5K
hcNkKrQIROqfpLCjShvKgGnbonROGSUibSEGUaDAzvAlXPMcSAtKRwPwE1iHMP6c77p3J5W3lDU1
iij6Ij8hSMGJrPDCdrss0qb0qjYlZEwRy9HEnhfVkkjY7SwMdhVjrLEQHgYHa/4yQqvim7odCMr4
Wx9kCtDtqZZ9i+DcreftW6Po75nZT23bVluPWX5xvSXpKcoDfJuPP72fS2J88CA9jvxypmsrMSZd
l6gotjSZ1UfNOs/1rQB+37Y4NwLCOId8DdxPn0JsfnmcYjas06iN68WN5A6QFMM8wFtDdeuEqI2f
R2uY05e7RHSKeojfaj9otpCp3rDgEm68fB+QYUK4JZEWliQkzESppTkoVTK5gR1Pv+0AvYHsj7N9
uKBaK3C9Ub7etke5DnC8FOTsBAhkgrsf9gG4I741sbRMpS1Eh2NMGXGTniwc8jb/B0KekBXjCXxe
auWctVzDBIFvmHqzLRoeUO9rUrow02Ok6OYHrCgceo8CdTHmrs/0qmm9/cSexRtLJ8mKHBfK9Vk7
WVLKP9z+BWFOKxUDlCGWF5K0UOw7AJ2Hbfm/pMZ/TqnoeWDHpYR5SixOwZo1WtwPgjWCYM/rNQ3C
1LxAP6hoQxqfoQcymP55f1Dk4HIe/AQcFQY18N5UB9VZ+QL95avXfEQ6OCAac4hQR26KS2032+4L
T8XW6Bm5VbzcWY1j9KZkmKM4z2XK8x7Fmm2bxPWeLBWr8KptmP4CxqanKdUnRdKSeGEeksxM6hNE
xIS0FON4TXQrhKLCLOnzQUpjebZJgxaBj1GHhytTnAkem5MviWvDKgGbFhUeI59m4Inn+V9YCNyD
EQP2bjKE6zpMXKwWzAmpJ78oTpAEc/TB9xITL9vAZrLDIEaXZ8rcaPSSel8Y2ppp662XvyaIZDzL
rMsvbEZ0vTu/7FJ/JaJM4TSuC7VcOrWaD87rfQCqGDPQACb/3B7Z+9LGEuvBpzoprW5C+/zgMmDn
HgCvwhZ7C0GI3PULirHSQkc1SuB074qLz6H25Cm1UHDhrSBG3JjWFsiPnLEMCPJ8WDuM+fuFHSJ3
0vMLz2A6lT/NrcRS7R8ATzXEqQBl1Rp+oFf+6khJb9BH9mQ998R4EvZF+qCxuxuUqIW3uv3+7O6L
IJtHrDqLjB9cNXNxEiwGpa2MDZCKYLcrA+q88vvCZ0iU8kyF8uFUcCANfKdHMqiAOSkjaQm/Z3XR
POPu6nPB0qn7MudgM+LSYsr4nDeCuzEPrX9GYfoCC5YldjbTNvhChCGfB46H0XGzRbKIW1dpF/Jt
dvlNfm869zC1rKscmRbkIrA5QTyleI/qRwE9uxztzWuUkD8WQU//KGusGVaEkv2Iya0t/QQfU8+9
3R31OaqvexSw1Gvo914Her02e0qVrto2STGgOY/OF0FyQw63udWWKVyHzT+T4vISK74oQTsvQhSH
vcMxe51gkia+TaWjhKeqwdZupTdj29H1/BCWD0I4Hm/burdVON2G1ACoySwsSLCkJ8fy2x0N54WC
49LhwKotWfogjKV5+zKgsNCzEPqcbb4xUpHtPTXCLMjmBk8OTP7/sPM2k1TgtPkPsLHueHEotNFL
FvjNnhqiYhBnIWQtd5HXjogFOv7KvNSEVgTDPmn+9C1hlDzAnHAwEEDPT/RVwBq71jxJ/o4liyCA
KlRN9iN7OS3i04h3ld/uiOfnqKY9VI4HxF3xhOMSBdeMioTGX6BVu7ClOw+0mof+FYCbb1L3B8kL
S2DyfhOrydpMBRv0l6xgmG8oYkJ95IrJmjuBu5j6evy/lhkASPvBTB8lP5TF8sHvB3P9Aa+48OY5
074mIpHBVKArCHf5CG2SliFHA5uAsnqJrAkH0DZWOY4gzK/F4+zeCMhLtIH2NSDnkvnljZs/ogiX
sysPWepVMXOr1vp/8PxD3WrEZsyk8FuCXxFRSiTmsqxQd2hYMWLljX/XHEPdf1At4Vprg2t2UvaP
vcVRB7UOvC5vVPrYsOH49sHmYC/D4LHTLtGo4DH7QE4cxyBO60uL3M9NI1NKMnWqnNdKFlXGMz5+
79xJAUeYBRsAv9Tg7mTtiqaxdZSQhdxVUGeA9/Qmr4TKVna6AVLGQGuVn4iuV5wUego///4j+aqS
uf3zo78nHqftyNAc4PAFHq1nrqhrWYWIMH3+pkYS/Y26KyNvJWjCr0fcVNqfUqCGHhKQNq35wYYY
y8xsFJgezGSkzWccVeKODIXpD+iUNylMumaAqe3EWzG7H459sSibLIQqKrzHl4TvzI6jxZBK6JQ0
NiYjM8tXz2J8uQL8r+CS/pLodtm/inOgVIpgUyAXo8w7sxQ9hWl/I9R8w1PkkFWoXDFeQ0jMujyy
1vRb1K85Qh3S3yIP/BDuWIgCTASpUOjVBpUMtsNws6bRIJ226tTy5VWEOs+IjIYUBE+Nc3iGI5BN
i6UN6OGuLHKeJJ0NvFq9NpWILs4chcDBgmQSKYsHLjpi3W+UMLW9L82e+KQrNUmXeBHS4A0qP6On
TduxEURvT24qBWi2hT/Ht/MgcE1yYbudK+YFBGCCtqE4e5oRn52+XUic17h3D5k28zhz96pvzrew
FRB6A3MFRVqxv6OkUsNWVZDZxiy4oJUQaf7zrdk2sQiQm9UM6rwYULEhRUh45WWfHPav96iE7X3l
9oiuoDMZuZkedr444ivgnVnu4H9kANMe7KF7PJND0wtSSHfDy1ifX/fAHviCRYFui0xdp9O1DKq0
gC5g75Wd1HzvfImcFMC2uD1/ujc4YgFspHwIxld07Nsgl2eFgT06I1b6nTC7pDUCFglgUysgpBjC
vOlsos/UVEUiQC4NPf4SqAXQT+968Ew5HbMNLXWXRuJe+jgbfWVbnJ1IVVMAKo87taJNIgftJyUQ
5a0teUxfBy6SUtHtxMSideZq12gXVwaWWmo3OKEMUE696LmcO+uVoDi5a7XKsb/kOPZPotUADdl5
/5Wx8gWz2wC/QC+/COTBUWkVulZKxBAlR0XvrHI2LOLZwh50oORMFS6uyXO2wTKYrE6Jv3cKHNci
rt4n6Eq9qVvkwFrQtQix3bnLJPMU+zLJbLJ86c0LObCan5DdbQ3tYNnLVdCAsXk8IWGS5YpnN0qo
vIRBJxS7c0xOtSzTMsrqZHEs6KRdW7YS5lUDwtexTFST8nE7UlRywBANkCns5QdMB992Oc1cpUEQ
L2PRUWND9Ucc6J/vVzdWnkXV5zldKaDLEUw3gBj/LAlKxK9n/3ntCMEpLagdbiB/Q/ALVZTry9r6
ZDjsnya6xkKNmU5m6S28CjJdu8L6vEEjZy9O273S2jNJzCCzhD/0hRUG0CLKCz2JhczZbURe2U0K
s9xSGmNeUgl/fQDCDlx+zAeE0gaMTgCtei4AINaoKuxSiDtzOjTx+8yG+5bBrUFFlh/+CbQPP8Jf
WlDLiENBm6CVGHaRsVz3wWh07L3VNXYI6F/h8ef/gVUMyAU4rxg0QwRtAEXFMBLuJw0fz/4JNqlC
QMYlAA7uUCUqlBcMfZYBnHT5jhStmkR2ta1vVW7RPsajtN/BNK1mkFi15tGfpkPryOsOqsmDjNL+
wu+rnxW5Ez6J+SX5/R/o5Gu+C+o/o6nxmDmdWbKnNnpJan9MIoCrgP/KK1Ekd1NDopLbTSmSlrGU
x/bvIxoui7VvK8QcPbP3rM9mbYw9X7GTf/Weqr4W/pyWgLjAne0sqOMhDs5Tn37mv3hicFIHsi6T
HB0SO1CwYsB9XpCEris6x6uMH1MThcNlq6CZStihDllnQCfWhizROTzM20VNiIwcTcoQvMuWXUYc
BQjSPOfIFo79kGsZ2n9Aks2j5vFFCGrVkGkocqUixg1NkE2IHkGQ2Rw2dKpruYNg7cEdXl/M97rW
CaUbXKzSD+KIa5oE3pROI/xKhSCczWrqQvJK6/rrnJJhujh+kFbgy4VJZEqQ7rvduRfJjKfzu3qU
yes+cC8R+EcUBiVVK/pUydZCC3IWPh5MCskobBnXwEuRYNeFDocI6KTblXKB8TtRYfShAa2+lFZK
gx53sK2OtvZmuowdsTC2OD2/VYNKEAcAT3fXOKfJUhrukAYqhJedcXNKGqNH1tRVKoqmVvGMeG6+
47vCiDd+cLLxp7ImTBHBg9gF59Ytl2hZFF1Txii9NRRkb0Bq/u6/IV/U+if7DNxoj25Mf222TQbs
1s6TEmRdaCISNu/msWB2LynvCwJNW2LaNGnQuYt9KhHDCrf+wELbbNKGd/DHSdgaSzdjcIjxRR7Y
P1JNR7nN2Oo1gLAEEreVyMkaF68Fy4F3AgXxPKAU1SZlEngyuwD4Yw16yxUXh6Q4N3cwwsADcrBm
qp2W2oXbBN3k41tAJuVB+hkURuK49De/8YNw+YPuUJwcq8Pqgjsp7bVJnADJGSAhEJA1LjYT2w4Y
JU89BsarxUYPYQ8MsiOKnT0OAOu/TqOtgvGdcc1n6zYlLg79yXaLfhg9GmqPtaObyVlaK0bzOOW9
KRvFd8Fkm6VTrrFL3YbNBvLqHuL++THC8Hfsiy9YDhVZjVbhz7UJzig6ycFfuexWt2yidpEcZ/A5
rdkhJJjChtlGdFY+bjW0nDr61KLZPN3bcDUaapjW8FNPjztF3gfb+e6/bU1bXVHsdIwDkOhZQbbA
JkRpfakqdRcoUzA8gxan2vQHdCVUlDwWLbp+hRD9KsvFeF6UFDjkHFRayerviYB7P23QzMvQwnAU
wkjzp2OghRNN+iYmUF5ogTA3Gg6UJ/dV+VAvkSBSmCYUeNjutFZ+uUkksO7q7rtyRsk9+ZmDr9CX
pq6bLEMMQTD3YiBOBbkZWE3oK3WDYfoHh9Sou/lPaLv1FdryU/vPHQYU3PHlbnn0mBo+l6bRtKXK
2dlKhouXCUvTf5uXx+jvmmYCn760HLrcV5hM8sn0uRkOrDgcby1XXu80nIS8mKNUCfC1Nfxdnf94
f331edmt9h6J7ZQUdHMP52eGl5xnMcw74KTwdF1xqYn+lZLDB/i+rJMMLzVkXeh7POsDgW9VYsba
/SBGzQLve8rd9n1zQYOUJ3+ho/qnRKMesLIW7yvV5wQ4CTxXN2OCJ1AjqCPw3UA3V9lQ0H7bR6ne
DgQnE4U9yxsSJ6hemOxBd1CLv0ZDpB30XkeLRG0ty4R2pnDCgtsZ2kFLRx/EqUZJ/rUNxASgC+t7
BFLkrSBeZnwv9qaoNWHxI21D+ohqS4jIFeB+2IRAiQWAMe4RL7nvTIJUWdJZ/t8/0wV0oINyL3to
0Ylj4pTWQTU8TmlqhE+7gdLulSVfrhAtOndTUZ9h0hnB20RlhwZWb8C0UjNmvy1KtJ6OfYBWs6Dj
h6THsbbtPwN34OeJ7SNnplsnVhMEdRSEboJTrMfdNsBuAEKZzuD5KKHic+2CfFWpzGDCup70nOfn
XyEQcMEc4/nJtXX6EaQ4ueh9pCZxFy3PQC4+65AgnZvoxjfhfzoiDM3+zz+v707Y9dVmnrcWLqSo
DrT4SDpTat+V2B/V5IsNKEdiI8E4mhfvdcmNmveajofDOfnfq5Pw5YFb4sf0q/x54X98BV1m2QbW
Jzagz17lYNN1Ql+SnOI2GS+/9flDNeDLMwiWmibzlapeQZG89GFAoRgfXQJfN/Rt1tMzzq33sJ3G
K3YW9OnGs5binZftVq0sjjbxww/9BzPw3I/uCzQh4jmUDi+4znuQrJBFN/krHt1Os20gAG4i6FRE
MXAXML/Zs5cVEbYrEg6Vb5+ppJU8BON+anukIdkVYdbxVrWXLyY9On3P2iojGCTAOB4uWV/F0I/L
Bw7mrkUwjBKQczixOsxlw7HvtpPXbsr4vDZZgYhk/a9u4vGog2yJ6Zs2BAfpCFrKwoXZjcFs9tFb
Y+v59OEa76u3FrLiD0ayTXAmY7ZOjpodKLIZji4dpGvkSuws8e9/6ibHDDmiSocl8m9UmuhxUVZg
6hFz0vd1ufHlXgLhAzl0VBPwouHlEWPV/QWfAoRGUB2FDPVNSy6ydzGnvW+F9v5b2zXhDvE5F3Nb
E9zuD2EAx9DlMHTVml/El2o6z/Kb8gQVDuBFWDjMnkoLCpvZmCpUlTTT+A5z6C24707HQAhf6XW5
m3pWy1614NH65BcXKW+JfBxSJSGmQDeHdI68Hxsbc33Nq/IIxX+n3DdQFH73cC75Ac44Pfka0xJk
CDtVv+ro7j6qlgteR8YiD4/GA5TrOt7aXlF9UnCmWNjAhpOix2y46MUXYo3kVyvAdEOW4Cy0R49a
DX8icxJYHfBjOpsJ/MkS2x72avvBmJB6xEAoPxLV8z8xGJeG5ACghI2JbfQnqFfg3Mey1sUTtyfx
X09+rWYZaBL6oxpFMIuvPnIdIjMJXwSnvzzSoPYTiFDifpmokPUB+D06BpEBgVf5QZoDl6ZwldnX
1Kd99CGazLdJCe5r98z9w1L7dfkrBJJxTHyqztQBdh7R3cKbMcxEAbm/nPvgFjYHvptYzzXau7bE
9dAf4vbaNZZGLWQpNdNL735g0gNVxgT7pNwd8XzHtJqi4+efytZufSGE2t5kQXrY7rBEyXSQ4LYj
Z18/6QeGuNOXG2M61KMbmFyLop1eN9dSjvXaDY0gbjPnV7xm5Z5ojq7wlsqviMW9OsSx0mRSQlaF
Sv9D9lVfAFe2pIfDS60pkiCTP/vdBYxgItsMkBSCdKk1CF5UbhPENL9dBCzNEc8GSyJIls1hCKzB
Qg9TVXIvRK46Bz750UFjtidieGuDP7jGzif+/5aGd9A5C0plRTU+WQvL9mS5l2R4zOEJXqx0ZciW
M9XPcwLZ/JAsC68Eh99O8RBMGQ5MJbjy7NT1fhapwFBCL5FF3zhPP9HdIy7hK0vXm5Mw3PEr7+Cr
dRXnxWTvCSnIHihPD9sWTB+45igHLd8ZXFpxswGzCc+2OmLcS9IgsrcZrD4ojS4/dOjEE8nGIJGC
HmlHtdlNBLvqh/Afs2Qwb+InNX4Wx6iBlOA605apJVnsUvQ0Jzz0Vc/TxBvVxfI8EGDzUBDZI1q5
DKOBikP23a9kqPiTxI3XhFe1OeAiBgkM0e//kRGJg80LVzFDOJGYIgl5lqaJV6kr+NPf0BJruaf3
I135ceDOTTzOOug6eY6rHt1aIROyGVB0X9eMb6JWksgtkU1FgA5y5M09oF2xtjnPT4FlgpVjJjPb
S1qU7QhCyKaUYMKx8McmkycoiiVXREEufF7DRQcEeL19o2BYZM428ywTqt+fpbQLnVg58PwEBQEG
Qn0dSckqtgXH0Breq5qSOKwym8VK4VOBW8YB3USHVIxiGbE8ISp/lPHMUmlYsl/2lIJJyX6Y9e7s
LFukhmP+Rl1vcXBpr+Yt379pePa0AtK0DRu84zMeko4xBKMlOlPREPllqJECyEqVQw1S45vwu3Pm
Glx/I9GwRleD9ItDa+ytk4VbHwg/RchFzpv1w2vxJAxs5LSXz5fsIigcRQI4VRC7jcXPsPKmy5Tu
BO6rqCvNs5w5PO1aycxvU4NfcbOfBOhM6/FcN0HvrYEB7qgQ6eAxR//snVMU4Y28KgFgyk5e7kEe
s4pr0kdDJwI2MC/HdWTJlnbBbcN9mK1YIBWkVRFx9iihTi7G1xFSDJqjEF8Eb/Tli3/4dQqlJ+kR
z7WFXzFSzY91tBXgdmDr2yu67fEADtQDZdXaltPJF9qZzfcJmvyxxyEdjv50E/LMFUOHn4sq36+b
pJsH78beQyTQ8LuwqJp1ea24JlsAXJPN5KHRQ8p08BlrXeM/2chRMcaowvIt1Q2AwhBbsovpbdeX
K7Vb7TFw/CiNeWIA8yhc9lbCUbcdUa5Y0l0sF71YdJkwELc0lTHeN+QEP07zz0ilCMsSnEEMFXq9
UFXjS3SO/4KqKGkNsYnFlmptb5q12ab8CfthX5vOB8Osd9k5v30DV3gO1kSvIyyYkQqV5m/XXbJ9
8luaoToHFGgmr/Y8S/2iyDNDDg8ASzQuZf7QKosiQAoQTfTNZd/VlEMPGvr561VLHNiVm5ruH6pj
gJnoKo68cBmp3XCom1lLedMRiqkujUujvR4aTm/8lWcqtUkINjCwD5/y7S0QtRVVWEA7j58r4EcR
RqLyM4j+9NkjQ4b9G6DLERoh2TT5CFEhcmYMmyyxnDVwEY0fbY+DPqRuP6ScjEsvFHEanYWoQGxa
PQFmqVbk49pYzrS+lAdr1QiJBXkHnN7OSCGtt7wR5H+mpo9+Ufq+RI3VIagTeZc4cJ8rxtu+nPxE
diweOkB9orY8Q7q4u6Qv9EEWOCUJk4xWEsgadJqKtA3yrmxhQ4Mr/uYcerEg9ai4eBUPijrTqYRc
47ZdyMjRUxBDWywIfMM+60IlLgaCgMSibDgNMmIHb5u0QO8lbrHSmTEgwBAqLf5DzVnTVEFE5aKs
j2pC255NQPEjHT/U2GS/aSO1aSAZDQztoS9ohjzWyDUfWgBAkJ4Cz0+8MdpkFkaqXfxaB212RMK5
h1Japc14pvbr5GogcAC7R+gaDIWXW8iFONWnVBB3SK3UewLuQJFp0ekav/OK/zOBxtkCUaEvJ98P
NYvkamMYw886kc9/KTxbE+WvkPMETOOGnG2XaCR0AcXuo/H+Z9A++b3mVpkiCyroXhIR8eCOPteV
wWRLCH+ZmDCxY5OfukvJ2azA0gNQvXfI8OHwSPqpXAZSXJzzmPUHc5AkiDfAmAKyNuO2wc9qaN94
83fg2rozTdjE/ScJRAGHSolAdIqhQrAA3ctO5eDfz8UdNgvIZDIbcGcFgMHamPqOSuHY+E7SyQzk
+0ZqnnjpV8AvfHUvgMJLIwonrUBDGF0nB0N9FmTKBFuMM1MiwnVa+0xYqLnKsq6isLl1ZXsrxJSE
u6ivpvYTDco/ocRtjFIicT5ePpa/p9w3/kG2nFAaZnly3cggJMrQeUZEhGkcVoCrwTptRyGiB1/g
JGnSFPeaKD30fSJZW3PHf5J3iDSFaSTI2vrXNyUNNO21P/iNIklf2smOiLGuGAALF9aegaUmC/MH
w9HX9tHjh6la9rNEBxg4ciQa7OIpzjM+iTTXEdweL/XEjGPo/dO8o82FD+T7g7yE4+9jwA/GvD0M
hDkMO7BoW2+qzWn27KMRJhbOCsUC06Fk1Q3k/S+Tq3BnaKuJbhJvuDNrPC49ry/cyXwS3KQI9WgB
+gEW/o0Yg7n1aN2v5HY9SO7qf1EGYqjSrLn/5pCfVNxV3YdWkzcztKqDVhwaWxyuTe949HyNH1+M
WOO2ObV+xmeVdLEhTCyEDdKRxOUzq8Xe7hS1H8PWPs0RRSEYmmYT1tfZLqPj0b68JmouN3Jgbfpf
CIt1f6bVirobIHpJY33lXk0v5koSDcrO9rCFQvOeKpPHruARxbASU6T+Cu3V++lHg8vfBW7n9nHd
oLvVzg6IneEhr/zR4Y/2EMOJUZdZQKNmN/BQaA25iDOHaVaXfD0DgI2NFXc2pgqBwuLqwd0BnDci
XsWO9h9RQhW8iQyok133kAvBtnNVgtXBP7HhsxFc7nJaRuhr/U1JZD0lnqUZfnSRfXvr5W05hdTp
WnFLjQvAVP6nT9uzSh1lJjVhvMzw93PDGBo11iF+55u7Ph6HvZ5DnXh8sYEhyJQ1EObjPOZnA/4r
GsEmnhfxJL3EbWh5ENlUsDlPnNuJI8nHYlnlq70n+5TiMbgGZGLVqslysiDEqW6gwEo1e2lCVJwN
2S/6sESFPV+IIPsoC9sywGd4o4xbpJUQA5fbYdqKmHyvmXya0gA82zYG/Q1WCVNme0eUQgDCLZ4A
0RNq7BgzJO+sRpt+mvJv9yWrG/MMykDf1bMzSEAAYwNm+YBMII6T6z2qQbS1P76lA/RaL8b1UiJa
feOY4lYLoCd0Pv8Ad3S4bgTZdrUTvnu4rb1bQnxop7pyj9eLsgmBAKNKEJpLDm3uScNLOouuToyU
BrizS38WfWPLeOPzSgyIezskf1U/F1DIfF6Wi2UDMk6dAQZxNcT6W017wxxstwF8Etszjmjl9f6u
XzQnOU90zTPpdpOs/WsLgiZXsqXeaiBmUzQmIfINfRNyGxn4KPA9FCXjqWJlLFeiSYDJpt32dzzt
nH7RABS5Bh2ywzjmtNFEVRnxfviU2hykZpwR0y3hOThBfaqkMh+Ma5qB4pm31pS7iecnqhhyHttp
cvQo5AM6i//3k0vor1H5PFOdQsxnp3ou7dxRh2EO7HjY6eEuP8VaQ5u8zgLNkER+oQo70EwUTc8t
1NH3jsHS1cQ4GBVQ+fmt4LmDpEDWBoHGE88hJpZfnGNjI6oVwaf+7ekaFj+KiMgI99jyTWLa2F20
d8ubPgBEIfIbt5HeeZ9S9VWpIi2VavNCm/vIAXSJzuYN1gJ4Upqs7vMeWqyRGe9dDxM77rpessHz
2r+FbgqctRfacLIQSlAP57SiPj0ficro6hoGnmJYwtCh/7CD4MXruY2uO/SLm1RNYXQwFiU6X8yz
CoWcthC1bfZXeuguMJHprXOU2cC5fBV1XW+93ncSEM0ALBXC3eZFJNEyLLhIuE9ZJn7w6ONffIis
gxMBS9e+ovXCKitT1KId2WGrZiCxvSwiaDMJOxQfUS+/xHn6r4I40HDnErmTSNxLOftnZGBSG3t8
r4rmkiJ1nLrUIk2xFK16vK+2dJQOHn3GHIX7n5ZBC/No6adLSt73Alm+meETKidz/6ivqs7xfdSt
DoiRBQOCYmcKvFKZnqtCFCgpuTXCuNzPa0kwPaDuuUER6pkQ+Opi5ISO9VreF1ZFdnyE6Hpk3+ps
4rs5hqa/Ap5AXjTTxJTxXasaj03BNsa9IXvpoc+Jg+52R8j0OFB/qwe24gNLg9UWGUSuEy8MgHsZ
SkyrKz4Z0X+Km61ZoopFOjbwjbswgyYmgcRQezXgVfB9U5PMCJhYZxCrSiXLfo1quUDXl+FkLcwp
7wW3O3Mrf43cyq+QSyIrjgRhX2/EY/mlUljht+CCwVcwTTO2Rr5lqWMhiC0S7NiuTfQYS+cIXQKc
SZBOL8YHWPt+Lknzq15Kr33nP2/9MUNXd/5RMNNn22ubJ0jAfJCSBLf0nEqYB8lHiurbr2GkzoRa
Y3VkcMFwiA815AgRYN4S3M5XI8iOZFgJkiKOyMGimJh3Q7c/NPnrxLSLA8N2BSIsbkCRr2RVb57y
VgUzmErx01PYq0hziAj79SccP+BAq/RCXo1b0rcK3Q3TUdBuXIQoXdbQlmomi5ckLJZSOoLxFvNi
7H1VRP0oxoNKboyvCMMHr/QhxBCqwE/StcOaZffQqXayYo5sGUrDav7Ln6KdtoPpZqNUo6/npIWg
aQFte400TI7uh0BWNX0G143BsA6YTV95N9gtwfyC/Kxja/TU6iy+mdAjnZP0x5Gk7tCB/eTL21sQ
2PKi/4XEAfhLwANydduJTOcHh9xZGgPTeBUWwIHEu7W4aJg/lZy9dCeockO2PIVrXIED5yDJxpi7
3yPZcnznmmdjwoX8VUpea/xY5Fd8+c2ffu8T4TGC1K1eDRSg9oDPJxUG9RXIGtTzN55lOCoFTOb3
yieutBXPc58KInwf2Ral7Fx01zB/jSJPkZQrP+2AN1uUQBgSQVHP7QG+xvH3NecH+LK1C686Omqj
aBqMp6jIV0TfEdtjsJjU3Xt19iYtw7MoewHL96lKFfhn1reuce5FYDs6pdqTf58x3pimw7qMK/nR
GW6vqUlBdCeIYlx8MiGm6cU5E141xsU07FpLsokwPO2WDP7cx5gPLBxW9busCmXdMnsdiRSDUZdl
ls22C8lBnNjEYNrjZ5gL8nnghuqcOGBbHyfmn1FsFk0wx2kcoQnpp+oH6f/cP9em/p11KBjlGmAp
cCsJ67itNybbajngRTdtucnJRXrbJIrJLm7tuPz7Fjq8jbmwRdDGE275Ioe3g55QvpnDL6yKMuwf
/vYPXo6D2/Jl/tloUVhHs37vZ9wT3VZReGdzrTJygpzakGVpS/gNt6S7cb2ZWxjKQJV3xXhI4fDD
9W17KfDDO6xEdUNO5idZsM01i3HVBreDbsmZFWRjznxGFV9iQCOEBgrkyIX6/7nellVH2J7Gn7tv
1nzi9+a3zhZ6PHPcXGj3C1jATDuMxdBofDvYyH4iWq4TZ7x3deMg4h8snmMhoFTtucGYvefmEbN9
nu1xqTzFM9pgyhPVX8QLM+R68osFRdEFyVInmQqSeK6s1gcrW4fslXjpuRZIeEGx5UyR8iD/ZFKF
YoFxG7fx9mMEpNXeY+0l8v7tVDBs27xfVgo5viVSpiccAHQB9BOJeokOwY6gnlAnBHjsACL3pG0I
ZL166NxLngwQYx1/2Kgb8RwsLzOmC2ONWzQ0GdhWF+yXCGMPGj5HPlYyyFIPCNdEqpchf6IR/bRv
lAAy5NrDDu1O9gsLjKLHQ+5856HsKwTNVAJfYbpPTZtKHPFHrTQ3GqPtZmZwf0SxKLpc9LQdU76M
8NjLZgRN24mc6yNzJ0tB1mv14KRdT872Kcp6SDnEanxXgEZthtuai6T0qI1FNr9uw4uMAiM1isI3
oegIJAtGxGJGzNGx9PRv1wkrIVoN9Tkp3EdquSlX54+roIO/GH8o4aUuZk2jekosfRzoOzhmDEjo
0W2eqnzvajsx2iaH91eyxyip97fKi8DqYpGB+7VAuC6y4Nd1M7t4CB8uy7i/mznfQjVAAe4yozHL
Z89yfwRirzF/S84GlpSEr/MRSsSgSHwxm8Hpkjt9Bd1cBaYlILt+hhXtjk0w1oSQlvhwfML9N9qW
eE9wPdEtDpD4kuLuBlnVZrQifzdOSk0NGUkQcG2bXpkg2PWiLVth9G2qsPH59myHkrP8i+axMrqx
CmdaLeAAwOCqwx8Oeta9zoog/rlWdMAIXhQKHV/ypBIZfWJBk2wpWgHF4j3pabU4vn4hI1PIUNwK
ckvyVT6kCijkw3nZ4JvACXbqJoYNkARZpoVJ3XcaDXB9PBik4MnVbv+kG7cIEwrwf8dhG0myJIfb
AYEkcY/U8EuwSEPr5AC6O7+OGyhPIsWhGs2BtxayTb8iHDoJ9QnBRTzW9uqJvvt1uujrS9TwMz8a
v3Y8ad2ftVO9dR1gviszus/jqzgLg/C5IKtUpj/37jrO0f1Pg5lIYxxpI3erGtHdaLYVoviweg1n
izzM9s3EQLZB8zup04KHasgYY693vFrAf9uIJV8vOmE44+HnxtMtyqhW944sGTbBo/wdEiu4si7I
Rlpipy7Ca3rxxWyMdvpbDjoZwaZEZmSL13m7xK7m4gnKVT8g3Q2Eo+1vEzQcccKyvmihKdslez7H
i7QUKcEKk8+WWtYgpNbHanJB4sUuxD3fPyTaKOWpXpNH04e6AIMSHIE3GVo0FuPMretTkj86aZdA
uFNO++sHrirQy/AS/V3G3nciwBuGGAAfKTxELBx8qBlN2xgiWfMZHHeEDzxcahqv/fSK9MpjScvg
6Z2GzwlDuw5Xo6r1/alylF/0WLqR9NwO/P0Sp9oU6n7oVSSLInyAW/+kLfbED6qUbhm9N2xV05Qy
Qht1UPVfYMtLWVn6Dkzz9d3DYCZbsSCv9G5/s2sRXxDnPGlROAFIFIOpnNcy2pgK0ZAOT0WKs9Tj
fMMQdk/UoPT5XYYzsxYNDrl3dG1hE/KXUVfZsW9XgvYkTsli/w+wMDRs/4qyUQ48IFCQZMokPQ8V
N5ixIsBuc1E4/Igl2W387qTGcNPzNTQ3Ke3EF24yOaefNXKPu64cVutKHrL2rXwWW6JQ8GZSfNuV
4LbTBzNtrX/3MWt/+B6DeDzCmj4aVTvT9ndZgQogBpqc3O0QolBUZlz1Tko8qtT2qjkShuEnKTi5
HWQPd88OceaPC+ljc76gT7+QwUoBb6oDUn4tGRoa3tKaLtInhnQYW7BzjFN1h+PbqpI+PK8YUtiS
K8Yfv+DocPeDUAOZEmu8jlXc5XwU1FAqNwGP167+zXXm6Yg4VRssk5MwqcbopPriEMB989qIuOga
M2SixddiFh9lRlolS0HZz8CNZTTxuY8ctB8tK26hYRc2KXe0YGBZOx4id8UkugrRF24/VVzZ4htH
UltspO29CU/WqkBiHpfci2YiU1OpTKNYf804ONWbrNvOerdRo8/8wQhUa4nZg0Y7yY5TDaNoJ6VT
f1ARwJjYxv28UlKdPB3pzPWptUJ0U/63B0W0r2LJ2kkIx9D4pXpMGl43C6/8u6fjnHFvI+2xQRwt
K/bgs/zCW9JSXr6wzNnZ3ZjhP6GjPIKfjoAl5lHEBuBhpcPb1TMTQUX7lhzdnneTfu7Znskm9AsX
qJARP04Ee4z783pW+6tbVWWpr6J6JNuEKRnlmCxG97nOPPjSnk8v9RfVRSvN0C12oSKm5hyB8KrY
4xxOwbH2nLAH5Z1Gng+xRB6/OGRRNbgUzFiPQjdvIW/JOaAoISd0L0uLd7Ued2dzqRgvxKNJkRWY
x1klIny4dEizOGawXKmheHeHuEpWery+DzxIgivN/w8c4PN1pngQp85sW/bby3vhl5ar6NmlwgHA
wsfT01aGymvXVM485du3YmBoBMNkRZFBC3esNyzJfiDPNHpfbxOPWpRJvCQwbuu3oshYIA1/KsaP
6sqcO7eM7kb0kRdwpYn89BvmU/5yh7Im2Oe4btsf87l80HyF337O/Likf/0aC9jBgj79uCNTGBhK
YmGvpoLeoY3PJGSY1SEuWiiz8psx3AHEA+7rc/xkO0RNikbV9IOgujShN//wAT27t4NCF7gwkMPe
4EXM1RmfGMiHipJUFZjmYbSs7QJ8X9/FToWYFg8hjq+mh6cUIZuhlJkAtAPbR61GiBWqY0sR/c41
ccfwSgQ4XUGfzBHpArF+QdjB+7cqDwJXAevtv+g5G9tjne705AsE09GJUQn9vlS0ZOTS9mRoq0le
G4/dd2OJPSYgqpZyRRG/QVve+kFORowIrQnA1MsA0aDaFHEbSJWV4k47/EJyZn4GwDwj9At2gJ1B
iMaQewEmDcnVA072SwRSBgGzXs/CdezswCejhpD/y+ckHZ5JlP4cAcRj0QymRKOQkcNsZr3Jq/N3
L2VBcyeXZzoW85KeqZ2NN8dphwPtgV82ljpI5/2KHIwnwhbaBURjPfBYCfjTU/5mQch08nX6E6eG
Ccwm1NdYL5Hjn0XdPQ/5CfBLwExNzo/AIZ7zESNBGVWtSrj+kJ1PJLnwz819cEnFZDCQK7U2css8
2v2vxNyvjroNgWM7xAG3cmxr8X7d+7Tt1EQJD/TVey0oxfNtmRkEr4HxspksbF17Lq7CDppCT/e/
18QwqcTXm3dNYItywSsWns7fmwiKgFCf0CqPaPSDQhLwYobZybAzwdKNfGykcoIILG/OD5bd31i7
y/khrTrG6wND1pOmksvrxPngZ+nw7bfql8iKU8Pd+bcsy4j2DWWVNdZ0O0/1Yj4iEu8PBlJrEG7W
G4fUt2oCcxAX3RsuWXXURkpBKWV8e+8UM/FvRRjgJNYiegqrh0NqMi4wouCSgJxVMap9NmfYUq8h
uNjXFlKowE/4TXJkUok674HzNLRkbXJ80/G2EezsMB+pULPvxD8fXTQvE1ldHPmDdZAYjiRMEwI2
tvTWPcdOfgjOnGM4fPxavqoh6PnVGk30sUVJP7eX7vK3jo/c8g1KSz65BHi13+wzZZevky1uQdLi
Q1XqJ5NIP+/HxkCLyo8MaqSGWkWf7psrzYgPfW0zaVbZF8xV69GSxUiEAPtRt33VO4hGDHFPSgxa
LMkGBgcSfIjaIp6wio0kDmfFZrMbGmHw/9xR+qTJPBqqQ7jB7gYsQT4VOPt3hOdkGkYELIKU2fEF
0SxRtHoBVjYEi8mUqbJIyZ0r1B/8r69bjZg67aEVsiSejFd7DkSVudzrj3zqTp0+ZnYU4I//WqMr
nU6Fchnz4GEvk9bDbl5M1vjq+cyS/SOdKB8eakUA3r5XysdEsHTJg6zePoPHzUntblgNskkohdnv
eYmFLkh9arThY46a3PE3DO7JAJfgavusX1NXDm0xF7QA23A7oFQx0oLlbPZGJ5PFaqenv9Ykkm/X
hNf9U9B5fwTiFmuQplBAS2EXvnHYd/1Ji47xDPeXPj1JUzh74XQBa2dQoi19RGibtupxMHtBE/FD
rTkRBuMmAu96/p8U4RtNDQ8YePoaxIaVNDwSwnpow0Wlq4ucvrrcXSPv6Dp9SLbUuwueyEtL3miq
juNrsu8Z5Nlrx3+NKrRM2H8vWBxuTG2z3SyOZq3wQBqXmhUmkUzvxWmutxubS7LS0tXpkrPDl+Op
yUzVUW+/+0vCtj+lI0qxDeRyBuMjvlqIhkec0mUJkj/Nj3Yn11W1cM+0jCYuUvo+ffOybb9eoiaC
tknoko0EcqLrbFrI0+biGnIVPW8JmOsKMie+MiSKYsowTdo1KY1BAy7+8DD4OloDUzNW1Kn9RA6V
JNYEKd8uvbjZ3aIVGkyOtbHsY9cerJn+5/B3bkqYRrfioWdjmdsXvA9WjuEm18Qpq+n1Z5nV8Lig
IPAGzKmUfzCxRAkoui5fe4fvSvLLUH/UScQ/C9AMnB59kVYqYxauMHXhd2ffd893klgWIcggKto9
8i/JR5pm62u02eMsiOh0mzMG3omp+wwfp/fc+sQ1PkcDa8LepuLSBgtXP5dm3leB3SWIy2/hIerM
48TLZouzj0qjTVROxa5y2FU38dsK55jacf00bGsgyKueLF5OyVuf4JElyGC9O1Uh6Q12jbhE0lGt
PhNhx2vz1NJPZ91OXx1O9SKO5wB68FVVSf5ZI5O3qrRLiZvx8vJIVUBTej5ucQGxvvuJArVqOT+W
y+hRuWKs7cIALtuHjED7M2zy1P0YeKVhHF52q07joGzXwXuL47iqSAjCvnLsqFc5XC9Lq7E7FaEx
I15iv76TDgDOuH6v++H9GRJRz57pKMuKWfJtUBo9uyxWpDYioudj1rUHMYNEzrqWQkqDLNNvEeBq
MzBBapYd98hu9Hi6OB5ujB9FnzcQriKuM622ic3hkQPzoi8EmSHUc0GLKcQIpClOzObqmw8yp1yS
/GwD+5X7vWYX0cjuXhZ+ODuXB9JRuM59M+4vVLZTFQWmWtnefvbQD+0GmSsqu8VxBWkTt3mZDZto
mP7Wv6HIes/veNhUr9nBmmW6ISvFAkfX6kLYz4H3WatxQvuchzRxejJM8F2mnIY/8NnBez6M4Z9+
P+De41mFducV1KY4yUN721QYppU3AUxPw1ncPKDLJElLfQ76eUGpXpj6XZLb6I5s6/pxlOVLjn4e
VCoQy254yuatQqhRKnOiDlbPZAgyse9FpGa4XNputNn5cjzkNnwpPIkkdofUvxVBl8okF8+IjxtK
sf5QDU6/0sBzLeGbw8xBfEjgiymL//RjXo7Yw+3C4AMWcuZQrklarTeuKjTteQGdzbrtcNEzx23S
qtSq+lOJ7Yh3ab3ryfzN2+iDGm3Iw58AhPv1UxwlmpPIRYKjKg11ipcTeTThf0NFTiEYa8yR/qsd
3q9YicHbneMdPiTlKo4cOherXnbwn66WAkUWuwrt4D5mkxZ4IJ0u1vTe7wlLyMAczoGtY4SHR7bQ
srfVDktT6fKXmFbE2lyCp02v9fMFUz0XGj0kpzwpHtZVwylh8Ajlw99tdHCjwaz7e+9GC+FZmzH7
d5uRnMcIHjX1iEug4LUuAraBpxFTI2JuIXP53hYAF/sgmlUjMhvyPkVAw+W+1EG4Zy6KMBT6tTXl
30vpyTFv2GADZJJyUAgcWjqT/9CCyQl7Cppensoj7l09mKuH7I3xLZmqtWQJXilHWGzmkUReEchz
0JaASkyFAgqF+VeoZtbAThFYhWeMikDLS7clWu8pXJlV0l0u8wpeEYMMm5ASPqvT+aEcxgdH0M1S
HrE1msV0RiKHqu9WDlfFlQm/FRFlcLzdX9oaSPYYwVrVg6qCS9rzoMIQfCmwJZJ/wnjT1ibBs3lz
Wm4qSpefeW6mavXUSU6VMumehY3tE61ShZ3zRpG10zTdRI7Du8fYEOeJcyhJmEBqj6QD5M73Y8wb
OAcBT+G7QMsA15HDjdFo5W2/A4QDR/mfJ6HpvrdtLdXLl+IwKDPfVwYpvzLCbwDvEgyjg2A0GP6q
VNo+Q5YHhjsulVjkvn/b+U+pl1mEP7z0cJxgJbLBT0Dydt61LQib8DOolAPJIEs0F4/B9O3IwA4Q
79QhovjWUv6qkBWPOyjwM8KvTKseKfQo5pGHAr69jSIdM/TSS+/GPnZYGKhLx5JhGbyn2MqywB+i
0ECnidDsxdx5s/OdsE09Ld1UHV6vHcNDhOz7DQqei7bOeL9ow1l/R4kiasRhiWdJDPP0GWIMb012
q9PYHiFu43e66/z/6VgsL/UGogW5sHW7BCBwkICPxCzWpw7MEs+/XKigXyf9YgN/OvRqzxfxJafW
dO4hQV/4Bh8Ct/R0Jek98dFCDkKIs4Gd1Zbw2ZlRWNeUXrtov6u6Aqi4phhCxlkDzoau3w4naaLv
/4Q3kQCw4ma6gTEBLL8QBwcpm9tFe5t4ZUNDlTFk2HSYhsWWxRvzbo1l1J0pnBDECfELCuQzToRr
MNOeRv52hJCwWPh0TkiakAx7n5Zpkn7+wULhWVt7VgRZfHpQ8sF8ADKo3tk1PsimR1q5tWVoVmeH
MiSO2BXEeerCz7DVTERdzSqIAAgKXjxNjr/WrDdVAZLjCiRhn4ZPcuyBjaXhzm61jBCdU5Ito8zp
AWOtHZ4xMTCtkI8jnafczb6PTWlxn3TP2zcujqoHK0+GKFy6cgs1qKoSGBZCF5IgzEoqQuGmaGxQ
Rza5ams9CArBLXO27FGxY3AAvU5F82Ic9GEkAFCldqjIIN23ECPgegX/PHZb3ZQtQEZrc3A+djJ9
2onSziX5BHNoavhssfKFjDyTL5sh+6iiduWqSmhLuI0QCgloolEUWf07Jmi0zl0LN/gfC+7/95Xs
gP0LS4QnPJHUy2juiqc59wYeJBGBnURdJ636dUsKCiOPNeyNAWVqxOm15YAODQ8/FuxRpT56ap+7
ElbVIJaIFK99rlSP6ksKa9xRJpjMftYj1Ze9OSj7vc3ToAK7RFj9a1QfjkhdHtIzZ8UzEi4BoSfe
FEaYKZJ2NJC71UyWMY5RNEEECrxbc2MhkHKrQUXdUGA0/A4UuRU4CRVRRR0eVGxpILpJAX2xgVZR
K7F2xTC8B/k8IRBTcyWe0gUrvuedSg+Y5JsC1YbcAxrJ6YGucK/MmQrVAoEhDv/6ha4/DvhM+jyi
dGtFVQqWMJLEvX6IIhJQhoGhdrnN98KaqjSbbx9HDqsC9IDdxynAdZtlyDcXGZfgcaPOLKFuxLUj
anJPasm61iUF1en2mWFyhyGhYbBoDY+xZVE4H8xFr2yFQfkvrzr/XQZ6/8ET3jPZBmxOvU58buc1
rM6bE6jpBMtmG4fxCaMjPVUR4R9GHjjNaoYgxVW5K/MLjrU6ssk5LuX56+5QEFM+Bsfb7aHQZNaq
Tn2WOZ9pkfqlvimQeA9DMB3AOYAkwRSRyiE80UuzQOMjkf2KJi6HH7UOhJdyOKhrH5fO/8pKOn1+
js/hEklXdvVmxZjqp2mahS4h3SJcD2TLEx5AX3KDNrI5nEhve5qIvfvE6Vsykab1IhNjlaOR5yF2
OGtxmEWG5LwNn7Cr7tVnSdnLDeouWdv5VZJnjwqJpfqv9xRHWt9Dfhj+zSqzLP51UmepGhVmj/Sp
+dD5AP/cVoksL95O2rmJnp2680o/efj2pJT/0whwlG4+OQvFAN5X2e7XTq9M3q/2X4ixnOqsK1sW
prBAGuoswWhXn72w2q+lQ83YwUdv9AS+HRFt9yCZK2Ne0IjPODZQ8kprxHorQHQLGPyV+3jBfXJG
uzQ2dk1LJ8amp0xl/hXpvSPjbKfBmNGvRTFKI5Z5YAQsBgQTWSYWFiUR+dR09LC2VS+jR/XXL20m
FHcoUjcpgxwTG5fR4wR7MCBevQw5fYuWit77w16UgLWjutPWsIzlIhfhU0so9yb2gOOsEH7r5frj
+t4Xz/ssjg9UdhAW1h/mt6tPDEEtdCLHJ7fElAaItgcwqKJfzqOIxq2lRa0V8iPXMbnLwcdzwkgV
2Ndw5K0OUWZXxzZdxjS7C/cSKThmoaZuamBBdpSc9SVxH6BIspdW6FYSrWjROs8uik5Yak62Oxfb
Ntu5eFoQINKC5Bvvrml3/XjVeWd+HpLPpSwQ4qoXKD15sSfJaNlKZ8eFCKUnM7BTo6vqlWdBgXad
5he2SX29Nr+/awQeqe0f8xW8FRxgXwaXbyt5lYhlMflX7eWV8mzZap4ljXFmi/IBSKkKU7rsEK7O
e+dioDXgzNcl1xmtpCKLVa3OTmPbT1Xvj3q6megmcPKm0Lx8Ri/9bD2CRagcOQsZr3Txk+zjZ0eu
5AOetbp28ijA/QbKnyA+7dYZlpboh5Lc5+TZars0vgbQn94lgbOJXafxUUlaVUaOWJcg3xKXCfLn
H1Xb0Ze//qD1uElTA5n7xUaKtM2VDSJDtS/5luJvXo8mg9Qv6dzv9344e7QxqxQcP2JZIxGTQ8v+
B7YeS1mD7xjAS4cabXprdnsizTh1RyWGLWX21u05XA1UNpWxcPaJMYoUD9WVtcp30uRXENxHB5xt
bZ9Z3vJqybju+n+9av/CzvQDNxyqXKL2YuJoSbyH46A/Ip6nFCnNwKTibZNOfXWzlueRWLwnclCF
t3u4hVesJPgN3lvoof3W18xoxkRlOb+abMkH8Dl+pf0QS10JTy0RHwNYaSdMfRfGQzA7km10hLwV
1L1DI+4faOShr9i41W+VK7Q0nTDiSkefiQdtqg1yKRyXxECFWbRPdrxGx666QqzIy/h5pZNievNi
nDYPsxtX/PdHULsbdnIWRVnFx0Ctfp29T2RcINzqmdZBIn7jtjoQcZM2tgAhBI2+UDiNq3Cz6MRh
Fv4l3DZujQ5n1pFFdTPTdnkvoMedVAT7NHWZRL6PHcJiUtOG/HdHcMRVJHSF3yGQve/r3vUTm5r/
4L5ITRDSqWBjX9+XRgOevp4M7hIxLpm4xPr1QhT1QdYvB6izFaifYTDXh6d/WCTKWqDZQFnAM4Tg
tOBQJ0j6LCEP5mBvhdSqpN87H8A4i0TWXEZOUvjtBGjLL03EFsClCgqYmSLim2IRmRHIox37g/JS
zqwZFjQuCE7L/RsS129b0VV5mVCIXK5nU7QRoA49BrnENLI3jLrW3Tr9HGnyf4m/OxH0HgRGrqWF
2Y9oSjHAxMfao08w1t0DoKr4Flvrnesa0V2JSt/Hwklnk6jEU1jPenL7ZB/ladJIW+0Wl0Fb7fkT
wQi7nXKPLfIYFv7netiCPWTYZ4kp0G0YK/FmZLUgmxv3SfIqGTjD4GK64KxA0P463Lx0XYAy0CjM
wWfLINuNiTbsF8xWiM2kWoqcWrmnvO3G2KOH+40d+jAU6VLuBJ92dCxGEXoleDz6UCk9aw74lNg0
N7ubU03ONQmuoFIVD20/n5RCxN0+f0Eafar0BQKsYpvWLDFFonoUH9mgVYbSJt8O0R4hnrmaUcBJ
6oYEoo4ctDJZsjKgmJsGt/SGHm9W0Lh18Xk91biMfisj3r2jSh5G/EpYdttb7igQMvpAaRA9YxWi
UEmgPLZ6GUtJMbH0An2/QmO7paC73hD7teGEjyj1ASEilOzmyyOOI6NGm/oCD1+825jbH7SbPZiA
RCHnhSnKOSr+mY25Zd8HILxYpr332NK1qdOw+LoV4rI3nBQy6Ut9RkpqEFltQLgJJzFBvlMVUhQZ
iS10Uzbo55WJMzVRnPXfb0GuWaf4ts8zk/CgIz6a6rdBE3L8PzKdMgoHHzKzJA+ct0CGO9lehjej
kMjbWp7i99Xv0VrA6Kt7twjHcAFDyIjTwNiM6gnUKDjYrr3cdmYo3V3bbpHGwqMKnxH4R5BA577e
pBHynPsC7hcA6Zlv944raEzgF92IMn9hXwTm/rwbcezLYeD0cVAbTNudt2w/LGcJnYY3yZb1hqEX
11T2GVlnQi1btbvIj2smMf45qkqGk0u1iz7v6BCdG6wXS7kTC2hIKMHD5qgvAX22IdFGjnCklBrO
j2ceiyFsdLtn+pFwldQsLUOfG/rHkrfOZuKek4hUpt+oARSMZUQ4uk7UvW5NJYlD0Alm9Qq4mD1s
2tpuzP9njwOcvJSr3Y8OE0YZIqiC08s6qSEyptRxySALbydvBnXDVE4/2JsAVdVWRWIWl3Z6N+0o
TJvNmUlK6e0fgKt4Z4XSagZ54gPqVuiF8j9T9JpxQrypz+vIfd9HHVFK99ojOMFlyNCzLJ3EjvlE
xWvOVtB4Mpertr4zJfzKn1EynYCFbccQj4oUpIDAg/YKmiIlHdqfDHoST1SuhC1ELAARKIMoIgFQ
DX5CxS/S6UFaeHK2dxKDMqfm2Zy1L52NYq8xkxSNc6m0AIvvPHaIab7pL0bRoomSA/OvBcOElYv9
e9YX5UhU0tnglVIH7k5UORNxWu7Ff78GvlE2loA5cagGtndhzCCtvKunSY4KvrIS7qyRAXUyIV/S
SkFVSWai13i1RnqxZ6Vz7trjnj/a7UWio+A83wuRpSoSgwthgSQkQlIRZtFzXCWC+5UpMYyIvlDl
lgbxMqsnQL62QefeEI3mza9W7hIem2gTafUdrBeBGluBjozldnCP9dLhsiSzOjqDxz0A/30RQRq4
evY5TLAB0M9xltmtPaRmRw8L1mkWH2V2oywo7cgMbWTz/D4GunTajz3AH3X6FtXhpAEkdBoO0bYi
yk5OLRF0jQEvR8RWo+T0m6FrsV3E7O/B2GNYHkauDjNHWPASjawceUT+8TirKzt1y+Syl+L+YNan
fjDiM997W73NvRXHdjRjcUbhx1TrCxiWVlaiI0o4LaolQE8+lwE7yC05qYUAsfPCSc95/Mt6Govi
FnxSwXE9rGDeXBFDPFpEWYQRxw4hCytuYKhXe7w85HE9WWtzYZxv7LAblhJ/exmcfiw7xVvMbqZD
f5RNREZm2jYnphU63wCHYBWM69B6b46LDgR5X4ZWX1K0NNEEOEEs6VjJwulVVCZahNfwjjewDskH
vP02gvmrOK2Rajg2T8h6A7tDjlQnrZFuNc3DA2pypAAIiddEI/fXU0CDNOT0Lj9B+VE/xvw32gd1
LxOC+W5Tcpzz/HWBwZ4bRIySyMg8rKdmO8MuVbTEqlqPZiJ/2rmjddNCBW8xi68yvzNaldZYYBpZ
N95xehnBY7JCO8PFDPhZYkgH2m9CtORR8bjzpODkb6iURHai8gfZJMTrIDZesz+rU7iXwR50jv6N
1sqAnq0UrXpVqjYQgetSFh/qJyJ7N9l5cvcp6uoI6dxjWE9fubcJS8v6EI9sXveSybbg2KDUNhQ5
uQZgIAGW79pQ5MEstKE1f6l2jJ65Qaom5VuTCW4Ugum/yiAPEw3r1+TDhsBIFsqODFcvEplSGy1S
Ced3cDdaRvHZEf5Z77zGX+SxTfT+93UHXg90vRa6NBwoC4bQD8K/jXu/GGqvVfCW1NRzMpREb0dd
S+SobIGUqPwbpKVtZYsffKIqwpEbL0WXEWziZ6GB+Mlrckrb1ho1GpdVbSKouPobYleLQn019jEa
wOw4Octc+MwjrCudYoAlwCatCvKM8jybzHvcSZ17si9v98Bq7YqBGkremmK1vLhsOFp3EWn+KFdt
H3Dz5AicvKNAN56CVBNQ6TZHLHwBWXGStVkwE+fn0xcsxRpBvGxWVmtmefKeKtBiwDDp+ioGFaJb
Fj8/bMjw5ZWZMvjUlKI93jNKQbeU/oa2rsUszrn+hITumMkh8/79O8ID+zWnzBg8i0XKn9eledze
hEk0rpYhSRm9p5ODOMOELqee+yELizETZZi2XbNzLzVehmr01qwSq2gDfBNmQiXOu33GlPJxUhoH
4enIvfjUxeY2azNDClu2cxIb5VrSr/MID/gvEbn623aCO50ZjoXHKPx8JCYwnWDd1sgfNWJrbbMr
fkOF8jhiKCJ0QsYL9fOEJ90LHdDL1Uv83UbnnFgwlOLiS8Sp2Wasup3YXTa0JFFn1drdKmk1cJGB
GinJi5ttqXqV9cefxClktwQ7Ux0ywWOwhYxjelh8kj3O7Q8Kb7E0yiahMSVMQAagzoLoCyCNlVRy
1FN6g/2Rv/7SbNzU8+asDYMUzd5rIBwHF45fu/TGTIxCWlv782hr0KmmJ2u7fApvEx9jovhqWmPh
EmD/qM6XyAv0mKdv5OoyeK+sMLqvZipbn0sTVQG4TvBae8x2thpkH57y7hNf+/WRfhkNIzCTW0fJ
V6vgaGpr8vROmHvixCrHUw3jeh97nk0iNUcSCAccaOYPHLhBj3d6OSuWLhKcuiPoAKB7qamXa8Q1
CC3HCIsUYZYD0oxfUjnMuDnl6dvY/IWzFJEXLWDDH7imjP5B64f9Zg2Hx3hJyOY8dZMxeE+uDrgr
VhRshl+Qs+oeuf8/K7S93LGhVWXfWY4U/VMy4GRH307n9zEQSkvKxa62Hjj8opmmpbmGp+Ysmvdh
gtVm8VA326qrBlycLVj7NUSns8ZpzpklYKiBXncRyajheRoLTPZNGFrQ2jYCFnDWPhKDUQ3LhUdX
MaOogdmuQIZi7+A2XE3JNoefUJbkMV67IE0619sdUbBizj1f/48fYl4uMzS0looq4+SB42G6h1Z/
Pv7Uff8RWeAYiuSoNraYe5pueiNuWfwwsvhjOvm8amMEGbr8hOKgeNKKjltSK02E+OfsoyH2tOdb
GITeuHfoOtaHCgcH/I6K5nF69dazJbZYYXpU43XCy7twkRSO6B05KcN1/TUROp1+0WTkDOfZXXGE
dzqgzi5XlyRhhZ9GuSEP9pRe3Vcy4lR9mpxiiS3Jn13U6Lu/tVgPRfv/wzO4p/KGfInMpJ4geUAq
/bGhxz0TApoPjTEhsSAxYPcTUz9E+k1LoTuwz1rR0Bmb0qr5P/8UylmHbmLbMYLmOF67ZgOHZFiI
FpZy4BnVwj0SvDi5fBiYVCQy1luRKjYyVSDCjuH0wpW9VP/gEJ1gTUBPxUydkx0g2kg4AwL5KzWJ
tUtoK0Hz9sV+suhakFB6AHHIiKSRku7qLKjd99CPyGP2tSSuIhR7KvqSLpJR/90RDre5euap6uFx
mVstc3mkOvEpYDmcYqDGcerAEkHa+2FTL17sZmORu3efRrF4ULg2sugj5yVCQtU2UZyIA6zAxcAQ
z/x3hYX1USRmb8YcWwYrpne+ya5I3jh2L8wtUI0GpKKBWcTUzJnJPUg8RnNGt64bAxRKgBklzb/r
1cbs7biMsMB3kSKZ47UbC2Ym1UKJhzeZKKGV3pPsIOizkKF00lPb/zqGTDet5W6QY2PpZrO7++re
IU/9xDVG8JZylSWbtlMi5DFKiZ+6/+m0dQ0tl0SVFieQGwiJ1Obceh4CsKpA4Vo7OFC5P1QMi61q
fraQerTKiHUyLPIYXfm+ycEzpyirZ7oOQMQMBzOCYBiESrXAqDUMfxH5nzEm0bupvfrsplNYLJKf
McnrzEmeTyafI4iNUR27qNm3Y4y5xNKSgUQmibnEFEE0xvJQ47epG82NHNXy17lNer80Q73RSKjQ
iIntfNumQrmTzj+qHEq7UxaxQLMmP6V724ZfIRAujfn4Q7sSJwRhl+Wo4K8kT/73i5RhtDMBQMW8
p2u3aKXpYIu2V3R6yT7XpO2ioyYHMKXYk7aBV3v8E67xDk3EQaQcmkS+ruXM9pb7h5JeKq7lh27D
bPWmSSSmjF9RB5ET5CJz2OYuMsacqFgYS19K62Qog638lfK/Y/xJaLaminL9Cl0pyS5DOIJk/rQZ
/wyQCK/JmPSOeycHX7aI7ohZOfCB4Q4vS//cXwWPrrIhQWcucB5EtuqgjbLSzC0Cmnv7dpUS64BF
cau5UCxUrbvaYF4phMl9F9GLU/+mibUKh3qD+/5W20JJCKNAFezGPqKhC45213RM6OgD4ithnAz5
2TepN7s1GAvvtEkeworislWioeQAX9jZGgybCHVKO6NCXf43MTKQE6fRe/+YhtWDonWASaohlHXy
oQQ8Ww563jMPZEgbQESunYjqacywHMou/sx8W0rqbnVeMQll4hlYMglEQKi63xeMZq+YPE0A55b1
p/X0hVvlHJnZQNAVzoCXz7ZhVd01auF/BAxAurrpTdp9Qr8isKjiYJMqjmwRdH3ufqoOEbmxM16g
LNGrQ4qxOtQuLuK42Fevy5duC8WGi97+FHFHfag+W41gJlSWZL345mt+uIVK1OPIwVIBgSqPbHdn
OSIGN+0Tb4whT0Mz3RlHOsY4NW4+ivWVH/Tb6p/iaZDZeVw71C08bfL6PlGG+4eBEdqGQS0zY6hS
z1p7j+p0BLMKW4uWji6D8WVVa2eQ2aI9Y5aPz/6iUYJvzUa00Sod2nfIVP/+ZTMQ5yA1r60Y4xl7
jv0w8MgI2DEEzM6E8ApsMckYOHaQluN4MNkc8NJ8tmTSygOGxpWSYbm8fZOjdYHEJ6/d1oknP767
lXIaKLSwmyi6Gm41eowDTySY+DI1ZJcAKH5ttMn53N+0r2Zf61pQ0mW/hUpSERY0EwKZbEf8CqJ3
CWIrAfX5dAP879/4j9lxE6YB6so0jGeloGyodri7GX9uCcLs9My3tiNvlzWW3AAishX5X0RD26PN
g/hFlQI/+p2+HB1v1YVv1xieDUMU/ulT0em2/U0Ze/W6f4KGu5XpncIM6Bpsk3Yqmx5gYaogfwTG
iOTLu2SeXk58ExiUgVdgkp3WFhvE4N4Z9ujBQWLoZi4eavvHGIfbHXsjRV6QxGYl3VjL2Bmz/R2r
T8iKDZ1noDJRzWnrqTL/VXzqmeD+qo6TCaBP9S2qBHfb/CQFG/QCM25a2Wig9hz+J3qllpIvI5FB
xZDTgpXFZKKlenq9LZgCc7GjDwYpCTj7+ezSwpEmJvE64RyBh+dlHYuO14UCUR9HSJYNZPpxPMd5
TjYWLvBHjpkvKMca2ewKU3bExdWefXjTocO0gartv90dHkvsucrDzwsGNBYN6qgmqIhGjThwlU56
tT6xxRRxz8uWIN1Vi37AOwsmzwmAT2G2FU34PJI9tUjccKdp6UUX/jHpa/OUXdPQ4P2pwgNj8H6x
XUbxpSDEeTwE3ImBAEgSC7TTMKAW43GXLXfLZcv++DGs2iZnlvdF8XMcPLBkyjNOa+4CzfDSC5rp
SyUbAjerrWJ0OhGRSfiFhDNHxwR9n9r+zRw8P57/rEq8yA+XOa+QNmccmjc5IrzMselvd/BkhSJs
RgSanY+b5Fws7lPXPZiI1LuieXIwYdJta8LLNnyB9LkVfHN0gYIPeDoIteW9axKHHqi1VMdXhu5W
ykPHtUx7mL1Ee53f2Wp5wytx4nKkPah1+/McaZXvoglvXOIdMxPnT6d84NaxvJPEZeQ6ALrQuGMW
HuDjXg2Hfg9dRuA/YqhePSGf+428aKcuMCtsMRihr3Wx2G3BEly43Dd0rAbjObxOK5ZNPhGuLv7x
TB4CoIjhQCnl5RblAytPk0+roZGKu1AZ7oPfU1GgEgUuO5H8Lfu0qr4EZogVrZfyPaiFHHAeb6n6
kJrONov4Hj8ic/1tLXA1fqzE7SDmGFcJsLXHNLbN/GiVu8eqwJFwMUfEDziRczq+w1heJfisZrf5
v+VBK4CQSvDERD6UifM7CkpHZm52MPUuxv51bUvyi6P2drkJs2xoHVWgz65cfoLVnYhizwr8T7zw
K8389zYFzEaZOhXfKBQ0YE797/pZJ2y9AEqK3la5IPydNsQWOJoIDo6Lyoyehjv3EjSArf5Z//Tl
Bt+RXfyP07SyP4a1gUuGSimd7bpFEZJbinJ9uFYO7dlks7BuABE2X1e9uUcOAYHN3b7uJVlK4T1o
JXFIRzs417G3xRJmOajPLG0k/ai8yzhhsEhHvKDLtptD9vlhjdtNwCFrh2Viy+ACsUDRGT+TOgEz
UINDwzjTTyE0+kBEdkLEZmlTi3zmktgMRcWHDAWf88otMWMqcySrL0vuzmqXEXLSTuU2xOUzKGXq
lPoaTwekWHBHmA0Jk0paPYteRgRY2oXOHBqAbGQhDIOeidP3KjCYTmzWl9WmaLQwr4s3y69pw6cK
kCPOGjBL2OU8atlxBnuPNXM1UdRV/4KZnDbTSIIUW1wKY3gDK/SweC3AVeohOYW4o8Jr3l9YUSb0
nTxB/1rBmuzfFoUSYwAozl/XaaSC5D4eau1ZEOQkb4NMz5c9Yw5UXrgkkiKvo/89DVmGHJUjs4m0
vSULYbnRHglWpxms5pnDRyo0sL5euRVvVErK/Brnass2P5zxm5rLkiSMI67RHBbIn+LxR5vXG//6
byL0YnPwym+VceQ47zWG1jR6lVMAvOr+aToM5ErM1pGNhBfzZHOWNdr+uQ79Ff//Yi+gLK/N3wn9
4GWr6bEEgbjwTkABYmR6/ffj3VcVvoOfxPtuqA+84jVxt0J/D5gqNRUDiXjDwLbumoK+utE2BZ6c
0DodfXJNDUJSF8MCyxChoo/RjoYPCTjP7MOjpc7OQE25g0flNl6ZrxATuKEFH9ThHUX3FdHdneIx
Nf5mqFUuIEhSs0KnsvGLKxLXZPO3LzdplG8pkbSOqexBG99lyXANvRlpiNTUuY+Fbgiz+IUw9TWP
1eBAWJjzIokaYrMsPLlGgV1Lg1dgLZA3wImcLXcaRfzX9BQ+ay/gY0Fazt8FK7qp7qWZW41O+hJ1
sc3tc6BEEeCXZXkbkexC4U1Z8NgT1IMgynUj/cTyjjUbnBsDvcmk1SpaUl3sT6qg54klbXgibyuc
ClylsbGGeJQhdMqUWGtnCTvPdikfXnv/7V1evHyyYafStJtplCVRekTuTMuzMGLWRICWrI1C+2Bd
McawcrmcD6590TMssqfMJiuH6fM49DKOG5QOQ8hkTtvUv7TS7Cf3wSXnuQOoYqfO3YAo9P6MuCn7
T4OM0mTwpefJHryTQSehs8C6Tuc5P9aaCKyuqSYOGkPfYHyTkicMYL/gB9oMmGTHwZ5K9r/Lq3y0
TZIp0yjnHPWsg8YZNm912NzPE2EUrbT4tDrX6MGOBGfqbyjHsckht4hS5QXCSFN8sWdZw0yShbu7
NvVQaWdIeoZ2nWnWQ9WSHoOQWq2c/jdrnmA3dZgPI4lh5Z5n2SioiEtk9EjwrWB7CzRPOwBP7cKz
8KV6FK0XWXkdobZyyIoVKssxOVM9CwOYDhOYyu+2xnndT6zSLbn1/FM65RzBbBXHepz1rXWyvK7E
i9zryiIqrWtjxFMiHpRVFQlUqIUS857PsxeAQMODBMY+GlbqxM8UrBGQCoPYrpEkA8TxTlgP6H0C
MumG6WZEQ3pTMlDa5n7HYdkFy1dzM8JLa94xhmZrC5l+Pu6ene541LRNCaSzvN0BQqJ18p3nFnvM
RhA82Oxs66nlst0QoRHP6DAz+2coFV5Eodl5ninClOnLAJG0qPcRy0HoEeT3i2oRAbrEkrKPKxJg
SyGFMwOCjXKQO57oG/JRBUwm8vebdyHAf8ka9KGka2nCttA+bi8n1cen8Brb/cbrbfPBFIAfim8/
sgl7XaEGRHza863e6jnbbkUc0vZRBQZHck5VMe9G+bWufmjW7KvNQOXtFhsZ+GgvspZYEPdtYSfh
7S4azmUK2X/F0AyS88/RWtDZbUkAzMm8U0ksFywyfhtf9sOKVMASVF42g3Sc2MaL/mTGhT5dO2oR
Hg6q8xfacQjQj1KKPDNf0BjUzaJ0hxVtYMynhqjimoIYVNZAnTCg65xsRgwHVGs8UyV3aglNPSFh
J8W/v8Stqd4cMjoYC3j7ckOqjaYrcHBUfK0FbxwNgBJ4TbodfZbYgT0x8SbnrKIBolSTUv1a9AK7
amKBeo8P83PcU2SGVCQMdFXz6wztiDKjgnoJtvd47uEdT6ppap9v181Zy644D2g3NTDnGAbgRNtN
BjiTryDh+JlXZmjr22lxzpM7BRPJt+ejdquNFR/UGsMGDi57XORpBm7DeHL6/CvfYNPg/dAnwNnO
T+2EslPFmwvZk317/o8yJGAAf+H7G5x9Bvxqc08650TfBttCiWu/WPxBM2JZMQ2N04BF+jXO2QCk
M6vYkJAwUWbtu5H/7IqZEEMHFksLTKBu93xbpM6AKCefr4c8DrVwAvfFfv1WX9N89wr6vYOUOytI
guqerErZPMj1k/uvzI5VstvTUdsNKkE8cpnIvFdaeFjofCT2AeDbcBPuzzIPKzO+3GPv26UZvdHC
N9Ar4edkKgf1StbTVU4Pnb/4ef/XRa63b2wVLP5NCmZILQNE+Y3TSAMj1qTKOBDFmnTaoP6UcVC4
fMjFAHu3WT06LalPnK3YzUSs1qrkF/PzYq/Y+wus//P64MpUXXeWOK3M0DEK8F6Bwdr/7vnxBY/W
Yq485t5DGyYHlxl3cSLJCN4NZH6lJ6tRFSN9xKg0Tvd31c5zHZ8wg1i80EEwKUAUzC/PISeFT38h
zWHw+jUPMYMMCerhf8auiHRal8yCfycbhFKWRrymgZO3CXIpUuRQ4bqbV4AKf6mxkS3gOGeqtEAs
WIIQvEHlnAkIlA/5rplUIjxPkL3zQlFtkbNyuSwLPJNAkORvsqjylHt3Cw64kKEQtyNjQ/bFxjoV
clb6lHEykPKDar7gO0MhqH2lVpanfZP8HQt40Q1G9J2V86A13eQNbob6LuXv+1My31gXIgHohH+q
KGIG0XeI+kE+gBZSiKfCpMUbwb63IalreJQyvgXdUKhV45yr+CYsOV+Qq13fTQcFam+JxTl6U35+
sS69+5Ys2p0Jnj7UzrIHzvHSSNu6mhNPzNcH6qS2EOZQ/zk8SUXmaI+FuBFzpKvEnrjnAVryt4h5
7O5iwgPmtKkHwd0oTgbaaXwPKu6RXtQI3kzopPxl+WCQQppAJh1FqR9gFQ1Iq+LN8z3gQKRl4Sfg
xwYx38zUpfv5CfVjx829SYhNCGUHfqgb6/mLv7Ez0Uf1IkQ+cNC7gP90XapO2CEtNkwFTOl+FGZk
MmkpAtNl4WpJg4CfMaAWVtAg5OmaHXW7fJbcvuPaxkO9q79r0NHNT5yNuVuRwHQ/BdPVBMqVvRUT
RYXFU5pFAUP8DQ/01WZHvF/umcJiwKfGbsLcdXh72xN5EpBc7Sbc+EA0I0W1aWrg5MeIS2B9Ir5N
MWjgBeXp8DIfj744G5Jux8bKuOKUUN9xJqLRcBX+pLVdlguy30GUBz9g8+GQOMqglDry5qaDR0KA
wMX53v2R4u7wyDQBe2O91OxGykc3VfktkWLPVXBjy7pEBO58paKgEqmtLG5SwXAeN56DHeZEzP6d
snnZIqZkpn60MZ2CxeEuIoGEPUSBQPfboaxz2n5KriUn5IFKjgFSMjJXumLo9TXQt1oUcTfJ3sQO
D3gOnlKtyoLXtcxroEBv6/SbQXftkB/1s9ayBF5XUkQtM5pkQU6M/Pl0suvGt2j5j27GLd9THR7M
zLH2h6ZAn+TwTUMY7+8JMA5/vUz+3gnyUVRb5S8kOTUq9qbT1MACT+YF+wJE1ffkQk3c0RuCbL0e
+zvzJl9+Ug8mMwjADtyAVbBru9vQschWU75w1WSU5HhNraWP40Cz5pz8uuVXRMDuygvgRDAdQ/3i
Oe2gXsTPJemwq3/qWdMxepPIh6WtTPVTGLdtGCJaNaIvigzjku5nYA5ZWtGqXIcnycj8Z/mUBLG9
VmEcYrjCKye1vMDxTWzdnMlihPpf/gGlU650Jutx65gPFig6xk2NZdvfsfsnL+ot83XLAXxXG22O
idw3jZ7A93hBBJuvxpSD8qbuFMdP9sXMJ1cMPHeIhvPnfsMfSxTxRgMNkboUYddyOejcZmD2gq7M
9yblVTPDDxKyU3vfL0H3fh/Go8JdrRWKJV2sppv5atVesQglKMSJcyswoPnVsoEMSV6k2Y8cIor/
INtDoFC2G0wuZHHY+y+cW4WXlm2mILGz7frR9c9xRScN20YFy1EXDvFLSnGuxc/y4OEAgHV2iWwe
EWWRC6bWxIIXJERYhORKp8jTkgAE3v4pVL6ZXfgp2/y/GsmncKfSuYp2HYhDYxt6iXKTd2XnI9oZ
5DEChd4QrDHKXiTd+e/fqJmnKmgh6mAzunViWN7Sn6s2JMn/De12Va8JgRixkMa+8MwABKlJDxji
sH2oX9MrINX1ix61C/2of7yWFrccqwa4Gf1jaivYPj2zGy58riRtHhoZtCPJWaW+i3PAx6jZKblq
R18RpejYu+TRbjiFLubNukiwMjvvHLXrXDzGeimEow02SRdOE4NINNoD+dt8DiBkImAT4SFUWMBo
P8Kj94qpleQ78q5TrHiDqmnBKtCoAaoLpX+md8r0mwIHY7ym5JTPQi1e0Ci/xyM92/fboKG0EOTh
sPVtOkkLTdWghGnGUofr4mcHCrgGin50ffImcSg7VBtkotl8OVKT8O/2ns8ZfiLbypOxA/dTerMY
cHeGnr29/LjcVeHyCee+8SqaWkh199af11cr7EA0YuIU7chkGdmgviLyqZk2/VG3JwEYsK9/m2n5
CcEM2F+Ju9IR8lyJTW9yaWtRwrRYc+WI8yXHw16dUpLSfxiB8Id9jt/NU8VmtXeiyxrECzZyvv9E
u/35chhYeavMbAw+LOB4dhsRmRQ+ekRRZQQQN6yxNAkEGtS3BxZxK5SeI7dMlJo/nmC1IR2ofPG2
vP3ZMwSgoKZdYFsgY85TAFkUypDXCR91uP9KU2yQOaZxXiAjhdehlrbBVw1xmLJB2alIzwUDn3ZS
VqtpWz/SA6nOUiqCZ7IhffFhOjZV7ZpQJInUd2EOtOD+3nf/+ABjxIFLnWKRApBFWRmi5OMIgzXU
NEc+sY62lCC5fPU1mhdB3fMr/aY3v1YqlvoLqdQ4jdNg7SPN4DMVeKWYq5aqZkH66ctx6BAtn9fp
qtxk+JPmwKgNAvHBMdtu+mlbjXBZQ3fLpgSb5NHMRrQrRO0RzrDRwRAy4yPfafpmAGXcw4/ER2ND
RcgWY/yTolgJ9XOAg8/2dgNDX28YbjFn+u7kByYNfcPIHXG7q2J6gF9wTQU3fhWuebS0r6R7cfWv
UzBgfYEk+fLix1EMYFj45OdNOdAjI2fpBnGu0T1vR/9lSOuyinu4ag9MTX5QgQGGBFY1QtMBbqjm
m9JNbR43FvSANhHCSXTL0kVlbkXFNegPu3Jbp6/SHodtG7BMtvuf2EZdf82AMu+R7J0yYMPGVH00
B7vemJCjWPfzca0ImUK5w8Zw6FOxJbFatb+n8ELyGysqo35sQOmhACZ1GL6ZPATK8Txt3adLc7ae
FsE++ZaQZQhJxN/aQ1cXWN5uHsHt/uwxBgQsX/ks5QtxhHUpd736l1RgT0SdEhV9Fp32gTqPlwTd
FCX8E78t3Um0wpltw7/xsR/HZ8+Vlh6elgzG+lCBAA2IO+j3CJ+mXQk5KZoNg1WFeu3UKqWUSGH5
qT8USulaILYeXwDeCAxYm5GxVoaiB70oZKiotb67Lq522f6xKrRcmWmYsoot86+PlMc0Ij/D0gT6
mbyIUe2ZTQl16nt3v9VGArl+ZPCM1xlcoGDugTH2XsTtgiMs5dUIYi/dQrUAFSXzA0PgwpaYwiLH
nvZGKLc7fryt6YGHcQdEM+lp9T07Myoyz/1ruypKQfV6bVSCsA6ZPwRXxKzYFXsdKgtG5ePQjULX
5CsK91dTC4/ARvt2inMJowOiummhHIg2bFuVFSw/wKnGpBGMltpF/lP16La56Aa9reBcj7nzuV7V
M9vzVoUC3jlLM5eACym2sd7lk5/Fzz9yrqmMNWphh4VXCIqzKniOhHQdlW0n5RVeSQ3/m3QVs1lB
7DFkcornog+XN52Lc0B85m9u4kYUryXSeDZJivWVKstTTI9ESjBhZS21vzCAFDS4lEh99qA76c9Y
kWW8nztXCfaSiHOseL9jGPWY3gS71autuWAJ+T33GplQtzTi73JR7v7mLgyiWVl6PErSJw1Ej/vs
QqW2sMseQsvPzYOhJlEpwvQC3+4Csm0UYzP3xZT15Xt9tq3Nk4FoWwqccDtXBrke9SC72j+CiKOS
o6jVwvq3JAdkN/p2reoYkFX4T51MIyLaIBG8XJAQ71LIPAjoOQIiYLj86d4iQjUSQFaCCVlw08I9
TpWl7MuNdzBNuP3W6Pu+hsNCzHkA9sZEROuz/pcy+paiY9YHmiCMBzm5QvNljVlevLsk0jopamQr
xIqXKD7mhTd7tDCnYYmsO73XL/q8+qD7ETHzT5rmG02C2x8Je/kxC7f5U1/PV6e8VfAhB0b5qhxS
GBW5PxWcstqet0JsV0LYhWwyOAQ3LCgK/xV7QfTYkcML4/2Ca5iQia+LsRv/BTSowQFphCyPIFTG
5LJGKcLEBiAP41cXwwJUWLwpAcZfMwbIwkauMUkT3j/47uDOFr0Kc4My4R9st3a0pcBLKLhKHDz2
0OZo+jI/feEM6eCTl0ktSft4YDQ2gurfyQhmF0IaHL8s9/1QoKjGUeP9w4PV28g38wYnLjEHeL90
IPBUN7F+Y6BiVFeNBTUi/8kXxUWxiygt4xs/DJRsj2r/TOEODZj0N4Ol6pymfUp5Ss42FJRNbMHs
DBJv7+QKhlRZoLCPFJBlbLppCXL8cmle1qy+JlupU4ZYO1ZFLaV/oOvh9FQm/1n/PARDYfZxIISF
WcMnnMkvY0nSEU/mGMJDbAyhu80b1PNlb9ugQ5HEv7ZsCInCzO1qvqnZc/YSkXS1c/36k5elo9tM
MKdCXkTE6GCtaeZ6JJlmk4Hw2EBgToncs/RQeiay+b5j+7k/ioFXFm9pkm9w0/Dg4zzd61C91/VT
iIOotB9ZLmawJGttNsfWYrBN/tGuo4l646mVfPBWgcwHeL0mb53E6YqjHSAvQuzcwI7pTZSC4sEg
1jLL0WWS4kHXwrTCORYxm+xAzZnmkdIwGR2bmuRQQbyQDRTaYcfYRe4g9wEW0tFPY5M8E0rn75O4
VYJdg+U0cMP5aWv9yigANEpc6lgUq4rYeZQ15d1bXLfGKhS1jKdlGWPiW6fbpxZ1t55IQGq9Tbji
NMHcpynKf3aC9+9jlxnYPu5XuRh4BG/GN8+trEMEw2Gfbzjswn2pmu5um7/1uPMY6sV6rruDj3Cd
sQrHhnr1jx2eR9X5iJ5eVjLpts1Pvm7BZxhphqL//ulhUraxduVRypy/pBCcTC8LjkPlWPF7oClg
Lg7ELlXenf1lTJo7FLYEDo4AT/rXBrrNJomQWNG7n6uc9rdbZolwh4ZDxkK24vkvvIEvTPQQW2lN
2mtnUQmwF0Q7L6kQ/T7DQAHyVCmrw9y/iLq2DMHWDTCU80XrrfJP3LchkpMl7lU2eCeUdz8zZMLy
lUoLxIekiibyYFshG5924bswYVnmcpY2kDgsAJlZYiXNQgg0NIqmzPnwCwdYCRREB8xEYCEpBISG
cSj7Pe6R5sXofHmNuCKal6dir0PsZTpqI0KLCVcKj5ObnoPvK0JDkHfGlDOb3ZvDBgiqCKbQ5uwu
OfmU/b0gzDX95itFtU9WvSlY6q4MW6FOul0+G6TsssjhQ10BlsV/bPY5aM8QSw7ABKpLU0SuFVJJ
KkdT6RypAo76CKQ3VW5jySmwpkUczJYNyEBgyOKCmsFe0Ds6WNP9cSqI6I3MzMggRV4ZYGvMcSIx
TlKMxmBeLNRXpXTcdCeJaMCgacHVZanN1lr3q1eanFyj2BvunKRd4aAMMRRUD4cy/x8Hu56XZoGs
peDVs5d5rO2n0S3FgzbbeucOQfxW+/0T8fXKI8gY0a+ZRqNpzhM74mtnXOjQg+DHztwDls9wEQLC
spJlSW+jShATO5KulW6iTeslt28ACyfuQndc+wNwkfchnwyMMI073ZMabiUgT5T0iJ+MMuTQGlp7
ygRC5RxkIqHt62lcdw+kZsqGFoLnD6nAQasQPo9YOHW1rOytAuYmuXfiAB6nXjm5j8InqCFSnl3y
8LrigtaNWs+CCowXXG99dl4ho9KQRy1uY5sTG24jwdys3rl5gD6AjnTVmmidrWVDWpH7HHb+YODc
SO1HJcc26CI5uUPUVUX2Mz/yjKKIZxxkOYT+X3Y/K4Qc2R39aptEwcGVRdalk0kXWWSNmUJhVa6A
+xU5dCJDqaxBbk5DcXtXf/Qvimrm35BEabrUoRtlP5y2hNXyFeXrX18DP8vsVdJAaiBJccLKmwek
GJTxyF/38MSFDVx3CKiqbxGbYfDOlwoXaEhfy8hD2vNBhqsD53tyfvyG/K/MKE4iV9j3bM8pgtHO
l48Mu+NkG2K6DsFirLb1gsHh4cKvZ5VtPmpBfltU8XZZyUPXQEWuucx96QFLiZGfbqVmDL4Yaq/W
Omk0lyegxQzGRxrTlsnedxJC1aQgd6JnxlP7IoTQJg9hiR1GqfWRSdTs1PCIXKstnUs0WGbG526K
tnFjacd8G9fpWmkdMfLwkHIWTj4p6182/+MS7JWBdb+IlteU+l1nLEvmFpodd2gT+bmfVzzzFjHO
raAuoLlstgSgBxEhkyL7dKkQQwJN09xh2+HsR3oPIG1vl6GMWAogp+cGFRMUJU4u91ygUvIqz3Cz
KWtpaEESs+b9rn7qTCylzswhX7djpY/DqhLmH/UUEA8+57kzyxxUUjzOhO9Xf3QnOesf4TBhBXhL
LwfDJpXV9ws3nVfPw3UpzSe48oIVdTI9T/AeayFysj7ya0xdQQqQsCPOj8j4cbLANkqDrU39+uB9
MdO0po480O3Xr5fdeeWwtknIVGushm0Hpgv1CA0KgDrIgwENuzbLPmVmdpNLwt6wF8Q/4zNedGJa
kiR32Hyt2LEPHRlX1UW+sLR7N7Egh6spMXziZTl3xGQ0V8rKFkH/nr4XZDeAAvt6zz26DJ06LjOu
zYxzpfODYT4tmib9/9ZPme9lb96qfa3dqmMPwlb/AHCHWM422rR/PbXGfq2Dx/lKM5shSIDGhnCB
DIVLHfvgkxh9WDGc2R1kINWo8XoPPb2LwD8HOZAu0H7mR4D6oPBR+AWYWsBmKQRSDa0aDOxt2udb
IhBVtdbLRr+nf2ECA39vNMkAegxqOmXJdbg84imQpb2uhgbpCzq7Bibb6OYbxhGJ1n9soGjoFE3s
xDoU/4mv6p48hc5Q7HDQY77ifO5ipTMio6b2ICBIs0ii1DR8QOR25aUVGkpFAzEtno5uCOdZnMQ9
GP+XuePwCO8xE8Ioq9tilw84pH3CeR1Sm/q904O6OKBXtOo5M/WlT31CYUa372i97RipVKaBd0Rx
yOuYh5REkLkyeElsdUYh3WNasI0rAtw4L0fUkqEbI8jorgaZfDQp6HoZpkF9ApuYXayJSLVEGeBy
us0dHiAtPn6ltScmxugyzF0FhbrarifICWIIxhc0V8CUSBwiFnbP7UKb5oq6DTogaIjgXoZcUqZ7
I6FJTey6MakYUOIUmYGaTg4sVg08Y0W3U7u7SkOUIPFRsnDgUJXy6vdmYSI+K59Fk/woUc87mhhb
XA5HVOxztP90P7/jO+0GEveDvBEGYSm3eqdXuX5kIzb2aslvJyDY4klXikJ4mS1iGcWmrFsf8wyc
Hes0FXQZPWDwVRkN2GHYjKUJYr0uXlsGKDbIYOWqz7FgePR/MgCwElk+/dnyaFEDO//4mOiqKtTc
8GQ58HbxuduP1D6IoavJFseXqBLHf+SPxlmxSWHodKRgGNdGXgzLrxpcUKDiq5VWOVfZj7bOh9aL
9nBS0rHxTRz7RFWU6rVp7YvDZT4dGY1xKHDErAQRoM5WS4rnSsufVMlwO2u2WrhhC1r6PXR83bik
/3W4kz9wVj1N748sm6a6WurgE7Be6o3u55AVlyJaB7Qu5ILcQPYF6vgOoLArjFPa8idacp6BjxGi
HBAVNTB5RujnBvMoHAUeGpI7kyc42VFPWMMB/8NgaHFe8SWOGi7MLa2TXPYVJpg7Xgb9CKGpZ63l
PA0ZpFGC7YnLAaZcQqYb1HTdNP0GLFTVYGCloNjj+5tF7zhv3S/YPy64j8ZAYaiWZCCyQwtBuav9
C/aH0EOErYZwpBDwWY61XNwLxFiaTc8xXSZyqd6sV0+rsOqtfNRGccEXmPtJsIXsUPdMVb2V81KF
ySD3yK5nKYmmMOqI/SV5jmMyLzQHeLMEV6RLgnx/vCZEog5FdwQFPC7ClXRxHKG5SrckcSdDCR0x
XzzRavqTomAVqN8tYRpppJuYbikJz2GQ0EmyUOEpFS5S/Q/mCkGTI1VJorwC9QW46Y9Lwtjq3FuL
qxzGStJfZW7ru1G6L3tMPRHqTgBrWbKTDj0DWxxaE7sQwGlpLppXylc8YMpmh6AuLSD+w3YbRsaV
XyAMe7FvI7rU07r/XR0hDo+AJvJoDzd2OXFsSWmQ3JbUHF2smSmjy5DBjUR1MsKTNSrpsan6Cez2
GsWV/oa3PnMKmE4yxWITuSZ7n08JQ1FSDgwQW0OABltQ7Fp7oqAEOkuVrvuyQJ9kww8Hdch7Ot7Z
gI72VQyXSxW0bkJnT81d+4ou+wSbe5+se8Iv1Jb7jfkPNQ57nBbb5tdyvjVtiC8VN+c69Oq21FTA
GCgPm+yuPPQL87MEdSZmQCZIZgn3+qnz5C4LQtjrUB7va1oQb3roqxQKM24peG2AaN8sU6wfWGoY
LN1Hu22JbdrU5bxkq9BjQhMIcUO3hviGhec1Q81SYggVCwtLcCfdrVJz1Y7Huq55DWLwL4LT+WB1
9eWzQf+gyWPebP3mFTKPAi82JN+5NTsnggJs1Xekx/NBPYWnCjDYheQpzQi34noFOGw28S4x9z+6
B7bhlbAIcaOp3A5olBstaxnkC73GAJnnLStVFf7hvE+kuCd0k3WrRVcrSoR9/PXbmnMfPxeRchl5
aIJxSoQsc+m3Nj2+sBohgjh9BLbJ11xqnuPbDgsX6SZQ8LuxPKdHd00EvYFR48uhbPQ2g9b994wQ
SiGdt0Y1gtpC0kMdP3soIWRnWmfRR/YUmouJeUwB1xvfzQ8oVFwMMMTp1EIF4NTe2FUWbdzybdMU
41vJcXVv93U3rU+VZgdp3WP8LTBO6QbM1eq+Rs+C/KjmoNv9m8YfI6U1utVKEREd7wc1BemWlFpm
mi7jU4W8Xkjl3VzsJt/Knu7PRJYj/P4MT4ashiLrcEDyxThL7m04y+wAoczdNlvTTPmET369CrCD
Wu/dlBameLwzy9uAfg0co6IlbRxz0x7gDRJYzKLxtUr7HnvX+nhGmhD30AqfwxUGhUJbm45IjwEE
pfrhpkQgF2LjbmBIcwkmkrq6gsdJpiPac8XQXkk2dNmvgtUDLB+sFAf2PoExZ3MWgx4Iph2KaJHN
hDdNA2DzwrHn+jLhQnwLwXlTOf+3LTM8gaBAmlIgUCmroqMBm9xQJ2XvntkxlQA3c9HLu81JEmQn
2qis9leQLi40uurd51nZTSOrqjpangA4LxFFtFt5oyuqwZAtY4unLtYz//nuR0BrTl7lle4v3r4e
YsRxre1l8KSTX7T72pCGu0hveKvzCtOiN5ZeyjqMBB7Vgpz9X4zK0jJQHIa/yuELfmRYTV7Ob7uY
V2lzJ1bk2U6D9umveS2KiDeWM4rBLj+sGUmCl+NHxq2PL/Ep4D9Wv+yh5VdQsz8S6DLQc3snsH46
JehyUU1afZDPWM0XEY9ZEXsoNP9i5yD49Mw+XvbuZWJJ8kyNGPqu98I/fnTogRCW6fG6OaVFRGe9
TECy7SvMD8xSh2IwRY+iCfRNeI+Mi95zjeKuBn3wnkFBJYlcxP65f5C5sjYaNC7y7drSuJx9ycL9
Mm4SEix+2nr1NoHx6XwpQQcQ/QDYAJ+4K+m8ZPP30tScviSmG5xT3SMumUuwC7/q0wlTZx/cOAII
3N/ZzdKoTct+6EKQGqbsVnhTPR7bseDTBGhZbpqKd3G8ZwYPy5msCO7mj1dNGb7hpLlx1SIodWvW
EhD4yOgpWoUQQgW6HPb+O6zhPHtVaUh0qLij1+Mln1Dsq+ONm6W/RRZkP2JaPOlP0S3HJ3x5Unmm
4gIK4py645VHX/Dyc94B7oSnLOuMjaDTTrNW+zdJyWi9tvNEZKea2L0z1Dmfkug2Kd0Tkp6zCVPc
JKOSfOYL98sSjnZU0TJwLbE9oHhzCteEMSUhRX3kzph5JbRcbXlzGlJOqYYLf7RoLaR0WXGxrCG2
J530QG0MlSoSjx5HtlcFRdfuxwYkSjEZ4C9bVxWG4DC30kFEZfcrXjUhO11CmjHf4NBVbpT/Vcjk
rg0KI6OikcDb17+/ZSaFTuNyKFIOWM6QsmoC3CLtwy2JzPLUVDr+eqAvAgQV0bfkBGERFwHFCLxd
Fzh+Qg8gl/XOUeKiqPTTcoWAVS5FE86Nqc7mrdc8Q9o7F8T4yxQ+UcARxscTtsmhKxyuIte9aBbY
ftt6fOIPnV6mLSDOe8G1gsbOMPbUeZC9zvoCHgVmOeIQf1PAXLd9K+pGR0sRj0LASElCsgH7/GM5
REMMpHuMSieJNT3TfLqZcv0sYqu/PhKze7HwTmhwReseciFLVtXhiKChRTE6x9pAvPbS8/yznJXe
fjYeuJcUZXJ/HTSAFOF+X7UxBGMXK4JdFzEaLyslEjun6amCY5BSWe+g/3ty2aq7ajStMTsRBFIC
7H5U1RYW+acOKLHSkDF78k/f7SJ1gjvzh3Erw3TZN+6ghmqnHjzYTzyUkR2zeCvPa2TvfYSqdZ1g
SMpZRCwYEvKs8psTO+rX9F6yP3Wz0VXuPMkZl02e0tJxO1yY6PT+oKBTbpt0s/R+2T0ZEVzT1c6/
LYhN9OAI7D2antz5uVzoHM2FcZ+C2ZHDkEPL1htsmyHn7dbKJ+Hq5RHpUBv2y5kKtYlofsDCIrL5
M/tVRDMZmD330+KlrQMGKktvZKSUZMxnlvKKqGzsOIwqIAipNK6Qb4f3XTalUhFWb2MbgSiKtHce
Q6Q/enOQnhxQsclmM4U0IH3ISLk0YxmoQJs1zKaYMcTdh/yjT19/VKo/B4REVzXfrRBF5fZjSoR0
XdA8vOm7as5U1+HgQTlzUN6ch5HR45OBd9GsNzb0xNm7gpZwCSgsn5uV3LHvRA71bDmEviw2LFYq
RuvtZMuQxdyQX0+wq1IxziN8mbQ3Rt77en5Kc9BlsmWbTKuOwZGGki+aeidGT5EcU/eXLwhfNm8I
KXwt3R/zNSzvLmIHfIFQvry8QIFe49mt37TesVrSviSmyrlOPMB7LcI7FBzEOoQq7jVGiPn54rb/
b/Obt4W38vFxEE1VJW0TqbSM5EkqlUAJ6Mxw416wtkjky6p21wonlLZcO/96cbRHOQUB2pXDQaiM
ipbXDqFD4Ebkzr/C8JoIdKcPJY2BPW96jSL/WcAz99Tt3UCowiuLjmJPJBQk71fh8xPDnojv33MK
MGJlknIlE1lM3sAO4FQEzgcBF4KPVF/KqG69F+bx2S2keRCfVAdHTl7JBnVhZufZH56SdlOi56Zc
b9pFN4NpggB6TdtXdkJGUFs0JgnTKMcaYd5a7G6Mx7WU7m0s17PV8Szxr2ETugJMYV1m4n+ttPlS
fVtscIAN2TVvoJgKfM0IGI7DeVxmgzwNmjDxiFmkOUXdDUUkM/xKH0KdLARz1ELd9Q6zi6OPZche
nI4nouY1PtjTEWaWh8XhxXkAAhjk/cOVKRNFkI2cIEdN6ngUCeUIuBammwOaIGSbXF0nrSAeGBaT
Js7GC+YAui86zj8B10d9dzhEtNtIsHmZ5vGy9ttQbwis6FALBE8uiIdiiBsp1NOJYT6JRVVT4nyd
9NwhQNUWh5QRL3AxTgfduZImHkMo1A88PhvyXgufWCPXihLojsMiI8VAz9gQ+IA77sfQdyXXAu1L
9RBt7UdEq7QZhJxnYmUkn6J/9pAwExOB+fqo8t3YOm3U6KtrtZqProECl6ZFcMUwb1LL7qryd+kv
5nK0Caq0mPyt4PHjpCaCSIFruixgCvZJVz/RZGqckpNbhMnjXD1vTQR0nv8OjXujrx+l2yrSbaWl
WpHY4SWDn3W98PumwHEOM8vaAKgrce7bcWbVAvq3hWBeZzCWMLmN82PcV0ilsyyIVWKCXrMqFztL
HTvQoAbcZt9Fpr/K6DW8Qo+qev+7ykNWLHf4Ev8zBMnZmtriPZl4zR8+53Ax0swTJtW4CACAan+y
hAqdoh1VIaqeMKaX365/VtYa6ZFc0BfzSALiiUINFJ4HypRu1gE8rWJYtas1841aS5RTADGVam4S
c0D5bFvzQRZAJU70t1HuBiq++CJSjX8G39vmJrToWVF8OECPfA2z5ZrssXY82HK7ReWwnYVJvyAl
JYH5qXbdxnQrW7BYwKZY87b6+nRvTaAm5KPhm+xB0q2mkXWSMZ8g0K3IZTYCumdWxce4TtKLa1NR
qD9/SMwZr+6flkwRjJhj+rBBUdQXOPKoB/r1xnb6p4te+ephoPMJvatDdx92xzY/H4SopojvocVw
68oyStk7pbwnfx8x7JgS0bD8duNcYa5L6HbDKCRkAlytWHEWWOQH9hdRb6Mjy6knMwL8rceGO8Xv
gFB3AX5fAkQlyJkNTYqNAJzD84+Ds/yUlLEMzpk0jggFuZA3/UdjmzG4HhqUVA7/6vq9lLG/mRZm
AyVidxsMeUDt5YfEoQCoRVk6ut+k/wfnzJvJi+srouTAI7rePxA9jMdhNpNcFICn5n+7H4Y9JYXn
iHVL8iyx4c0mssaZh1ptour3Y3a0JgRqiK/cuuwBKgmLi8vvmPv5u1hZuB4I9sylxbLGP767JUTG
4KgE698N749d6tfN7WXoym1krq1Zer+7OHsHpfoyGwYXf2hSqMpMKSKtiaHEisFK8n/T34EOGeaK
XRtG7OLQP/FGdclEfmoZg+KLN4BwNpZuL2Ie/TgykCm30WWY1AANU8+QMOo+jlCxfg++U6ctLzKD
5e5+7haSZv66TgC3SGNdSD9UQjOLdBulYQHHcZ6ujhUOkuEgRwOZDLr8bs1+MlWj/8DYPiRcdA7l
Eps8Je6vohKupX5psa/TO2a6tTNnqYf2Bcehevei8QXCFIKFJqijcZsOJISBGvVQUH2qxGMIyIS2
m3zypI5cNq+9Dyq9wkDQ6liU/r5DODVa6esrVXyWuGfUSXn3IqtDQwCV0GoZz+Fn1iu1CLi6ij+1
fWlNxYkUbIvwiJSbvo0G4uFklc5YJ4FE628Hhnzj/IaL2+holpRYoh20AE5Y9R+Sio1xZc2XaWj+
5AIHP4ehAQaE3aZxn70yJVoUg9a5+GdSRA8iQdIdUm20T6Mkpb4O68XA/byMUQ4nAqd/DJFmqHpO
Vyo6+O+MRHtAbpmC0TlsTBhqBypRMIOtS3weDLe8YnMQtfO4+IMkQ4IXcLQCXYP/xRjrc/neVeAd
OA0riwybb9BphfHgQgfS5s0qCWkH0sszYdowqxu964rgVCTAHB+nJxZSByl57cyauQbU37yRxk+U
LC24MSEcFX/KUsT0lmcXZ9EBlhG5hGbujne0XPwrftBxBk0mRslE50V777+Jl/lv2iuRf3OnGq6w
vA16ZgcA+y4fpi15Z66l+nnVpK24e+DK0CgHRlwMgUKX8TVQRKc7/5aeMX0o8tBdj3OwF7kiDQNQ
mzoApbmovPnDwVxQNDwbcsB2fCxhPDvUvDbR3oAcjzP1w1D2WZdNK5LReFEYZerb6lhh45NIcNKB
b+SrH4kCQKmojNlsjtd79OPFXOXHsGZp4L4OKR51Qb+PDW2d4fIXcD2+qVDI23rt/GMrqMdMzIGF
lKvNaVycfhJKq8MPGzxhFkfHz0sTEbEEnSoYJHMxGpbWWYPeHGlCz9ibpyyEdENLn9RSg1h5waQ1
frIXpK3Sn88vgLerEyD7qz80uA5B20iZqKNi0AT77/+/kP1g2iuzAyGEWwlidvVFWpRWYLlhxcVb
GodT2lfAzrVqlVOjQghVFjg1NqQxu29v3QjbNUslIuf1BPtdo+5/VuzLsRgMPR9EGobc47sjD+YO
Znm7bfiH0lLVhMex5IUSZb0hQipPtJkUWr9azrs2Z1OVgwmMhc4JrtW1Jhcl0tlGaIwPijcZDIGN
JhZvUDoC2E+lWj2tL4kZQi0C4aRGj9zBfJ1EYoqYBhnWqUwHc25d63+nkah8YGjdhTahgilzIo+C
LfsGftbsep+Dh5T5VUU9bm+NW4vkE/sIGq76pwbI/6bIiEeAN/gO7pGG4l/7DIEyTyLdVPKD9KsO
cwTUFl1rQvsGqXDzdB0iA2bYkAUc0A595Koh4PDNGU4f4H+NAFug7xnJo5SuM49+tF6o/IA5lAwx
dVgGp75w4VvtJh18uEcn7VCc6drvI/sgI7m2bYsBzpxnD/6lXmPHNhSyJZoJyyH2Ot0qQ9cBc7Od
NUTLy8Kfd0trkpyUZvqEh3nHkmFlGDGW0wq5wMwhujhMnCRVj3/ynvqhd7Oii0oVdpHTHqsOyKz/
fpfBaNhAjwuERdX7B0Vlv4/oJbN/m3Ld7G2x7V4yGz4D9yerAn7E6zTfdbdOLvEkuAM7oWUliusm
lMo3J6Vga+6YUDbNdcbowZyfqfZUyhHqEM9gjrKUTiMvTGfDjtkzSA1wVHzDFp6xjnuSglRQeCGQ
EgttIKAmBVM+ek3wuxSRAVjQtKfm5nXDOgWoKCP9cbLuBptLrY9ePwJ9xolNGN9eqTEMmH8W0LmQ
FQlr+G8KqfOGcuS6ucmoAynAoRpmZ/jFfysJZSrLvHUSOnyeiHF8IrwuplcfD6YlWpupqhtYBkMr
z93zs1H0Ump5jXvASv2zCH3zVeuyqmLBbVfD8bMJb/3i6CDZEh8rlP7boMnhD5ypuZsnZCxGphnc
u3NDuGNRp28POzRgeM12qv9ff5ZDFa9702aGAEW7hAB9okmP8Rl2nE/Ggdu9xCwR+84uW7BtcKJI
cibfR5YOyVDYlwk5iatGxHqvQEBSvTofThjMimK5jbjt9qNXzSO4zXd9Wy3gipq1vUOXgjXp4d2M
WbaSo54ChUIyX19+QYIJmJu3Y48uICiAt+mXvpz849JAzG28UgxNOI0E7dWqMwhF7+JiPVA0Gl6R
W/MWd1UqwSkH6FQbBe0ciFkdn8oHWEgVKU9g3crUacZkkmKRtTuQ9tk1TN6OPJL/a7NpXLIczfvj
2JENa9hC/vDc2/6BzTK1WErWQuPQd/u4NXz3layXlSxo6k0NY8c9DAXJScKF8ygVR1t/B7PxE13S
qeA2H0pog9dwdGbsgwfebAFTdD+ooBuBIjoEadAmiwbkg0Q85v3ISwc6R/eNZWq7C8wUdVWgNGpy
DdT1/IlnipfglvJvZRKzqsTw9RD10PTgG9gXrMYsDIfbkIT9dw0EnI+oRbsh8D+5SftUdTmDFnoz
K4S7iOXTTGzzcbmB1lgzRjDRoltOmq0jiTeTBlsrDvq7L7s3zqp+zMccOxK6bWEGGzYh0+Gr4D3C
OAvqHOU9Q7+cMfOvQ/HewZlYYoMs+wHUJqjO1btQlYQfLzy0ecgdC8BTCXYF0eqL2uF9sPNwY5O6
Cp68lGiNd0YJcXJRjhg3J1hHM8WAnxpCLctBQad4XDvDbrj9LP+S4QD1eSHQLCk2F3aCMvVA+axA
5GZ6RPnINEWHJhTtT9lqiQI2SLIn8bBoCgYnwVc0d00RTe3Np06fNFLdfS59XOuQICxsqUWnd+iV
aVvl+oiyAim2eJhgSkIKjk/kFq5ZvU/s6DJqSs8VNy7McpoNy2OHrghv4V4WOE2nXir+ZRaVGJs1
uLwEqBhUbMzOeUrTn8bpstjvaRlJfavjZChKfpNrwU+sMYzXnNGOb7rAhmR2gXUiPIg5DR+GL00K
hCE8BazeM46+5eqzVssjoZDNEKYjPjve/9kaBqGx7+u7AGaUCZcQXs62fPJQYXH3HjpChddNy9S6
/8IM7vEqJU3silNCBgcj/iJDTq/D2mDK/7GTtbwGGC7tPq8uSDZeKhJb2QtcE/3QI1A/qTYvU2Bw
kaUml96xuBla+/CFbIJ0cnjaL0Z9jozFi+NJe5lsuYe6zlenNC74ltRnqJvvMQ5Y8/A293v4YRY4
s1OsUw5qNUb7NdDwmOlrsrUDHpq6USO45zaFQ3+gFPGWE/KYdSWJ8uyQF4fDb13LduRz98y3MyN+
+L1adZeTy9mHK00rU6hSR7s2oDNW8nUCZAKhjUd1yISv1D7YLTkJDIlGwT2gJi6vmi7aM4M50KcN
il4eAQfw2kDsxfCX63xvlwY74efg59qlofXVURqR2zP1+7Er44aXghlSHB/aWcsoMYdNqQzl9S9b
dD3bQ0FJrcsqDCid9yuxBKo8DMvLGV2JyjSzsoZQDlO1UhlCS/FpY3ZkRoXYfR1s2aO909MxXGy2
V2CZuQ98AJCgLSv/x2lmDRIjf0SXo7cEMcYjR94tj2leITy+ZwwKUNO5Ff+PYbRvH4M7+ko7YH/+
dkpIUZF/FEu/3Ek9btQXcHOSaPG8Elc5+rvE//o8+CLD4wPru8xFyD9rVfJQSMMpYUcUjttr+rq8
Sdr5/lFLz+A56hd2WA/PQvTF7FPHCcrk5OtMuONpsVe/ZOjouEtJASDyiu2hjbvEwBn6F4J2Ll4P
VuURhh+2a0vcDKNiu6qxGvX6aL3WC/747R8KEuxGNgdfcmrJyMvrBw1EQUsvd5Rhva8GFPlmK4uB
oTxM76Xd83u61VifIy+uMVCEJsdDM3JgGIO/Ian8aiM8IU0nnN6HQCwFF8bzZdJFB+UZaJn1hr91
5q0E0ZCGYSnNsps6cqY0xrFLZWIOHszT10cC+/nFQmUBPLX+4F9YFx0xQ+0pE5LTKOvwcnetcHYW
OuhMC7l3ykWek34XBz+ioetskwDbCmsUxgZqGBTpzqh/rG+VED+Uag2tDpd8CjPztb2SRZ2wP44t
fGHgT/UGWth0iKNyiXZkee9HCUzMLWTethQjpgVoWHFqtru7tH70mE4EQMLRSWcxAI9N9j52mp1N
lEjbGbsV15Tarqu+99/E/YhJw4WLj/fAWNBC9To2ro3EpQxmPpfzgz0CpzoeHtEJNbhq7yfQdXYo
hAsmAeT9iKOqNdBGYFayo3+Vla2UzTZwwvGxgqs12tS3FjuLjAtu0XZF2e648rQP/AA+np/zErLA
om1FJVmCHaoO7SP4y5RxxYdcqzfi9Iq7gICP8dkDB3S8+6DCxEoRLkrNjoG5GUNS5OyLJNATC2vo
AeoJspRaglPzqDUrNnYOsjgo1u8Q5XlBAGQTaDSjwPAs61Z2+aUa3BOX//ez+z0qb+5nTvHk3LhL
Hkh9l26lnvZffIO+Gg7s4j7dLQMRLAUUsmbDl8S6xlGKcFNkInXfP4FnHglAI82cNrS9w37U3zFA
BsKdSyzOVSK5APkH9nJm3LPpA7pmreTdXQbTPFAHDfsE7CFECqsSUfSmB2TeQvT+z1+l7HfRDwJD
rlqAlP2JuwWJ9FQu+9HuGa+IDRbsS8OlOpgaHV86UiOJDuLI1GUG51HCXw1BIc9X4qQi5QI5LD/h
fMVhTuNXCRLht6PwrqEhVEbX6dEa7T5LTGk+gNDfSKbGfoDf05nBGOwnEh4hYM3AkNv4Uc6KwWQh
pNkdbhfYQQ27Bz9P1IlsCK4Afzn/XCpizQx5Pzzpf6LrHlh6egErHrIdS5LPT0ndhAC1mn8vbBc0
cNx1G1JYZGdiF2nM0pCkpv2v+077MEKa2Qg4P5zhCXlct9XMtzZER95nrC9fw4TAJVKHIHqYEFXq
DRbqb4H/nXJLvwphRLE1xcOQbONqzJHGRSQPISSTKm1jsCxS5MqRBQwxtEl2Gwe67bmiU9zVv9Nz
pTVNikz6soEzSO+UR1pOEZNGUVMuUAVs9Iq3qFUpMgWbLbjSZgG8EYnattZqP22SMDIPto1uPrIZ
pygvhIZWqj/WcVUvnSTb4cXGJEWBj5Y8+BSBY5SSGaErlqdVE4ftFCH8MNfkMXjtIuGucVFUt19n
jyQUH6/mcjM/fiMIvuLB/C8Wv6J4vN5HZxhWBf4qqwzOEIJJ8zhx1KBQQ4fuI7I00SswKa19DDCg
gcky5TwsHrQW9LhwYK9oZloMpYhvk09uRUOkoune18CKScjJWdgVPBOu3FdyINNuGrMAUUxDB9td
oGjmA7W+YE3QpEgsSEJRIob12V6yIDOL3AO3c4HSTLLEP6M9UmyeCKLsmH6ZTnVS/imR+1YMZFUM
vmLBxOjL2USvaZXpv1RXSlOwQ0jniLU9PKdi/pnuI8ood0ZYtYe/LD2XjFaRSHAJ+a9/jmLH7Wvn
QWyPRsXGY1lRKCupaiVUJNolW2R07jSO6+J1kuIjuzlNGZHxmUAWzC8Yez7m5omnixt/lAZj2GHE
wxZjmduhi2sft+EWXQPNlEltXiI/GD4kjsJUOR5l+6mae1PL6QUopLZ2uKy6aBdhqUh0vL5/sbbs
SEUC/Fik5pxnhfnsE/L2hrWfQxVSseTcAn9yliBuuxw7txQejfJfhyMho/ht/MO7d02tfmBp+v1t
+eUqoxGkyceJYFG3+vsT1ME2ZEnYonWY3hFR2x4nyIZn8kFtceeNwdr9xqTMs3PbocubX4bY+3Cw
iJNj94oKIYnZsG+VWeW8fjMXZfcWwku//fdpDfi3iGxx/JheC+F0O3w5K0YD1dxyN6OsMTy3wcyX
fe8BZ/hU7nQ/io5u51gmuUUkBuidRbWKqhxdmrhy4w9MfZBJg88lp/JFi31nSHa/aN2QERKefFo1
usyMMzoBXjbiqATrgURfdNGvQi16J948ZlZu46qEY4t5e9lyfiFxQIbAq8XUvgxnUeDd52B6oz3E
M+YKQZrsHdpj/ej80z6c151b66vWcG+0i4xH8nXPiABCd/02MLXTVxpRQqTgCJCHnUtqGejPK6lb
iCkKEbB/gox/GpAuthxywkKzt0IGUgqO/68zjot6cW6L6+xiMliy2vNuKNxzK6B3eYhWgVVsHTUK
KU9V7rsDl3yRZWDzBTcHYxTEfECmqGQuqEnFKPNBkxmvGfXkS+glGc98gQUf+9mrT2iO7aw0XIEn
asqLvZoJvwPjONDI9GFsCNOp8EW+8CrPUOodRQVza0LxzyLgMKAjo/AhHtDk+OMJj8X3VXPRLCKo
qypeu1II9EJAkA6+ZmGdc7bIKfBRQx9V2213E8HLghD8xIZRqXbJYW6KxKy1walBcjiIWof7URIB
jYsUm9gYtgoWu4S/6tEpAGQ/wgUEVfa/2V4PHGMIcJGGemiL7UauTgwxr3Kfg5jL/EBoLYmf3RD1
Bgs8ZKR9CxN1qeyTEMvdQz8T/OZRHnWgZgQsfnwqqtlJ6CWKoOk9P5NaxRW/p788FQLMbduqaE0d
lWWSVSr73AVu2aS6zb6DedGt3eNbM7DcQGfiIlS7Dl6UIawCsjZaQ7XOjjjQ+joTuxIZppMdkwdG
p+khI0cV5CpgSSgKP9fQmyQO9aDGBQ82JH3lq6cgdUmTXh77SoQQyto7n0a8qXTD6vBNfrUjf+Xn
MXTM3qkDy51m0uQzEeAmlmUMNFZbmxY8DiTvqXHmgpgC13r0R1TuiAuqzUq5Vzrc9RBMNGXzHtXp
vgBxc/8HE3FwwrewC849Gdd3vdmOPyBal0l235H1EmqkGVWxyQKaB6TjPWlTAorI1Fb/v91dw7tn
mlnD8fMRc4F68VnADaexk0Cn+wnSiqS7xD0rGEx0yaBmVwLVEpuwkR/o3bnX2Qkkg2yVpQEnBcEC
H3HUF/kgsiENSsK5Ptm+ly9A2f4pMZivY6a56b72ffaRMrrnzd8+77EgnybmM+Mbh3Llwxsgkqg9
BN1TAWhfNxs3QCpf/Gezf+bC88ODUzb39d45sZrsu6VdUQkO/nwBUaFcfomVchO620pYgrfC44nF
kgjnoNNjw84XCLiC5Q2a46Tw0cdav66+cjT+MdcKAFgNHOEPGpY6gH72rqSmROyNE7rSomj9BsFQ
YBtyS6oZCf8wmGm3uH8gKIfV+aNVNL3OGXV79sigtwuE/xAFaloTl7p5WkM7ROccHOVyc7ajhvaw
fNtBILz6H5FhkU9AscTov3WfuNPRVnHEKCDVysz8+2nbk9TwNUmUbYtV0zsyoo40wDPqENwQpHKe
VQUxm0q4V2ezcHvr1GsVNcWBqECpZDme7iNjRTk60prAskiAQ0KC5fCiqQF4MkYWIxIbNByTY1Mx
xaqfmn/rRWrARkmG0e+iU2feoimL7AfkAXbSntgLOxC+nWobtMPK6Ez6mH3R2lyR41qThcqnWNNW
DZZCnXXA2YoDg36bm87wRN/yMYN95Obl2PvTsOhKgtir1h4zmpYNh4c+PjBZpcpHI4kkjLAC8Ajh
55M+cp0PQuAAKNFNcyJ+RzmsoPaUAtrFnVMsetqzp74Z/PH7JKWxWBiOV7tCYPh7ErvlR3Q4U8hA
hNYz9ZpSFppOrsBLY7oMppTN6fUw9yMZ013a0Y3mhHhYlxdIQyNQoNIFTUfPu6p0ocsEoqRJhHQB
yDmNSonNpMISJ5H7epq/JHemUQ3apZHoOxhezHZDVxgJyWmP22Kv1p6FfIghZfEKJtVVK2+0tCrR
4XzrXnUA/n2uSZcuTOH2HCr9O6YFzMgNRWlxtWYL/nzhaybOVOVH0naiDpqDU2gY32k4T2KOTgJ/
x0S0Dyraaqdv3u3WGC+0YEArQS75bU+ESHRAemDAB7xPFBcZvV3iZpgPxHwSCJIRy9q72lAlUyfX
bvYcqx8RLKER6AyLUM9lUGXHQnDc6MRlIspYECQIPExA4OArDeMJPjkqLW9yeKlVmhsqHo3UouQw
MUXFiAwOuAa64ctN7uCoCGHGwQ2PY/EOzcChm2yVc8r19i+UEVNbfoooi1lh7FNOVltVjiIyF18G
Rymm5x4m42s2KSW2zVKF+OhRrRksP3qjd8K5WAcH3ttoQBS78/LttgdkzAC01zeKIkYuJpmH6gew
lI/ruCgs350vFWzcJIFPBnDg6QMVlFAovZ6VtmiraBF6eCKlKEHC0IIX/2+CHNFJHP5LzXg+e3gL
qPoMG+AhKqDJalPjeVhLRAvBaSYmuxi1QW+UYsavY0y2eoqGjCI48k9YPPHQG3iZqYhuDZwMK2rP
/vDoHF/9zYeDu9NiOX+2RCeGU35KzPRlDNvthJivz5g8Ht86jzVcVmqOQsEKZjypHb0iTvl23psQ
0by0o0/hW3PByU7sPPddNfdx8S7kfbnEeu7PMMvdiAKbNqdliYElRYIQr/HVWlvJten0UXe2jjBr
uiOBxWW1+cI5HVGIoHvHXR7bsmNKIkdMWRSLFoHTIKDyB89PT1UvyvmDGP96ZOwo+HzPO7Ieskj2
h20pC12IiS3X8PlyW+B2pv+JKVVy1/yyYk68/IejQwdzKUowXP0qz1Sf5+5PakwNI16+/rRwYLrI
fHh4SWhBfRhEvZ2yRJZ8TlDjy2acpWQpZv/H3Ti+9O0FUnUf5hxPfh6YSbyB+bb9UXNfhIaz3hrq
rFE5mlV4YBP3iNIFFL3BKaTC69JOwps+S1n4g/kX+awaPW2oPuapyCdoJtB7F5tzLRXFtkKx90fj
nD4/PZcSI70Qyw1eurpZXZSX26hX/5UFLUT678KBlH2vMSyCUMGWTaXTfUovmLj5JCg6vdqH8bFX
LDp3m6CSJJHYiDas22Q/LTprhustStxYXnOxnLei9SipZFVyc9fEeIHmiJqJeOw4dXOPe1FyaBZO
EiVK9EbQCJAK2ryk6ct2oB3vf1fMj9RTPGMfj3nnMMAAT06SGIftWfGJLz2vYpZVsn0KFronkEcq
GmSaqSfoEprvmBpSQDols8vYDKhFKFE/0APMzXwLvn+hLi6MKcFV4C/6Yt9YKiDzbnfPOSmSdvUJ
iMFJY4e0VqtDT6VSqzvQ2+8en1K5injMHUdLpCrumdANsyjLQCPRBDtpa2Zl5OMP04ds5Z9w8PD0
7magCiHKigfChr7YlOJJeSvHtHzKk/aJr2h19R6GZHnQCLrCdzw4JNvFtUCJzxZj286llyvINuWM
z2QbqsgAjydkZfM5qtL5e9LpjDKIlQOsK8+SwamTv4K5tzcSDMNMBFEVAxY5ww1p2rKTXhC/p5WS
ukL/nM/+gKsBCoHpofFjS53jWlK5wVLSVPHVU8kVGL9JEfDU2q0y049eUO5a2IQM06LZgAZAa9dq
A7R2xnZHAEu3DqMMBrbnp5HQ5rGe/TPe/EX/OCzigb+vohpJHayBc04cKwf/4RZHsGuC5y2aMelB
lnhtG4ecOVhUKz5g2xg9rGq9EdsimgK6/Hda4rsZe/U6OUaT5S+LD5ECcVsc4iXO97cfJvrjBtiO
/G4XmhnaTz0fLtfX2sMWtbBxB0CFPYtgtO/9hvFi5XgbNHCqUewvg6o3GzPDCuGy+Un5FNNJ4a4l
bfmVaZ6nAr8rxUmQ5aJ3E+6rUlFtsdbT063+Lnl9IxsnQvKwHpRCWoEclOB8Z7zHL6BvKu0ev6hg
gwtK1EclpNczIhcuuraubRVijDTZ54b1MU5vZqmbnc8EMFviLExoyAwldWzVHS2ZYfnk22AUPeQT
cUDIrUwX9s5WKJqRQQ0JBMEXt2nP5yQ5npNF8LgiX7ZjsLbTp41VJA9jkk/wz3fZS8qHNjbKU7P3
Pq350mwBN6gmJ9jNlPUQyTRLGvQIDOAE8Ma1aw9WL6BoY5iNkq88kBFx0VQOyTUr1D2fTHTL1JHZ
1xEo9OIoqzxv7pK6pt2P+b+oLlvI09MFJ3cQfJbTO6Vhxya4ROIJ226HMJy1m9P4BFHRYnYDEqrq
VKfzo8npT1b1o340MwvGj5erBI02INpBXrCLDtyNWTVpR9f755RMapcrW0d03FfxuYgOAFns+TRY
nLDApTSbePUSRmgyo55oeb4NBMIrcMhq00lM9ssJzVytVTTTD9MyI2vfceA29YkeA7gSZSBOcAkV
kXdq2dgS5KmGveD0Yw2d/EFJLnoDT6Q7QFnjvMkmpSDf6BeuFSYFF9IbQo9DgpMv3MoZH4Odr0w5
1WG+SpAuAQobY7DJJ3uw1mFnvN5TC1NIz9RGCu0w1gN6/k5Y3Bm+ElgZ9cdR+crQuIi6XahcSN9d
KBk43rNVN8ozHasxwWvI+LL3ySYLrrL9+xwSiA5MwYaXbESYy7f5izAguS4aVgQxFcTCT2yy0RyE
ALAjjYX3kCnTmKKT3TJLGmZdFbLxQMSxI9jEljxwTqhoALdlJ4RvYTp0v84iUOqeQDH19gFUR/dP
40v9t9Q0lB8YyW+JKWR/+9ZSSwVIfwO0U/fN6ManDvPCee4BnY03huoSTlrvK8OI9Ca5qPloknpm
2O6lhvmap4L34UhTJaa721Qrexc4YNsOvN98j6Dh58hsQZabxWdY8KsQLd+8IgNKSqU0Fw3S1IUW
lIvBtyNigyDMpiUNA5o/b2udcxz3FXXS0jmswo91TuIzJuXQTaOy8ernH+48i6rYhaQIWaP+Q9PN
J1BqGVdOGPuymrGRe/IGFSZlm8rwslhSpdQcumDrWSkpHY7xloxyA0HNkhMtpfkCim4Rmp/PUL9U
7KjhOzw78bhiEp9AeacoVwe6yz2mZWvt5VO91qJFgRL5arDcf2fRZ6S/VlEYue9tE5OLwmrcKlZl
HX2jBM8Qo3y7D1DpWKTNpRHl0wmOpOuo+DWdPbUbNPCn8plQV6zjcu3dxqn7uo0LU1xkDFWf3LYJ
ap/IvmCEtAjhWue/6FImAX+YDjH9VWdRf4l22Aq6rtpR1T1OrI9LPsZG357Efv7wu131MrhX8dhW
NYoKmTH09TkaVC/5o5jYr0r0sc+wbstf3Z3xWaV4O0P3wYtnKml5nv/Q1d+U8rb4zGmQHof7jjvy
k1VG8ez2vKUf/VIfPbfigXr46phgXnQkqkFejiuMfuaS/T51lG5bf+TNf9rU/Hij+WQ6vxACCBSA
1Y5IxHx/Zq+v0yAX1SVQRNxKuo2ngUFV/V2dqDdwO7O0EyuqI9YteyrBtxf2W5YEbNZ0074SauyN
/x8X6gUI0dc0XCQ2CokYDIFF/KsEIPP/UeZNt5HSQ80gXG8iR0VVNRf7rr6YnAetQJrHj2NyaaOq
5SXh8D2QJfmDwSWNlz8qvxqGDnbc2tV1jo7aay5kQ2k1pqI3RrtRD5v+ex34fEJBLajiYLuqsu0y
lUTZ1TYmes/zuwJ5+1SP1RiG8y88JtbKC3KvBdB3oahZeyZLGBmk4j68gsV1OW82loqpOqQXtsyT
oxK8FkVxePgiyYlAWIkxR4pFt5Eg5ANSMJIaS3btAtP7sZVT8ZOAim9j5qA8P2u12SFihuVFCh/k
B8/3y3kgkFPwhWLCK1CqcIHFSlC70FmNm2BUiKwUf07cmSI+CsPPd9fEt/OqluWKvaFc+YsgbZHO
lucxVBbM1iz0AI7i1tedO/UiEkzhSJMpfV5+1okSqIGEcUdRWJ99Jo1WynxL0y12XSXyFQjh28Xi
RzynUl/gNlc4EHOXJRMII6NnLseqa/5+qlsXtgoAgyKseC31jnlRp1VKdHwLdKv2zTnaXbqOX+b4
bZfQ/D/bmlcKOs9t8VbRsyKr4AejsnnnV1yCquR90A+MuwQGBh30MOt23ngXNIfJ/8s333r+dzfJ
D0HWO05bNEbOlMPWTvMiCEMU6xi1rmTNo/jHwhIh1zmB9PEc+egMpa8AgYK+Pk0o/j5pAoDNWjGL
r3Kk/7PCvYEGqU4FvJ2XaOKRvHPnJfslZ8I9sMjyPGXFyHZeznLR74Bsheae/8HeCreEYRHVDBbG
mK5Lj5hT3afpY+38belC6Nki6V6qtJkS8x6MQ84Er1fhyumzjx0rVPfNAEd/kY95I6hnoBUud6S1
jgtOyt/fNcWOPCBT6hVDGFivuTSRSP40IAonWGaITh6k7njcFr6fXSqjXovn7tAH0uGs5sqniJPx
F7EJMYR5uN8kwCLTKduBLKs5hBYA5cRXoIbdJ0RvzegWwhb20zxkp5MmNV5/MZyjmc+0ra7wiuTc
r+jl9+HycT3eeNxEXqxtg4K0bSD7zeGhsVtrXf8PMNpTlc0H3KkgOUcllsFZ6jFv4O7pakxclyrN
fjJgf5yQZ13ADEpo3IPs2n+aXixYRTqBn035px3I03gYATEcIvw9Wpjp0k/N/wBNkLzTYjLruGfn
nwOFhesDivfQucxv0cufI+GdC5y4FyKuzaqvkEh7v2W4bLANeFU7LqUhpIJRhgvuJ76R9xoKEoRW
ixoMrNlVDjOMJspbZyJ5qPpQoCBZR7ltVPy28+MJlhe3ErxqBRgzpkPB6eNyLAX5NNcVpZ/5/IxJ
DUjH44dZPVu/iBnqEvnMa4RXe0RHpA70kOYV+A1EpQN1x/b4heimYUQvKfeWViUjAftDMl6d8V7M
/WB51vFKfWhwVLMh1BFsNwXoe9TdaTIMNk3dpzZh4ccXG1ZPrGoLiY+lqlHUu+OXBrr5++I6VgZZ
Nf1ZzFqrMTSvRugldkDgoL8wdCFukHkfEyDXCYleRrKM1A6SnhBIwF/aWuv4IH5VHnR3iMi2AjFO
7Ven1kIdfM82SMW0wUP59isBMfm9nY8ew7Y28+enJ10/WzDDYkjdM0EfG1670sbAIvLGFZHM6F1r
8nEuFY2DO7HxrwrDu6JDthlFz7clZ0zffadI6X6LufxyovTTQtw8kHBgE4ZYXF8FH54S8fY9PDWc
x/iXJMrAZHiVVwwTZZZ1LjsHXhnHHWdzscaDHq1/enRtVvu8B9bPh1LOCbuHnEHHroNHZeAZfCbv
0pcCeJjbkuEgAj/f64/NWgNaGUqQDmKYqSx4R6qMHMiJ3MkOt4uJ7HsUFQyLv2PP8Lpb8z+9ugEQ
DKYE5AdAmqhUHLuuHzpGh1rPErPTqfyz0lxyAPhbw9cXndd2t0Of1Wi68eYtUjzDQ+vZcQOq6UqJ
ssSWHQ1+ROTsJouEqqN/1mKnQUrehoR+sb+fbThI1Vj4kcBCtJu+ymQqSJMbxVbCp/+Q9Ppm3CN5
vy3USQJRYfYQK5FaPkbDLD8CduYiS6vCFhZWpNwlaXteI6XS8+8stMOR1yxJ6cL+aZxFDgi51N7v
prpphMuG/oCdwdFsM91Dt+QzBAxZdApQtviFBW4RsDHeoRgsUP1SNyVnVP4pKgGNSAa8l697Gdu3
8HvPa539EV1xkm/I7iXpJrd90lovqqJq0mOucn6AfLb3MaICmJLwzI6AlivCHc3of2v7Qt84//JN
5ESvoYjMQJEW9stGW0prAs8JuPIfiLxKKVxdWNTMyjTy4lFciicCF70Fs98xoVLPUo/1lMOfj05X
DcqhGV/uwhL4Y8MhDxPvadOIC0/7WtcdMCtV/7SZoSH0mLMn7FmRMgdYD5lcuOYJQtLxeGQuIsxa
XgMVx0nuqFRO2JneoPC6qZ5o66U/qNV+oYndMeX/6gaFWo5AP4lXEFgoPOJVzNllkNKmx1vqx/Vz
IEQqoATnqqv+8By8DFfgIi+6FIBFHmO8kTdxXpuukhycbEhxufZEfL6EEw2FiHatpl6FEJMqxfVN
0OjpsXS+wLLxpvwRSXPZ/5bVojTw1rgh6dlY+oWSTxiBBtW8UdjUPrvcDRjFzs0kcQshDzu0FVKA
kilR9V2KmueZFwcWe4JYSSfPEOnYb/V58g8E5fAnYBrXOFmUKZ915XE+5SCpG0V4WmwyrO129t0H
0mJn5cGQbymBJMXA5gDgeMa7WY/d0W6FQo0EJGy14K4rH105nENfHM0gHMrZbifSXUkm4c/qCNSj
hTVk86cQEaHAGKXA0M+C0ZQwczyTElTE6BYuiFBNjOhaLZm8B8nHVzUFw9vPwljJcYdaVajZpY/2
viSAKwXHpGp1waNFcHlR8uoucgOX0W3+3VMgX7Sj1TMPCNT/lAENJfOHmiaJf71YPROvtirJFC0/
X/Gz2NREhAehjF65tI5Zij7swmwq332wGmIDNSTBiotaz292RJ35VWWDl6JjYeounwbgTtDtB4Eg
pCZ+Uho+qrRO2EbLXWVbBlyXPbrTtWTCDT1suzmIxgZCnlx7+C0hMpzMMq5NsIKiKCtHXS8gdYly
qFTVX5uxHUoGHT5oJIfP+p4gk3Npqe+eNqyMONQkZ09XLS1/JXCwrj3DUR0Hz/OKYmfJj575I0Zi
9Ll/Am7OV8Wy9GXxYeX1RKTOkVa0kaqnL48SbChCp+Vry4agnSt5FZq1ACkxVUqP7ap74IEgqKf9
21MKQERI+0cYQ74mALQYR59rMDYnaplHePsPpjomvRfzO0MP2frxGkb2fWdwp4tV0jE/nInfQUAK
EKeV+yo1WJCFFkdCN+BKKAWKPbLxEw9L9p496MVBoMVvI137S8aTeWTJtzdr5UNFDAdTGiXOlQYi
rOeYZL4JYL3WlsLxtSREsID+aGZM0GTfmpeluM/D4WHTs/IItNJwbqWyBJnFGzkK/ryb/NK3CcBW
VhP0HMZi1QohNGc0NgHli/qC/gGZMsk3k7wIdNfSq8fCLURFGBT5JguP/RioG3zvSPm3ixeapv4O
uimbE6aDu6kjKzB4pe1z9fA59Q8odbxxr9yDa470HXXtc5NalzXSu2OZWC2EeSEW8KxoE4hPM+yH
0hIsCZ0+eXQyYe9fcxBxtmFWb9+216pKDyotMhGKHj4r2JxnQPS0vLn5qC/EvTq8+xfIRdOBm/DY
cPrW38Nn3yPG3WqFeyBaSFDcXbSnISMuy/D2bIT9QjsakrehyCh83l4ayT2+eI9oz0U3tHsrxJaG
g1Rr+HUOZcN7bQic3UEHgZ7CNkCRcIwE/+SdueiGcV9Gs/QZMkD1pMMFZNF8QD5mCO2Pa98Ib8MR
3k+u5VF00Y6NixJELqciVa7kRsVvGAg5uTHK9YCiKpHD8dvfNmRGj7zYksw/zaWimhf33Hi/3GNF
A2OyJS70YG0fnL2F+Zs8URf3z9sX0uvK94jnuvWnGz8nLWYilnGXO/z4pxtAwbAxjVQS5BIAAZoH
yX8OQLxQgu4ZOHRz898iI0b4wQrUBy+BZ0VA1EzDKzYUfdtl46F95YIrQI4zDYqSgzqzHoR3D3Lb
1ZM5B1NTPi2yHT8feAH+oc3bxEVIOqp9Hu5wwvFX/RvdCNzSHSFtZ3eY9lAfQOLDywIrkTxhfQiY
o8te5kW7eWzX4lIDgfYQAO60rI8bnmg7x4fK9SUWQ0jOH7BOaR0ONKNf4JWBXIzX64Gbf44FY9cS
zl0Wms8E/RpGvOX1S8gOkTGBVGh7HxazSeCMtcnCfSJEx6D85amekqcF6RkUiDvZlB0ZNBiHmsb3
vkbHdFrgdLg+c1VAajdRkBwlajKt58HyW/oWp5wlfdRanrJyyMHGita5jm4f4GsfmNBkagHLkkT2
KTMdnjChyrY4oYXV6v2N0j5rMPdWjxGb+PdV89M+8DiUql8Zek91yf4FYXp297i6EscTvSbJyDct
Pn52N5cNf6rwmzVmymMsAprKnO5sPaWvDCxsnGRg/cWi1yEc8PQ7FsuH9DsFI9HOKBfD/bXB83Il
OCdyDGZxp8/rPWEZ+qUOKIi17UaW+2OcLFcj9ZxGiZOP3TPl9glql5szaopRV0vSYT6z9BzROA5t
2p1UKF50U4EATaDJi2kiJ9dvXW2v8FzcJBwFaJtGujF9Rl3t7EBtxVrDLQi1BEFcpXS5iR556VTt
+cjLj9JorFJscORpVCyhwrjzAE0YdQHXk21QeMul3+XHI4/c3U1NBFxNEcStXHc01mD8+73vtTmQ
i1j5DjAjsuK6rQFZ/4eGM/5xQYrpZfZ8jbHJIrw2omMEKrDvxAdObmN7wTxsre4wH8Hn6L4CDdEd
l6PEmNe/uVdFe5QVJKqweqLC5RitBlOQTAC3lt4SxzGg5Xop1W+WEhgGOTjHLUnTc02vYnXypkrP
PdspA0m8sfmlx3jPuAhkZI+6IbK2aEDv3tXr8j/HRwu35pmVzrqjk2XWIsP6nxWinxFwz1llX8+Y
UUCZ11u9VagL1FkS5JjT6MFzR1CjeUrsTdA3PoZKOAhyMxlF6AJXyvgbd/6TnvX4Mfv0fmawff+m
8KvWk/CKO++84GRngcTQd6QLxB2/ptrFx4itCdXVVbXKG9NXJy4JELoyoUAs+cquggXlVBDkPeNb
NjpJK8QBbKGVZk2oqAhmYGxcfpvNOpWo+c5jNgHGBGsgSY1uVxrtD0kZTIZmKGDg4XrBpgSqqcFo
Irh5A9ihZxHE2SX9nyH6ithMjwhb62sEo1Ey9D76CVOe8vrofxqIgjRnynBzdo5tBmmCdTbA+D2B
5vRDRYVRDK4VomqcU6YeifKBtVAO/5AkuXoFCNFbHe6KcQQaVqi38nXGsxMVRuASxJU+qOtie6Kg
kkYg+NaAcn0O3e4GU8IqeCVFY6hCxrm41lSrWH7TiAiS7KGTFD7q0Qz8Wv13wlO/lKrW7SEiD/e9
n8qd1CFQxTbB35RW1v67j1FgFvkkFxcShPiR1YY7ZQ+zW8a89a+RJWhtYXyZCa8AqaxkQq4xrezz
/px9fz1tVYRdaSMylT0UaYrJjR4YmXd/QVtjrnJhYXdNtisdEDVoCgmLSV9uPdRTCGqo8fPcigDn
RHJow/xMZ2Rz8Uxl5hhbrbYoqibuB4iFodIW998HPtf5teJMmZ3X+/Om2nGS32eb2uDUgWhJQ6KO
y+o51om6+AmKGa3eyt+nLUBkdmUsDkL+X44DabAv7lUfpG2T+o59uwegnbTVVS30CCEG8X8p89mE
FNWAHj4bf9VwRtlobuwxDB1iHzS6JmlWXeNgginFpC+CKID9Ezzima5EMQr58SowwsuwbPNNW68G
ajwqhFF2Y+4W+KwpFomvufDcfcPAmSZ+xHq0nWzIX1CMN1yadAalezOor5YqAROV2N0MzWOVuxTo
UAVzaPEUfMHjDUPaTfU9YXcGvXvsie0tCOaOu8BS2BKx81zz4xPR/XLeZAwC2U0gTAMbhn6GUu4q
7HP6slxfQC91m/5FcfALNVFcmV0gn9vqpJdLHnEZabq3Rfc+dWAG8Tesv5pCXsABjUWFlD17om55
ipBtEjmZCAOqY6MGGvdfRKsJ4vprvjmk62oWtP3PiCf4SY2496sDgWoZk1PLj2e8cXzZBd2ietye
rIDXVJtD04G1jt68BqS7fAPbP7770nAyYG4g2E/VaO/3PAgspjNkh1E2wVShUhbIDBt3H2UIu0vM
tuhogHkx3mdQalfdxt+JqWUyQi5rAyUrAS4s1/f43qzzD6G1LXrWWBrsPGpMq9RdlPI8LuVllIKh
F+p/ch5ORGaWQ5GIniM1wVrckOuXKNsy7VPr3+nMhS8mOvev4gxATk/h75q5+vA28otv1e/QiBdu
z3yzTA+7NxJdRXvE7LlMsN0Ezg2HerqsvtJej3Q8HDSUt6pjy/ymKrv+vmP0X/b74lBRgReuIQu9
RKZ5dbWSxYDgKtC6GM25iHV1JOK/5lV2DwpEftPT+7A+mlaEmdV7mmlcKY41IrxxewCwdT0ArjEl
kRYZ96n2zHHF75UXIGajEVhvRlyQo5fjqPKaUhNXvpIbi4jBMwdmJ78699N2NcocyhZBTyqnEAFz
59vgiZOMQEmY+jsvIi4H9h+1LX5/HLPrcEiStw4xKQ6ogGRP/7OQlVSzVykzsQvDgCWIHgAGqCnZ
LwrLEEs53LgfHNAwVxynF5bkU3kTW2ODzCG3iGQQ65xq1QOR9KawpWfNTTsJfMYkIiEzHzfo/we/
ZGMkzxxWNl0rutduD5TsfF4JN8uobRU6IETVMWWtZXdcmOfA87wst48UZPe8Kp/UfNkXLrrFQZyO
+OAkoi6y9S0m24Yo5/d+rXd04P5m7OqCjsCHF4sY4VbA0PMdYIOLN1o44Ef6nNL+c1kajUQ6i7UR
DvxjuaeV0Zeb2b8BKmmU/8B2mSrqFJ5drNoQ1vNjJF3xMESK1fV7OtfaDPvdh3hs+2OuJAbf182R
nDHf07p4bBFFTgEEsl7mSdtkp8/Wc1BuAvUG7Zcj1IyTgTsVtp5czNJhWbDTXpRW+dNXlYcPTpmf
clDiGCJR6bu5aAcJZQ9nL29tIXRwQ6OYIFar7bVaGf7bddLXAU4mWBXWFHFZFyN5IZxKYcLKcWQl
hQwWOOvxeCACTVDE0CESIsOjs4c8BbYOhiV9RgQQr9NeeUVcAZNIEGBJLhmSYW2zzWgpS5RzVKKJ
4qYu7e0AoaHHoliLKdN1jybQiPzn3WALMFTXVamNbGUjtl6m11HcP/sNjiNr1CDvPrAFC5hB18Av
E1EHL2hN/ALQR15BNqTljUUVje9htindAr07y93CZ58fUAIckuJ+DgA6icBX//KNmNedcla2UdHS
9v0KkvplNL/D8BQAak98qehT2G+OLwRIXWUhp9czvwG3y0YpgcMQIFiUbfCUfjGsParH2gUGGoS/
fXr8QB3FFrjEOAENLV582YGT5HeD1LnAdAcLnW1+w2fGjnK5mbf1Ny4esKTjb3c8Gj362ZBVbnYx
ef45s1lA6hUex4yFoICAFnVxAizIAF99LZXLO285dy3pJSRdB5P34cWffFJ+GVHC7AVtkWBrtjjK
NsgimqYJcfJtLAOMCrphhSvgpJNi1T4ox5o0T07j61RT2lC0zB0kjFp6+BCrl3W3iqsoweT6Lhuo
0GjPKdq7JsZvo2AQOVB7RcIYZSzLhKZLFSGluvC5MaZ6mwseZ2QVDip7ZaCRKcN0nbO2LaXNn313
ldiqjEGi0SQ6YN2f77JWcrQFERjkGz1TU4UpYWyZJH3MOwsxJXmNlhxPtYmYDZmfF7P/Tr1mJgxK
PIPHdZ0YO3mF4241k/5B+fBPF44f8mn4jcYDzMUzp16z+XOFSiIYShKu8QGEbu/BjIZ1UfOw3+Ho
yhrAOXvTxI7B/6UnWNV+EzWXq3L/PBye+eDJTvQE1NDBKUbR9u0IfnQDwdWslmTYJeXBd9n4M3gZ
e3NGUaJIwkUTVR1/7QXD0k9fnEfISx2smpGotMh0tNIH+4vCBcH2Otb9zuXdEG67GteJqtxB0FTR
aUwIEgx4J9gmYW2SMK21EltAa+c//fCcbyQzFE3np0e3RoUae5Iw6ddpjFYeOn+Zt/oUBE1ncR4J
Tt3zvGHcBwho1OaQBMVqKfssjdwKOUUChGY+rizS6TbY4e+f2KpYCrOZZyMbuHjURmXbszQnCPRr
mjrXC8LYDu3Ox2Ncy/0Mn6h9S6QuDgBQlCIY9ra7fjPk5KW0eLUWC3nKBp3qIKPOkZPhaFTqVn6t
q1TZCC4smG5SfgH/6X7amD2xPE6xYJkQGo+PIo0wI0K3vKxlNTFXCl2Btp8cbh1NrP3iazHaxQmi
/fwHgoj8u+VCSXUP4ayCFv++2gdkVdpImE6HJ/3abK7aoR2xD3Wl1Jn7P9MeLCX/GLNWZSI+moqK
veG8aEXEwC5vkNY/WxmfxWKBPt/B0wHBofkZrTtRYGpOCqmrcBD0jmcbVCkQQ5R/kHYBvtx2yq2R
fIKcB1b7V3Ne9I/Dk45Enr88DkIsfNYRBW0wuLS4iJbzYeZPyMmD6m3FYTHMSrlpl7eEdTRdh5M0
rfWDyA/ZAnK42AXWm6ce2AhX+XtTqeJq0cZEpYcRBweNtg5eXzuHJiVdD+WCANZXJdqpQ6JlkSE/
rWC+AimYKnW4/agDvv6VOq6a3uewM7KAtWCu3OSWs3/pWRCir1r7hZ119OjVx6NGtR7alzlXsDHW
TlfV//eBtiAH2DSxVX3JXVuugARs7D645Jop5d+3yA50sJg+g6z12ihErUQBOu1oeq8Mh8YjsMXI
Da24w+y4ur6P3kkH6exzewJaLAbgrljyPC9jJ7zu+mb4DuTShUp5x2y+1HMglZinzAm3BAti125S
hbnsTUlfODh9GznxlU99jekLRpTgG+n+Vcf9I5D40AfAyKU2LeWbd+pLYD9sWqpXblJsGNXWdNne
pml6tQKsAQuhi9ftC97Hh13GWM8X50k036GuOIdealr3sSb+HL82ktMh0WLyGulvcDKl8UDbXfYa
dPAaQYngaWziMVbciCDGdovAfTRymwIWGQy9o9ATH+YiePAMW8mOkcaPLMowxQE+iki969qzRgOX
e5XOLXV7QzLgnRvZGrIh90ldkuNIHCdcUOd6yCWz8Kt6DTXRR90us7zUdAF0ZNb+QhkPJFZACP/u
Pb7ybhkDz5mJNaCMWi8D7Xr2n9QhaPeLzQUZl0wRTChkUX7wwWfVKX5ma+B/wrZLh0xi1Y0ln/k6
jeCcfmQyoD9qd7jX6kEH1Bb6c2Jpcq3WqSuj8tUCUkykJEYpRvt3x9jUFQQaeEQiC6mnkDaO+ezZ
rz9jD5b+nx78xlz/8tZJ5KIpfKLVqXGIU++d0nRPQCrN234Lb8cv3dVzkc/UP5uC15cdF03gb7Je
/BD7mG/kg1czRa8BAIiLPPsu2zwpVN8IfGTmEgHWWpKQ4tqwSKOp9YTaxHulKfWzzCFSx3dV/5cJ
8q1U5cAT6r6E9i4qFdKe0gHFQL8Dr0tR9NyyhId7cy6VCzV89jmiPr7a4HEqD73iRipC8GZhgMTh
qaaWaJ1B6zgzyHsqpBSPZ8pbV9lBjkn9cGdl2ZvZfIM9/t/AIyMl/LduZ+YGllBDzO7t8WTl9qp3
x30xrFQtf0AgdCBhBN8dytSDa+uhOIn2hwhmjiF8ZfLWBe0tQ+Z/Xp2LX9fQ9BlA84Qg/3a8zbFQ
dbJYeZDOch875aF/2P2Dj8Jn8qCTHU6A2ToVra/oLM5Kbtkl2nYjkz1THn58pofklFwonVbCBVr9
ljgVRfkxmoVftTQoCDTKpX7pBcLZbncoYK74ak+OQQD0GJ6rcxE59RZn2gfwdIM9TG3I7kWOr2VM
O4WcZyRc3kfni7JKtpaEKjLPHpsl11gw0jlZsJ75hFl10Cd9oAuD8YqeXQIEu1eAl7X0vlOZ4u/g
wY2p5n3ApC28xwu+1ExocgEydYYUFdJQ7qaj5cuFtLODEFkW/NuAbU+AaGscwuc6BufNgyTQ/Yml
cLISmldvkIjIccqSPSfrYOynjA/fDxMyj+D4rzgXabUehgyx35RR5tDmNZlTlB9VkNrniIq7e0Fq
wuqhn7sXB4m6vid+rWODSPpnZzan0x0hRQNw+IWhO6tQAcZsWEtuNVAT9H3C9KtQTaBjjNysvkP7
j76clvEUEj6lwa8hnUQZnTSWoy2PiHXT6PgkoyIPVYqQvPobL5ucwoz2aXhLGq927f+i3QqoNvS7
J88Almd6xydEex7nc+G2zWY6HG6OGboWueDuLyZoJf6jZ57gK4TgJRxDfrFjBkVgiKQ9QvHOXO96
HnPT4SvKc2EoXq4PrtmcImyP0IPmBjPUzZI44vXEMMm70Dz0olFSIkFdNUf9YLEzPCM6RL1mkDYR
Xw8BSZcCmkWkroKOf55zE+MJwN+NO5PV8MJkEYB2ljmki9ZVy7HDZKGhw0m/qKJyAFo+ESEWI0UP
+LlyF+bxRj2QB48C80mjjPbLTZrHyC6Wfygh6A+jvJ94oZZZu/2ZnyxGwBcujNYrdjRCfWTHJC+f
Ps735O0Ns5Zhb/KyyV3Sd3z4KWSIDbuIOs1Ql44eraU/LGBGuIOWUue7HRtLR+GgZZkXZB0JcwRL
0va0FD6dC1qRPGSEd5pIniiNYGGL3TG8/XwMWrlX+1ntuNguYnx742oFHxgr88hZIySSiMo3bg68
HIdbBhWSkpKl9HHjXv3fI8NJ9CyrwqxMsn77F6pquxC6N03ncIKLLytJBvSUrKcvNvEVeEcZQtty
0FqKOqB/4JafJt1KzTb06IQkWO7sDmFIJTfdrGKKRiVrH/k4RU0y0hRvA/2hC9mqjIQhzCwnZAh2
h9Txi/+2PYK8sy9XRbrFvTAA9IslQ161AegaHILh0G9aQUtSleu+pSB0OGE1XhvcF38ZzCSzdLdx
96her5IlfI9Z5eH35TWqAPn1A0GrKjMTOB9sNEH7EaWZYjSM90HMo1HpLfTwfrC7VwgSjg0bzVWL
iLIo/cziI5NVyUirBPXUAphJ4Hx6xZrWzAbHlOp4gL2vL8RdGtitrFYb2IuepNVjYUdNU4Jx4g7N
lEF1L1twA4Pc6onD5iR/wv7eEyuGycEIsi3jtCWFyFww52NtdHbp8SeAi9LpI1uqEOSY74Q139dV
F0zL1BupKvDHgfYURt5hVkOW/MDgeyecXMOj/qbiGkNEttzNhCRnPcPKKCgT0aAPVWaEjy8pFU42
KiioNu5DjsmlCJ7lxL7ZBEzcz8mVKZhQJtUsZ0o2pUIjdV8+2n/TVwn1kh64dqZY946p3/kBuuQK
j0vvkiIHkZnO6RD+by26I7WYgS7biLLqTEGLwYAly1c6hJxAdprvBJw7fURs4ntVoFx6ejZVSvHb
bqXC2GN/+ruNJRs0DrgGyd6Xi2hLcF9GUXUZDlutxbM0A2ZvXlPk9NYltpBXkG+CzkmEQt9OwQtn
FJ9hFKClttI5ckKzFLZbTjpuBsG7/dVEBWQ5irMC7o88lphucDhlNC9AiGdvgN2ZlOYH3JgdHjqw
R8IZpBkGXSe7dbEBpk+acdK3zUeCVr8PQ99bniuvXdhJFY0/wyNEMo8rQiUglLTvth6+bGH2+xik
CJWotTjatX5T3ou28U9y+wk6x9e/XyzrwO8qR9iu0i2L3xtt3FgGIzeec1E91nevZpvJntaB1NC4
Gk7ALk1zUT6QL6i5iJv+1tA6SHAH0hPNphzuvnLnRvIY2bIQf/5kRLlGbmQ8rwiI7f2icvymoUS4
FG5rHqqyOW8PxmJ2jRWiP6QoeRVNWAAG+hFrgY4Iqvg0L70hLAP00rsm1wYx6+79DXIt8A112RW1
AlIUQkuY3ZxFNzPFvICyzuBmVaEcWS4GK91IUUd6wAjiYHr4JFF/qkOJ1KVS9qxf8Xnu3D/b1gZv
q+beoSayoRiguX1pNHrlOBHx+dfLeQr1vk6QFQXj+qDw0e0jI9ScXguAaSsthrRu4L7JN5gfOXaD
zgH1K+ls0K9MWoPQ8Prk7QcA8qYaDzaC/m/oY1eAQUREDPflaPrEkinOg09WiQcJVU5epNJqFB5N
BY1WqH/5qC8KmKLlfy+YCVeJ/6HU+HcJ4RfZGXoouoRlmpGjPRrpizncT9zVbqEBkKfO49zrBxoR
jJkMnhvpxWQTLmi9A3GIkynDW4NRQb1oFRBgB6ji/1Dv0Klls1ubWDJlFsdmPu9KrPWRuKCAEoyk
eT7OVh1KQHVhr7qPfTssWhnXQBV3L7kAPfLH8aE7XJHyEMKLdXRAetyrZ6K++Dhkv1/B4bz0B5DM
hqr/qUbSpwbhtZa1lWQF3Q+oT96AFjetz7Qk+FFknJJoXoEMm1Zfak6IsZHb+svNFy579B6wNOKZ
QauxYkAHzpt7VYH/eINAPt7UGi/dULSw3cISq5jKLOwCTj5iyTtQA3HIoME1TnR+0jGUBWJbbrwf
cyndLuRhkOgHKEP038mJ20Kc18ZL8wYNOOx/QLMu7Y4Sg4u0qRfByUg82cJrh1MsQR0+oCT/hObx
Tz5urwEgh+F3VULyIHvhNqvE7+WFfxTRPxeB5KhuhM/dvCCoWAL5doSYAlyZcnbN+letjv9W7+Wu
dUbicIbPoMrdBg4MVCY9v3JCPVAi9hCy57BygUm04HPoc9VC5MOACsCT8RN1U43pAgvbVi3nhylN
9grVVg5QDqzaTfd2e7vg6C5Lcj7tcc1fk0WexajaxZmqFbB0ZyP9uKP2L8VUp1D6Uu+biNU1erG1
8Gscks3qYRvNbphzjDhBB2TaidTAdr2n4hW6cSooL8X36uovkvrYnSV95eVabmhhAPXIi2qForTN
TqHrfP08F+JZFkNHwn6X0Lar4onB5yHtskZ4TwF7jcwnuNZrbCBLmZ6H0SQQFDjNxuAdBdk9xnYc
Y1HacKsFucq5LcKtawqnkBt1nAvR/Vx4p+poFyqzd4eJnu8fee/tp7VDFoHw22k++s0l88cB9hBa
peH/6Ke0vDC6Hp5nf4T7ab44p85SHe/InGhP4AoEQu42dtPNIikBW20sTF+ReTxoSu+lCOCgPojw
Fnu39LbjNWrnXVWOXlELXKN9FM6mEfWfj4xh0xMDSUYROYgMMvG8u4KHqh9iS6kr/NNYdGMwNSxS
5ZqhKxbBrnVzO9pkT+6+tdDE0/6D9y1DmZ1a7Y5hUxCzxNCi8bT8rXhBVeCEcBOgHVVUAHh0Hfof
RwoIwEDOGxhHkNhKDW/27a9eSu2KiuOqjxQAZINpMYOfPqY7++gUS+oiqW2IVHcfBt2rNHzcgIO0
ZO9xjoAZkeNrlwwg4++l18NB1yHp1VYWTPi9CHutWHb0cBYBVOBmbZYzPqoGkZlJCLLH0Sp8FhQy
RS1gxwJ63JIyqqqGLraxYI3FiTL7YBo6oouRLigqL0U6UzhanPvCchponEeXI0ECr4u6AvgB5Vz6
dSL3o3Mehmiv5UGLiyiJGNB1Ji5B2v393ZsV61vzTwJufX0DBTIq8Io/h0h2Un037kn4JabUlj3r
gAETzNdNHXaWmxfdkviRTs2rHqWIzUfTQIlOzsHOQreeNZIfl0WX4ORUPhaVW770QbeLfYk+hqOS
hjEZA+EHKuMt/WgODlSTNGVWHW9ddG+T93vlIjxSrxzRu9YMgcA+aIqd6224p4+zWOz7M52GI6dk
MIhXnTK7McZdTiNoyw3L3j/emdBQ48pMcxayNhrjxjbJzOkhzfCnarqcb2JoxwyEAYgSKydO42FD
p/FXA7MbAYIMO48WTpm65P1AQzmBtrrrn+hdv4zzhnzqrmFfU1pfGqG5O55Ma+wvaoKJzy8fTCth
j0er8Of6dM5oC0PIRw2QRpo9IR3KIKK5y0AwhTuKmgvFEvSXUsy+Vy46nL6eovoCMb3XyN1xAMVU
+Yfzkk1OW4F6MHAL5Iqf4Y+SdY0QKQXWxNWQxpspOOQ+75CSPfpVnfnrDZW6S2esUbdTdGSIoaYk
B1ow08FTsLW3TeCHfDoTHjQoh3rGU8GHJ9RAnKW9sNOsZx7FUhy4pMXn6IPL2WMy7Xn2nVlztocS
zWjxawV/NKwghzvKXCloQz4wFe8mqpyqyn/CH4u+rzOsVj9NP9pB91UsVGJLqsKtDBuK/bjO3mTc
muUPMqdSZVE0ED6wYZvRoiNnKWt6m7ChaPmQ5YMaFYzJjlI+52/aPNTRGw0KwsuM1wbcuqYzGGan
5zlQmlPULl1VoJ8ajpcB6M4d1b0OmyJWOb1veVSm0xpl/U8RqzXG6ztOrUCY4nGGLgeVrKVrOfCd
YP5eZfct2bY2n0I95iotuEMyMJy9gaYznkcXOXTkckizaeu00kKJ7xnBUITPDCToPWiZ6cBjm4pe
bY1o0xdzoVplqWd3RbRrMbuCz+vMBDJfig8Cy/cUXErgm6B6I+6uGU44WZqd/K9/Yv1vMmGeVvt/
38KD2E4UK0CFI9kXIqprfD9XCAp6QZ+Ul5Iy2os2Mt5OT4O8BrGLul7lFsTX656RXsV1vBa2ZNqC
v/9V1SeizznlJMlniFTr5iHCt5gXPiezSN33824JwFYxW9LBM0oTU7bCfq16PsHrED3MD97FWwvV
8dU9diM94aV0YiIptU0eaDL0q1FxIvmHtamJ/zg2RsfrMIUhUtuGzxNH/6Fw6fai7h2ZMy/xpKgY
rjuwHNyldDi+WCPpZhR+M8x0LIRBxv80yIQc+pmsXzqzR2hvHuSdBs2O4lguw5YWBU0XiJZR7zib
LC+zSvIhtiX6RQUkrgeqbWr3+C0kqbYQtVaq8WHsuczn3gpnba/MgIEyjtaD3XU2pVmKxxuWvAUu
ee/5pFSgirCcPaehV6HiUNlHMatEMPlkRVS7wMTU3T0KNGTOlQUtv1N7LxZMqz0Out4mHe4u3A3O
BKxmNYs4TlQKGEdrv8pNAsrPdxlShWG2RVJzJmUwzblPfgeFn/u9xrweXjNkATF5IcnJnjQ3jIDY
A3dtR23Fku9st5I6v4W/90ebT/4Na4tCKSq3lmjCNyNh9ZCN2YfDroVgtLswkBK/mEvsnBhdrhGA
b4Ip8vq+AAaKg3iSA8L3jJ50CXr0z62Fd6yezWRewSY1OO0XBMg3qsW8VVf84YAnTJUJ/APgXdDF
2EzVX8+2s0UEHNP5T8oXp/ctp4csrK7A8LKA8H07EsEzTX0ge2eGMEL9kFBdc5/ukFj27EpHxxyn
oew9Xvo0jPe5/GAkxO99VwWt5mVwl74MqbsdRRLo5S8hsFibEHY3jXB+Ca8qhTm0P0k41x8TMkSl
8sYFWPH2bZNVShNCy26P/+n34nTII+uXGsNa0bNmYxntspfT/dxtHWj4FZUce55t6ikqexCvNuZw
UR85xfKfCNcVguITlbt4/1pNcW3/pMXJPTrLvT5j6lsDL7uk5qw7w6cROXmd8zkwLYytixeCWkhQ
yiyjRSmZBHWv5aSKLE53fPLL/MvSr+7gZdENB/bMxC3nqrxMiovrS21aplXNWK5TUzWmcZtqilrR
kdbvFWhur4KCH1ZRJxAdRJT8wv9aHfVtGv/MiTC8mU+hurpnqe+qEJYuR5Hn47giu4M9KkROEvhP
WZuDJRqYlX288UCjmD3iWL+gj+Dhwk0nBWmDptHeQrtkcFh56oqjCbIJGm4dpmLeqA56T1oZ9RQI
wbemHzXN4vusZWPhJTx36yjZYX7wMnrkQAUOWxtQewvpoYnAiMPInPoHF3DsNXZzNHJXd2M/GAOG
5JyGNQtWOQD7sRc5OSwQGZM3YvtixrXmxe8/SEcNItE+vk/szqF2f/WPqFDeMcIuLKIS6YponymZ
oUyyG6Ru4LxmVZpeaSvg6/SkSArUIL+NlqwL732x33vfOelpsoGgjJPrQ6PAVBsn02wsd+6033Hk
KunkK9+2B4WgN6Ffi6Esy00DnboxtYB6daybAzMQjSNqfkbkBK6TZe3iqPlGNVjxhPU0q4Ln8Jop
ChCDK966rEHHXeiERqYnulMfR2XRk+OWLXq4nalYorGy43ioFwW7LFCM0NjRgMmE5nd546KKPliE
lhzLxaxb3hDfsIyJmfwkvtls6iS7yWACMWNF5nIT6uJAip9PDFpLZr5JF1ENdwDxyHvTVFuILVdf
evt1i+4OLFGW87dzbjY2VpW5oAYYRAARkT/jER9OoWYy92wFVC9QA+mGU9IO8pg50ejxfUQP+49o
I8Z15i9gOvfBGqleU6CcfpiUyv/qyxiK8R2RWKVEDgFONrKht+nf9E/W4T30GNZNLJ+muC/USEU+
gYvtTDoiPpLcup/RyqxwMUaCQha5NFtjlEAQQYjvq7EqHRgwRSapZ+ViXrjiyNLOCuPdQqOueEsn
CeYcOCtbiacaNHrU/6jI5zZh5Bv6iGZ4uoJM5bEqeb1CTSp0scjojv+FK7jrojV+3v5tO8Z5yUux
r991w5ThAoz0ZI9dr+Hfa/S+jsxJNt3dlJekqrsSSHIhnygRI68T6dL3CVPtkC/W0rjGM1QRjAoJ
wL/Ghj6Gu6coWjztUOD1VRFt4ZJ142INnQoYV2HgQnpkk6/mxiahl3X7+6mkslK9sXZEI/EuAhAk
Ej7x6jDLOsZGDD153ySiRllBUrreHRFZ+ITtRjrNC22AWzmvQOEVe0mZFgAqlK24cwfgbC+WINUQ
ngdiFRM5CPXQsKCWC4yvSKfZszEPhi/Z6KZfuqEy8Rvs2EQcMd2ZBfnPlOXYm68uQbUKQL3VcTYT
56VXcO3W8tNEHMlZT+YMbSJWgqvfx+VBbG5DyoFjL3tBzbyaItB5qbn05eF1Ts66S4fjtddeKgGw
DFIA5dOZ2mCWLB5gEalMqN/MmA4NH1LlFuAI8+YaAZpno2QuXnJB++VYqMta6FqNAszqn23PqiQB
h2ix/Mczx6lSx/4QwvVXfZtGqIjNfpO7FnW51fzp+70qphZdQZbXullgfSkGoPfqCHy8JI5ZNw4c
75PTv54uZ9tfZsev4E3Fvua1zYKnZY3duJt+Dte+RhpQ9pxmfiyOh3TGba/rui3rOpTysJio9NlC
v88eHk9x+GxSII6RTctVSr3sDFEiLIfNX2ZAR4i0PSxjgXBoitjuapst7VWbcG4ONaATN0UZAQIj
N+mAdpZgCvxLPU26WHoKcYROgsKfLv+fbB4tJ0dUlSpHDrKh3XhtBAEAirkfraXvhcLGmmYJ/sbd
o1hfiBxAibr1LuuPiUXFd3smo5D9Xgr2U0OiuyhlM0gAeot1hamsJO1jS9awPOWH/QQVgGxC4bmu
U1AODK9+bxW9Pjev80w/s8W8nqSQgWcZlrsS198e87z2cCxZDCpuPH+49t9bPid5x3lXsndKXJuD
+ltJ52zurTq0sCp71UXjsvYVG5dmE1BQvN/T98F/nN8uLEtvGW3aEnbwsT0NCqTpD5cqJyGaJW8I
BZnAa3+ltvJZX0FGmNldsJIIALWh38WuShnjqhYmgKykDMZHN+DNRXSziAtxgFRW7uakI4MaHcOF
aCtirDTEp+zskP5jPBQkDF9+h5bXkpmoXcVU4RNEnuPIhjngZEPlFH0lTnB07g9sj69sinRt0paG
eApsIMefYAIrkA5tOQ+7hiA4FHsBotWhJrBRYlJ7XS1Uwt9eqHNZOsQ01JCywZV/fLl+/kz7vQDW
oB0sHdu6RRtFvzLocgzTBEphGe3DwxcgCPZV2HvdN5EARAI2D/yjR0MOEDEgWmo5i/cCDpG6yHnO
BcfdXF3HRarBXJvB+f7pzPucdMNLyDshJlQUi3V4Wogunw7c25nrvwxaD/zS3EkaSLqRrWZcV7aC
40qH128v5allbc5evZmBoOBcRWO1OMXOmHmPHmavYvyrooUDSg65qJzR8oYYbSgbvytGICFbfo5b
5c9aFS2FOou5hAvQoQ5WrxLM6G9QUIqi+qgaFPH3SJMZogIBcDcEIeiGmb6eSbv2+/VzQj44N1/T
YVbqEkXHpHgZ59EpJA6RVvDOpWe1+eprEWvWzIqOvcCl1d9709qRZYZDRVB23qaUVYWUFNIuyRp3
ZfuhmGbO4BIbn8B0XbFLAETeuBmUusHU9IkXcPV7NaAdX1wbWbdd+skEDFNRCkberi5LJRnsALfB
ZUfxhv3DTceabqPmO3I5RovOytW6VZX1cL843ajpP6AoDu7TLuiH5EexYtjCPKh3yLwy3m61XaQ2
N2ci3HsjnjsU3ghMuP6AE+cv5IvZkq3PptoN1zCIPPuEQKfo2URXhutQ2hc7yNRkJoWNztQnBZHD
vcCMio05Oin1sV8U8aENEARaV6O4GqdO05iFv+vm02MQhl13EhvM/ssZki3YIyu5k4x9gAWSikib
ZdVuMWyvSc9Xor2gkNBEna6huMxuwcD1BAhyI/Ong00H0Wo5fxZYCakTbUMqkfCeskgQZWW/+pVm
rdiSJquYgEBi+KkjTOxI8oTgarVuTfseyVrOoxlZXKonYmG0rntVVbvtC7VCrTKP+EMe0PEeSbFr
Rxspop+laYBEgXUJUPNV01TL2wH+eVIV5OfD9j1p7YNGL+qgkcv9Yo2z2RPKCD6hFPxsCS88n0E2
jpCuqSF87B8t7I1TWJ8cvF1Tqhol4IR0d1xhzc3vjzjw6eojCUyFrJxpBMjXKsJIaD8UG7mC/3Af
6zfuM/wllJ8WuVB1EesnPXilcA7E1YGX/2eBKEmeXh7q/qi2t3aO7/TV/k4OJMvfe+FCktR7XMYN
PQIdfGjtWLGDWtdfqx5VJaTPqfChqtUNo54tmXIvBLeFbDki9A4Tt21+mRS9RmzubgmQ6eyf1T+b
HgS40t/Xq/790Wx3wFg4QDSRHf/ftKJIoBAeRBUTJAjxiyvVxu6HmR/BOxprReazOnDFW7K8WPCE
aFZvhiaSArIs0M8LhxtvMcU9qUxakEHqF75Z1Fk3tyQqzQ2bWCzwzTox1nietLv2uLgQOtuh6mQx
KoN28v/6mR+Q+4ttsDSz56b2mpheNobSRklthlLjdeZ0UwoY4Q/MRM5qnX924KDw/f3r9kajBgg0
LqknqUcAQmMxkGLwnhnCpFCWp6kozIBNjv1ZIS8/Zz4KTypQKH3jqQDV8xxnzcBs2jBFERRM24zG
oVoJlOqiq+x4cdrKF8xev6pJo1NNIyoyDR7Ur4zsm/X/tphYhVydaav7wn8UJ0CVdYgc0Wdj763Q
XBQhzAFCnWpXP2kFlkdEGR7CHLdSw46p6Ju9tDTMk2POfgy18DyEFJ3K4gTjGXe8zJFS7VxBuwhr
SLaLZgfWHySGsVzzIJWU8M1PMcx+qiP7HjF2A8qA1dxwZEBS5oZto/vVIdp/vy8fHL3uNLq2on2P
HU2aDLo+AaBep47zQnsughLN8ZeGMCMOTG39e/eDNrFyIam8f+l6fpt90v1zQiQ7SPhnkxYRB+e+
hp6J+gdLLU2CWMTnrfdltDCmuTXAo4B4/T/FJh8+Xk4OQ/bFPRuRlR22/ElCKZ12/EKTqhRDDV/b
3RqE5EaDf+44RiqDDQczAOP0NZRruN968ugvbrRCZPPoUDAgPk2HPetMQYBcnAvJHlMUdTmQadG+
6QI/b8WzqfpRK0NUha5YTWbFAlY1WE8Zsim2c9lGuYm8MFt/br8uvSmMCQ0U2pmqpY9dBL8JVvqE
ERZOQ4dLda9gr8EjGEf08SCj2Pg8GzfK47nsu9Ob/GCtTEXrvoo2bmA1VX6uzRhR7ny/Jn4XTDFg
mfvbVdQCI1QzkZe6WsGyoAlayS1DpP6/9Tlp4C+jpIT5sYj1yeuCqqoDWLoZcOxOTJXzfuuEYzTl
Jm6w2bQaIEhoqDXZ865FIHMD1bNNlDtHYzpeRbCvLiefFLLfDEnV+yHGcatcG8U58HmhJlZcho9k
1SdF/OE9z+T7nEFaI1JT79DO6seP1UFsOF2EkjGDQFpIWQlMrPD1EqaqD54EK4OxK0FuZ+Vj4Atj
b8FLVLx14wD75LZgSj1pW5cLSRwuAePOhGPDEOVgiiEgniNH2mE7l477QV3m7Af1ZfkCqnRFx/Dr
1Z2EGbVPblxBI4ucPAgNVnVabTo0/O3kWs3h9Gx2Hfja4Z3vkuJCirWtTzEEkLBCEbZw/44KufWw
hsA7pqimM7KFrHUGQPYMzs+SuPesK47AJI3E7x2nnAjfDLck1l29XsvHgkvWk7GriA/N3ca/GVa7
ddD424DGDzUWjaOyleg5WLFKxG6mAiUE5aTvuFOt2wwFvVRStCIawBmVmzbAIqtixj6ng2XETZYs
MOUPIOiugn8iZ9vz2WLAA2SXXlOsXp6gOwNcZ6lejbH30oFYOq/HT//6/SC7HwVm6L4Sw95Ruo54
fwIaKvsf/GtVCMOM1M6u98oTHzlLdH6ZyZBzXXWROB+Q9YsEuLNckd0yOMWLodO0O7Eb1w0iJVFV
SZFk70v9FYcTO+EpE4UL9ers52X1OUvrjV2fOmjeYJRf1BnUJh22hfkGPjrfNZrqw22+oCc+fl+H
TjFKeBaa9BkX3qudLe2UvYyJ5W2TtTY6ni75YLmQ/ozlsh7osA6TR2hRFEZ51lQfdOn1NPWY0h3Z
u4v95QAeW+dM4+3XgSiXzcp4BDjPdwBQSdepcXkrpuUyFiwkRVfwmPomgIdDWFK3v2PH/hOsjOtu
927QcAshSBmdY+un1/zhrlum27vbV7ZOofS1/4huWItctJpBnOnnPHMLZ/DJ8dCNfCDpcnd380zO
09PRgwgMLmgNN3JG9dzGZC+jPEvBQLnm2SIPWVXAQGpV2z9etCqXJfdIAO8JGdbJhz8kijIWuXHn
n5tNegfPoarVIfgOJSiBlp8ARC1NbOd3xjYtjVQALRFT3K/FCVceHnOVMCTBT3HHNBmBmQaGuofx
QzaFL2ifT77bxenmU3CyPcxdsUIjENQf1jXOeMrr+snFDCiwqEZQ2rVtwUvrgyMrzt1HLiw7IJV9
a+c22mHv6WFQdkMTFP5RcugNiMrbZol4/qS+57TfgpzpKdTMyTGpbdBh/Afg3IKHXbm+WLLY+sY0
+qJoJe/xfZmiCk0SBsEXzMQE9gZX0460bCUFxhCwexrkJnXXKosPIT+gVBDJp9nGItnJWbQZivPo
/TK9S3lGtPjglHvj1atm09yxQI3FLNDOzKH0APblFNlCuSlZpbocQRACCW2uyBcqCmqmzl7b/t8x
Fb5j2xHnzY/hQmMlu9PE1bixNXK3yoPX1SraYNgyK6lPMQGAdpLJ5+pZOQj/fb+ss+E4cmfNomDg
AZ/CEAWSkH6mutMBdU/WsfGj42ULJuiLAFKIvFGkXE4YSEwavQSSoE+VCXZ4sqMi1qy33G56188W
CP6zvh/QRRrWQw2adYHLYWdD+0z+tcaFlqUA3r+eBX8fL4XA5y5hfG362lpFvQjXOeyK1qr9yrIV
IwZhlxFxFxwHA1EFFPO+Z4t1I717sLaoGN7lO84tBpbylRSmLdnNqGalp1y52TRWjFsCV1UaohNg
XHSmCiZ0AlI2TnANwDHFHLfpEaU7+TqtT6m33PNUcYhFiSd7lOdUM8SipBClnXmMLWrmQ3zgHq0H
q2Uc9NLYCCLUBbiRcHyJ6poGNz+vsFJ3JEK1EjLPwFW+dY1QTXVVCEFvkCT9P+cBUsrc3BxSGWOV
0/TVhxF4pgcznoSvHosPD0GalFm2PSJKmZ0ci8jgmxq8GFOXo4WiXYSqzFXPkFl3KyjpmQVpHwZG
Mlvfr4Us5O4znPMNOp1Xvd0Gyq1SSyBMiTSEklQGjXD5W57BIbroaLODfYLI/rXN4VuTB07mT4+C
QXyGhHvGiT/ZY4egcUXt1znBNZSN/RbeOoASOgLrHI4jx0By1ZEWQ293X3YXdeg6IGTBLcwGWL8T
izomj/OUFeYGwL+Axl5XOlz2xTF/jQnn/GoU/Hn4kvXiym2u6MTz81Og7O+jSK3//aNDY3IWpGim
3UkgvGqTK83ryPDCd4o236lfjS6SXmrgt0q9HH0UW6Mnh7Z+Rk4JyRsbMfZuOqNZNvh7BnVAqkBa
15LSl+JBH1sgWR9Kmi9ZFt7oogMvKmFWRWW8cgGxSqOTLCxQuDL8P91ym1csB44Mc29SO75OZWMu
GM3x9O2jUhB+QaM1Bc/qxpM0lwX13jOTCNxWuFJ9qC41T7PeO+T7OfPiVbr0fMVw1zxf0tg5jtku
B0vdUiyR4gai74iGNb0pD5PJA8NwLx6yPFNGkNlVmvaufFNg4ToG8FbciD3f6QUgeMe0qf2nYsJG
Y+6hfcmSXn3mZELD6dimT5tAcRNPZeDzN53sjeR0OcO0ILRuCJKCli45JY8L/rBtCnPKxxKxFV29
iTI1YgY2qGKkdBE8NVwws1blkD27qrkUxu3bsCcVGBx1bHf3byCWlK/oC01wrUJkyZJiIpIiagcY
WbNUf6KYqdMGprLvOPCRnwi5+Gw8couUIJNC3w6o3pDTOvZqUmOR+g3hzdEXjsb/5WCLlH8/BwV8
4Lpyy24VADAYelF/LWT9kd22GmQCVf57J844KiuCEOZ9WEwB5kNqxLDbeETajxV+gduMF+4P3bTU
sPmwOAJWqnXqWwXiNH0nCOccj1vhFVhd5bGRIrLH6UsPcGPt0pHVaatLN43za1uhHVaY05W2wfqN
GmElD7MXVcV8dlDAxZ77eATz1CH8T98N1Li1b9j+d1KnAqzGBEnQMd6XiVDxlabEaQNSPxgT/Hfq
1IMV5NA/4xVE734N27G1SnJ9bfifCPcmG1Nxp9GfOhWtjSCk3BMWt+8Xa0nLTL1HI4ocPChxcwx9
Y8gha3HFM4CosZAGVBjlovQdPg/WL8n125NDg0eIsFBiZuIonTMwwzGbSpunqgSPrR7OVwdFmA3u
F3QD7laSYg9XSsnnkrHWsbi62YS/CL4jtr6qgUy2i8xksslcZE9d4aySIMR/OWARCcTihCc/OEjO
eyp4V/AD23qqBRsJCKFFMxYKDh4xWOvKhUekRWHYJsYXHNrxQqHewy79jdGJIq6xG0vX2fLSj8dT
0ZcrHM3E+4a6dwhSeppbiYWCmCe//P6tNiN7S74SzJXLMsmOMAggBs55ytjZ93E0iivlKU8dfGFH
IqjcfbAOsSw1DW4Gj+wVwopEwXYWwW271gjH1BzgbRsWs3xlE1311IzaScH84FpYbf8sWgdfHOOd
Y7WOVVEDbeqrgZ53zoDwsW/mFoYpZ/B5q6gruxQQNO4DqxDrLbwoHjV9LHyQmS4Tds19n7un9pV1
hv6M9WrHbvdKcln2BWG5HzcY69HZwbaeOBtpwkXkOFtk+w7PEkTj/rgcBYjHu2mkowaQklNC0Jx3
uO8ezP67YPrCZtjQL3uc78PLxBoHoEmjIqIfF0QrfVOFeh/szWkvJ0izPpqJ+utXeLTbhZs9t9t+
1ME4O/nOBfVhvXMFdDehxZseWEFiEadjdU3o48OhVi8Ro4RUXOonzMQNxDmWa4CHae/u1fR0uhfJ
ciqT4tj9qOZ9Qh13CjlloC6ZEzsjuTKK55a6VHlOZ500//Hm+Kf9SJkw/rJzV16/PibsLw1YloP1
ALzmpmcEYziJcrlM46YcmOz1hS4yh2GpaBPSp0i/Q8u5DOqdZiipRktdgOiQodJfjJlK39XuDQqr
VrVmj39tczq8FKhXRJVOb+f9R6ZcAoIS+sE0cgiGtriobeUg169YRsHK20V9/Cm5OcC7ubNenSjW
f/pquHq0vca70uEea6w8KwDg02nq9Wnpx0S5gz8d270m69DgSiDbwzj2Cgvfsja6+eO7Wuj86HyR
vHBL4mO0l63R/ursRnOpfXaHHVqPfW8SMYzancBrnqWF25ksIr8E3wlxuMOYInL1AyJy8nKghp+I
icO7Bk3Y7O2/W683c/b4m6Sb3kno7KDmIJ7cWxIVST2U8lilukTRO/ybwym1ZVjbfgTnBrRYHDcg
XElBhpUUAFiApcf8aYiFdpDL9LdIQo7W8ACx+U6++ABMNOFO3nqAaAuhxRjx407BlO7sgiksZggN
HB4m5mzUUskW2Icw0vo79/tHLhhgIlNfLAusWZcGBsUe/DSkyTvgF/VIkeEOAoGo5TL+cq0o9bTy
arDBiVFaYIKfe6yTtazXaHmvZ7FzThKVyRuke/KOk1Kpomw2ZwIS9iJyDwhARQIpdXRMA3Fph4cv
tf+C8rStywpxEcOmxBhr/lA3M2ZNrAHaE5hNRf4sVtkaipVS0yJe6tmo1vERIOV4XKGcghg+rDji
Uv32UYNVSLmUU1DiRAADSUQ6mFaLkbbisHJc3TdgaS5pkuzbo7Bfv2DIddy1C89t9awvaWRP37Gn
wKA0OYfBWQRTgVc8r4UFb/m4QdojMszF1iu8k/F2/cU51fZlQ7VAlQlRG2OHWaVa7G6ApQK3jqS/
DiBLHHTeSpxDu9hyByaf6wI20kMwNzBqmncLKkcuyB0V9qdkzo9e6d9mVvMMI9BdaGWY1IkIwRic
h3v9jDYpg5YBJkjeR/dJGRkyk070K79wXjgv68f0LTTxAJqPAqNJIXBqvcvwywtyi2LR9FNX7k/s
41vdvjZmIsE/R843UHfbM4iDm/a6UdUwr9kDnWUIpsjuvO7+7ix6m1nznR3b51B0LFeySxGkBFgG
pxW+o9i7SXQyCVLGj6G/czRZGYXTZ5u55ocz8kX3q2vlQxr9J9lJ8NPm00XZ6AziM6ecFAUXEzFz
MelAI+Sm33vn1Wev3LcDn8r0cQX900/grjH+MEabm4zZktLt789deMK70nP8AnMiaTyyEhcmZOOt
K0yMCreJbmeihgNKM9I1X9wBc+UzTO3mBgfq3LeY11vx24P+VRoWHgr3PE8c9e3rez7iAdtpj8C5
35Mc/5zhegQM8t5bhEdZoC+W+SqIRPNohW/y7KvBwa93iXqsb25fsKcTPuijfbf9r73vlY1Ztbiy
ln+BbyKJ/WKZyq0GHO4jC93T+nAVItfQ5Y+rhWndMac78phxWwZeS+W5+9vzx/vv1kUkAH/yN+II
0EHop5bkZ8UW5DxflkpKsEhzH/1ozQg5GcZEL5OvHf9zeFsPjFqTQHOuJ0B8ir1W4onTGGIPRgM2
dEXivCgu/D9X2gW+DI1DC+9FWbOwkQNqdYyJ+pWXmFjrU7s7ywMQDXxyLhQfEND9ImIo8NNzkNvz
kuhrGdPEyB38+wvukdCmPMKWpzfnttny0UWxiVshktYqDCU5+oNzA7zJN2LUPr+K2iQATwSj0hOG
/pAMSgmJdX9AkQ/iUsmmhpDPo9G/RPfMSetfdQCmNWZgg6a3Z4rqourn3ZbhHI/Mql0NIpj0EVhC
ymm7B3kiNWlrJla5bRBD4k0BtjASdKwaOz9G2WDQAKu/BOXbpmH3eomYysIDsJDWYXorme3XlsjV
IJOseW5m2jEFwX8LzHz/UamSAp6p5oxvO9fD1VljuH/saGCdhnUeVaDBLe65LDVZ7FcF7QaL+jC3
Wnhaiy6VBCcJXkP5k5v9PnKsc5ZA+U8d956z5JSCu5eaBtEdwwNUitzJIoc/6VxQeVm42i0l2c6M
QlHfRv3wCuehCWJtc8DKx6/tTfS6rIN9XeHhMgkX8z2z58MkiO4Cwy3iinTAQb+2WMv2tvIuITZ4
TSPV+mW/Rgv4pBnYfZoR9GgDcpcGGNmlo10ivcN8Yy2rk2z8xWlbZukk3IDtcZON8A3GNBiAOepF
ll7nIMSpEWHn7Gjj5NEThF6o788/MfNKgFd9dDerN4C4TgpyXw4CP5bO9G1dT4CHeghkKk1JAXr1
CtFJNHPGg+oLSHjjInNfnWajnxswEnvPbhZRiS+VayJJK/P793ZdhNKh5ZZTM2lDY1u5Fy4pf0Af
86sCBaakpeKIcIBDlYDHRXP5Pss6Qfxd9qd9A+pWJReq5kvaHXCnkPONm8xC9CBEBUoRPaTaAkr4
aEwCeciR7pOZYjl712jXVrIu3UKS8MvjftuklEEGyXGVKMswNAF0Ct9mEJKk0mXUnEG/YgZyCM60
Erv/3Pn6FDig6s7bwnoXkWACnwzvTRYpdYXgtlew+1oSqqITN0Kb4VcfMkB1FJO+5Z+zSHcdndpR
bCIuuyshV6A2f3euAI1XQ2IJtyuraIfUNjjteKC/kEYWyFub9l6pSoiwu/jsbjP9nlm+2ZUYnojj
TC+IA1gTLTOOThYq/txpweUFLIin4xhFGmXLvNL2xhRaLG2HkL5UgeZBsImh9d5DRerW6aa21zRR
PO9sD1VEDFOJ0y1U1LBaDc/Wdmskk6gLJ0r3kvtVKzG4WSZ3cZ6zRhzYP+EoHwv+AQDQ6mfJ5AOf
tUt4WWAclP1tszN65gTBI+K333yJ4E+UhgyFGmA4PN5vDO12xyjnFDZWB0u17U525ZfCE62ytB3w
cTkc7xv0shBBdlFBxReDCasHUZFvmizqLU9zqu+FOE1/Wm5Sc2+dKgIjJzSDGom9wpXcXuYjAKzB
3DQkobrNa10L9jYndcoR776JdpMOSz3Za8QtbheY1clY9Nzm6287/EDleO3ZHxbvwHYYgL74FE4A
ul0Yj4UObYx//6Hje7GT32cwaxI6HFNVnElCIWU34v0bXs4eobkwQ7dG4ciNmqU8eqxLqu98ZSxj
tHMxa6OLCf4bGwuy3vu/i+MMNlVw16AsrOqtDIsSRravkYQAb3GPRZLmXCWtz59ULzS2x2WLvJYV
0/LbNtyl5JXqTFAFAmF/BQaV6tgv917Qzj5V0tZ/FYehr5wexRx9ktWAYwiP/LlwuCO44c4YvL1i
qqA/GcO28AiDYbpMY0+MxeCbznmJ+CpD5AbY7aP1jsKsr+Px5eJKax/+Pa2ntq0ExFn2yILC5K7A
3GlQpu/PzG9Tqq4yTKQukH8t115DOUtztCq79PvbDjJqQXvSdaD+5XBQazsS6Cpbbwv00Fvt6zJ6
BTCPJYq7YqTwRSEOJftEow5Aw5+V1DGqzuvFD0DEqKflocQ9pL0+tikq/ffZQi7MMAfkdVKVP6O7
YaFFU6Uxt7oqvXwWKShR+//MYBwZuSNNejW45tBdns8VcL8zw31EHLmeldiPxa8ILysnct3omFOs
Jp1NJQ2WImPsPbb0p8DFT7ai5fRC2PpUwxJ+L52lwwQuLXC0SIGWVwWRups1hzuU6SvLQp/W+hL6
w4PZe3AzfIrPkqM+CXViT+YvzYBq2rvZSjxqRaIy41VVTrADn31UtJ8EZpYnxDEAttolfqpenqX7
IdToih4auYaQNqsvJzStGDwpVdouYEnytA9fLm9INmJdS1XunJxH+TaAeGiQS7E91xT5Y1dsxqm0
27iEOIo4GAbhBEVjscFae+pmloXWwwjRsaKtzCVimK1rGgnPuJ8BZP2und1z1DCgqiPXGyj+bjp1
33bk/SnbwOoPPWRKxwJIGn8gUGQigifQmUM5cZXMwO9yXDn1Zf+G1ZCiSNB1Q2lTKlq+zKd1LwbQ
QxF6dLKid4n2IRir2jV+kPVpgqERcHU2hsNyDOz9wkkIQ8Schw17RgkjylO4aFP/e/NZmzwJJlfO
x0rEL+3jP5iefr77oGN+3F1dtn+JOFUZJy/S83jmRkw8jneBDQmMXlb0D7h21B8cGcZpQ7fHhVd/
llzMEPTJzNeJ0qUD+HrXn9gx5XkVjSEBL0GIwHExWzTfprbtjUiNoPQCq3Mj7soXYh6/gMouhf79
qnR1GMKrgAKIwzwBEVNTtGBDZacrA2OvDLkEgwW4GW/lfQmKwUmKGmNjcCSmcOBGzHgzyvYSV58n
dxiodFfqTsWt4yY/GtwmFU/beCTPWn5h4OACe7XgteUNqtLWlndVw3JWcPoqvqTq4U/7WpAYYFlY
p/utllIQYDUpu9eu/mYVwPK+/74O82/N3/AH/f6EdA/eAZL96r5TCjaGUEJ3b5VyNPg3v2kFVZpA
vQQK7uhzOjiokHTCspJHE2fePWFmV6pcdHKlfTUrWgwqVT9RIHWd1KJbia3Q7xOEdiaueXSOjnpc
sx2hjFhMJWsEFalh30EPCbfniguCY4GBg80yBbUvjQrLk83ve/GZO4QLLqdLyc4ygU4FQ9aCaAwS
QsV/4m0n7bF7lkzn8ro2IKxsenZ+VgKIjlgeXffn2xepPcIQVCQg8kyO+7PNp5IYzI3JOp1tfZZ+
DTKfyY3YSVqfVSNRTsbZDZ0FkfUj0tCaSxnCr8Hp7tRytRFxKp5IVXG3aFZkyJNxuGWbjGv8wp3I
LMfx4ln/hpvKt38Upwymhr6gn+vl9c8osZwcmzgGn+51EERXZ4Agpq88ZskBqJtIAzPmPJn66I0F
0PpnvJ3wksv8RsBwAQYKMKDQOOBm6r8Y8XI2mOmW8zc5d4UiDW4PknCOYCGCFN8ETM2zaV7dWJwX
dqd64jE7WSx/4Q0ZytA4TM3ijV0Dxbdi0zciid8XT/KvsN4+4mfQBTWVfgxka9RmhERNiU1g1PSJ
K0J2vJcOZv2brFvhtpnqTb91bqOlah7XDpcSQEhyQsrcuVazGKLoMoPai+c35ga8TZngeg0wSUUj
xFyk7GDH5eYVag0AEUUUkLMPeeQW/7w6nu071bdEB1TKK6JVzZ2T+0WP7n6lF9ThS+veilOoWqO+
0rduFK7D+bj+QxCEciyMm5s8i3kciJQmapQdjiFprEDXan9MMZ4gghEsOcH1jjgiijQR0Ii/g+Im
lO2oTtQ7nNZ9/aXp3WcNZq8TJ5eDBK//aoYWGAWxTN2mW1tE0MevSGR8gvaMZfXOPK2H/h4GyYMF
c8yGd7Qrg7q87Ja3Dopa1ajfr1N1gWaUvFEOrtjvA9hKvEoVnA897uKnbet9H1gK7mObO6mrSq/+
whnkHUrGzo3xS/9oWQbi+fv6x/fKmC4u6oXN/58YBIEmznDQBTuvpQQEQU0PBEL3YcfDE6JoczI2
G3YZr+6w86XsP3450LFcNt0Ka21xxmj5QtDrXEcVorV0L6KOEvtVMe970056lnHHeh9JYT9Uigal
C6aEbgymTpFwOX/FAbAIon9VnnOcqueWcdm8xm/Oc6K341+QTdCfdqqY1IbWnUDsCe1Z4BR17My4
lBX46k1Try+dncx0ayOCrftvZ5l2f1Z2BgVOhzZ+oc6doNceBPN3asIqT8FuuYki9wz+EPm9/mrq
nPSyz2i8q6qiflwegyqhDnsjdH5lCEf08VVBV6MwRtjCsMh/5RoftsJebc6jdjj7xhe1hVFJegFF
48cpoD8mXybtlKr4Impi3rX030g3K7j4NSZLpCihjhnFTlkRFtz32RBh/YxUftV//wjtxvzEh8qV
OMy+5B0UwhGxD7lgMYLr1bnz8ntwXVrWiYEgUBz1wiYPDOeM+279ZgT6oFMmc/9ZlE6ULfitrDHw
e9RHsKRMWA6qowukjwzECa5zEvp90DQcAhs51Sdp3wauM04qkZ71lNbt5BQO33UzQW4MfwTCl4k0
b02blL/i/2m4v+8BNuwUqqMXGB4twOq/qvVsnnclPzv6ADYr941jEIzvQS01dHwkoh8Se/ixmbS5
OpPw9vPzFWyRstY1VgxCKeOm0vZNKMT3AtybhkhYUfMY3VsRwWyoDLArq7GLY5uuP4TJ5YxJNOyX
UwMAJLEwfiH7oWa0AlB2TrWtMn/rZ93Zd/nxcUuGpCFgCPpd1GRSW73jWQJ/KNj+Y0Xl6rFDqWaz
V8mlz6nfzJaDzd+6MKgxc2sHpSrFcir9/CNavgfTE5yXzyHCqwFl1h1pF2hJU53oUJCpAUszgMxN
vxUucLM5BX0o1hjEE26Zl6PHaFCtt3kd7E1fDZZ70AO/ujoXSYCS6f9TmlgfAure9ByHe8fsNvNx
L1Dcho+U1qtl1yI3tjWnlO2z8Mxoew5IYwi0rt3Ou/DIlAgn1mQDDI4982tuKwx9A5oxbQ/s7rz1
8XdcPhvMcBqxKEWJbuterBi/hQ1X05pcJt8RyEcxtNU0ZSPptmY2JMqGGxYZYBTrQXF61nJb3P1r
1baBuhaIXtjZeIyQgNocCzP9JRAUQtApULfmrQbERCYXn/SukwS7ODKtYaxzzFyJ/XKARcbV56ex
P2Ws/Kb8wasFZ/InVCaIqM3mZ/DDGK8k3fg1xpifyPQRkWc2SsjFYRax0lTpaIZ/zbbY+NcpYXKo
3i3ppKD5hNnfGe2/abHfTr0E4Mc/V4tsu4JQ09FiV+06hWodGxAlMo5c53aaeaXjcX9OAjYx3XHq
aXpwGU+bFPW84p9b/8rEjDRuYeYclVhDVXa2KfSWyT/7WF2ZC12vmkRy0piNd6Wqzb7Z1qgcH2ig
UUxdyl3pa8APITkGbmLcBig8VtjLLh/fhypxs+Yrm7R7lD66Y9eaKSDRzoiRm1quHihWJruSt1N1
1/0vX7ho3ytwdFPHhibT44xMd+3bUwSjcjouDX8POZ1upvq5sEZHYBW9Jq9DI3y5dNcZW+hvVjNd
qbAWiNKil3cF7p3t3TCQLbn/X1eAo3r0pVbgUfzkR5WK/kTrTIzldXrJkl+NKz+rgfg8X6Ms9J7E
1xaTZxt7as/cKrQ18HSYesncHS2RKbZhmb6nyJUNkP+f/dAEsFkuHA94xSPLLTh2OUxctmDw+Hir
OFWv0+E6HB8nH5WcdUi3a2mQVpU0L3gCkfmcRRmQ/av0l3bnL1Ix6cKO7ZYoL9xtR6q6NGDB302z
77A53w/Zo3ynTSH2CY/cCsdrzGp2Hkq1S+6whigxg9RaeMprXTRWVw4TR3KqWAgyLsIwjHl6PCdd
zO9juf4+dSb+5hivt9oIF+LvCMDbtKFuMN0tvKcSe/GATYH87seFGj2EzkKP2cVRhhon/nCqLFk/
QnTST7FLIJsrBTIAoJ5Zmlc2w0LgFQ45J/1zmLcPCW4cVvr/NSEANYFT1Uc+sb6fB8J+xl/x5ug7
cf3/k7Il1YIoBF+s8THEyRUy7axnjQi1xf4ms506XCeFss4P0DsBZYseNsmxjcpM5iBOZhIOsrTX
rGBnLyjQqjJKhGVVtoK5bZ7XLZSCowcl7M+AjvRCTomnIs1xDCImY9J6l5CMEwv1fcrIGTJNfwQl
WRTVIFInGMyjck2Z/YTKorTQrXGfcLjMEShY1dFdEunKqgh4/euoPnqjYGnuObjtT+VhFFo9ntwk
r3KOei8URgdvrsLRts8MUVwYd+WAXKip9CXWjmkHDgtrthcF4qD/PShY3/L/j9pC4pY2xSZtCfoM
kXXBf9l4MWWDpCl90v7Nt3eS20wjayZjFtURjvGShfzjvaxlmT72Dp+DgSMlnDAQtIxYbLZhFw1E
lq6agXbLsAzpKutCdGn6zn53Z715xmXAhcAWOtS/6WX+1/HJzo2iLM7mNVaCrt4Sj+Nhv0mzwlzV
GnXuPATXwyYLN+BJiwEjd5N0mrg7lPhseJAWqwaVncfWgeKiC/4YDCjTm0y442DSudSZz7XwyhzR
d975A0c8xo2qi3LHbtQ1hglDq4e3fCCle5SCoskDwfAhPKmeo4nSxEU1QWoerBAAsoFYS+ApRm+x
C/cHCTHQ+2sq+MFSV0mKd59vwqSMduYELYqdwGAsAVW5ciFcSwzrGqxQ8AtBsVKT1w0d8NUukPz2
6fJNSTmrwlNcv6IhhSkTlz15GGGq71Q/B0JVm+ZGpowDLS+O9IFgbO2kIui++oE5MP7c0WsyzfNl
9681EXhPe8BEk0xFifKMs8mBZiNQgbzjCpUg6WtVtz+VhuyN9Lnbh0vo1ICBxy7lXalVAeRERDgR
SEoa+I+t+jQZRiMs6iAV57PdJNRAmGIviW2uoBf6x28j9ZiAOKRso2yb1DTBKViFr4PLwD4hEqIS
YNMN+v4Nno8xitz41E+fMPVbThfncmAMUQhOxAJzs7N8YUR8NNhSa6uh9EREFTCEs61ZqK6R74Zl
Er0Ggf4V5Q1rTOzCoUWqfFJWoKPeA97/bYXn9WhqL3iFEWqFQc+WtsbwIGQ3aoPaIGt16ntVMYrP
Xd2FNfUcQAvHOy05I2xqUrxHUJEMtiE38/UqZHvMHmnWwL430fFe4DNdVC38PWyF4pXkBROzCXl6
JuyAgx6RUw5CIc32JcuyTgqFTk7MttPhRHCZA6zFYnUz30VVKalXM94aaTjCc9wa5q3nRaYM6jVO
znSYAVIgvzR3eC4g2tQQDbeXUcexXXIU8ERparRVd7oAPp+CEnYw8bwQbJ73um7H5glh4PpBOzC/
SwRPiGLXXi+HJwDy5Byr8yFpR4s3sKvG5bYSLbxiuhVY7tm5yoFsAWI/VpZ+mNC/kC74fSxbTEAe
d8M+KSyyhWgr2+R0bkx3ny8svLlCjPpuYfKBRXLYZWYGG1sBk8gbCNuTuXqnQjAZK0gnjfVm/Pjv
AIhJk+udFpUTgmp0e9kRNI2xHlzm9wsZAwXVTNIrxiqiUBXxbevZVHlVX7UDc5vj2v/ZNUDEN1oi
4ZEDHsY2bNs7GB9aQxVx/cUil84MHXcjEpucOVDYlSI1d2EMFvLHlmL7r1prqTuCJIQeQlrdtElw
X5GTGtunxGVhh936c+LcKHiMGNbBHnUy4K28Hmt5PLrGuCkSIIE6C/ZALsMLWo1nX2sS5G900ey/
pLJisf+IaYqfE6OBhM+KXw3/3IS1rqlOb83n7tv5gbw/IRw1coqKCF6uZX7TNqzmYNRoXSIebXLV
KtaKv+y9rJQK/9Sf8xhG0HhhjI7j4iDjIjVD7FmL9BPecXOZV9VsZ+hQRC1FvaZ0vHD+rbF49Ekv
QmhILfwWQ9WaBLW5RRjXxF7iqVGUFDZRa6xOgfr5tYcXyPE9usl+SbbXnW//NNWuLPi9oJdkiG4u
m4ousYbCY4cvB1/OCvp8PgUezkW68NFqHs4yC54G5kx8QxAbm/2vBgeIn6THtzEoG9Nc+5mV2OYB
7wX5PJjhoml2Gzlz9CSQi/OHlaL6IpZmrzRG+ZfMs2+UnB8EwX/YyK/6R7XKWqjFXe58CGGa3r6b
2/x4kgIQpWQRlmg5prLr7wohwm5Bx6prnpLeqK8VGwZU9D5jq1L7mLk+F8C+T/b+ORm0HH7yhh3O
LcT4ceYMKCDOg8iv9MuiVNIDLTzhtlOIJla9p46c2dMRARP7r4J5b6qPW0up640aM3TmRtocZLJn
66BVr4qGniFpahCWHBBgZBsPt1X7v8ZXJF1vP1yI7U6HJAalQS5Bt02jdtdFUpOIINqNZHnfzddV
ybBjim7cycamP34/a9Gcwj5vhSSvSiktfnLHQO7GlkvkKV1hWk2YlRzFzgakCScbvrK9u4ptw/Vd
tRg7YHMUujUy2N/brbhuCCPk0TcoIOBh5TYwT1YeG2c2+/V8MpU2hUBndCkmWlbSoG3o64Is+zzF
520UjbVevHYq7IDFcDJxCaXHSqZsoCcZXe+LPYWPwdsP8tZoPf9xU5UkXaUdD6Kgm11bxwmJvpMY
WvhZotX6Wh4eagI8BlDb2ryrJJhC7KR9esvOPkydh2ksERNmsTCsUL2ifV1DP6mf0LrfZBocn1Ow
iBP2h75bb8NxLYqFJ8PhF7jjsm6ZjVVcb8h2bDBLTWoLHPRZ8gTjJKkPCgnvALxE8WQjCYh5WIQ/
Oo1KrJ0EK/+SH6v8yszLAdQqELM3uJFYrk9k784fZUx62xSwDjMqSkY48THJkWMQjxlDvQU6cG/W
vg9dq9j5S/Wn/WnnVjJyUPeSblEUtRcRzM7iYcQuPnvI63emXdSswdig7gLYbD7TklQ/XkMQNdw5
fi8yLPWy2msCH1icvAH8BdJ6Cc9ZnPToyHzjPP5PhzIncpux7EPscv1lmcidQKn1/MbLTinUgd/J
rmz/TeXOxQCUwEs0ehxvZ41Lkk1IJHWbP+rdNnKCNM0WS9v7kgPXQykComknyKeylHZ7ncGSShL3
JFYI2opHeiPB8uMQtoBz5+izA6GCowcZNwrebgvZb2iQ0C/S7BcrdosE/gjQXfN4qMyqtnD91G2l
sdBi6+v2ysffzSkvkVzRhpSrTTijBD3bKb4mU2JpzDctXgTxTpnSPHIil1uLoVDaEi+HJOKoDtzj
wODUOgVSvXrsMbLQ/9GSafrdnOZKehB3csq4BFpO4w+vB5F5eglN3FFH16pDUaeh3RjG9lCYyJXN
cqKHIIS12G8SlyuSMOt76OyFQgrt0IotPRiYMdtqMHE18fVZu36Hlpuvp4lKCdnnP3PiPK3gznBz
FLnVWSPBmocdzoIWmS90wNA3ytmz4WLRvvMd/FWYTY6aiuL/hHmltkIeZsx+/FghD9cDuprO5jw+
cTRwYk8NylQBfze/HUIOdHgwL646WurRdmo3Swn7nceE951p5nETkEUs/C/20US8i8YoO4hbaROP
QuNZfI8od8Ubek6lt8sLFf7INp37RKRV0koYsDuFKHSdKt3Cj8crXUojw1X7KNcqq3LNOv+t1eF2
LZ+2Z1LSLJ11GWnp3vEbokN0b6YpyHCMJXJH96Ws4ouLgpuyKDZCvNXoTItB0wczMJ6FSq12by8U
WZJSE/3+5tD3Acg0GdViZqhqc0yXcZQlz3FLvnKV/UMpXoq2LGiFoHH6u0uSKrzWM3ymAE7WfKA/
0kw6btt/WsVfv2Fi+W44RwKy3HXZNRUHdBcGJ1pl/Sg9PW0Xj2cQM9DDiUG6Jwsihauv77ztISmO
cD8ORtNrYfWXwZ/Qtp+PFyGcDi6DRiASrois/yn3uwKATjGmTPtEnIKf9HTOmW/AUH68fhSa+xwu
WxxJS1Jq9I4QFwDaowBtzbMQNRJpFI2iGLhEQLyJ6DrpoPhBjiuXntoTArGkouR9NIAGk21krnK3
J60K44EO3DfV2PcpQcvCIZz0+Do0GCzO0eiOsFaZ92VJmu8nucazZt8lHi9EjNGSIjZQgmhdc+io
nh3gCYoX5DxdDDmiRRRtRPZPvlcDJZcitgeMobCKx57+9iryywVeKx2yXl1i2p/Tg+wXYLJgS5Nr
EzYmpbmEQSNdAno1kRqKTAFsE94/RXpfIT0RVyANi5hycmVXW8fIASQGV4MmNQN8n5N3Nh0sNEn9
P7PaLEGhKSIcr/gp9cDKsfgVdEukxCEsYzHaaCqYMSEG9dWgR3sCuvem2V3Dp0jYOoHyqicDN47J
sljmyfrvgjj0PknUdj/MYnbuCDOeaFET6ppkNQULX16WHn0s91vxFrUR9KIHsQIZFfruP7TLkkhy
Mi6WxAVKYdcjlooF/w9z7TzWBXNwTrGi2LBsidImxsSXvy2/9I0eeZpfLDvhXZgQfklYfXlJABd0
YHk7TnuDj7i0JxSefSNSY1Fip/d7f137f1hfZZynGy+E2xYr+HIgaO0LzPMTk7opx8/6RNi5hag0
Nh8jajLeyvzZpPD0TdsN4BwGP95GgOYlJjK5w68ovom3F6OBcoyQjULSZwL8M26qyrJzKt+tak+x
dWw5rcgh0juBGQVT07YLUUFL16wjm/I6meTGNhci4wg80hLVVF25Pq99idoa73Fkgnnk5+T7c8Uk
DIhFQzWmNPyMDJ/ORImAH/DhiwrLRw/HO27QD2fA+0CdhT9QFqQnrMp0p6uIUvfALUetKwDyrRbS
DKLTslcpV8kur3/Tz9GpSCd5u6/dVdSR4/1m5Sw1V8drsA1gSFPNxyY3NlIJD6O6hCrfRGBbvg6F
/EfmqXbWqfJqjOkRztzEbTShh4HU37loQVZ+jgCkMDdHaCdwOK827UZgaJNxSv208oKW3V8xM1iN
W1tUPW4o6bzTQYXv+mP3vICN1MvdwNAtACWRx720nTFZcDYYaD4DRK64rSIL/R0sEFMUhxymgrnn
QtUjXX7cqB8eI8L39wScQq79tWmbfYe8lALWhBgRQM28NaJ+kFjIckjnSWTqQ1yDVM7ifBxkSNPX
uo8pBWrP8wdQWHSxrjRtPe7cKx259Bsa3PP3xo1OStmSyIPR7ThrimtlW5smXR1Et1ExgIoV4Fcm
so96VdVQi4e6II28FPSpgmD+Awi9uuziZu/Wp6KCkX/HjDr/gYUk3SKrIK5IAxMehypcWSPXGW+j
4dxNTGPAzs2RNohNG4CUVxzBfwgMBBMiBIcOMpnWz7XDaKjbNbKXHT2OkZVQAgzuAAljeJ/eQuWN
N+pVjP7bQvth3pdq9ozltu849hYcyZWM4NYeFhMm/NqI2JJIhmJEj1tSzqcNG+tEIDExNfey3Th8
gTlEU0m45gtedLJC+X2HZ/qEygWzp/Mk9nx2a/KUCe8MFewPCqWnsZOi975Rc78+oeAGveRXqYG5
z+69hc0HsHkNCrYX+uHmnRrVql2WVgPazuH8kpuzcxyU4R3REX7jb5kkztX5it6CQpJp4dLei1rc
y/JyDclQIelJov7ZKej0BveivVdS4Uvhtr06/g8cH/4UFJlylD1OYUdHOGQBjVySJSZYOx3IhahR
quv6J4/D+wBpouWNQl6iP92MAoIp+sFiUa8CQQJ8vYGhy+Ss7jiFp0Hj3o/f+lrdI37kmIgmFjOn
evxdAjKSmuUj67RRXFzyWkC8bqtS8c/+0ufdCJ5XaeCEgRiKy0qeDfvKW/nrLa87ZCAUOS4tjRov
Vf/WSfXIXPGTIofPYU/69dIKVF+TXyCa9vS25EmhxnUjSkX0TLDMHL+BKUsYe2QyOT4zvaVmAuwx
XjS1D/KqxnET2mLpKvwHX1dge3wljbg1YvLHmuI1FjGbPvapsIgic4ITcM1RZS/ETrw/B8V5bwBW
Y+eOf/gdHF3WJa5mQGIlpqRpVuZ/lbTj5kRa1t3UHHixNJNIhtlfY99knnOzTcu2NAixGJy9kqj6
PnJ0477iQbhhZ+AIfIDwcgYP2oJInVE9OKIuxfNaWdqjC1ZtFAkBxqGAbss/tvqzfCcdYypoNXS/
FAUFvDBg1slV+WkHqHYQzT/x2N8iaeYnrSUzlaEmukXQkkIbtB3Ne8t5WNc1Mo3dGi7mWCFBVWy6
5hsWpYjuRwLvcW5mucDJPKYP+UewMQOPsgyX8G9Bwz2XHoD0e6X4BaNx9lKezLwokfP8iANO+ipc
PXcA7osTanRNQKUhq3cztWLpJ8lVuryZ/sXzoy1pbKKncMZ2CihRbHlJ5ec7cG8ZQPcCf6Y9M5Jl
FDW+JpN4zzp5Uo8iaZ5P7xsm15VlQHyecK/nZ6gs2Xjg/sGL7mEzxaS9UpwunqExnZ8fP3rnN54v
ngxsuOB7SSaO8NK/joB0Ar8oLYWplYToqxgki37o9PT2YMjScUho7yj4rtZC2C2PbGb9vCMSzZeF
AErbjcZQF/FUqjnDfFPalY+vC4LH4cMUcGRoKopgf7Q3xOGQCUxiU5xaJhAokPM4PrXQr37CJtI/
91IEw1fLG+xcnZAb1ERqBOsGnlMsJ8BrchJUXH61L0ItLfasHtW0DFdWTpw3OJ4yWiP5oh5mD1zH
B1IQSjj542mjnx6D7y1i0dLpVwzokF/x4rylyZSAjRpkq7QbyXk0fyqjlelKtEPX9wo+dQqT/fjU
uF7NOCcLdmo7Om1x5Z010x1k07asRc5AL2VnYxi5mO3VMSlNcATNsJPQCQdLBFkqPYBojif8kPlT
ukTQnfbEIGlqILRXOiPxSOdwocyj5nzWJ6GWx7xNRfe2MkcIO8OBa8bKzhpcY9FURGlSMyc1kitY
cWaoKh1kFp+7eKjnPKcn9u6FL/0QLBtuIflIuJCA0iU/JmS0X+pSKHwIuimC6fbqbK572GIq1QF2
WvkDnmmrbKNNA1h2r4n+cnc4kcw5ef4FYw0j5EoOchubS9diVtDAemN/tUA3q5u4d3Q66i8u7Xf2
AUsHBit6ePGO33ur1W9ZhBFKoCyv+9vE1cRcbJ2BersazLs/lSnpiyBjV4xUgQzWhMsMgkfDHO7W
fW4ncR/y561l8e74v1wCQfvxik7ieWZXX4DA8RPiiCtEZuuk0Id/ckZFV3jdrCIMjMKKtcHoYxDn
2SAbQYS5ALIRf3qo7dyW5i1Xc+IT9w7FuauW4Gkzl3U2w+3M5cENYHyuMWUxW4SkbR5oyE5ksgpu
IxGABa3ir+c29aqIpcomotS5IQvmDjXria96kf0/4YlAWpgDTDKHk8UIYmJCMT6i7w4HdUalis3N
FdhIBN/c2bE4X6czIz87YqzaKbi7NVyOtkFbpj2w6CR6IV2KCn7TrOJGAMJx/VH1r7rJTPdybiQb
0JUTyiB2qdY6F1hh+Ja/od6EIv9tfJ7frc3TpsY1uFfGUd2ErPlBK6m7TNSdSSeTyaGHBt7hq7Ty
v/5n6svq2/EassyjjWcrz3qAFZTr1eJi17KKC2xGLX6VRgUl16/pJTVkNPYu38X7s970lU8or1Vm
dJr2CI02w02Kad0TjQaadIpoYiY3qgEmWdBPnRHkbYA7mCzTWFsLTLUwrMNT9vlTFBqTgBGA7Z5Q
lCuKh02u/KacdoNaJSG2aewKnkZpnkPROXXEiYT/F3ypWxY9MX6FDXPHxlC2HoSIGb2IT5C2KlJT
VKavx/6ay3/1LPRAyXUYkWlJ0DEQMsgyroPQG/PIJOInfN7IUb7qzLwV+o78hITjdsJaxbs71Teh
oZnu8r5Qa6dlxS5C11GJmECbbsprWiBTOnr/8OgTFicltPrB75/JFTEJAm/o6I3N81i7e7NbEaVR
syLrSp1eOTM2qSFf/0eeLfIyi9pmvo4OgEQzEfrl7rUQJYhUzr06uDKW4A2U4KDLOyvtyu4umt5j
snWPeQ+yfLQ70nKAFX0ANZT+0JQJgZV5F5VdEv7pIHssvLXwCsYwhUMg0qf8NVHS91NVAiPDR/Kr
V3wN6GQFvc9YtgxgXeiNAWv9yDFT5Vq+6l91zLp48NQWFUqdX9Mt4GbYtuKThAiYRhAEz1wA00CT
pdvvqG5oB7ABfksGg0mOU6D5S4LMFqbW4ETVkM0gx+oQuspdRHYmgNWir5CdQDNEfUtY4LVdGNxJ
7ShacDOnx7yDBc8ojPc8VZzzGKMLITeejirIvVfcAFwj/Dbpxr6XbiFXG0aY2WGMFkur+36D4AEK
SbaDSS87Y9a+yjtA8PxZxc+WSeQI+69I5CiK1Mrp2KWbGW72+RJuNajaAnwQni7MXVvnO+BDmUxg
k91WT20uRj4iEMiApLBKswd9aj51MotresiIs56bg/7ETzpBYxaWx+DC1TCcBQXYFtIZzKzW/sVl
TsykU3oyhMZVTD8OLkmhIIWmoKQnKsG0/ukapU9n7/5pWx47n067FkknRsccrCKL0vDGimPxIABm
9iMhrzunftVHg1BFX8o1dfTdqUSq4sWlLxzGQ/aGdN1bJHM+R32JhCVKUN2G2oHNa0Gt0X86ZJ4F
EAUaNMcCuavOGAprlWDe/DG3CEWKaP+HqcNFY/81q1vdWFI9t6mqsPKcR9Un3eQ2uX6DvJkfOy1l
kCrTIoQ3IMlX1W+s2E0QdtclrhsULwuuV4/cz+/e7cGE0RZOMTPiQ2y2rJuWhPifjQje8JW3BkEt
7ajxWBivvY/b9tVqVVMofw8gyjnKWFRbzZTuBxXbWxPSt+0ai1RVWytlWs0hYALOvLITmAl64UFf
FtnIAIUjRR6Rh4X05GmqXU05S8Eub8xY7sCuGAA01EeeJsVXwa3MjBhV9NdM3SJ4xhQ6sahzJeMU
1Asaccqk/kwYYX2vSoRYq9qs8edivDVEtAcjJE4zOOZyuK/6qyFyu6QeRRtg+zSY1yRfQ9Y69TK1
lenwmMhZZK+5av/RblKBq3wx0oEeXSViVoJ/q4tDrUCx3WvxJFeN0qn3yygmMNZdeZJXQIVl56hL
rY+5l76OptVwUjVr3HmlfaZq0CutvLkEVd83QbS6sOTf4pZRJ6FY45hinb7SLHLqMnmLfPD41eNi
/E8ZGurRHuHb9Rp90LUysuhYfGUZGywlRWFLkbXlMvYtSwZnleL23cwr4QtapgR8qE0KUlE66epw
Aa2dPoKsnGmT3Zy10iAmJTWDlz6g39Bqtaw02Pq9OjmgrZm8oUxsg/qkIB3Qq8WuVnOX5ytT2fKP
EnrJMhNZP20vSp7XG30kJTpHHTRnWZbuH1qnRT87l7wcB65jDF7aP4epxui0/9pkyNA6ux3jUtFg
2FvUM7SrGdTjDsHjPjoSJCRujfD9rBkYBt0Dlllp3ocQPZHEVhdaqHSqkjTUSpstub/NKcFnvejR
JO3R0/NMnbrU/G9u9r6O17UAeK/HuouaXIRc5Y7sD1HHsGfo7SS+LaabWrGDb9sBoZE5Fn6BLSoo
xj+BmQHDLewFSQiPTSCBo4/eOU1t0v8nIiyNLlgqdpa+Gd9zMyBNx9RntZXmJQU962RV54WfRmSN
XNR3YpbBUq7c8C2ePVSwitlKacxa9RoIZqo6qLH6KIVn1sZh4WrX7qQSqNZJvG+NDgrDspQPwszC
lIjLHu6vWVRdvqZns3J2ftL9TmsyOVW9dYxZLmlEXB5J4PdcqpgKrBqvFpeJu1VD/RNGtgf3kCAt
O3QHj1kw6PfyazDB+hwT4ck8IfqBasNsFjMSi0TZwY9MlIIBaMsH+fZT4UQyprUWXAooKBtPGeAE
9y86Sc6xJQ2X1bI+E0zlgnknJ+LIagyOfIUprMh9ZIp4NyLu+2oAaYGp7CGRF2atPxUk58abOIJe
2iNd1eU6MUYNYMNOJTnvowtR1jDodpFqAVQrPxAPA+XuIBy+pE0JFZG8hD9bom4atsY4v8+2loVR
Pw3/HshzDQGil9NiNkLNAa7yWK/WJgEoa8ejFRX6s7vXkKA154K3kzaXYbd5KDYIZVEfIBzZwnH7
mtiHjbsyoLGyCKlgYFV3B+rivvYhAZG33Qpof0YMB5EFHtRE3ROwgigaiMnkKZ7BMXPmV0NECl+W
ZFmwXiUSMuWwCKclxHuScDEQMNMfucVMDCDbStFBXns6ZTyZCc2mtusDTsUSnsxq2Dx5S7vzf9nx
4y/yANlT3fkzqVZzY8mY89pC32Kac03i3cEzF/OsddF0N2FSc6NY8v1mpgJuQ4YpuvsbxUgdEzh+
T3hYlu03PBc6oiZiUl3tLLxEEl543AprUH2/2R0jqSCvJuezObaQi/RBvrhViM5yMrsFtVQyMfMZ
nATI7MGprKOnIcYrf9V5l0vmovZs+N3EdqeSSYoxqstVecozExIDdoYx9ExN0O6bRYONz4rkduSX
oknvBuj3knizSWtjncpCceLJHqjn6ahDy6GvCAKzxAhRRKye1YRqtTmNE2NYwRqBHCVvTKgzW1JZ
ldcp85txMeJHnL3PVgnlLA2lXr0/PwXi6JJK/ueN+9aj3y62QLFylaeRG1DVh/fwKa41IXQDESnk
nM7NkrMgt3pI6ycr7SPE5VfBD6+0ISaDDpDOZ2zAnxaWGo629ZtgnP75Tj9533IXmKXPJ7qgTbww
UBCggRtlxZ+tR6/bUiHFxjY+T2P1vWY9ncj6+2lNtTQcNEfyGSdZnZARq84dkoL/U7+kZKJ6ZBMq
BqQ6m+h3UOAu4750ZfDTNRo4iNrr6y20qs5R1QC5dP44K1s/37AkOvfq3bR9uEubJlcrkafKw5Y3
KFLcftUcu1rJ7Q8B9rSMhYimBc8TrIhcwJK7hd3JJZb9LlKyFVvYxsiT5uL+r6TTQmB9ilhZpKHf
W1dbeghgAJiGb1bIHjXgLTmMPuHciEh443fSk5q3edhRg/DEHHCZHshMtqicD+TsnWRQsMsJB9R7
vW/2SpRg+IraezdXZaJqKYcGcPmznRdqmjopfvOk5yIhX4K+vk4Ekpg0KphL1zGUWd0krb4lE7ar
glURicY5nvg3noqXWQePQGXjMbjO6jkPoZF+LzUGeAmEI5WuH7/HzqxGM89GW9hUuH0zKpBQFNv9
pF7Tg7S6FIfrLZrUqGiYbjfE3ajMjyxlp/XDkTpZv40qmHW+R30vjGZ0O1zKDUTBPFREJo6Cq7Mu
31iIWbUNLiS2pLczFYiwD32vVbaUN9ouLugN7heeSkaZLdzrnW1/MSlKFN1ocYTIQUI8JzSrLF4A
7/XSqr3lB/+fDn+KwfFPHiVjleI7vsKSuOphF6whNXvrG/9+5PV/qj3iaAhgHzH8LnScLzEe2tuz
PqusgI97UVzGQ9Jyup24CSvDelMYOFyf+m6mA7+xH1kNFYq3dQYGtUcK0y15359Y4KZS7i4X1lCs
ohOusYi6k4Ty4peMgcguYRHQa/IRLvaO8EePey4aFwjPBVytZ7R7FOC1wTNuiILMuApfVsy45xeQ
yy96m9w57o3WunJWXnydqzPVk9xGIz8ACVSpVNoskGVnkmyzXJxTfa6caZo5yAIG/vsrMyh0A8X/
pf4WY3lHt3vI2Pv0k4gd45zZmUeBTzrspbAEQJgmuOz9vu8t5js/dETPSBWve6Ag+EDqU8qWOQRf
aNUNKZcueHFCOhmds/uc904TdXIp7YN+VU/LPZwPMAi4fIu7BEk99UqIWgFn3/WEnshXs6dCDsWN
gCPwHktUGi83JKnT1CPVWgzECrDFuducWTSw4aQvMhxpOSWsZCUePnGn0xW5gKQC3Puvyuc8F6KQ
cMu+HAiTSb+Fubx7LF5ZrhW4bcOJ3ty3PzMbvStK8Qvu3EHqbR+6dd8zchWXnUR6IBgQzsvwhAF+
0dvZVPvWV+I1pS9+iSJP9jHh3eMmKRSwk8X5bqp2vUqCujG8bdhp6mBI3GlI7ff+Ge7IhGS354e3
zk/NRjIeITA2Tlv830sVxGL7l9Gv+H/rhGZCP8+QPu3wV4gKFvONHS7b+heav2upJPQLzfAh3vHM
Yd+REWZ3Azp3Yy1KEj8pjzzS8NaKmmWAJjw0k8eIVaLVuTItN8AmURp1YDcFiikTYExV1OnsX2EF
Yndw7oJI/sSuTDPyqztpNpsijErwjsuKLrU37P0B6D4WOfDdeJVcCXXgMAT9XoI0/Npy5Vg1xsmK
hr4tpZ6WgnvvS69eLS+J+9cJ7QsApb1hrKMIdx2SKkC7Aqgbvk6HNsCG8tyINSDoQXdood0ZGygz
DR+cBsaLaSw10ZlKMXHGjQxk8Ip1RDDcfhIMYXNXiM397SOEI9nt0wxowO6rhIbz5PfCtemzcGD5
ZeAZRBLnUkrfwuBLB37Qo0WIpCr/wZmvb1FtsfLr4Su08JTdGKYOD4WNsZgRRqhHQKkGh6g8xs9B
b8iaJ9GJzYCTu6y56Y3316SrVUiEEjQdL4F7TU0Oq6eiR+Gj0GvzmM1nUSE6cwSsxKHFN8e2ah+k
zXiQuGy6pkmQaPj6Ttr2z0d9+7Ub2N9FtdxYBUA1xgZmdWToMLM1MWuSdqh99xhVZfFTE4VBrYPD
jLNpziS8A2NoProKAhuPCMRohIJ69MXrQavBu4N9XQx9t4tGRwrxI7zxsEPNjBzy6TIUcmOrLFQb
hC2bimm0b9Hld1E3XJp6uE2/AqhQLbEUXX0edGGtfm01LlsjGCEjT4WPp5N68lQnl0SQPCIPkTKd
LXTGYzv/DKMmwI1amOUtM8kgN+LQ6KT4IN/QHGGpi+Mqj4/LXDs11njqB+IuNUSJfbM2A0wtRsTl
D9b1Gs6RS4MzrIDOfypvi9JfTiBJ9UQQJVqJbgsM6tr7zROQA48WbnLq7m6KG3u45/M/y+rQyUx3
UXTigFX9YdS0jJ5cSbrITkb0HRhWF75DXkbwYB0WYBmx9frOlxs9Zl7CePXxqtA2KDZ1/CpAC+3s
rqFtPPrcm6t6Ca++xfXlvs6RXzT3JpiSsSMXvCXWlI0i7VGA4w3bwSDKPEhRvfNlkiFq3MEuSzHV
+NyWhZ7otHomhs0i1EMn7mtEE0zOM4a+U6CvurwEYGoaY/vuYZ899qnXlNGFip2aJQxrbOdqnYFL
4QNRoWzpRPoyv3A03qCsczcw8nNqTJRHn0dlITtXgFZ6ybLDRUEmSR16vmnwkPUJi8hhnLcRsRnY
nTgL2PNAQOY76ZOw9GjAlbL6S1VTBwWyl5wAeEhm1//ZkqKmo6p4Tq1gabRKxvSWViWXidTEGaYY
BWR83FGhs+I5AwD07sstDQmfkJz7IRrd5JIqx9QtGvbzO0NaorVrnBaatQ/RZkBbzVP5ICxcwQbC
HUClGWWnkExiU0IBj3r9OwWJ5hUb4JHh0CxXSFqgYq9qb35PWK5hV5K5+LiU/st9LdM+iCPEuKDR
LM7lHvHXWtbGNsNKjDMOL7Zr11L8yCl83wTx1RXhMD8I29tyt55LmOs9YRgv2o5N3QSj1gun5Nu2
NmETn6nw7UaA9m1J3dKxYBul6xM2FIksMGGNnTmivISel6kr7ZxpIUWYjB/sxiyXSMi5NbvYsFc9
bmT0frHOv3YhhoAezvvc6V7axXfV3d6Dui5mljtuvaDrLMJAeWIM57d/h1P64pE0qWytL8Ttt4+l
TnwQIb4MFGqXKacwOwoWX+DnIOx/S9dljop2NZLgadXPwQXs+jGc5LFWt3+91NrsqsOD5qfuoQnI
8YNwpG+llnX3a2xFbSr4Do0KQ5Pad0Nz+rAtDHztFUEPJrDnNL/YAXhUMgwLFAs4e1uXowZ+kP2h
WO62ef+57KttC3FtAQdCRbznsG4k+hA8EcIjiveg66Tz0nqdD6slkiuS4c8gCP3Nx4uXKcCtnKBZ
9oA9ywwOXLClxC4/OLLbjoq//7ClybyCeV1uiEnH4TRLoVQGceTVrfMGo9MiMJaMHRSnMIBT31ou
MW6WL3R8j4kiXZDI6tv+1DJ37fgQvOT7NsSg0YoHZJB1i+Rqw0rrYAnYjAEf3BK3V2ESvsgFJC6B
W3W82S6iyZvn6eZLgnd2s1vlT11n3yN7OklSv5xRsq8flsqc+wMyzEKQ+67a/Hk3ximb2oTp4LUV
su+57YV/AC9wfzsGWxCYKKlLPm2CEPQe7FXQToEJnHU5Vb2fJFHNTzEh6jDLpF8fx+43DIkflpYG
xg/VmgJcDO4qH8Rno7spc/axktoLoxH+dCV3lruWzfK23cyFD5kt90OOVbcvhBm5EoeSyVywhSAs
G0S4f95KkCdfm8Ogg6td4wawpHj3Q4i3qrccN1Cbe0JxvszHGJO+QRvnf62a1nC1DEqMDss7OhWo
GvBcv/s68DzaTjD2aDfpwxKpDE/VWbF7Xl6zRo5JYJ/8xuDXX+/qx8bclib+n5fncR5zFDeDlXC2
+RN2PMGhV3FzQuZSME2L6arC+xwXbdS+il14n/JcvghOZA55Blh5TM2wNLonoCsvr9IbkVnA22WZ
AUVZ4hXksND7tnCskVxavqcLfTCmkG9DiV318WiUTLfKastMrtXMEg421y5GPze/TrWbKi/A2ehS
/WhitHgeAZ8lPbMdDhIjsGMBH+09RIC+7B0cLHZCkA3WhEqiWHckIr/VHJGDPPfCzUI2h8e3Iahj
OaQ+b9Yu01cUc5KLCNXbqdHO6elpz5l2nheqCdikI2Sw7ozRilUzTk1TMpJGQJEZWI5KHDifWsoF
5gyhuHzrjFHXez+s3k6GvFJqtm98uVMCmktjROmuMIOfLan41MTPJFdtdSTjOVRPbNIGaqHFsL/Y
/yaDvP/KJzX31hyATtXUN9ovQTD1u4OpTKKJ1NFSThOyA7GUpdU7GlbSA4KOOT6AP+nRbCpDTH+0
YTz/6QghvAqfQO6atAZiZzHv+RKVJ18WNRIgIbKWZKesa8KWDkyUFIEU+3LSQV0lJuvEVms3+17y
/BhtQhy8i5s5Ycy3h6Y9v/Pv3Qh1bHrBv/uJLu5522HQmSSzPaFlIRo8eetk1nIW0W2fADy/tmq0
OQIh66Xjy6Har9zmh2Kw/zDEnpI/YqHSqKQI/CyV93FEWa5GCaQ1BVA57kxQmuDVSA1rrgSWI1po
4k3QfsMYHRS/mMpaMEpQjlmWgTxHxe5bhipBfAk6kknxdK3CVsixalXfiHfVT7nauHpv/AVgB1qG
oEjJaToEINZdSkk9i+4/59tLtRGPLwy+pavos9Lmd1dmxHQVgj2RXNTMkvPFVhD7NYGefFHrRrxd
4/rcZKOXpUZDEKsbzBRhrqe8mSNjoVLzHBen7ZNFY5luBrABBOoxEkkFVLiYfro52901kO6Iima+
4I9RW4BfOpYKbgHMnu9TR40Y6A9FD8GtIkLtaz96WfGLpXFi0OfGbMFvzXyDVrundhfhYkZt9lGe
mMsY2HR7JKnOPLaSlX6ZX/uZBk7iVuywLKwQWIovq+kYEY1Y+PQ4WlK32WKlfFY/gR2f0TPZdMcJ
Xigv9sB5+3dAiM5f7xAp7eQQSWbr0/sYk2nRZKAHvpIWp9cbPu5tCmyIOXDIuGURo7Lb3FDLuqjZ
FxtzfQBUiIHNAgp6j85OpCVqj7bhdnoQtsN3ksVPK00cF4wxuCJAye4fOYKUiYfyI5oE1lfhJa+J
krfuWlW1SY6E7rYKj3a75xt2dw3Ss4W6iG7oprNmS/E/imb81j+GS6FZxOvwrAAZQPoC7Z2VuQqf
/nyYrddj18ngYEYM23k/qltmY0wr9GXKkx0IuY7RteVj8LXaKeTSBClueXf+siDWDxDCA76WJ1cA
vshtN47KV5tu/8jAh7jyST/T12Rd/6AIPO9+ajyv0jqbk36eY9sf3GIlwwQyTj88ILU2pW6KgAbA
TX625H/BmAcsbBX7jLNwDYAMFZfiu/BzNqMWph31Fozjr2lqL3EVg+OEwlDHUmfJYhZg9+Cmo1Ad
N73nKGuac25c9V6XfNRUjVP9zPC8p4J+ckVFeF59DD07nMEpgv70OOZHhzKttharcd1iVOIYHnrS
Qc6EdUYuMRHvVY9EzSpQYoUjVeqhMopu04KquZRRRz7AaGstOlqh2OELfiSZzalWDSvgG49vUSgN
4DS4CdAh+rsPTxyWYSSedoF5/8W91T1fBCS6WpAhuhoZoFYXor2RPyB6bIiE+pgyNrnkTDVzWjAf
vRKjH4w/OpEb6cQSobhv3siCXMqjBO/vLWKOeroo/YRoJHdGufd09LKrt+qJpBKQXuD89YV+yaOl
ww7SDG6FnGCWziQEzY2nDPFd+C7+Dz5NwF9E31LaPONtFtg/GVtCReNJJfnyYYWM0qVMlU7mKs2f
qDE5VJW39lAdEbYNcUZfRckuEzP24QI4fXGzIUjzUGSvw6qnECaGMKtSTUpCh36RUaw7sP7BZyUN
zsq6Wet913YLqu4wZJPPegHlyi7p6OGQsfV2SEcKCNeTKzvj8WofTeZ5kaudXwAJqyQE8yDS8asj
DFHFBsZEq9zP47O4MADGyt41qwqKR/UPo3JoDf4MyiV2vUJ7U/gkIlzGY3AmrMdWh5o3/x8DTr7Y
jxuK1HS/XzoGC11DSV8RDqZEugmHXoDLovSi7WvgmMzsTLQ1+rY09URHb+DcZ8+ISau0fMjLJ2Pu
drMbGQgPF9LCKyGAA2B0pBGi7f/thLZovF7m6feR2caXnm1AzmmJL+Oq7demKNTsXBCzQ+z4U/KN
628Oi6XL1TzVMzwGN9N7Mmg768QLywCeCEFEfTn+igl7cC4m+2zWLOFqHHmQMT9o1tziZ7vs85YE
QnKKSLeAAdc9+2i/G+0bgIKoDX0JakBKoV5785UX1AobtyI5uK0TEGY50rERnwxo6SCNOuWTsu3+
p822aNrHDTUDiGHN3k06unPBYHU+mvRwoVWgZEFH6/BZvDvGGhjh6YiLXQaLIyJKeR/OhacX0AIz
GmXbw8T1zmnbpgyyHVxVcoFKQ2oSh71I7ais2Wgab6oRj/sTC/qCnKr6aY1FMqhlE0HQPFpXKkPy
CE2svUMwuxQ03gYecFiMj8Xv+kryXAupPQ5HfuD6hWdZsZ9r9bfeyRrYQb1SKB/gq134AgY2yhEC
0/a9jbezRkTEzkxh6GuwHCFOFyFKGCuiR0rcQ4pAaET6GuJhLbJSSxCoooxNdRyDrMG0hee6kmO0
DZi69w+M8zm1g8lqYMHwsKBaw07bcudJDDCGM20pwOpJT1JE+ptP/K1+cbOt5i2/PN6m6jWc9jZX
8Jxkc8sh/gisveTkzEVxWe+OAEs6CrFT2akAIMJY8ER448ZP06n1vatdSDq8oBJd0AX6DPDClzrh
haEVRd3vKM3ZxtMcvypk78amklKjqwzJC9eLuXn+yGEWD13dbQ4ORx818JBUPoa2JrrDYhnAftmg
QD9kODnaA9klfXjJjW26TYilz1OeHpORKiyp+K8ujh6yEyYtLBDogZETtfHXgMckdhav4T/Gldux
dH1GqQj3XgjdzApUSkfY3xTyuVzgQ95vCEDuW1FYt1hRnYW76O3IGBc6BQUAOPeze6XUIUHHrJGn
Gl1u2mlL/ELfb9CXoLlsx/a5No2hL+OlEkD77kB0pUsvDRYdC8OSUwOrDthvy/eaEExk8/iYftet
lbJUFRArzNnpnckCXtPQN5u4kS6i/wmaRQkT5lZxRu3aMHg6sUqcxvhIJwffkZj9N601cMh1oHVe
BwTLzm0qMfVSqSKpmbaoPBwu4vALae4Jt8hWN/kqap3tOjJzzqs7REIrhXwqScjzFzzqwpHqNCVd
5anXYZtP3cCF5yylnZwCC+is/Ea5cbXAzsttX0a9o8QdlUxnxp6a2uhv1hNN5sJVaGFSYc1SMWiu
k1pJMrmLZomWnq6hT/1m9XoRAJ/wrrlS7lP2eJUJ7eWhtkFzRtJoeJYtbaHSctiafWYHcJuhGdWQ
EdyYledpEZ6QONEozJ6q75TFiZpzsWUauACLPFlTeUufg2hUsDIwTYXZFeICPSi+thPBUOIYcTNz
uxqZrU1aBz4PjW4un8GDwm49xxg25JDtQoC201Aw5CtdK3BiI1r//ILUbRyuiinSB+hlYqPOi32L
vpZIAJwro8OK3lUhnKJxCYkNKXEmZjgvccrkv3mdfjE8BxpnQPVcvz+8qj+w/8nWHBhNOjaybw5k
cEHfikpUq7crFwivfa+SwmYivMug3VHmKifvEHZX6BDRs01Ro0Wk/nDUfeP8gpYqu+8hfaReeyVP
IzFY3iE1upUrC8ut18FwxnfQNFrmT8H58tYPfeo7g+u80Q/GmNjJy6UZCbYzSX9LeTwaCtw9VSkn
VXtKfFR7T2mwTaYhNyrBeZNhCZc+RKHZkjm/uCaVEo9mOwzsCNRRpnEGRhg8pOTPxOf9aIuzfEAc
6XVpwYkx8PoQ2koCcPfH6/V7TyHOuiAF09E9oY+KD87G5TGpjDO0RAvSjFemfCSizPsTomag0MjR
iybE1cT2DKaE+4702r1b6wZqNBSKBvGT487OTpNE33z35zrI+RM2oGmXdptMfkO4oY1DsQqoPDwH
n0ZkNPAbsH46JgCuURBM7I1JMPUCKwkzVcVdTCGjORXhdWAvFeOeyTZiiy39RhuDCBIPhm1URoPo
UPwEiJsQ5XGrMDFUSgyROTKcVFG5pCCf1FXJdp6/QuHtw7a2XM1IGhW+y/XyITlK9qaXsoJNnxbC
qsNZ8PJ/LAbhdEiVF/AxTSvFqpdQwVO0Vpy4zMl1/BGSDdGdfRQaPvAYPwVTAdfa9K9ynzcZ1yGD
FOKEH7mgEf0IsDiSWPjXZjW75yGTscLmSLg+p09LEnoxbg//CkWPPJ0da7wVsavNpu5Prbe1SJQx
AOJGHMFACmPffAJLQzqHA/ZRrafM5RqvS7a0hIjrsmvTTbr0B5SOPrZFeNCjQOCPXhAy+6XKLgTF
ECfFXM4O5eTlo0B5OSQTJ9i7ejMKmRbDAQeS0QG44uHyM7Mp+qerj4r0xakEX0pUi6TJnVSl5T94
9snqiotguQFgqY6w6AEn2rGcoMZV0r2gBqZtKezU//p4P8QEvZmfKhh4dac2doqXCmXM/yYUwx8y
r6MtuKiZ9oVxEutEPOXQk+zW+PurqhY/CyRaTEqiagFL41qhUWor2zbE7MauNj4/ksKLnw9spinH
/li9QPzIxJfRfo4w4qoPz32QcOlWbpnDVP96sPnMs9ldViPuW6cs66IiTMRxg7MwaGLXKenp7SpT
Yl+JuBc9XzGQw96b8piO1ZU2ruApJo4qzXYhvUvszWoCsUnv5Kpe6G25zy+4nyDXpetlZujDqpAm
2fD3NLVlxkwqt/DI7flDBZjhevsv8HY+vWYZ1WMHhcbAvMWiY2qnN7oBmmRdEgzJayhOUv4vFiwJ
4RafDAAr4OQqHqIXhhXoppJ9zEbMGW3HXQmGwHmjocMnZZ1j9IbANks5VXaGd4guA71GAcvcdl8Y
x/9GyAc9UbITWFk//V7jqFSW3dqtpbH1Xb5kfinwfRNAcfqGOc9ugaa1GfpcA04rnqbegoX5CzAw
1i3uRc7V9GcZvi8z5avZ04jhZCLE3hCxNuu69WTcujd8xN7wgChWwQO1FLkQw5BSxEpSfpDHhOki
Ni6UTlVW4em6uSOMDR6jbejquxuIvUEBs+tuNmqnxPcIEVxeS2WlrBJYHxIr7nCNa7v7NxTQEdw5
4WK2AUmjz0d8yaWA35p2mdq6j+xNWVr/lMpuQN3/Lne0IzrvN3s+8cLeeP87G00WTVzeAoqKaQEI
58r9velxOETIDJXMQMCr8mEEUV27MAOS3GWPv1Q0GhLr3oT2Re2QWe6ZOUDa5V3VBhaumXQJf4ZQ
m3g8Z3JsFtwOPDO5W9k2tqSBukFpDVrWY5mPTeoiCnt1U9xrh/1DWGxv6E6Y/jqNX0qho0m44iBs
zE67BcuvZMg3wITr2vRwwQlbL19I7KnLAQZNoHB9LiuzleccMGQkxq17MhcQJgVRmAoug+zIcQ+p
vlNt2+yN5UzJLGA2D8OurUtP7y17i2XoYprlMiCaChK26KcuSU4ktjhc9G8A0PhFpfHQveGUWp0a
BDn1bSgFl+piRxELwPHGCvw1xecRFmJFN3e+R2br+IxICtW2tG4oD77JF/I+m4VajJ8s6/cbwYhB
0sOYXSYjki0nuAxna2/fgnk+V3V8Xyz9tyxnrDq/+awjPXBXcTvAyUxcUZqOzXbFyvt8ogjRtBBY
JO+VjqKXJQJ6cS+hE5jWwB0exy13kmrjPufvPQlMwWyg6Ctz51hA/BDsUbGoafawugjSWsLEWEXA
fBjxQjE14014Miolx8DdOIVZD26aK4A6XiOAZMRk7IsT4UaQ5E18DJOzwY5LaJMNM9YQSywGhXXS
2k0SteU3l8NsKa24cVJog4APS4MAe5jWvp6qhpmf2scFyCrzViX1hknZ3R8UCxhU9G2cBwUchmWw
OGig4nsDimd6xFnknlkioQnCLeQ6SBEy+l1fOPIQ6uNlTMmxHXzEi4oweHKHZqbYIiAMZfCdn8AL
R12y6tys+/fIeKkHM4F1lz0Mn/ZeVZ/M1xwd6WCoTH/50mssBwhaB5p+YvB0Ek4Kgelbg2B7FH8K
xVZChH07rxzL2vTij/ogCFwW8oX8MdMKxTsqPC4ZKlYL5u4895/zczWcngeUX4nYcsVqDrynsUy2
flH5fWfTmEedLOCE4M45fcPSHng4VvLN+VdKue3cZ3roIYU+l6rfsKSCzSImNm3anrb4wNQlkj8g
k5gDQ1fzcX++vXamus56xOlnPamS7uE5GRHj47qcJsnrzpR5QFkFnUXy3qbVGCu1UmFgfhRrDrTu
c+mzKw4PrOsLrFbATBmWXq1We7+yYMbE6LOWGx9S50VpyKbkywLxFTQEn8XGqMCC2ayqsT8NI66j
w8zzOeRjUpS8um3qRXNq6CrLaaNF/mi9YBSbr0RJdzZWM2Axuj3IWZ4eh6+SubFI2pnwkvTvd1Zi
iS03MlV8b2Aeow/7Luqgw/MNhKgEPZAJL4ns/8QEeugInqoIf0HLHNZTB+s/L4pO51XOH8Nvfz8e
v00jUxeM2zoJleb77hF675rZ0CCY/eMfGQg6kTOa30D9dOpcQeNfVdAcMICE2biP6feVQP8ICtpP
nzJiCQe81irdn4VYA714iyVS0Y8Waam+2K64I5Eutu07OS34USynMSQPFzzIqE1A3cmGh5d1q7aX
t8iU0xW1/pZT+Zjxy+qxzJpEwLLAeqojIOHU0lFQ+M+V+aIGNLMsL8WaW2WG8V5bnLbBKnJxzh93
ImqYrTLdXTW4h4VhrqZe6pVPb/vJ97cNfeFXCW5l9w1DIZalHG5Bgc8fG3v6IhFa3vsYcwzM+Qz1
zkOtE7tvW86D3INwYgrC9ikg7z1SQsMlsl+ksTOScbR0j+dA8rfrb4W2sYaPPICgZRyqHSzHGow/
y3RtK3raxuxXvG6K6GI12mGG4XU1DZPpeQQ/mAbbKd2Pr+oESZkvFNmeUJYNzHP/fPDOYksp8seD
c7caYQBSro9hXiF+SSJPDY4bx4qvWQRDcz7THo++3Yq0MQI4X42eF/2z4VayQ7zwaDlGxFg5vfS9
INTaWCMLNAr4iobSHHHyGEe45KMOJkV6AV20087nDjsBre6ACrXg4Dw+zyID9XbKnBcxQnsGT/37
TQgHlffqc+nlYdaa8PySbigaSxxCocrbeGlwgGPvX+dD/EJ3hTE5zTiHfxoMaxuuVz4vvAgO5Ru2
IUInFpcuQN7ap9uVlSQQhZpWGLhehMrobvOkSwhjQhkdaQbpEFWyiwMLf9nBT7yfHpCjabwoCXba
EKLJckoTX1lCq7o6dOrtFJJ4/1u1eX6JbHmvkr51bLvx1/SwR5X0+i1fbxKm/yywIO7H3dTpIWIF
xaFXDevElpf2hFrDgoDLkNNgOOQhL4f7FTYBVNp2kKqeEN5HyvFrGyVl2MVGQ+l5jQ1xDiSvt6nC
ku79AKtQzKqOQcKTzj4ERYtcCbkM+A4pApiGspxayKxVEK+b/taU8iiLSMRxW14WUHByC3Y0sA2z
O3cm7ug4vtSyAjd8MxX7DXEnBDzO2HXirXy/FOodyr3eZu+coZ0wb5Xs669OEg7lIKjTO7jXokrT
pnGFyHb3zm+7J81eOO7smrFwdQ5sRDLDdQluYOXi9pWbA+EUiOtbrBsdTpa/FCLWZWS1OFtBiakx
pWIIHMeUMxuodBtwvQ9nwndaetYJpm4WX09IVeLXDZE01k0CoBtg9Z8eTtloppDBEQoR8sRqwXy8
4+Q+4JikqBiVL31vhVO7hw8ED7yN6rRdgXTs0gAMZwj3G54RsyvAmX8YSMFWRTEMs3Fi3IRsIG4/
4NmFzhddKQIXBNVF4aVeCnRCMjoVy/ATdEOFo1FlxGfN4LNhluqDSfDUgxWYo9zHGSOWXBNISvvj
w1oPtLXm+M6TScnoYPgq7SW2lwK6UEsYODSp4yn6eGV0lePb3WD/cxBxX7wZBwPYUFTW/NiaN1iX
98LO9/JhLuT38dr2JpaQMd57WV6ZQBuMlEhU58KpXM6RVFDCwM0C0HinHA3qlP1qeFBHf9ROX9BW
FzctScap5mCfbzvkU/NFYDTZAScv7iZ4txiEjgHjJt8zBYjLyr6D0rxTKgSEpt3b4+rfxrsqbiEu
H0V8Ldv0H+kJXFnMS3OvNyGF2tMNHaLcuhV7ia5XgaoTlVfXV84HOAZezf1FuF/j+fpT7nzsT8o1
soymnjuNC57hZjuABbjPN15keErNswoWhjApSwApynsXZr+d5R8fipu2qKIkAsMMWEb8s5TLp0Pc
FqalIFQ9UCLJl8vGsC78z6wzmbyLslIt4yxVl5ZRUh28gQ1u9jQY9PQdPxX6ghBgD/Ex3PrnTkLO
4wiF4+hxRY4x1HLI5OZMPb8dC3XR0aU+tqzeVY7BuqLDbLeZ3jpmx/EeMiatcdadK9Wh46tiktLZ
e0qxqXPeTpi++K+H2A4XD7a0KFBtZmlN/WSZjYijv8ivTL57kwgaMn3KKP7loIY2D+SdN8kWNdQ8
5adqlzzEBO2X6h7aw/BP+NYdB2Uj6tg6ybQ7irsSL7dDsJ2KaEIMSTG4UESpv52uh073lzbQfb2h
C3tTDmC6U6iUH7m/FrJeRmrIH4awaUryizlxfLWBSlOP967QR00IvM4oc7rUGN+0xmnCZL5P11v4
nrjwAouCmqWykB3xCbZqF/4b0Ad0VldtzsTVSO9noYqsEDPNrcekqdwI9Mn4WwHZsK9N5bklfqow
J4tEw4yzDyFqJX/jvVEDV4gxWlmJ//SH++BaGhJlyfLZP0T+BEHHcwgUByri4I7+/lMsLC5qPFJ2
b+YPR429iaVy49xOsvyqceLspl2yJS3mzDV6+Od2gqYAcjCu8A39lClbjyg9LxPi0kSIG7wqVH1H
vEcB/B/TMV+V4J7qWp/3WLyAOXkeDsi2ca+K1N1qU2+1ifnoetMM5p69AW91Et/v/mKcIqiFzyXF
zhW86v0mJOtmExMGnxSavYjE0GnvM3HBRIlWwYYrlXSeRh0rYcXAOsoDbeyaZWZELmB83V5EO9AT
756LXNktEf16x+Y9TucWx7IHbV2j47V5wamyFb6x/D9N2qunUi8tk5//5s2vAS1YUZwm6KE50XP6
RV5H4xKKeP0vhtXoogxDLVX7oeeC0GeE9EVranUODLaRUiH5VaOcuJ8IWFRw11A0gEXSetnvR7zR
K5/gbIkXPakLfAh8K9cImqrfSCD+uMWRMGZWVijVKSA3n9rN67c/1S2lWn8I+5l/Nn0czBeHjNr9
19PgfKYsuMYDSKZxejW3Z1aMdsOGue0XvFTo3J5bMXpZPwezgopDwAPZAwX+g7A8WFG6XWUYZN2l
eG8e37HcG3dEiX1wOoKmWYmySopMW+AaD/4xZ1PA7WxMMix1lGfr4KAer2711OPOXJTXiXGZtAlM
Jjbv6rhKTce34C3JZRM4JKSZNOmsDSewkq+u2GfQWaW43Kx8aJlyqELO3CIsu0//yOVzWJW88t6g
fhsnZu4R+0LR+WGRJBuoqCpAEPtj6RX0ArTUin6cPdyh8NOzpC5zW1AFqCGwW4sfKkRm1bnVhC6x
aHGiifpXvNc+KzDJYDqqi1q53VOiiXqrIOWm/JO2PUqC2QNWrF3HCY/24dupQU3kAl+XS+XotBEk
xMxerr0VVl/rENNJlqjXAlKMOjJwpikgYvDujKyO2yx/qOlTlabc2vhZU/RjWQM6BKtAKaJMTlKA
0NuN06Tn1jRTLe/ZqSP63OeAj3Mi+IHoYnfmn/wJ9YwxxGnR7h73+X8uKMjWn5qtjk7dXi4i7+ke
9yS6OQ3+jkG+rP+MjLHucJyzQ4QXlEWs7HlWps2Pe3owMc4m/gC43QrY+KWAhsbaMGatOTTb3EZw
x1/UImTwxkrxWK0WOyHuXgiLgulPUUn0mLls9qHdY/1l/6FsifEQqZZGqDwpWH/QKxhEqdN3byko
BNVZe7oEkPBeEYX7/JdyDGaMOYH4wC6Rn29VTAGil2kgwcMD9mxlLMt4QwMLWhQWk8rQH3bKylBZ
ghxpc/ejlJcadJWsSnWpsK9h047GfKGxaU8X+gNEmhLiyY6P4YGh9/xiBIkkE1hWAs8fXdtv3ayj
/e/q95p93V1FN9UITaMpNZtC0pDU9FmVH+G/H/F0rCbQb/GOOGx4gHE0tDsxB5Lb8z8wM43NeT+I
OD0EfF2KxHm79deCB5iwsa4hWtCE81qD+M1Tgl+T6mZP67ZQYSyYeL8V8LrDK42vZ2lk1WccNoPc
VbngCBuYzDxm4yAsis4RsQK9cYm5o8xB7H1qdc7qzoNiQLoMCOHYIBYpANTg9iVhwc1uGfEzvtEr
94zjFThfagKfQe3YXPorW5nG437l0j2DWsbC2TodYr2j8IBD+EpB7phKcCr8H2cSfScXeJ2GxfG/
gXkVyj/+gjosrEFqaP3FFjPsWvkvI8HwTp8D2TygdKNPV+Knsop5dJMtqyRC90HZfd+KFOmfjMxR
gtb1hSmqICGy59Sh8CLcgm9u/qHQBqgrrLXzLd0W74nKfp2fVmKWay1Raoa0hg+6agIWQLgvtqvq
YcaOknF22nGI0HAjJ6lm1ZNiupOjn9UvnzB/ibAlEPx2uoI9NyX43eHv0t9DWWpMB8sQJ4SjP0BY
sGX8KqalMbOVf0i6jcndBJdKdK0ku52Ch58qYCfus6PNHmrF2igh8S7tsuDG7ZMDBepaVp5jMf1B
FvTyWiKZg76hWcQ7kk0u9jE65q0ueo2s0+x0nmIIbYWfhPklPfrmLleAKI6b2t259LhdOZNSQlzG
8QdYdc12Iu8jqCobX535pjiViOFxUhzPKaaJrwKutTEW+aMzISHp2Jn75klrkIsSUUtFCVGgU9dt
Knbe9fdQyJt/yfjLNLspJk/uQubaeQcU11HJ8+JsmdyvoK+zIuJhmdKiCK2zWRQYkMheDYPVDcKA
ZrJYA1zbRHF3Xd2pMyobyt/4BpvRjv3yoYA6JNtG3zU3PsbH1ZcPXqTc9TP9cDtyPvfn5e/46dc8
Jc5xVCRB9u1AF2DETWhw5z2eADuEsKQljHQ7V427gcW/sxAOW2LCbigcuZV9PfM6sohjRGtLVNx0
YRQe6ypR0M8Thw5N2HF6Hjs8xSp+X3KH7tga8bONHniYs214IZDhLr+AqXzqMX0LOJIPZKi0svWA
soLIuwEFsoQeF0ltv9nlGw9uHU6o4V+xYzGvPnbG9No5xQS/KLmtk3TsiX+XiPyRSrBKnn5S9hJg
X01w8KfjJ44vMLT86lbhh4D+yLDOL/53dE6dZSi/ywGRTOSYJvLNdRbWulY098kUQzodIw78b8Oy
YeeDMak6TesTXeXqVKy+mAoHeAq0xk/xOPPidbttfJ+f7YeCFDsVjDiAv1bBC+jeC67iGkisokU2
AZzGVkkJR6HXrkz29XRNh4grLQdmdFC3u/xmtCOFkzBICoMoO2+mXwO5JqofgmsOf2yeNslem6a9
d7IWZks4lNtoiFzFlkDk37ar0bIhUFP/8rkg7hkSVLNlST0K/13UL9FBHhVXo/0gGPkZJyAzdAv6
+O6Wb8lRqtL6G0fGOYf2pxIWO+TrZbS4ZSBN7D7vwS61BNBKLDGTOKcD6TKWtMZxn3p4PPLZPXp0
LZsTtFIJd46iIZ8JRkwWa5FtVrB8lhSY8gZtIgR/tm4VCkSt5b0t12qKeDeCNYGDG0cIHbWDdVt3
MgwqjqVqEkAeitfNHJAWSx1duWGECwjSc9BprYGvcL3OJSBEf02TZyGJJz3IOCkdEOe+Ks8TVR2Z
DWno0BxXgUOtCaX2BCdwus3E1AN5JGL4rcsJnwydKZ45W/gGfoXfK/KKWDcCZc+j28nRl4oDjjby
4YN915DbXEBKAiu1ZQT0WHvw6YVsZH2oizOZ6Eat81YWWzVEGVh2VvYCIlFVBPlyHzTlCByzIqbu
nINiLwGINm6F2HeF63BSXqFrqOTWoy/oy5sx4g/deJ69hZsP+E2QW8M0M+M71aLM4Y6cV2LcnxZP
qLPsnGLgHQivTF55j0y9C14j8FW2sBbQ7Sv9JKfM15BRdQ8eXNATXP+8Z0oz18Ky4OoIy3ZSiPpA
HaaTFUv7fqOhnbBRi/kahCGCq3WpVtPlAd2EgSq7kjSrhQKloeO9wuR/TnfxGOUMlzdAxK1NMUyo
D0PHdWxLAQbc/GlwRPPPEOMbWq0uQMNQ6Dl53aHAEUd3pWJjsk58W7UDFECLO6t0NZ2mg/BioQ/K
6j0gdO+ejmMKl0UnaeNC9moHzWcc7A8CpAnrhlNBg16dSJjqqwpQVmIQiyEJ8X32h0McDXvRyCvb
Rx7BV/eZ8PwbkyauCd2CQrRr/H2i8Pss5MuS9Xtz6QU43dg90l8t9sy8SD7ewwIzLpO2IYRETXJM
W6VYWR/ms8jo0tcPg+HK3PTdIfpXjFxw/tux/CwjFUH+mmorc9R/RH6hlbP68cZhPv8ox8SOV+QA
Cns1AG1rkGO5QaK9sPFfc5eA+krZC+xsg5vxVuNxws+2g2aBkNGUJJ12DXRa8reiJpk8KntpLgye
gMhlMpPV6ugmZxydT1MycEwrTSkAMZHXJHjAt8dkH5yNRdZ6w/ywC8R6Re3ZI++y6DMmqzWedXsY
saOfu3MZu7GZwcuSf/mEYvb/F/NE51rxVL1R2rjXxyQYq5LX4RGW9OMlNLaJKYuYAQMYnp42mFoj
eErUOhJFzPuSALTM3/bDScuRdtMNHIleMFnnPUJ2VdqIEGA8yjH7pFNzToZGUwT/fpLrIfT+edKM
7LYV6M8/BGWz7a+1LwDzrBMC4HiJrLgGRj7wH1UIzYGp8dSSqhc7Pp+YZAECxYP5ZNLzrRGFE09z
oUHsfDA+Z1RgO6Cbovpti1oNQnTrt3ziDitWVZEFjhd48j9P8CMraTFpWkNMDgSLC+uwU0qRri7q
FOu/n9tc3/xjSU4Bd3cvCdcL0jBDChXL5N7rLNWOmn/zciKWNkh2NTbOl5TsJEhuZUhxt3oK0FUo
phSZc5M0JvV++OPpM0EINE4nA0QGwx2aLX/q+OAQJwr0mLLAoXWjfDWArMhwenTN6dQkOyGzWSC6
n6TMTIrQzfsIr3oeOXig/OzsGyx24w29xC1TsL2rtkOddhBPqEf1APb8472TtG/nHIWhzgF9Fbvd
1aXo1P67DgoWdsbczrXkTv2crQdYbBYvAlq/shNTOeGCpAdJi9uViFc8TO08FLa6Wb1M3BpAkKaG
IDx6GJfkRFFVw20R5rI+SA7UHHa382csFqcq4kyIXGO3vvEfNRoHZ+1Yp3d7FuKeI+eigcDGQ1S1
eJnURyHxCZJydV/O3akRRvWKKYwiMDBodAVPrR1DorbpL7Jht2aoPsDx8LoAtLiyueUiiULBd0ex
oE5PJDBqy91Xjv95IFTcV8Zh5f3Vj8gX/OwWL+EdeGWDXzUglN/3jnbe9AJxchn7zXISJ3EVMsGB
JVYKJAjVme0hVQFE+XWMKf3s0R4saFpv7q+N5S3gaqnfyoOC85hzyR4CwQEaL7pMr+eAdcgxe+BM
4c+CBIY5MFXaFCFUE0GgvQKwRHsjgyx9yC4bp1/OgAXNsmEAJ/H96SneQZHHixs5C+AjvGlwTren
ZUyA1nvYCH7SfQC7Woi+J5/oB/9PZsC1bqBnyWPn+rsY4fIu2DGh4NITaFbkn4q/z6esag+jDGzi
ZxYQtgkz4mcJgvPxTju1vtXHADXlLD7f2MgjaAoFgNL6+B8SzwCM6vO426tPSnWTmsm7DoUlXsnm
TpNWM0deRVvtJF5C7kDiuaawOX+kr0o6mc169oLQpxl4CUcET7zwd3hzv6reJ2kNLru4TVMHQEG+
zQ3NgdYswJ1QkgNS0vWTlNNm8VRd+msf6WqqmG7GrjvA7K7M69Q++eNJSzlP3oNN4gDhOMxe4CWx
Lf1LSsUgDgo7EB+WQvIm7f+s9DYgE9K6KiSfFrRgHTaodB1vP8hBCt4x9mFOmWXZXMCuxXPAvP25
1eFycea5HgFv2/78bjjJ0/JyJEFa+r7NepO5WCi+N9Xv72/KoKnZL0w9a1oM23YrDbDfeRLyvi8c
82q7J+K/PBYBS03xKhH62CGF9xgvS8w0niUUtxy3Wubszfv1Cv8M05cENEYU4jXYCKIjBHTTe19L
cKfdlhcAEqS0VRR6PkU91/Q8IDiHJkCHtUCV1SYQcJDxnrd6sVP/50potqDqH04QKWd2UoqbtSYP
8RRggf1GwxTlD/yEVn1lUoMp7/IBj/4Veyxx/1cLXjNyKOFQ69Ak9ohy3IpSZjlfMQPJ94zY3kEH
PqitJpiKVLs+JBwOoJViWIkW+YNQIkwq9gouRh+BafyrsL9fsDTgkSp55KJ3eIUBtDY/DM1cRmlH
Wm9DeNUUZd1Tq5vCHImQGAcQb/pJmdd9aM9X+Y2uzxD3miQRzv/uxyMazPFJiuv64JAZsNam6p/9
/5BhAR+r4q8s5q1CHRYDPOt9XFn+yzPs6NmvSE0KgBxWjVk8OBFwv22hvqJU1Cf4OZJOpM+zukKU
QX0AVGiVJwDaGH5hs3chSr0jyFNBUsqNJnv+gV+pC0dMxrT8gEFmp6fYVxVIWCeT5bksPAI2JRKL
3fvNw2cykjQGx4l1D8z4hRMaNm32Ib1BzIru6ixOLx0mFcgwehoYkcQI339duvF5gcMQe+4ticFN
ETBtBFcb/FNykBGbXBxdkV6oAKuzz4ASPJA7keKCxu23YkVEXxGo8RWnjLzFyWwTeCiLcGatZsYL
UYLNlXuj+4/L08ZS/+31wjCWa6TyGz52N2QouQN/vh3yjck/pkxrnriWX7rX9mLBapkXpfbtLW0m
qxyc/zTrB5YwDY1y/H+fj/GqqpeM4UKwciksV9bDCLnYTtto4DrWPfBXLv/XJh19PXkkVwX+EJAB
psur8/OWywormy4R/Oi8Sl9DmJKmlb0o4p0wQvKQOXtLjxTsbKmnFQgx8e3Ln9R3jQuGZeMtXwio
j0F25RpNvNKosEvT7jMnW4HNAtVtjYwejJBmOtuWyTL7jsVOPgJvS64YcIhdKBzzOOKAkrcC3cxy
GrpNp02rrKkkur98dx0ZqAcJ6ML1WkuLjynrr2ECAET+CclDEA+3ROx4Uv77ccYIKNv+6B0HKnAE
yjKaSwaKTN9bxSqiPffDR9sBidEDKiYHIHpxOU7wiNG5Py0SLQxyVMJ7TjXPQY4SXiTGhEk6fqXK
Kb/NxLyccQrbjbXjDEtCvcgiGisubkukMao/ypQF3Djs6UB2Zl0Jt50j2n8Jy5YVmiyKMXJwMe6V
G1ZbyHZyYXmAa1I1SArMBHNTcRF3OWpbyB+XHqPeezUiXHpeLtrHuIO7IesFqU9Lt9B4g+8MA82D
c0Rf4yj9b6xV4ROmUj4PQ2MD1eT4k24Z9wIkXsWjTBkqS+yyyxYjEEuYEJ24Z0YvqCAtJiwjGmRA
VZDXJ1l0uCyN/1hTnxd/MncdNgu9f3vh3iykWTm0C4FNoRoChzS7rXnrOeTp/b8SF//mMcaTD8/E
urQ9AJxDa1u2cnRGVtNzuD1ftVDaWBCjlwEf9m+E9jP2GRPyb5zG7BS+Z43XU7ckfPXvx1xbJDVH
fJYDkC5d4WNi3iCiay4VOpYgaib3I4NZrZI0UI+g6nAQ4fQtiA5oyBFuVa4hK4UFONNvcq5tpFMQ
rc5jsWpt9H3I8ZN+VQK5O0IWp8q8Vdi1XSKu2j7vU1tn46TOPe+rNlu1zFKSbjQdWFNt9rXEnTdO
IsKNJk/UI0u3yseIXdEeUpKw6QpziT6LH9cSOxI+q8/dLp4OkPleRQXr8cQQSj2MlyWv/9sLav8N
Iwz4g+pj/pQ+Vvw/lNuVXsbtdEWX8vGoHcyBmwwygLYbzxqIgJgJc5BebdIhjhgqKmD1IVbUjekQ
UlCKcszVa+uygD5z53gl+jcWwzDEUdVyG6QH0XoHi2ds/V99w1mhv4Spc+ABtVY1NfQ/2ZSwEVYm
tUkx+eCOvHtvbIt4FRsEVvU+GUBgUDWexZnjrC9PYZqiFSvSbtm7HCmcxgz+3T+A6xggtnXKdOn+
tFnBMkNEWJ57AkE6bTuOHyhyo92I1tthMlkH9tkqAbCJGAOS/VLp6JAiLc4e6jTWHwQ9R60JR7P1
D5hqr8Tb4qIPW/ZLv6PwvH4qTqx55snokt6UZxvnV795uGAgJvhweMEgseM1uW2cH7iTXtdJDaQt
SFLga339+iIGTEHgGCvgXqU0VQzTsfHUfLABlAY5bGsdeBDn97NHwq/BOihRDI/XjjltzMpvfM6D
v/3XEU/S0sSBVfKioPi1upa7kpSZ5xirQVy0OPWxzS9y4wpSEVlip04BQDZJwpIdn1B2mwLxXWLV
olx6P9rytx0K/7IMERMJgkpnlb4/POq7zlQg0+ttDE962Mu2MEsJ+dMXvB/L1ikUetvWIgcYENvx
M8z88x+wR8GqwAOqROODL7GPXjn7xXt1jyIEqfjL0WBYcB51y1bQSK5ZykJ2m2Oomd61BWu7exhE
CZNQXGwddwzN3GYHK/QdDyztBud/QJYiPDyT+t36b440eJZhyj8eFfc2Ilp8cMOCcBenl/M7w/hU
MbbhqrNgIIv513NIxy7ppuFNlPORUyzilQ95TdG2txN/M4LyNJHrTA2oe3Rda56CDbkvqXPvr1eF
qfblkgFFma9dxhmuTSaW7NOXZH2rCuG4iU7sWLQugx3Fyder3zLkivVyW/323lq5P2mzk2RxgOX7
mKvZ+2PK3pr3pF3ne81wHJjkSqp1xOwy7nqVNEly1N5s8t1nHXO7PqLSY3NR51nAq8MRK6hbChZo
aOK8sQG9owtvk1u5vyZCuKzM1QVY5JFcVK+fKaGnEgruNDTP6Ozo3fxuKs6Dt+mralthzxuIuMuO
onDPOtyfJtZv6oME6uU9w7btPTzxl35tOZRE1jSrkagTAfzaVCWcWB29Z+GwxDNouhImnvq4Q1TW
1GPpAzWmqqECUAb9ZKPGP9n+4nE4ZaZE33jE+vmCyFNWeB7zaR0RRQQnW1Ck6Sxbe7J7yOFZZJq7
Vj9fDUSRG9RIpi7PAsX3ee2EIInL/EpYMi6jcWAaNfx1Zmpll1+9qQDWe4c0wcs6OosA8kfGDLVs
izOw0TsFR4zmhyDOIdByFsYZXeeXbFbwy8JjCU5anQk4OShhjCGDfXVU1cqr3ELoD8b+HhgHF7bG
KCKrqCIywmbn+rgjEjsRF1wKNR+DYOzWe9qRf8nGbquMoQsYUiFPTwrhNmk6vCEO5IHTdZF7dZXm
zrB/MmeLGCKcJAnea0XbdwG8Bl82vZTbvPTas4D+UI4KVYBB2IfoqLFzaTzbyh4QEYrVWioktDK2
TkXS6CCXV9mKFoYh/9GJk7np6vqlFWwHrhG6eb+d24PwieG3Zr3PEPqH82S8AeT4gGOAPEg9xfMP
dVX/cIsiNl1by8eRO9YSxH0DQGa7bZUjyL/OwR8AbLkv5z5uJzEtpJrzF0IV7zghGsTHeq2eXae9
jxAZpXaAsiCAHtI+s0xihrjQWl1U65MEaJQXNvJKHigQG1gFWrx0zu+AaO3jj8xGlfH02Tm8+faF
Nusj4ZBqZpcb/ddKxxDyHr3f9e86XqTw7EAnbYLfndsFBAkQ0T9xy3ev66pzRKiSFtdbU9fx+pLL
NjNS0y97Avfst++0+sKXqfi0t7VsqNYQ/08VxBJBAngYowCm5/kKxe0IVh1Vcm84YTXWblU9kGzg
xsqwEsK/8/WUUf830FQaJQ3nBKi0Kl7Q8tHxGPieCGVvYhl4UHDeeiUrhOijdcXwqJj3o3HmqsDQ
n56oysR1ZPfRm66C/ylbY/8RXAlHynwsM1/DyorM4cJ3saFm4Ri0JiKd21jnCD+MamMWM6lJygVY
QJuaxlL7929/YGeUVYnNVPu9aXMBSgGwFpmkrXeEnOByPXPgBcr/0WdrSCAFgRPccLCt6rbJUOWs
yX4uSRPyeFWGY//RTAuJV9r8xbSOFJllFtqcrAxOSiQhb2+XoHjt8qe2Jy2PLB1rSe5VeI11iZfI
YTsYysXtcyFapC2+mHCqYbdHASHbq3pqCFgVHU7Xnc20r6Np0lgA3tRqjvcEEzrO5QOHQgGw32lL
0aZTzgq8LSNYP7852fHGErA6tELodl7Zn377NL5zEOJXWxyec9VHNt/L0sDDGrWv16VQ3IdOSqw6
ptGiIMinEZExKwRMNDdKhqD/Rx+wUv0bALW3MLAFih9qIaINnxjvVmlt37hE9SROc0nO7ZaUHhzA
altTGPeLvjnqm6asy5Ugg031qwyT7j0dfy3xsdf02zegeNglimKehk8h4A6fJW6bZ+xLdRYsafVc
aYQ11zqmhwH64K/YESkrXG0fZUkwA5DNttKc/9G3r44JK5CE97BRapfoPkCV8HzFz2TOwq/SmA1/
b5vMoY0iAK/xSqAwLzGzlqbp1psUS9+Qqkn2+F0gO28dH1oSJ1bwI1ByUnWC0bN6S9QqVHfoXIWB
43+li+f3fd7MmWikoYrD6IIZFgwqlBpNo9RooJ++wyS1haiE3doghTp3Udb/0EYcVh3B/Y6K2E6q
rKFI7J0sLRT3NiLJHn+L0BpERQMneujxu0g4+pSwQI+ECISHDH2h6/JVW4ZPog32BQ1HAtfBpfa3
DQ3L0JybBeZbOrG7vkxrLMSo5YPVo5a5qPZ/7XL88DnUQWLWls9NWjpgfRBTsWCueabLzgHlCH9R
bYzogMWi05zExeU0y4f07/GAtsN56puvPbUe0ife8eRLxnKC48FEjToia23si3kCSx0PJ22F4bRn
ln9jqWP4K81YhJyOpRb7qfOrkQM1MHx13PrkcTg5gbrcmUZGT2AxTYnYzvCPOpAmQOkjEcH5p+o2
7CLcBX3rNz9zRnOfWEbyWIxOpzSIvXpS4cZ5Cxly7JH3TXaLppY3LImxeptMvNhJCmstu/PD19N3
IZlBnZRtJMx00lrVNdnerS1nJp5EHHr+UHRyigN1oL+NyEBmrnc35TSO5NoiK8lW7vxPATpV8n2L
PlPkqW8L1pPZDMtcGxvbEE1hZniYy2maeqcZKJJNqI2M0d5TMuAdArDdH15oUNX4qcbVdVtCDaTD
LJMK1U0Nw2BILqkoJii4FsJe1GZqwBN/vg1cknzLmDPzjMzmauC7lYueYPhlL/x0edWRm7lFEETR
yt4+mMKIXHbzlZSEdaCZxiSvafhg5hbjkdJG5trzduAzoh4N9hcynFDIfdovSfFbiojE8Rx8M3Fe
WpYHyjY5120HQcAG90K+tDn6dhPUP4opA+Tfa6D4nFg7vWc3z1Z7DDquAYxocDqritP3biYe0qDz
EE9ng15p8aza1damh+2Xeo4Q55o8ErWJ2M9REJrnaQRS6zS28AEWLhBS4YNTQ385cliOwqtE/cjY
4ob4EFAiNBf5Jp4+UjVYpOjSygm3FrUEt3MasyfxqErBg5xxmLBRp5bz9rCs5v0cHfFNjqzQof/b
QFltlImHHPSeSqVvJVGdrO7+WYA50DTOzmwDBAUIGudNVHFWrLT9HkExGKoyLrpTL/nOkpbOXpah
3AlSErXa9KxzQ3arywoC1AkQnbHa9/XCDI5aJgnU871TsJ9aDOQP/913GT82Bi6rhBiT32OYgNJ/
PjCIt79cxXhDTJqbJhKewSVCfNgfXwwJF672HDYQ2dhHkjtRj5Lb4IrBqcJ0I6gKIrQNPfg2uWMb
YSf7aP2vYTK1aIqqkWt6tRq+G06W0t027VmIpKSTXxXHCEHyhinL0JReK954CALz+b9JKmYjIXdD
i0kGrqKzaDrXFPBNPg+t+BFCFJXxjX6GiykxtFgZnLEqz0j9oYEc80pQNA/4Oqjpav1XcpcR97wV
8K5Xzkp2zXUoPXRI2TQLk20UAJJYxip7KN6HOb/i/WQCk9nYwzAHyte6i1crjH/g4+ZFl+gQMc2Z
QX4KUUnaXbMJyrsvNLwD0U5UHEJeIRaVSNiy33o2H4WZQlJXFhxm8nGbtcbk8vooI7BBSyHRsUbR
6GPdgw9Zeymtho5G3nZvJCuuz6sk4ANGhtCXVmFrWpe+TVe2zyNq50p2LpRsCFCJVhBpgRhdEBIw
Zrte5hkEL15xOzzGG4pWbzILdaWKcdztQBRVpZ+VucHbiYhOhx43Kp6zBTlE5onIttMCjerrMEYr
UczkRBPq22zuC7m/lKCo8aKRmhQiCKMsUk9UJSepRuRRQBkDbF2ofDjdCBkteBu0xMl4iODb+jSp
cHo533H6DlHRMngvd7iQwrfytMfvz/k8SIxeDRMGIO+6saYmCDptiwJ4VGG1eWaUJ/TAbwYd3d1J
PlEPhoHHAEI/wnvtoRrqwJyxrAKMifB8z4MJG5t/z+O+9R0Nh7UH3lSLBb8k2APEZR6t3lfsjUNc
l4QuXk9fuW8CselK/gAUE2iC6v4ax3ewqLyE4h9HoyISawQ8kzPqDBMa3pQEzAy6BiMbB0RQk4Tn
k/MCy3AtsAIoKB67v5FilsqW4aWst2xX1kI5zqwf0nmS8OYvISNBThxFjVjDdFgn0iMgEVb116EO
0cGf4TIvnvq/b1Py9BdXyJZ7ZRN1FE0txz4alz80mHIhINQdrr4afDlx5khytBOMj8aMVGCopJvK
3m4EpkFBMmY3qGtn3jqlNYGbuuBX1HLtK81aFHZJ71j2ZzZ3dxPLE/qzE/1JL+42ZReJUKFkl9II
EOpeymJ8MmuUmTk9rQXSXMU0iNyGqY0o97rDhQUjQkGL0bIpQ1HMl4rJk+XhBCnaZue3+lhZvH0Y
SA26CY1pjhYaYhu8/dkwfDX2lTJv7L5ooiYcQHBi6lMUY+DghPbiP9QPhFXUik5QB99PP6csrP8L
sbQOKbVAYX9LYiBMlSyZYVmBSjJ7AuAuaLbSl3QcNkvIOta0Emgrqju0yaZKkaQb0qh9mkkb3+Jp
Dj/yFKAYHffliIK3IRf9+jheP7OCjw3BtQNsKYtqaR381jeAjPD0rv62DPtMezPcVfXb7h00XbLd
4YASfGzyf6op2CpYlKdlW3/cE54C2vNMpmb+i9h3+4KElx/H1FlRD4NsFdmer8oCFVpU8MProP4W
9MFLzfthhGf8Y0+lxba/nX3jPZeLVi6UDiTYvnKlaMR/0p8ORh4xm5F0rp1PVuPkVWNFxeuNxnmU
GTdhfxn/Fwr0OychHwkwFjdx1U2C2m6koGJ9MTfM3opJSnUWt9uU8ydfnYehPdz5Bl1pSoz04IPD
Cmqz5Q4W6b/ubMsnkNyx5N6wPhwA7G6/HuGe6dry0DZ6s1qkc2yt4AJ/X0K/ErWKubtRMXsU14ol
RtEOJsL8wUW71LjxHfmH9rOTd0DtuKQ51REqgJ5X9ek/cFjXcLxfhpwfb//NiLzUwXqrA6PXYDDS
SX7JBP58FxroksnedNUHm+RnOFYuSuzqqlDzjtSfoImvmX3bpRsEgcA8W1pBKPmVUFgX0R2WN1wg
qG/sMQyg87QuR1xWQS/+wI4K05iu9t9/fwK2hhTFii9z0T49pZG6Qr3b1fAQNKWbXuakH8YJdav/
Is9Mub5KCH/FzCK+KK9inBT++wFLrRc/kyt+TKAkeEGOCDA/ytPMVmAvzbKptdvK4P4o4478Q0Sp
KeEyvzjUOLLwfK+ehRs8qUw6b8sQ0SArOfqCjEXK7e6IHsx/0VYaIm9MUMbm6sq0ASgUjZQdEUNT
C16PNT5Ns5yI8Itq4wMADlSJ/kUTClowb+8wMInGBWowxjilDlcNJqdIuanTeVPWo5KTolc9NFxL
WwNbFZ6chE6+LgGSOmAFLwvxyjGQd+h2MFvvqFGHkG+vayBs9cn6Tc+iZktLUbThKzyqRv0lCMBS
wZCYxvaBi2ETUf6GxR1FQsoTjjqZyEDV2a9JeDQ1hn+LqR6AyLLx1MX2cCsgtitHk/waT970SlGw
0Um4X9zX/tejIhjPnf6g64fh6bpkbeg1K/qq4pmfs6Tyv2Tyge/f9oERH+JOpP60WzqrDeNyOaR+
tNoKJ/RloTwiuLCKyUFiuL49igCaZtSDTFaFZ5C7whSiaTXBpY0O/N0RYuJOLNuTGvd+/baVTwsK
lZBBESos2f9CiQ4pNdo1dPCYOsE2Qwo841cPMlANPyVNEWiQJ1NV8bl13tj0WY/TTpDo7q38E2T+
p2qbFb+CJmAREzwN5P0A34XIHFzkYlGzL0P2D21IUMsiqiK8wWwZxd24HnjZFnf/wY2soOwgg1ue
IFLjR6dzZPXSUlT8PedxoL4OkQ85pW7hQdc3cXtj08Q+U9WmYjDY8WQNbm0c8ZzN2D6+Tl59hROf
ZdGvuCY6gz0H3WPtxQgqfqw4lsMi3s5NWp8o7ksxS2Hiuu2iY0+yV4C7dLGH1ZSyZX/MjrKln86x
OcrOFjnE8lYE+Ch4azBTs49eWIdm0WvyjUiLQzExC3W0FbYxq5SskpFW/lvdl+TwIQwJlxfoWkpU
NIrOjCaq2hRctM5yKJcRvmqZLnMgJLJ5WipHxxieODeyZz7bkv0+tihzxONkDVvCK876SNP1VHlz
2i1v0N//M2SCKmqwPvIHpWYwCUGd9vqln3N2J/7oW9v9wC/jAZfaVwTcMS3LUg+9sb2b2U6PqOdv
3LsWm7K1zzRpi/dqPUC7/thlYqwQopJezd8WKsN9l/oIlz2m8E6xBTBVESixO9RC/tFefGyotmst
MY53Jmnhk4vAKK0Ctddk2YO6WAGJqBF3YLgC7qPp8ufG+zMRRsiqI6XEKlJY3Gl4y5j4s8eyEb3q
3A9+Ln9zOCGwDhrohxSLgVgnamTJE0AGwl/1qC/XxaoUw76vfNcGFKYOmovPlYfUgMhDhQaxWleR
YUDSs56OY2ck4UkzquUftqxevK4f3s5K/y8rM3ve9xNhQ/pKjDGJpNXqVGuueoVqpAg0HvWE8BgF
SbM7S2R2tgM/x7t87C3DxKBqq6vxdbrSOiopRTBRrba13FE/UfjTTPgIU40GnfxkuiCMSZPgUKRK
ZJlEvkDaUloiuLQddUwhZjTnFniXLCKdxyufNQSUzOchj38rvkVMtXj3m6IJNDB/oP7lP/Pw4Gzr
5xDpgIybqj7t7S0zeJn6u7wVK5EZBVjf7jOdY3QFHnlvUMKMYtiqS919wUE1QWAWe4+IrGGz7OQe
VjHRkSxuFLWc2bX85sqDfa6iZgmAVE5Nzje+deMT0YVo7ZTT/1awCobcJT6ZWgXMk+4zl9zcvauM
+OsoXhqZWd3BMhGAmBYomzDSsaqM9uJe1OK3k/GtV3rTxuHzUkJIzSIYZBibtUfXkk8KINNCZL6K
o+eaRx1weJNihscDmFwhX7HgmllGyfeHz+IG/I+uQJF7NKP3RDrWKAZZxiM1HGcWoAR1llvhCf+p
knxhcy781XyzZVaDUm7/rCu1r7Efm8+7XHIrn+MkyU7nyA807UDSlIWy9WV5SW6f0NTytoPMUiHk
hYttWXy+YZXfibmH4Gv9bZKTQoMIwBxI1HUbnwCv8Hvjaan1n6sgn3RZEdC6aZ4v9YzGCgc6rD0O
tq4lbArqQH1Y6oSrGosU5a1dDpMnq+VgzDcceeb5NgtsBmhHhUCSV/7yGFcKmBzYGzI5EDLbc7Fo
2ZKWPvwEhTs/tvWGT1LIrK2Owc4utDJo3XGrhfTKv6bnjyOA5lJrcfWQ4wEee4PwCNqjscWIAUG4
h4br0s87cC4NRMFd5GFpjBkBljqIl7KvxPW6oW/laJaVhdR3TqiKZ+4QBpnKGA5YYpjPaGSSlz9k
6/QLAxwvyYQ9JX3/mSSgMd4gW2QZNJpTBM1BjEOAIbp1AeAohULrzIV9Aqqqs5KgUEgMfGMIcNsS
Rbrg4WwB/icrHiX/GsGHlUlxPRMVoLfAX+J/6M6ZyQd8K2r8UXyjagASj/42oQGVtQz2ClRE7cZ5
xXehddGS6DdoCjL9ktaUxVPjdyHQG+inFcxT/knb311Kw1lv8UW7Rd5zLdJeY9KJHZRp6Lkpg7+x
V5feZ0OG5Kj2Bz/06GQ5/YqcXHXJ5CrRlmfvl+xWwTugRyETFgDhm3C086SCET1y/DHF+EAoUPzF
/3WyEvAg14d5ZkiClPvchl3ClE3CSk6ptJ7C2tJ55xlOsVPsov0R0Nav+NOkMMw39PPOhg/luwPk
xRBGnvUtgfpXcl7NLl3+ltRLNLjjsyVvRiNABsFcyq3w3UXAeYjX+RU1bqjYbj0hTZ+HhGSiBBKf
sbfckVU8XBUhy5jUCv/GaftmeACydj70Ootacjc851HcF1MvdGv58Nthjs4K1kksPna9n9jGJetO
VstRoMZMuSMlpxZO8Smd5HcN82Ssg20/5YNnzRDd82jyLgdCkExVmIOvqlcwtn7QEVL5A+XCdrmh
AUs0SxloBbaxzhwYpDjAg6qButjrPOQJcB2kP7/aeLsgKRc2LZDxja7j0JP2Z6m3yJ8J5VNg4XVq
UTFFc83ET0zVwOZfTS/5c3yyYa+a3jchExwjvNPtb49XxD/JrDDu4jJUsLiO83ry1yI8GPB7rtOO
03nVxLtx3TpTihip9X89hoWlEg9hK7kOCx+30tB0SOWAZixrXQpB3voQ4v8QmAUBxsN9EjOTEnvJ
1VHIda7fI8F6H2I7RiLvU0BCd2lhr/ITMIqqGpQqk0Io/JF4pV0Lp3KwfmmuBOqfoRERQCbMFqdI
IpOXIDqe/rNvais81xQ/764O4qNo+pRVvgR2FHpIQtGXMAjEStyRrSL+Uyr2e0Hf1amjtkOsinaS
X0ouHF+flovgc0R8qqMl426yBu1NpVRUobDy7fr9cvLrpe4ptDvgsatbNh2m/BgpbhudWNXKxtHa
6/EoSipD1v1y4qe+V5E37lyHcP8rWM7uyPnRGU9dGvMnEscJht7m9txlzEfPhuAYl8jDA49wx72h
nhYKgbH3zBmLPrrtAIhxJotdaS1+/QdvG2eORsJL1E1cjyQfL4lSZUBxtfgLq2KwLoLTEhKtQ0iH
WCkLKHvWWZt/LlDg8cCoSQ8lMfk0wVAKYt47/afngaGWzLLLOgVZ97Nzs02mjRSxBmaOpffi9Mmb
bhR/9iqAcdBwJsfg8ZyddpcceHUOTtuS4Y0zEhzgRH1vGaifgmIdN5VIAMuBQEjqJd14Gz2Ys9Sz
yrbLykTDljl13Rsv249vLpc+rDLymjDFbGgzwVIrlzn0KO6QCWdj9FC32I1iUD9mxD6ztqoPPhIs
P7oQWcpbSfYB3pEnScFxWlWbDKuZbvS3DmriV8xxFucqRWT0IC2tzSlQs4BufkWx2KxP/MXfDbwm
7bdoDox7yxHKLhf0sesJXUCJXbq76v4BMaimoiIoqFBxJrek40zpLXf+PXR8AgTjMDtYZpN/Q4f8
IcsyL8G2bqEc3n8YPJKVTWJy60NcFUOCJkX1ZH1HWENK4f31Y+wNs8W7DUGOLb++jOdz+arPGSJy
WlRthKG9KYYD4f5vSe9dkPc7eU9KZpqoyV+XkERnUx9yfMwDb6XZ+h0Lrh26O38rA/8AYW5yLrOo
YoTLOt5PU930bKgIaVd7yKI3eM3RA8Zm6AVEsYOvkL4ldZ5oLwTsYUzaLdHPYyJgLsK3Wx30TpLo
39jdNuae7+TYbDc44hqCY58ZHAUWAiXfKR6o3fj4c8ieAbcgQQBFVi/Y7G8RVMkSgeAT6zr5kVQa
1zER4RIP2uOFpXmFXyreM+UkfoPGIATfnnUidclbIXm97OP8zHWDtH0e7YT+Chzz2X/KWTAMdJm1
YcsOlrXUKrYL6CRlg2ZMNyT1ggkgLxfalSmQ69DhUjJe5Eg+G9CihRRFoZojHcjE8N1HgaDdCU7l
pBcd17B14z8ku0h1rP+WbPKJMhhgfuFGuFMBnTnk8leDRJbR3yNmWDXXKIpeWWsTk696syUd6iTO
sg6Zm0UVz7A86Sm2gVW7AzPtJZUoF77ZLz4wD0J52ERcSY82v/Pkuhxls3frnEMoG8ny7nqexqhV
RPNG1NxscE03gmiC7GSl4Z+TRtY8kiJ6WAKluhp8L2yr+LKpFDRKYL57Vg9cnnm5JyxsxkEn8KsP
ouIp7SubERf432aiWLLEoz22CEBjkjWQgKHP5YHPl1ZiXR7vvIZe4uKXZJtQ0WZiDZterWFFfHGf
wfQXSKplrLN3TjnrPAUnt48MfltFUs/mAsQyxgq3snjnnQDaQCKQKDN86rmcs/PWurj4FDARUyrA
CCldtOKD1Rn/jZjWuBh3u9LU5NSzeQv3vSWKZwncRN4FQ6RGKMLHPnmEL4/eLwNwztbvmPCxPdq4
oNtDJRkmKVrY0Wjt3fEUtOH2K/IEDK9MV3NGJp7oZKcf6FufVJtmhS55gzR0EBpr/MvA09G6T0oY
yuDUnvOWaNmtR9XjTdVBgC+4HNsbM5sJK+Qoywbmuz9AC6ypEGBeKEs7yLd6U2eu2AnWwSmFoItl
JkwDeGCghFzRmcaQk00DV2QtXdUM8jtRYlj4dp2IpLxJR1CvfdSSn27YpNy47gwa4VKGKKOL7i2P
hJbFbVh1g/tlKxc7hUFLHzAoCcqFpTy+sPCynhzrteSUlrZy0qluq7QZZW2XVWthVn1efDFxnU8R
o+hgYZMqcvlWvMmdoPc/WQB0miPwBpx4bSCRvHAXb4Qkt9U0C31mAfYKJZkpdJOGsFcTO1M8TP1U
YG/Nxmdv68yKV3wTSFbp+F4VYx38awYxY5VDqeWHE1MQCRVeRYoLNaLVNTI0J8Nn6BED6/+DOLC0
4WVCirDo4r1zZv9N85BMoaXnDGlRyo6kF8LQrZjxlduUEmfNGaUwvlMRDyW3r4YE17Qs9DFfxvkA
F1dg44lkXSfW0T3Wp/L7M6EDNQ07PJKri9zEGVkHl28z5O6iw1D1YtSb60MZmkojQJwe9e+AbM30
ztzrL9N4cajFFbGwGBjQiu+YX4+ld3F4NyjMa8NXG+aK3Api/K+TUwXgN6tP/oqY1T8WScYsSwCi
+t/JazS0MOqznpk0YEm2ByfiW5p6resDw7VbU3NxFR7TgBZ50s6Z9h1V6kQMo+tumj4GvqJRl0am
lIqm9aFivq6phGQtgxdHF2LeR0EymbcQvWvV2Ho91tBGtRRLdWBKh7h2btDB5BmXQm0NzJQWSINb
gNylJt2ybkMnKqcbJl3SgJawJj9uhvPMq0LJ+LtftuQEXFVhTmvaeEWsAKpZowtcFpHTHN436Gne
t2HU2/BBW0KAPMnq64uTPCbDhawM6mq3Gsd9AEZAFiyW+Lz1AyDiO/MCWXYGggdh71RsQwDMGV9/
rBU20r/CQTdA1smA7xmdR2KH66DBKuI/4TKRBtR5aDiOXp5CaDGdjiY6Or1aJiNc5CdIo8TcKavM
T3zgWX5thlroLosZr0q2rFIJq469O2NwKj13GlIqOGTCJtsJZ2EhUYKfqoulBi5rdclmZqZ0c5AJ
Usasbs4pPe1EVQOry1vMcjGuk9KBj9c0adDSd8p9s9RkOw3vYUqsadyXDoXKh2FYCmfkeiK+rcy0
1oQBQoiGUe2VL+FFzzRgVfDZhGrP0ogqG/x8u83qhuNYkz8cgoQO+q3QtqdN+rWhVIvc73sNeXN5
twckYpVZxTQqOdoDeY5x6hY4iEcHdGcb/Qjy5aHOTBxVJz8cs1LJxc4B5BcZnax2gRBbM0hRtds/
hJGLe6GavXWcjkd14kmR7e53p7yBue+M0xYE1wYyW0H7wN34MXlNHRtyBZUplHQryXsmSxTD5oeD
OjhEVMB48VXoTF3rYm4zmPEWaOVQp9qoEGOaeYioUSR+Ztqc+xClpYCsAIKRFKbvWMNI4+fJPJi1
PBUDG958KEsPx3XrFekbTEn83BO2x4mvxO4Hkz1prdXOOU6kEpkd0A26445W9gx6Tq0WTvIwgtn1
exZR6qqe9cAehWXrburiZDRv4epm1ycm+eBVVPr49NJIK28KmJtDj3xPlD8d3Jw4ge9fNO4BvF+j
HdsxD9pFu9zt1dxmSE/zkhLtOFeQ4OR0OvoiTWJWlUqahUQ6wZuIHCBfIE5z4kmp4AyU0a5fB32a
MamnSDES5SHkg9GgRevMZaPE0DnrPr3lOyv8pllLCJXGCD0GsxX135balTqV+k/fv4fSmsnV1fvG
JvlQNdB0YHMEt6Avz48gNTjGN+tY/uByEQN03WlwlxSDJ8ycbVmnYz5KyW4MUZjArrBS46a4PtIn
vXF3/Mj+MG37UO4yHqt6+ecnfLpRxOdT6BEWN0t9hc4K4f53bY3vbM2pDNHtdl8XGos+XvFmUa/K
zEg9Oy0HOalyXEjWL5FCCmeXsjhYb6cVXFhxbkkLw4HiBctOhksGwMI26S06J3bsP1JCAnSur4ux
YL5gSe9GOMRHzTvnq35Asnl+8vs1eBYiSly2cpN5PkDZYMw0GUu9hOvBaER5EL0OUihohpXkp9Wk
NQYzVL7FsO3wZNFlQA93F7QDsMku6IbdP1KOC0NlbOa17azTOglgGLdTx5fVLKVgSdmPk/2/fFQO
fjG2ZiVo9+rDGaIj6N5/lp1liqLzac2Dgkcd5+Wev/yVC6JUSx7z63iBISTtJiPd9Cv4daM4URT5
RO4+AUiJetNvWGAGKAZc+voasu8CSLVtxcGiKpyLh2/uZbySvtzgBh190zdeC8ueAg3ZaBtxc6bE
bYWs8JshVPRj6e0uk0VnBupX2evfSOhPbeAJsA4AwaT1z3V9UuEKkmtPJH9PMrSTUeY1w7meFfQK
08jFbHUKxz5MgdfVgflCEZFItZr4ZRPQ7+kIrxx7sWyF5F1t8m1ZAJXmPGaR/YSZXOqfcOfJs8lW
EIpu7zcj6jFMiUbqccFG/iIBt65Lnb7riIljOoffZEISYmN87o4NC9tfL/Y5JEIxALUFab2/Zm3M
N2s5Per1flNSR6yf7GZ5hOssYVFqFQA+48aCYqnWe7mNn3brPllqIVv78wGMryTWR+fhVu3o37w8
Wz+QWFZ4ABrLPaaM+XS5dGtMU57HKhMNRHmil1bI4YxceHvVYZWM3ACwQiYUPZfXDMfP6imDiG8y
SgphGow658S3YYFlrEWsIluAVn9EquK6OtewngCp3QSEfHA3xVvoUJsXXQbUADukHNRAQlhT9JgA
jKujJGfafv6tckXhZmktU4eqi1xYqAQJHy0plDNOjqFdJPx7tMwHIIU9LJ+G33Y4BVX02FURDkbi
z/lAIHMSQnsGpcUfD5UjdzQK/q6vGwJbixe4ZD2QgwY3fsvzPRImVm+UFG1R4G0/MQClVijAfJiM
4Y64SVbTlnsAPDsdkfUKnINAVtWjihxmlKm0s9Gnz5rC20+gt8c+nk9RK0k/ql+lc8UFiyO+g81f
+Bx5/SpnsiUdXcchqs92nausf/6KVIh//uOA9XEK2eUaUZCfsS0JGXHFaT6lyBFgZn6bbM8unBVc
h3nDwkyVKGM+PjyxizJQe0/LkhU4Hsqt5yRpQs9TvU76H0cdQ3lIC8P+l17iD1wiEaiSuhvVLTZ0
mbOrowmfry5IuH8tKOQytNd1VCoQWw/SiTUbuZ5We5di3swFYydhM67FkBYasCm3FD6/bT7jwcul
BDkpHoi15WCHRyieALp5OyHU34amB3YdLOLeg7rAixKO45QcRudH4ka/anPga3Rx34ZIAkthz/J1
8AEftwlLC9u4jERDXXpOtbfHlSv2Ac6CO1YuMaKN94aYP9NOFcLSi88c/fIiNBUNEZdspXhGfGmh
QFpZqq4CWtZk3+WuVIqs2Izl6hAq3ARd6AfrlRBfvNSElGNbYsxJv+D1T/2uuUPJqQ7aY5PzCiQT
+l30ypabg+CYH5NRTiu9Xps6pcLOgut6fCAlr8kRbiCH3Hd9SJfx9buJzvSUiHt/owxDTWhsMTU8
XGylZaKh/oPNykxX9e8R1pSae9wEZtJg5kMbB6Zq5WwTcy5P9fxOB9kTkEd9wT0/x+McUT6f5gxC
TUsu9TDGUFucjXTXfundzGe7ZSRgOziI6lOaoXjv/tylem4pHZx0fbZXTVnrRjChuREZGUPbQwW1
fFg8vGp0drXfH5FopLPNkddBXP4/vOf9CKP6fKKHtiXc/w7JZ9nltUZvkxuIjz8gc644r1A4ZgTr
/FfAvccBchHU+l6bKUwfjvOGkXe8N3QMoSvjscwmjDr4dJiK6U8VAeBk+Y03G0c0MWXII1b/FTmq
mHJHYof2obPoIwoU4xTjVdVF8Y9UTYTEXK53CZgtU90mu8AcgS9Eqp5bgs9brsFl8vErrv7LbTJd
/aQ5k1FDE0q8k8aHfW/OEId60zwZspfMVSTk0wxMb/G5OhNeqjWrgGSEqtxrsHa07735/3Pu8CVu
yszLzO46uMGP6hJ8Ht3FlD3/HVG33n/JWCQUCQP9r8/dGSausIUF4AISNVb5C8h9X0f0nXtNGtqa
s3tGkxPu95OKb6v9XCxDYODC4KOLBlT9aqXPQ4munk+2lBotsmems/xt622vfN99LHQCTOC7Kfw3
khelwY21EaWAUKGsirKQU4iC4VK3wKe02TrlzUcnxIZ4dDUjvEzlqkH/c0ctYGAiqKXptN0H4WiU
liwTQkl7vkqS4dN1WXrJrLi9NiNtkBk9dYXZIHEbvSaIa2//HZtbBiCG/R6T0kFvLUGoS4ES1vFc
Jn/iFtU5kAZx4o8JjL6dIOIN/+1tus2wYwH9kXp/kg814kkadf0hS+L8CsswqK0osIAZ0g4ZucXM
ru0Yl0JHHkT84OmRbPuPfPrzcmIMul8hLhu1gh4yIn/JgDmcYXV0r8kngka9o2EIvUzcZsVUoteY
dHaLYRz87BLd53dFTGshhEOOeaWtbc3g/7NKAF2SkWlxguIfIkccvevLt5iRCzFdkJuMiwTLy7+r
OUxTxciHd3RP+V90vxLL/SUHRtBnmSjw3OGnuXnLFL17B+KNp4WIG9DXzYFqYY+B/OmRwng72pon
sBrvaKxNC5a5wlu4orMJVxeZMsK1xdj6d/xdRKVRbeXm4txY/5tV14CY4OT1s777KytkQ2CKl8ts
l/eqf6ubcJpb8z7npxDXMszPkTv7KzmxPx/kl4yJ8nnmFUe2ThPZ2qjQRlt54G2Le0SSk8f5/YMH
CEA9K5M1j7ETBy2YiiQfU7fcraliEtGIFydzVCU0rBkIdUVsl/GHf711G8ysa1cepSrQbF+UVt/6
GxM4aSUnpNVBj1DtBw9tMpF/anjdBmXeWrL4YavQzKdTq9mAUp9+DF2aRLzEEtQdGGieO1A9Wb0Q
6JaQQ5C6bqj1M8i7o0DkNnwdMv2JgDCt/cGp0gI/7lRkb21+PbRTfS7EOnDdHPJHCW07WfEvMpBe
bMdDUyq7ssKuihhLhHCa42MuuxMZ5HV3/e8dkM7w5ce7MzrXZucoGUtHn+z49NVVPiqeO/TOmBPf
Zm9orjoHnTOzjgvlRQUX1VLWBF6gnKDYqPnuXZL0UqLa/lwJcQPL+cvmr/UIunF8gClLQF7siRlD
DYzZddh0l/SzdkrcZT1APkL3wAxgWN3u2MDiNuweI3Pg31QeLddzFeL2nbIz/0IxVg0gIv1NgD07
+jq12oi0gf2bTMt1nwdxdP1PzK8pNEWpJFbIxVxzJHbQqxl1Q0nFexzPGCySvIDEKXo9gyHKbJdL
sgTLXVbtHKnhS8KG4q+A7dyLARAneOtAXo28NfQYUWjRrbOchL8FmPR3LhwSUiHtsusIAqlvKhq6
VWCcZi1gu0N/1mzH0u0RaPVwc9AMo0Rj+5zkgHLflzSwXN8LRqgCWzVPIgH4w9vOmTEf/lXR78QS
1zbX9trX0TpPdTqJPlpJAq/Lgfpa5lkhR+XvTGIpre8y6JFOm5iPJNkIE+DrM8J6XrAYYSQZGzg8
foF/+XCUHqvnFFWSE02PYd0WDrCiczEfVSbk4yA1Tm4D+zMryKTL9EJJdMAX8CHM8XU81KObEmBQ
eP5v67nrfBQyVLW31/wxQ4nsn8w0KtyDfMpQBaBwORjK1avntsfGRfpyDyhYnyrW+IaKYRx0z5eJ
GmaKDlXfKDxAD0jk5KzHkoeZnY9MEP7UwMmPQSZTA99LQ31dzS+Ydvu3s1ImgOwH6QOesSEqTX2a
oyM4eyTN+TWTyH/rwFV+BPqVQ/bNWHpFf0MrrXrNWNzbFt/U8vRuy4Kj79aEFT4gspneGPs+AMAs
pfmMFmX+wO+Nc9Pe3EYoAOiRWb/iIZMkVqU0vu+ZABmxiFAz1jaCjAEM6jnJuvz9kAdC57F5z4Da
XgOcyR5TvjJO+S+aPQ9j2pIb9/9FBvH+hEsu/VHLQfYWyQUeH90SCtWeZWXKw2t7Jg+21Az6Yg3H
jQACRfGkrMje+kiNvTP2HdUm+yKKKm992I+6mP3difOnd9U7Uv+hfdoKJpV6ECGS6w81SLLNjtsR
+8TmYBSIxsP78hyhL41drsEt1CV/vjHMsQs8LH3b5levtlHsprEIm8LNuz8I3a05U7DjZe0kGteC
LlUagwdSMXznEjxSInTqGFvsMjjo8CUqmxkJpyjbYr9rpV0jJ9tI/yuje5/MyZdQcM/Y73/n6Ews
9YZOK5oaEG09E3DUfL6Lc4M7wgeas3qPDdmVuLP+SM10K4n444O6Egtve4Pkr7C2YBQCGooISIGD
geufJvrmoda8MfwVHRqwp/7vSfJOmYlP2GifHEquB7+euhfuyILk3ZzWKm0ctO/umnBIbdLqcO2D
LwUz1TEJZu7iuYaH+C6dUHAL8PZuqsEf5DVpS7Ijd+4CAQciDd9pyaMZ8RVl474IKPnhddZA54IM
Bt3QNpvvsWGFv4Q392lkoxVkZXGyhkB/w8mS6b0dpF0B13p5R1VeznKlodxKkIULm7QaM2u2sa30
nKPp6Vfa/AiVSSzEAQxRUBiPUtvkMCOUELBqFpHziL6wv+KaqMzxe+VNUa48TYnjm+wmvmYoyNlX
fzom8HEZwoomp5sEBmtlyHw7MqehMIYs/Mhtv/YPVmUTe1X2VCxNGehfukAGVAg4vvLeAx2+uuyU
s73VqIzAy2SckiCU/Q6zOYSVefGC3OedL1zlmzxefUoEH0fQ2ttu2VNy2MvdKEAp1VpRMSEEU4/q
FmB5o9L92oEW4RWOE+D+fK9dAg2w1axzV79zlhPpaqOWwq6H2TupbTxH0aLZpv1oBFPtQNugGZVv
UzvjspY/OD/5hsqbl2n6hAmVWbd8dkIa8V+TP9+ClpNnocj5GRu0MmmqBmENGLOv+vuSEGMRvMMY
rgXUH8YCSKQxqMpdsmKh+ZzS5XqtAg1/y8mCYeWqfPF5lrKQ5nfMoNofUI3C/dsSpRK/CkvDIdxJ
ZwcOzsQAGtCpxeUIsv9NEUcQ3vPnY5xvg/bk4ZPymQkYs4URsXK/Z8a3hJvgWs9nREkZBmrRwyLr
ebZv6yLUWRNuCwIqPExFsi4g65gSy5K2mZQdGvAf05/7fQYOUuudCHPMesElaS0GH9o7tY5ACFay
vUyXuVjxG6Zj+ImO+TNvRCsxhiLNJmfwfLpMdXvTeRoIB/tskO3j2QDLfODgZyDfKbQ7iCIhrAxa
gQd+OrNnmv4jzDPAVur0Ecctg9+xH6IGPvGup9IqaJ7PmyvU0CPbgHp5s1ydIpOwP9Hgt12g0+Q6
BquzD/NZ0OQ84egLCYbWwC8o8NXdabwf3PKtoV52vfgNbBeRMeOzfUGTPlMF/AR1kTrsR0F4eHwn
HTcIROWNL9IcQkYkgQbXw0ZkCYXzcUcE6U8Dw+n8mwgy+JADN5Lx5JkV84RHS7rqJd0mR83/wSBi
BZF/sA9bqenweVzstHgXqarOPdAbXZ2xVQz3PHCDE1ilDA6Okrbo/kDP4nAZSlR41E1hCizcvQQF
GrlmziD2qw1gQGr9uhBUCc2imUj20eZzEH5Eehqfy17A0wx0iZ7vXbbZENhpqKBQNNY7SwsDSPsE
GaFPKzDzZBvCQfQeAdNUgI79hyXHyubH69NyDOFZTMl/Mw3AqFrg0wvemJXApqMrlnFCDHFCuOw8
ZDPUqoNa15ld82u6/xmIPQfPMIYIj4/y2k0f7wEmFkts4jcQi89ZkmyLJdfp5bCaqH/gLxuoLXb7
hqbxiRoiYXFX3g6TY0cQpFXwflL9w8YPM3awrJ4MkWOvEWfKyAhf3fV9GCUafmNz/BiZo0cplzUO
2yOC2N/MJQu4VjY6GcGS9tFQTyTeohKVOzUyOswwr8W7jL8uCDChc4rIIlukSvDkQxHi3cisvbFC
/VlRE21RcGZR9Zec2J3NRg6yiVEyPAp77sOx8wgBYQoAlYEuRxXUZGWeI0BapY6qotq1e8szLbSc
LSl6DCbEFygt3zVBBgYqexdeb1sDmne17BzPgJTuGzGOfR2qL+sOFsL4f4caaXU3DLBItInAP4qx
6ZalgmI/8DdmSPdnixsUK5mUMuLhLoI7p4q20bEJ3C29DUO0G2Ji1ozGgM0984VT/I47B5aIH1ts
4t4+WmcHmSKUASK5y94eY+gu3BVpqomGxVRzVp3Dsj7PrDhY/IDHZs4CbONwR0BFz1TORM7RUMUl
zjfIZ9r6MBOGuRkoCdYDjPKMk0fHq40tdKd2u1TMK7uHdBXxkFBBTr1eetL37tpJTeYfkI9fZNVq
G/849sL5L55NG2dWqdIsT/5pJKqwVeGR/nTgJ3Yq1koVgPKr676LSDjF/5yUbYDrKWlRvSgzDe5o
gtKko++377X6zJ1lNYDufryG+Ipzd16VwjSKl1agyPz1ez8KVEWe9MVjraMnMt6zzJTgDHvIrC7k
jC4HpwWn281rvPJr+pj6aVmIlFOWVIXbvuGhtZ9uzI8WTHLqkgLSgFRW7cr5Q7r9XckAVTGOwMeq
adI0geJpWasZzzDVgt7rQlUanGjBILw3ycIbyYNk8lb1I1lSnZ6eOz/UaHag9IMNe32QjHNnSZ9e
+MbxBnThhvS6o4LRCR1pUdFQwE2d3V9YI2x/HbUwFO+G1mX1PoUqtA5XU/PqCfwuDlJZ2fqGdVrT
HiF4UX0nhMwTFi4FKmIzRiB9iSw/Z6xpBZ+NsCh7458ytGBqDyRD9ibZE2oAhQz9Iu5jndjAQbCh
ypVqOM0TwsCq2LolDgz/tT9/zjS39HV9HWvr3Fdl6qw+phWNXDxMz9CkXTC+rbkEhTngVURlsNey
F6H8L09IbtRw0vUeQqjvGfgnNvWAo8oG2xItVr6ee/I2Y/KI4c9Wx0+7F3WvQEdJAQlHHRxfC7pn
/Noge2dFi6H1MB9RlS6VPxH86om6N+wkEZ+63TObF2uGwuZrRuXsNSKVaLgm5kE92oWf6nkYbA9F
MyxggYsfH3bfzCG4vhsurEcOcHpSHhWV4Pqnaffk9++k5x9BYJJPBtXwEZZSMc00gevlF1nTBS9D
UUJ7m5/RF37guprs0AZoEIipZp0SR2HnlBAcmk71kRXBeedouR7EBHTwp0JXJjBW8x5rgYd4LPbC
c5Xm3Nojh7WoxVcz1FoLXGjEwURajycxYNyDsGdqNuFjjkcdt40XHRiJNxbC/3Lv4emAhS+eAk0g
tjE+6qKIPNlaqRJ/rVji0wbwTZCoKQQhzE1525WtV2SlMYA6tmSqo3gDul4gz0bhiawYpyqTo5N+
F66W6XZbVLm7x42wANXcqmTEXKVF+3gbD2FcNP2pt9uRJuf7rzzzqAWwDxiRFyBYyr9nQLFgX18n
O+Uk/UFMOjNjk+8EA7RYg6LfsU+xg+JsEddWHzHFbpNrk+JUVxHN5jp5SBIJ7eVKZfCQe4xK+VCk
aOCOR/RJlpjGVHbEO9ly50XRwXddLEa/pOTAgiIOr5ofNKAOtogaEtHuC/WNth/W+bI7aYiFDwVM
z0T2g+h+RXlRB5JLyNoKJ4HZHkpAGiF4I6JzVzt5kd76inyZRzV269kxnwgVlWrBzIpTGpwUIyE1
hzDC/HCiBP1QJj/+SK9HqzegSGBS80BobkbhWGLSHw1MN5lXEROtE6gasnAoI5WLem0ZNbkJxG+j
tJGpkssllqAknwUkiOq6FtyVgMw7OYO3FiTpzOh1MW94aKHAxZyqWteIEKoadzU56gsI9N1eZQ1y
bodZppV/EP8hi1qD9M9nLGW+HUwPK8UXwOA12bjbKED8BgZWjJbe89w8jnk2cwdS82Jy1z8tzaet
vB61fGeoAI7LRVLhWEivFn05DkQj0luwy5f4iIijLvAw78qwBV7VkjPdy/SxpTgktRGy3kCfxRUw
84li6stnTbOdth4nH3BsraMVZHa6J9oUpTBAvfXoRrfV9mTbtnLY+0dZmze3o/Ov6mGnZXvGcNME
DqvM3gFRIOMzBkYhK4lInMjhvfbcx03QKvMZ8c4LIP+jIEYJQ45Pz1XcMSxAxd6FeTfaxqJHsa5z
csGnTDIWXnZ1X0o3bjS3wQgLo3NMDx+RlvEc3tWsY1+ecRXhhDtWuRi6VdjbozrGuEzZiNd9fpRN
Fm1hiyWmi0tkELc/sFiXKgvn2q5EZL6RZy9fnriS4RgT45vHIJO4CsIwzyVsgKN+mhknIjYNAd/n
YHouuy936RuPlz6vFbRGKkPk+B3JB8bv6zH+6VBuDRnvmMJuow8AQhBdvJq1Mp+PKrX4Ukoh4+hL
3xNvbx5bWrHcNqH5FD8D0MJuo+BLSzDPKjqhy4Kxq/Xu4qRpArPSZMsRF4rfWZZvH5bCGWcNySER
LvcFtyJExTqwLnn6wEBcqbueXXs3W/1YOFNbehwQpkIjZE4pGoRDYawGSx+OG8txB/PE5OtFw0bV
5mRW5XEgTxvols+ZTuQDgXutkdHSWKH8DK171RmZGGa9RhmkvsMiHwdMC5hvSqC7IR9WPiV3bgNK
5ypFrCY2NG1BO4RGJhabIsz8wZ6AHab/qw8muc91hqJuj/QzGYscbd5c2NvSNLFVKlcGZt/Yq3jY
xk1dKQmXsY+PMXr3m9LzbOtMbC2qAwVSz2se+bKQTc6Uc2eGkT+v1lBZCOaqgSSZZ8sdK7qu+dCH
q7FQJKfjKwQQo6E9313snnQCwD2Rn7VT7+zWmtVe1NsWJFinUs5kKmCAcoYLKls5rMgGV0fVYu8d
7SWcrOm0JXxOITlb2SBc1QET1bYjWoU7yTwUlu+AbpyEzCGVa0nzZhKyN3AT4+xhGGhpONZYz5xT
djpAoCadue35zhYsK8qI5wi8qKTOsWEaTiFH6JYKD68Ekl6RCMsUTncVytJrDlR1kUfmkccklqE8
bTgd+W8QMHTdWVzfhMZK3sDXkeHofOLo8dnRfLlYLNg5K2LmKYIRAI4577jv3d3/rLoRkjkOSxe+
uJ5vVkQXpwyUOHk+iTwtTx+sKPDdCRIbhfffhxW13CYEZz0s+msi7n3v1TGkunCIiVDrG7sMPp6m
aidFVlV6f6u3Qq63UZ7Vn1t9/OapEDZIyfesNaORa/oxWbQjMT2CaysgXjOioSfGi4wf6rqKKPqO
+N7NvVXFwYc1xNXW6b6KqlIIU8+SyAsBOdqDsWiE6Uel1VklsGKYA9BeWP7VGzyU7zbNrLGJs/d5
qcTAWOwV8045voV94eUb9LGJyjJ7yuXlaT47QgqXi8eOs10WGZNi47VkKLVpOPBxe794fm7PPvIV
6mkvaNnuw89TUCRLicMnw6Bwc4ArlmuGIWGYCABgEFEok1cMpRnS13ru4D5piaD1VDwueqma5wIN
WZsZknhKqfkaJTaWUPfzb8XHSO3P47sz0Ue8iStKBWACBv6I90TrW9KzMPPD4Y2nW0CsXqLL/fuE
/5It54C/3hC6Ic32bGhwuxKLmU7FXhgmV+AuBzX33OZqGGdLc82RKwj4XpSdCcid75S3qdSLksYA
JaPzjfS+HNiiRVF7TPeP35UtG2TxhDk/iSFyA2ti6IGvl0Ji2wf1fOYpJm3ENJyExGUouRBnesdI
iEmcvF9SP7MHY4BGCMyaEa806VPbAM3KBtopcURrq2EJ41new+NdPObVOJT02RmBcETgabD0yKYI
akKPuqJBJSt6suygeXc0Vrw6fM1FQUODchvjFmYD+iyuxOnCwppnAprsl3PyKhplfgR1riio/VVn
ALaKRs9mHJE62dn8oznmyppGTFED/Fx2Y5yu0vJlusHeP89ckQvMUMJxHCcubOVP9b8/MVnQLA1S
zM0+HC8NW58EKTarp8WGJ/WvIzZrTyoiC+n6iF7b3VDG5WbWSlwgBGDh2sji5vmiX33sDLf8zl8K
qfarQ0pYO5apY3rQkOevZS7E0k3XCPrh78mH5kHRzvw1Z9O/rwCaB4mXl1siO++Qnvf5YByhATjj
VOXJVNIYhx9Bn15Lt1Jj1S9jMPuBHCZhwsIxz+c5npaUH9jXR1SS8iIcrKABDlhvHJCy1gyUWAWT
NBAfLXiJXYUeJ6t+ZzOeLly7KQ2jHhWZbvN+1LhrjlBxM/0dmX54TK0sUqABolOIBbIlV1XTNvbr
407UsgmXrVkwg3f/dP2wS1iE0Qe6c9OOKl9tCNUM05qGblW1A20W99E9J1CuAvJ1pIkp5Cus53DB
iamU2fsY9+IbFKzOgCU5xbvacV0jehfLvE7iKgz8L05zoP5WVexQKLbqwl4OY/TIOk0P9oBCa/R1
lgiCnC9byYGhEnyUmgAOjaRjAKPkHK8PiE7/Le0qu3f7sBFZnzz3pkYX3V20wiYPHzeebFXOLFWh
TerKvredmk/OA3ADffSp8vBn5A26SAfiod25InciT+o+AqOoKU8VapiHsUNsnyhzlWSpaVkJdwRz
XtGYVxjJuobMz/h/OE9PtilLbaFJzYo7n1XeoPwEVEUVAn7Tpd/4asEkgbB4zO209iTz2nCUWWqJ
p7UZ1SZA64DUnbYzV7WTiY1IMlWaTJSkIfo5Bs7/P+9uJzAJ2k4SdHA8u/j3k+3p6cpza7erDF98
yRqpOuOtR5SO7kq/j5phiWszGy1Y22M9BvBOTmEGtejFSryzXSXEp/rzjJe17EoKeSHbZhXOySD4
FUqrI0JnV2Cyb03/mT+eLY/oulOhGA3Q2LVJ2SwzQDoCHnMPeSstWUoiyRW224JWd7OrWzrVYADO
uzowohYd64C25Jt1LILBIu5145p6YwT/0rcPEKK6s87UQjYLv7ELfsz0xglZrsEt6nXQm6+a25DK
YFJqr0hb5mlw5zyLzjyI8Qr4LW7m4t7dXIxNJ6VtCgX0A9eWTZiqXwNT3io+e+9wd0LF/XMmvFm6
tAO7Tp/OtFvtsfSvQfR3HFVkEpn5EuCHaAU+Gv7T0jLtkeZAKVjGW79KrY2LoGAAtPIYycf4fr/b
0Lvz4/Y14M4yKK8GLG27YU2/P9GpxAPD9B0dAPYNRzz6DotBhWW2Qz2oVnyttAb13zifNrB3DBHd
/tzk1kUFhLur9OhE1K/8GW1cJCULwTbkLWaLY9X8gEJwf3U/QxZWl84yC1YuFEIgxwXtOeLYGX3x
aknVHl/poJQUqzbe9Hc3X8eziDn61kxaI7CQBke+e7WrvCL+HLNhUHkLbEDPeXJsOFBuFbBxn7Dy
vNSbYcJFJEX/txB3qkKg5km6ScblUYrMR+q4MW6NH5N6S9s/xBjWOZ7jzjqaPMHEdJJQenYuwBrs
lXoH/eNEJx584dxoEgEFdHajNuzCzJNohJCkxM4XfpWBfp2DRfovmBG2S32GOyMuHQwN4hnD2wzP
6MiLFhCWH9ZCbdrS+/i5mVrsrDQEGILN7DcaEUlp8tJfYMK0GxT0OVTxeLbrB/RX9RQ90JWW6vT2
JYOyPKQjFlkPA6Am/7tQou/NLlPCGAK9ZqdQK4Z6dVoRtO0oZTlkR62IqIVJ6YIqrHLkAJzlWuwx
2wxXm08/O/7JyXqH1eUNDJq28RacxO+25KTtSLgXq4mmgLgajtUPV4r0yk6J/19HDphdHmBT91WR
BHvKOF8tegkku3bxL2ZoyIkTHLcPCHt7SOS2bmk8Txf33DTU0WOqFVscuxCBLBPFMXs0dasuKFuQ
fvIjQBfnwpC0L2q1iX4UmwGHpr1qu5hxEP432R5PiRVfPNtzXtDRRMRxlxPjI1UdiBdVBJQL22Vp
Xl+Dtv4u4QsmPZhUsupZ++1C2kECGGS9W6JHnAxPJ9HGeV34HIja0EBXXgnmQqSPQsTrsQ1rNUaG
Q6lY7PO7ge0nWyy8niPTIfial/pbCQkhzIPvLa0ic/EQIJys7zEjfegN9D62KjZqpW7fWSIhvDqM
qp69Fr1wakDRKQcA71wqX3GZpADEOl1rPEgaVMNTd1GHo8UL2sj4dSnWRErsAMQOggwHgolV0hzh
Wv0xdZ8DpDcEJc/VBL3x4RUYV75f9XJrH6qhpSINEnDMzzyKHL45PfcgOJaPi1flMg5brBpZX3fL
x5qsWZ5nW7A6LbMGIrvxM7H+v/LQ5MoLWVMiXAuROG/aL4zYVq+sh9eBur/dm5ddfJTVWmK6i5TN
dUdBA9pnGX9oYFQWXaHa3eJBea/Ern7SF6oiRVo++4YjWoJNypYs82hnccLJApdv+2FXhGtvTfVN
NUkmS5lOBCfoo+2gWMBM+aMDmocu6b6WmOHRL9qZfKK0dADjAfPX1vdU9Tv6YO9Fwx2lswRMsebg
YnPxC2+aNdAN/IfAYCW0uK/McBDtfvQ4ZDtknr2AWG4br1AMsm1P9Ovrv4M0WxCtzkm98NSWj2RA
kkelxzc4623OdN6CXq7K42H4QEZLsdrSzT26uPgaSl+YOvHNGpAKQiL7ezzj9aGHunxej17e+H0W
I6EVQEfd8k8TAwH+KQXlTh9G/QbteawiUOllil8gfDylxzy/Lc++jkOZPDKdB6w9jwwy1hGUk9e7
RgCjap3m6j79sHZsxrIUIGqdoA5jOx1U0K+SDL/VcG7K09tjUk8FwBPwOoGTwNE77c8v8BwrXuNl
4C/goqLDOfWvB902vWB6Am1XqFVazYQPYJ9zuh0umVJnV7k2v8e3s75YjIrVUGC67Nb5So/OBw5K
yNo/CR7u7vI8FveuxdihHashouHpzxGdglzS1DUmtjh6TGBn59PXtg5+Tr6T3ERsKL26sZgI1lZ0
6PSJT3/MP7VT0XFzv9oSherBpJsN1l5KUni5tMOt8qilrBTuaTca+Y0SIAvX0PR2s5qsDvIAgZ+r
jKa6OE4fzH4QnIoJfortpgpztuZdTaQS5D3MApcdNBt6HfJUScWTIyodrpl15RhqAkSOeZ3dP5OS
/F3+vD3mv0K8SHD3jlbdYW/spxkV2mOq3rpKQp1QAljNDqHXLV+PHNmLNzLWnbxRgeyFKOKWqHc9
kRlhqrcMq6WrkxlCgh1BN3mhxPjpVA95QS08+sspz7vNdktHZJEosN289KLlVwcQ51RJplosk91W
GwV9GVpKHFFFJGecburp96d3nqBBdNRdG6ZfIdZPGBYPIpZ8zPhEdV/JgO5xrXUcKdZ/excaZ19+
twzE+5/+piaIYJE7NhUeHSQPyxTUBAdM9fDmhIFOYELpE9gkIWYXyKk1sdFlETGkekQAOZLsueJt
PRJAArjTdX+qx9S9RvtTq7Q42Z8KfYvZp7OU7f15thi/omEMjvmyVdqhDM9U7eTdmJU6IfcYP1BE
1CoNZkgt8Dl4pioG7NZS6bRBIAlzvVwTOzKNZmV4UmH21PgTdCIOtGpbDyHLg7Lcu/woHy7p7UgR
5MLe0oZs8OeFyLvTm/N9GvvJgQqA4f5TANpO8NjZPXvROfz6gZM65r8TstitZWDsbVF5RYvS1wJp
LdjtCNjj5dUTRhFYosGWd6tMJQTwBVc86TMjSB5kptcS7eygVa+O4RKfXF/uwJPaZ4EsdlMk6b8m
W5p+RCjAaNSTLnYjMtmmhblnimEKHcPgAFe3JLtrDLob8gJL+3kupS0z+bSWfNSSdorSAA0BmD/S
LMDui6cnWZdPao5sfQ8RhJXEjMhWe2FZO3KdPT4QgQ2PTbbKLy0mYRsRZEJthIlZy9B7pTElvRT4
2/l2mGSxMWr2vm42eEQGS03ZbKHhkpIE0ouPyZIuJEfTaHBVwi0ktVXKRrlDkIzLubuCRWSjwk4c
dK0jEzaeX9Ap6AfAy2T+TnA6Q+apxP4xB566Wp9NZTfPmTeMFVbdiBgPSF1GcYGlfpErMYZboQzZ
Cdj3V2/l5fI4VYZjU2EHqDDVIQznfZU+n6sPPaqCgG7UKDene+2lMWrT3tCe3olSPIo9mW2KrAA4
nFRnk9Fwx6jDz4a+PdgR6wOHU6Ep1505ponh8Ledp53/NlUvyoncToXY6KiyJeNnaPEPyWpkTxIn
1yJOYuEUd0UCOhLo8tt5MG6uFwOs6GwWWCACoBSaYRaHAGWKoP25sqsot/EszwcGSJzfcoyMuUtp
I4tGsJOp4CyskUsG0HP+/QZCz0XzZq2qt+sKAM5V/KinB8zW3j1Ata6eINdEjXEAEcGbn9KihqID
clZ9jhLm6xyUUC1ZjcbIadg+QR5pQ6JG2uC+T/BoYG8Qp8YWFrB8wE0UL+mkThEePZebNyJ2lHRl
yhlAd2SZm0DO2XrB4xNfmCYJEO1HLl4PpbeksGeK+7GIjhbs9tuA4Tq/MCobCDICb4QFTem1Iudy
zfMhO5uIUkuqnaqAdYi5wjVt5wCIivIof7StekyKV0Jh84o9jevRuf1t8YScaRz9Om00s//ZtDfr
z8vucMSqO4QDwMGNP6CoOixI4WmDpvasdPNqmi2K7YfOe+GOUv4EIS9TrebmfUu8HS5bYjpK6nrw
UNmGD5DPnZcsos45H55UamTiEBAtB26M/XgO88UE2UQ2Q5rwwY8xJjg61PhgujXKfkASbB654z5T
STINEjGvI4es3emXPbFP9uiklrel4Gs2pc+/VjDbqrpCqJakoFXJUleTbzmIZhx/4pJqyQeM0m1m
BKqqXc6VZ4Hv1HuIV69Ls6gplhpyIKDtMTyfMFgD0Vruv0LdZSJhbROGC0xe8stO2pvDzmjC4Mmu
56cnBE7x+XUXVMIES3r4NgiHb9gDr9ZV+TtKUIIBcscX0qe/LdPNjWwmMc9R6G+8Fofu776gsoJq
VLuWyTK2qt16avL/uOrfld4ysYK8zXWHJjdyJgX3BIesPDe7NNUtgLrJAN08NormJw4Sxl6a46T3
Rqw8zKegGjPN7xP30V9CE8+vs2jG5VkR+GH4OPNS3e5wekdApXYF2HnJpOLeRjQ+WB5nCjhOF26c
jthSPlTMirKlheMFC05CLwuSs7wjxic6HkStm3YeAjEB01EoEfvVijXcSf9GUgK2ZsZIyn+6ZYm/
D9dlssdVEaH+AbejhjobMF61ut5V/pGax6/4gxlPdWO0c5TH7P0yVFtERdT8tHWlP9WtsTNUypdf
lAAkhbopNaKkMS8l1/myTs7d8GuQaSGcJJQpqu8YDLJHVuGWN8ogzsVKsIBXHCI+jo1uxxtQxwJ8
hO1I1p69Hk3pyQ8bNXmK/oTwtE4FnH4+qw3DXjAjl89Fa+C6DQAIht10qlzJs0F+q9oXuNlCUpEw
ntNAcuxSN9Rihm+terUksaNxoP2GkH0tVpkB+veodlg2OC6Yd5nMndofhRucqgtAGls/ufZ/knNn
Pu4ogQl8PpsseQAKufnwf/gSWlvRzG8SWIA+6stobAH5WvcfFToW9HcWaVdWL+hD4nJVrq8whZ7C
KDLtIW7F6kiSWhWMUsPHT3Vgwgt0ADuIIAaS583fpJyHO8SijPdagNELwZ6PCViY2ELVeCSJVkin
S6Ea2nqBLCeeOxsqBnPzWcHIjRLdUHCEwMETRXCJSb+4bobPhg5NUYGoUm5OTnFB2EQeJilwweJ9
98eqeeBcf0hrUMTZR0UKmGQbJmuknk2olpLNrXtT6pr/5ed9zAr/Qe6dJAujQSKql4Zxhrv2rlkW
GVTNF9LgRiDYx2yGCZeAh8nAw8YQqDcLXtDHS/WrABF+4Rri108YQfjWXpsBsU05++L4NATsndG6
tw4FKbis868Tcx6YDOeWd/B8DroniIWuvYGYTPZ/P/YI2wuRxbGgLW2bC2Nyd68POaisFdsY4uqO
Z2A9jf6hViB8ycDQNlgtRJm/jjsmkvYm/8ih7V1fxg4p1zLgFwH5qNWcX+mXnzIhGti6ZUXH2v2M
8irOpu25i96q3tJGr5+lVmzxJMQ0meci1S0VUZ8q8X0UjM/mFVfnQeDkFNg60SAv+6kLrNnZeddo
sPVwFdQBhEJncOdAEhPSxUY11OpmXO4DMH02Mp2Zp4v0EnR1mWi8Mrodl8cEi9WeRwih6FEOqsZP
LA4lPy5B0pRrZf4aUeWJuwc9xuoX3GYnu7VV44hm2VguLT251x8ZFRDMj8ODoxv1mGNQehD2uRMV
Xj+e+Ekrdwt60e+uyvabwcjvACDXpp9kkeYQIFpJ17fZ59CDXI4NeIQ9w0JaOfn0/UOUxe4+ZiIu
6fLX9QyxHKRdjg/hiZBBdaMKHKTFqtUAqkv2ZeRvghTq+vItgLfwD4OpkkEdnI70No1RaEZqRube
/6S/Ef2PFQtp+Bfg3jt57R8yOebqlK0zNTw2ZHjRKybNI4D2Y5VQPMBJovfZSi/rQD+ALwqVaYyP
EHFzx+mAkW76rneFH74/FWD5gLSxjcmz0ldolr6F7R3/fggducmky59jw+pERvFQih3N8UlNFafT
vlIgGjjOH53yps4gTl0I8ESsU+TLlvrAJ8Pwe6zKz9INF3SdkOZtgWhvpltc5vG8QT4cuXQZcjtj
9fvD73uFZhc4vkhgeKh3fuPJP4WlYAEoUgKl0QfsJNWg9sCTt1Dzyw5FOx2KHh0sufvviZoRTq88
JDT43D9+JDqlz36xWGUkccrxLjYbvdP1D0tiXet+xVe+RgTT4jyrDwfKo+88XY9WS8vf9HqMF78p
XEK8AReTGDvyXl7/UrnTc1PLRGD8f6L4zJ3FpZqOXQ/3Cy+lvljbMfnP4wOsFg/oRyP0xqtTSruI
f0A+If924sJK2McUsSMErDOEbUH6RBe2UJAUJp/A27QeyIdGGc/i4uG99z3S33azMorzyTtqCpbN
Vje5qW5PexSWLGaiXFu9Q3ht91XzxYLlliyxOh94I4jHlYHfcHXBQ5CQvuSetfMAPC1cRLv5YvZA
z+2wi7YFhYAmcUMS8WbaM9EAaKnHV2uWVStVoKc8nP2OpklO5l+RyJdfyvCBWP6JdMAmclNcKWWv
F/rdxnq/ZFJi3Va5NWDCE68IbdVd17+GNO/rhzZSoYjS9hs1NvK3eGkatRtkTEDUusH79BZONdkB
j9j47JnIqL6tq2xE7Y3KiGE+SmIrPFawHyyy88P+7jENhjb4s+0gjtIydO8k86UzGWSHN9YRZyM7
e2FAMOMdfdDnDxEv3xjd0xkSYKN+g4f7qX5DMM8Yt36EYxtDqrlehzsPkev0fE+TqQz8VIt0sgXf
6IP2h/UosbMbk0/uZk3BYja7tuBIk9+SzVWEhflYDmmAb6469VdE9pnIBJDQLAocfjQVa0gFstiS
bSW2Mrx2gAqt6ozcotBvbJgt+l0IlyrnWdRAoNCjixM6V5b9vnA0XZd55NXWGAEVD9R1x+HDvveX
VBElbGIKDCeKG1t+RupVFPdhASSG8ngxkCfkdXm2G/+mb/FvzmlH+k3xlXQ8cIov09Qh8VPyau01
Agq8o6Z5ddXGLgZZOgm5Vu4uYreQ8CLGaAq/gMn2QdoD8xtA18/LrSnH8JzW2EF4HhgdzTLBfkSN
en2pjpbgze0tTD8uKU0v6Qmnr0pwnhArwsKu7UIOn+Cz8qsMZfqNNpgksg1w0UypaCp8oxkrGAEW
mNH0is7EiNgq7v5U/jFdyG30uYXeWOgpPuLCD/AvV3+1H/TtlrM1pRHWR2Pgy6b1zR40eWM3N3Gu
KdWVM5sBPYt9E4D3uGf+sHCqSS6GGQxYOrlGz3XA1PKHt9sV0dZTBQjmW6UIB40S90IAyIDo4tXC
P8SCQMzSUtLvpHexp3Sob8yKMqBnsktGSDpwMsZGKWYkl+vms8qzaI0QP7K39IB8Xp9ggUI7Ge33
FCSNeRpWf5Ryp9+vOP0TPfaYkIuOqM0kdIUcqnvSe/IstCupJBYLXuGo1zLzM3Oh3Zv66g0po6Li
/Zj4FBmAlBR/iBpacWAFWKOnJI323M8KrGobiJ1dlZydGj9rhHyzSByg39vkBhiFSmcn/Y0n7J36
w/SdLHVQXfxh0gc1aY6dY5fvNohvI3EQAwiRLpf+O9EleClYtVfB+PbSlOIhEh4MOyve1Ojts43o
EKusQoEkGl6exbmOcAFPUV5LJ/vlyoHWzZZNYNOgxO4hCvqlMaazbqbT/QfQV6QwKCoESmLmWRDV
mPTOyMw0BrhRyWirY9g8ji84NyJVwYSgR+W7EwdWFVVTJxEptGE3uGsrHFN7DIbI2VeoFMN3Qc/l
wP1i1DtEhe8aa4faZZ+/UVOTQTeEtSd2QrAB5EpqTgshkLga0QeQ5dnud2jFVY1xCMeFL76H/M9k
dfaZvSPf/q6aFdNMz+N+C1QpgpN1UU9T2UXfwKFM75LDeJ0UtkDCiBngrBxjB4uC9DbmP3rrUx8z
UgoL1nNQIzNhDOAtBzlubozkx6IfRziRuRYU6MRuH0SD8al+gRHH5PL07vfN9CsEVWkNaM22Wz60
8LOIjDzJ48aLUW+J0iz2LLf2HfVJUV6nEe+b6BVra0kjxp1e4ssYoRDzH8iI+pqasUIazsu6HIRw
AhWkHJS3oa29xkLgztmOi8D3bTuodq7qEIf8XNM7uMjkzYbiGfDRy+tWTaXMzq2ICTfs1G3lTRJA
fXDCF1CMOzAtANtSOpkzat+/SpMJdjLHHx4NJAK+kDEQGN/t7igCEo6pwmQZr3+8X3+zkW7Mq7oR
XqGTcvxR/o2JkvNJYeihmb++533yh0BLe8j5zBQi86dYXVgSiDha7hfBAqeAVx1kSJKFu0oF57bk
QusEQuIF0HRB44DG07PIf4TmlE2JKUFzf3r1MkCMQugvl9a4XnBQTDPlFRz6Apyvgk5dpmDrf23r
aI9ydQdt5Daf2DiCuFWuFULXUhoGnAaAmFk0W1tRh4slUmAl1L8uz0O4SIPLrMX2A5sGYBWGN5JY
flttHV8uNpET2RTFRay9uOCKExR0tGGBXnpI2E6W2QOHtLNVZ+EF/S8qHj1pnb/YJ4RLipwJN4Ez
zBVvndgfWLcn7yI6G980bHzScdgHFrrvA+XGUukSEg4bFBg50rP8fTYLkUDXtcG/2sxk1tJs6MjS
CaebtJhuNZcsOabKRv+WxVo1nZZFlGFmXMK2lQh0OAMj5hef7qNrQaHiQHlxchrLP2rSvdMAoJ6h
xGIYpGcOqfGZ6iSePdqxP9jYY7YMYry1jqdRlEPlKBAfIEE8wZP4I4ETNAsyVkxusoO2cGbiJSoo
hMcLNL7eUel18NIfBFxNa6I0lve/n38ZsGzdAudpBrrYrVq2vmDPmMRQ/dMGB/k5At42dIHcEAyv
5fQoGKxI2zy/0ZNqtOZJkQcX8WXJSuMF2EM5v1W5p/+dSIGgcHSofW66bO3aVGf/UE7OFOrw0rCp
4lFeVRc4Y7MPQUXJ5GFTMhde+La0Bj1yv1S0ZeiURv/otbOpN4S34sUDNlmhN+EmDIfavFY8NHo6
nium7aFPDk263oO2hf5YBa+UmYwbVyxfxgC+JW3W9fu+vDfncCQu7a0IIrFW6ZAZXcIbvUAu6ZC3
3wdtK+W31QbFriHI608MxrE70bxiIuORT1FAC768lB7sxgGptaS4Efqh03/1mVVOnEGeLFPGpMWQ
skRPjEJSS1+Z+cE4L23uJ02AL4Pvorx1Bz4c9cP6ScirffUQyCe5wlsmaUgEa27/gpvcBk5kZQoo
Ia+fHGCt15SD5/cngqRKNwE3DPhZA/6Vq/wXQV4CX7Oaf4p/DOCsSs8ZKwSNmyf9GOYbRkIJMXOw
zbLlCYoZ5S5iXsTYaCxeJnxD3wCWnHAfOAWBGWOn1TTfLxtbo6MXSpaW7faootr3LLbMehxUW4ax
4P61e10XLMRPg30HeApNTT4mglQ4y6044irM8NxWm8DVDr0+6TSNlgcujDe/kvAJzO1bjlPWY3ai
RLVRtvIYilQ5wViwksph8bn+/cPh0GJv3wAGdWunRcJ6gTGO3LladSdYJsgHTJh4/0q1T+Ab6nDk
jGFL99IOli+VX/mY+4Uqaf/9KcGBLBACWjTgbMSNltA76vPby1hKvDc3b26bN+rwTIXpBobu5SW0
E8vOdtALEuQ+EVCPGpW9fK2yOEf7toNA7IQommWPIMHhGIX10rpb/d2IISG5eogVw5WG0qtVaLg7
ZA6QhlVaiV5QXzbkrW3WjzU3tpN3xF1yKA6sdLDJtsp1HYirWZC9M0c3uVetkz+0VZkXE7vyd/gy
eYD3nzz3kA109dNybmQvVlUWMWPt7AUMlcpU78hpq3iMGNipa3XxgEQbRCXo/GkZSqex1dSzVTHU
9ZhynwckjGgHziAFeRu5Dm7bXCWKTLGYbNngAS5+/vFLgbXpsqIZ6lOTErMfZmu3L+5ywT6NKumZ
ZlVdwmJ1ipNi7c4PQfAseT9FhBFvTZVTmoj5qHh6PwST98Agdl/+Vj3MunBVJEiAUwcco3vnzKAF
sgeggtza9d5fAjqOiuV/mmOwGt2RH0FZlyLG1CvjGxQrjgCGNjyeKwu8fDNW18OGU4McdSZI78Gq
Nlqct7/TT8v5FKzEDDYdauwzftxdfSaSYh0xRlWWNuAUccwhmG1EriemuN5DHYYm7KJBZeEzJx8G
MqJWKDYMf8ShIzJFjPi+FeDacgHx2P6kxb1so74mRn4Gc+b2F4DFiyYZqBqMAXUT5YWujZyLf8r1
NdjsaGahaWIsnWHj5tOCx1dHGnND/9BJKI7Yr3UGFXJ9vFDke52w18hLScBu8PMz8j0KevzGdFAJ
MC9oQFlBkWF0WYvQzQAVH0YRBqlbUie91E8OUxx7f0lPszJ/DyE6WdRXTOAQz956F+Z0H1fpv74O
FfPsZJBCZgIO2dFL0AloDJjp+Sbmn6NhW+zx3HzewmsnXEdO5+14aeDYZgdsGpKwHr6XLxsH4MYw
y9o+DlbgSpXdwWEc9C1IJpJ9q5ZDz96WcmnZaYYeJZE9DwJMq4r+/uS9J34fiStkzOgFhEX4ROsk
8mdQjkpRzZOnME6MbZslZqQMs4A4eAhwU2aMsRDxVA6nZny7+J9QhELiC70FBSrz9eVS5iBrBL3r
aLgoZ0nTMwmAlssLmX6JOkIzQstmhzkUu/l4uv63AZPGlGU2QTPCp9eEiC4VSTeM1FfUM4avi6vR
/Q66zQVw50hJbDBB8XNV+6jlHvFUhGbkBroRG8kOX0guYjv5bSQDWiyiJYjZqJLFg1VOzuhf4s9V
YFg5pD2nw/t0Q7Q50xQV27u48YESJPM2gP0Z6f3t2c2tC/+JtIy4L+h+LK/gSDJgZY/7ADwRb+P0
v9GSCX2ReTY2TkAl0vvbbO+R5nnfQX0xmSLL+zCC9/YsxFzruk/W59XoMw8J314vfu2nCBrHK24L
Rp8PbwrSvfh8aYvCsp5wKciZ1JyLj1gjBPKvumb3KHOQYcliHk4TTo2z+l4SRpZDdbwnunoAmhZB
P8FOSd0LZSda92Ky7QpGPk0DFvjkz8vKTzBgMLKncKbs8bEYEcaepwGfAJUvUzqj0YiZx9w8cc/R
5a1VLG8kmI7b9ULShbibu8ODglndreAycnrdcLHuN4tmqZCzzikmFhomnprxqD3CFACEDDvb5b+l
DuXYxRsc67Sj3Xs//cPhG7QEzxdxEGNKHjKsBJCj9+khEOXW1vv2+iviG6g4Ch+bcBaVzqwoGsh1
ZYerztAAeSCmtiZJMBL6BOUD53KUVQgXM2z6wE9C/RJXM0dkHjwd45CMlibeaJu+1I1bjMWRxPN2
NSL0g0y7CVHircpfDqcZfacvgh/7g1Winl4iRm2z09YpalVftgZX5BnOUSjXCNlm8Rs5X8GdoUh9
CJlPkKDfjphhOqwP/MqO4ltKIqCiTS2dMFPOHOew+mXEBq6OlzV+oM3RaLLmWjZgy44pCXC6VrVU
TwkaDA4OwgmRZHmPICc899Lh0TIe8EiZcYiOE9Usvw4p3Ly3GwmXA7oA2moJSVfith+gQU19p5t3
U3FZhbcBn5q60ya3S6ARIgdKkQemgeawAA1cm6c84RfHvlhysIMgyPqPsDmokwiW62E/zxhA/3QP
wFXXGKeD0kln9QQnj1m4s/SmT5m+DSnQ6LsBHhU51ZqkkybmdJpZhXk85M95Y1ebB51Q9M9u+pAM
8WSjmo5jeqi+1ClmJgfbZVn5p9bFV54mhFvQXrbVM0snMH7u8mBBHh3GUJ//otSj3GuiIYW5XRDn
J0G3lACYJJq1JxG1KHJCz59AtiFO2/dyVMlhvpQy+SEj86s6iftYv1u+e7nLnT8MHOKJUNdljfVj
/VKfjoJBNn24MqKx4Ut3fIEFjCXbT3U0VdXbyb8G73U8+ofulmiIPw+sRLK6FGjqbfBuVJt5Tjbu
g1br93/4gUBabAQ4DqC6OxoqA7G1jItC2cr8nWX347vUes8337BuLrXNL38PvmljC/xN732CLjKm
ki3aUnC7zn5BxIP0aXYzRVp0gQnduZqlcHSMjxN5X9Cw6lBQgVvvNsrXJrLIB3hltcukbvQkG/vs
E9YTWFB5UI3Knl1gAvDAvUIbjgFFSKtnYZEhP+dlFGD85n3uepZhMU/pwnY1qTW5fs1HRw+ATXms
S9vpYpKWkxZRRot482W/Q5CZMD9TpTO6bKtJb/oYWwbBcz5Ags9dEXM+zZSxg0+EyoWZ+nlbP9+t
b9gKChZpNLfUEChwZ6mAe2HKzLMo27H9BcBo2mHL4agp9jE90nY25cS1XGlfYk6FwozmXT5jEdn3
4MzjGtpU0a04ohJssQxsNutgDkGaVnfPwXO9fvB0gXlx3tzQ0tHhgtpfwzU85RJbP6USiufwWvf4
MOncycPzqfI/8WsOjJqzSuRxfX7UkxBTIY32D3Heia4xOi3eaCdVOPA0pJl72mvIcRDWQ7Wbw7Ex
MpWb7NfHP4Kcgr+PokucS9voZUf06vS3rJ6haF193aP3V/Se8V/ya45d/OIdAu5zuFMoE6KlCzQo
x+z1HXGFdnUtswQxV6DpzQEEgo7jkh4+NuufuKGOuFiUnECpch8jmgn/R/yadH06wM0CgHZWnkUP
ff14nOE+OQsUP8WGLn1GMjkFfjoLl6b6qYNY0N7S1aVDCkllhGcqJrvzzSkHJkEYLNaHfJzlHaES
9NFLB6Y1EMaWGWWty+ydL7U5gog92XQqgb6skEVyg9HA0pEKGW2tbVqUAKg+Z89TCRtz9ETZwCJv
0d0L2kJE6mgEkM+8WBab+38C5bYNxHvYOsx2MVehzrljV4TpgsEEiKI3irlmL0AWSBFi55a/u5TR
gAyJz6IYnYwxlaBgqCgumMctwh32m97MJjtqiB4odWlF4paw0J/k039Izc0uUvsNnpzHWUo/QK5h
hAMddm1KKQjPuIQP8rliDEIpFrE/Z445e35rm0XoSRzfs56jwIR2iS33iynh1yl3c6sFjRkG3F05
f22kqz7jamAlM+50SYuXdTjueEiW36PAL/JVxghQS7nwlqYiixnc/JSoRwoRj6/GRXMcu4xVs2TK
rPCi5EADt++coKxsWItvX7AAL9QamgaUANI8LmtZz9MPeDJVwXgKfh8ppN4jWVogl8ivCDT5BrqP
Wm9zJnUKoruIFj0Kz3373/H5SKCFq3L8VbYQln6LG4KEHX1dVda1MK8v6hqfAnnttHGmSzmS1RVa
2YjecI50LrfczR8/mU1/G3vudLJUIfvTk4VNQddKpxJDusZdRB2WjAUInbEqxa4948hZ9/hp0IN5
5wYOZA3aTUvmVcpPWZ+9ASG+b7UC3JW9/UD7u6QHDX4EaFzARUhZk/jdRJNSPRDd78nx6YAVLRtT
acVygQNEb4HzGDU5/qR/o/OFJy3LbiAAG1vaAUGg8/4101jcXImP8BaLvZ6DiemMGI38SxHFNY7i
fA1E+jVqJZeB3Wzzp3GqgsOHiklU4xDZ5yQjEBo+1C/xB1z3QkfIAYHz3nmc+AC5tUGQsel0T3Wi
cLeDmaUnJPkkIpzJy5H6XmE+f2yo8s1mKCjvHDzyQXqtGHlO5cxtLf9wyOmtUMrm2TqK0FQAD/Dv
ZufjQPd3h1LdeTkMOoPg/qCCbBPKTzcZh0/VADQ4jVF0EHp3woZ64xt3deYZv3ZUE1RYJqjB1dyg
zT/omUTNf/Rn+kUKqT0Wihq9HUMYz+TZbX6V7crlOlAHSaiwNecf6D6jdD8veraKiqssJZsvFEH3
QbHHJS4phPf2clNzB7sK1rT9Mz7nEbh13ledZcKhfZ7W4nyWVIEulnA+oi1TNTugZZ/+T8Fvgf9y
eeERy6BfFhh4dgMt/QKIECdLZcCL5D3mQvE58theCanDiPqklvvw49Xvz7TWGRmZLx9H5T3Eim1q
x/9t2YyORDmBOBAbPbzFj0+Y77jUHUaa7DdCfKPuPXbreOdjozVpwKxiiKid/sD8/wqmQP+t4yf0
4dCY3JdjAceZhhe6Fvj5t3eQn7P0JAJPvwf1Lc8A7fXAbp79+/Fta+oVmKxM1BYGoxN5yAq/YevE
blMvuEGVQf/lmWrZswJZ+pguVn1EfPgNk3RM0wC7zuqS3CIfUvCmw55dLJWWPKSH9hcQ4oyf7Uyb
f6/sDp37APxxPFTJ/W1cqsj1ysqJJTKF6uM/LLxYIA6e7ntXbrmHPuAEyZcgcqw82VU3Zb2jM6nv
VpiDTZEwfwxWg/6EiAm+jey+Cd2daOiKWjcZgrI2LdioFISLnkaWTBZIkC6dZkz/r6/PpQN3LHJg
4n3nTfcKiqNbIN1nZ/Cx616K+LWlFcAA/U8F9PV/coNX4ao8burXv3LUak1wkIdOTBrl8sJkuxzL
Mpgm6QcfD1qZ+mITaIi6ltJh+umQn40sr8YbM0OAKMh8rcQzJXswehkxgSi1k3H9nmqsIV8okHj8
7q5kyQYavvBb2FTTXG0hn7FiTWjJGfOd+2tHc9cnRa/2FuoHb48c3eMv9SmNvG5+A4xWhwvBy/0s
H/5q1jkbSi5CDRsR8G0AXUEOYH+kV6vfM0CqCgkQESJVykt4MsZuG1UYS9tpldT2a4D7RwExCb6m
PoYiXRX9WwhbrRy2O6Zyqmvig/RdIHdenHxBJeSoHc0SDC7GVCjQ9iQ1asTuO0IeAQW8F9KvSly9
lTmli90T2bbRO5Hb4uqlu0zUKI6kuEnFIA0Xs+lRoX96FRIxLwzhscN9ciHZNHMG6le9Izt12eIR
rF3hwCOCi8Z/rbGAxbNeY2Uk52T/C3z5xKRm3IVSjiv+VG+MnA21qOaV9l/Q6yvjA/p3N2FH2lVO
xB5kVo2hV4O9lJ9hjWKAz3ZJrGTPhMb/r+VQ3PMbaXeePOOPnOd++p9uRkbYPP3H6lbboWqEcsNq
NTHco3TkQEiMi3l+uRkwGlVLDs1/LKMY/w9ygVGca/aqinc4DeHNwyyMX6OpMpQR5MIARNy4uqeA
EwhVxZ75voQiGBqdDg0l1IrIl/SOBpap4yaX60xbQH0Iwb8Y0PP8/S+Y/tv3Jiv+yjbCFkntNIXJ
IXn6jXiOcRGORRT4qlRJUF/usjSkHBTPFjQOmK25mv1Qg6CFwwKp3Mk02n52Kw8UndTrBe1T4WEX
a8MfWqFEMbbN2hZ3uCw37uhfRetz6ta9dkTMb7jODCAFH8eSOras3icj2JJbO1jn1dfWhA/C5RST
/fixEFIPuIur5ybcGftN3B7GWHALBRt+yq0EMaiSPa7lPBHXUThNMb+AaF7+h/Ft9pNpa42/qC3L
0aNYcrhntaLjCPUBfRBwfOtBNiudctbulEK355qiLh7R9X1EM7Hivtz5d5MsttqZK7MCqrhaCSk6
3wDURfdbsqNJP2Q6qPAQuVzSIMO5rYCqGHztXXVkM3MKpfFNH95Pofeg92zsbolqs783aTAOsMFK
MzvWIJzBXTJ0fpQqwloHERJjxPCcLkEGeRwANkFvscs6l/mDiTb2AK6es/BCT1tFFwbW6YBNUX14
vITg9+ceKGKhSQQzuD9sxOP97cVOCCRiLgaDeBWBNo/MtSdf8mw/3awjNvieOfFgBQ8nNZlw0Ph2
2xsNtrtzklxGqgutQ0PYaoxAdkpR3K8KmEYBUq30suM4xSk590rKbIM6XghdqpbdlbbUBdNVIeIN
0XTj6Xy4reDPJXhYKgG+2Ylt5vKsyIC1pzll5cxXQ4J/PzJdzlETLnzGleI9P9RCkqs08KT+4ozn
pUMF1E5dx8fUgWNhoL6DoxoKZ8yvEotLN5iEt4EfhYkErg1Tn6BbfmgMiuLu+IRZ0O3Ys3HfQ+Yv
BYaWENRUqZNsoZ8mH+1VpfmycVwSCrgu0K2z+55npiXN60VFVbnUAWN1zEoQVMTic3T0FD3KTuV9
/iGzo1OILYu6ZYLR9y/VbOiEavLSeu4vsIKkZmEzmIiYMmta0nsgetO9RC24N0Li6xx5zf9OS4vL
pp1QLoFRO/Us3L6i6n1lDkaj124HS2t2UtgJZS9EIjtX4xXmG2O4Sp5f/QxkwVATsrdXaL3YfDuO
gZHhmjcCM6qyHkRNNayJFrHqd6s071WZECBhKXhg7s3blJ3CYyxjx5wsJw+dq8Ylo3tNbzuvj/pl
dvOJcNz+DN4khvOlAA4FD5aYDCKy+di17HJAfXAFYh/KSTEi94kn7ric9Ggev58waEPBGJlKxFac
RI2MBhSx1wrOOvJN4YJCYxNNnc2aBeibnmqdK6PVk8GfWbs8RZ2pwkKYupKs80v6K2yXSveGNrE/
LHp1Mq6AxDecYZdg6qZrLzHdlO4hPQFjF6gihwWhYMQKdeF/6ZDmUpBanbd66NKq0fP8dpI51VM1
ZMh4qkVK2Ecl2E0/b2U9wse/8h+mhSO78lDoI/idqzCXDGjDGJRBr/45gpY8z5kKlOHbBy8DxvKK
bnrrYb8DoxeIk8juDj7Df2IFylZxK+FdxirP9Us5I1rrGqA+ooPcgzQ8ORcojlqg5o1i1rZBYKA3
qy5aSsFTjSPjJjJehf1wIOg71nT+8KrekqzFRQ4teZWwFPC65XaZT1A3pW6yxCXMpSGlM//Xn+uu
hoL36F0em3fqQWvTIZSHCr62qoSq1cwk8pkyS5NNtb5YRXSmK5tRmTt6Uv8fECrlmJhI2tey+ZAd
q3vGH73Tsre88LG/YU3aSB+riizarkmhGE2muBuf2WgKamei5WOYkJ1Kin/WIhThG1Obp1BqEVL0
F91ttDnGAx3kmEgVC0zbI3GnOlE77tdxPSOurwsu+wgPCicg0OXLwEyWnLUXkPqFwpuHsOReudbb
0Odq8vjyHw4UyZ0GfsZnZIZmgCSrPNkLxvy3vq7qH8BmBUp4qSTiJ5HkP7oORrCfYfrx7BsAKT8Y
HrBMbRtK6lTRozsOOMyL+MxkRNkvbNqSo95NNz7gatu8VeOtYwy/B3IJQ6y3VloHwH2EH3cO/w3P
tZqP+9SypUgQeUwJOJ5laiViuS96+Z8G/2Kvq+OHUxjSQ6BucB0HF/pk0n5+0rXBQNYG27Zy3Jmi
8vcs7dDOtyBqt9qJv7eLR/KxyF3ymbgwRsd8ECmscCw4EN34XTrKHswUYVGRZbvOsm5srK3OrJFV
LfePLKdA2sqX+p5ceREtn5E7sECdxxXiJ6xXTNGSe5Z7zLOLujmcwMo6VvlcPfc4HnLlmYuNpMq3
0X4M8RCspsqvNa42FmFXmIJDsUqCQYt3+AyE+3PgvhPnr2flcnN8z8fZm32mPZ09077ppQRUpgFu
bcD7zLUA60JzW6tv8XIUJf4wUvXmAEoru6zcOPPEN+v2WSjGus+BNcQ6vo123MWXFB7b9uKXbWIB
9XVZ+musC9L46Zckz/3cHUu8hkqjKNhevs/qVcw9g44KZxjoADoN9MVaVB9i/PdbIHek2pSgCTMX
ZGR6PTQEVSz6M3PqomHDSj8T0V7grpMSlDmsfXHf0EIPrqVeL4h4pl2q9S1w11DxPTmXDG6/SGY9
Njow8MNxIq8Px5APbn0jN8+olIiONpuhAnfoj9K/kU4p7g2U6JwllQWHmEQ4BcO5Z+GJimfT7RS3
IBVQAmpnfKQU1Iyh+etJxA2M7luyz6wKo7FH85AV+rTmalAEVriYs9KP67pSilUOgmdPG+K6s88Y
tveaDRc3A/7yYGGvtOBZB71lagOln43VExJMxDHk7F1jJ5ZUHSdKc5XtzqZkyaV/cwkmRmYjL0jX
P1B7Vm4g5KQXLygCVAwZR2wroU98y1TnS2JT0FsYqFxBrX7U3VtWROZXu13hEmdVrDmKHqvzD57r
rzyXaKkWAF1ZtCMZHBBjSf+fU3Qjg+HbWZJgtvm8NFKwQ/FGDGpPBTfAK2djZgbf/co9M+RA/vvO
9PMIBq/Jg+NYuAFvyDCANuVqjHTzW2ISKeUrrIjZg+I1IqellWYOLnoNk0QXc7z61kTyLkLXfFb/
liHCpp+b2IR/9rmJZnuxeqG4C9gF4VRTn6GYYX/5Sf6D84Lpxpg2odq/oGKJLWxi4qTgULfkGihX
EJYfU17pj0BavGjIiHjAlbRRaJpZX4WOG6SGE6YAeG2OcY7qKF9MD4/Py/1u1scm3R8HwgdrHc6u
c8jF4O0K55i8DOijmTs+hkEy7S2+ltPznDYeTYAzq51eiJLlI3gp9AiATpfmxQTK8VzHaSTfaT9b
Ri6c4cZ3aw7Y10dGLimjflVewwA/9wYK37uTMwlHZKghPhbbmzXoKzkW4xfpnYwKkk7CiyyddnoD
fxPlClOanIKgEF0CycVlfs6oiYq8jeUIoM9qYClNcJY1NbiYav/MyjS0uwbKPSOBMygIESZ4Se/B
CKohVmxTYeV4xGdFlQuRBgMHbMonSMQvURgcZOzER3Y61WUTAdq5K9iTHTZjIHCZmUB9dkauOdig
PAd8XR2xA5UeEDtACdpdv+5SLlTW0ySPwg/cQThgvJ0l7JOXr29xyR/cb6o6Co1kjuI2F1956ldZ
7tEMCxTPHhN8Wk7DVezXCS33QJokmmgcIhyml42qs/DKOLvuHu9FR9P7TswgRGa5IXJoDSRS3xii
9YW6dEZVQKh6lHOGeEz4bsfXsyKDVFOG1OVAB8QpCTSQVOaiTTrAYN190W3t3/4q+CIJ/71dA5ip
re4RMelp/Ymo+yhbUpHNW8+F7w8GZKRQrn8stBdaCDBS9VAHzza4XLRnWDubfxyW8N7lOQ4l2LD9
3ycZ5lmCA1VDrYkxAGJTm+GCoR4ICyuFrTvBJyuduoIfXwZBASg0yitrLBvw/9ZPpmrEq+VkSeZg
VzBDU34XIHvfeoEInAPRczEpB2bBa0pH0Xs7mvOoEKWBK/7iyruwdRMyz5n+cUZoG5D45N9c2b5+
P8xhJc9b6DLg0Pox67XHyeeEb9jWiVeGWhvEnL4ih2pyVdzonrxXOFsktmvF04auYktcAF4Q8Zdu
ATlrDgLt+ER8Js2PwFZC0Cy9+F33lAhllG915FGgai7PggGuOHBe/LCJQgTOSk5C0sgYoSRdoTD1
UG+VfJEVw9zRPDkqozTtoG0bxz5H87pJesVeLffvttwelXQXpBVD1garAo1d42LlJjZMMI2ylLMr
grYtFFgepTg2sXIbTTt/xc3sVU2HAEysk8eEjtuRCbMCzx//61F5CUem5NmlxkBZB4cGOj0Q7AR9
hLeIJ/nSws2e2GAqNXG28RUTAXotPueihgFT+5rlNyZZDqEDZ6gQqQKPMhAW5nWg/CQkFEBpRdT8
DWUxdvavxxeP5TlX2ryCeMtueajxzCn29ut4E2xyJVqJ20l2Z51FQpL95Wdt27lS+yTLFXf2I1Mm
dox5VOB8R5sDBaPlsBIZz4s/l201vWsl4+lUXjXyMjw98iAr8YlsgotUJlUaXwRO6AO66jEzYnj6
TPFyEqazzdPGkZkZstWU2z1f0XwuJ/28vHteTFxNVsaGm2aGBJwNepMFyXbxKIH1BT1B3rK9XL48
DJ/A1UJtN33nt4882PMs4E3XllSufBksfGc1n11D2N753L8AtBrzDavQL2qiEeiH8dlp+pS7SmGD
MSvER6pNSydf9p+J9EIRCc2+w5t4DLMupgQ8UN9obUdRVydCAS/pAk0OvLHi0Yoec0FDayZCzCgB
zXXOQrIK+52MOiHNxYGujpPJU6+LXdd6jI0dc1yAXWzWJH97NSYtrmy6106GRR+TarWCSQifFlwP
aGx57Pd4CVRQml5mVWL7jIU1KDdayr6JA+oLauvLScHKVHYsk8Zs7Pjhwfxn4KpTy3WJKMj/uwc+
T6idS2UlEIgplGr1GlDNSFFOBGgS0wvM+s2rUnXOXfBGS8tIBwr0sL5wyz6qBuWFk8W3GdKV8MOs
wwgujHXeD2I8806xUtWqkkJRD5p0iIK753NaeYecjFtAJzcyI6Q7/xceZ3OTXIzkru/KC58Phoyn
ZxP2tIrUancveSQ4+goDPFaBh1BEZMUazLTc5U6/ncMlRjSDfKBb+1fLtmXlpx27FHs1W0c9YWhV
XLcS/4GSQBX1ukXzwD+lnCjhYKGG6t1DfhNsjJSaCpvuk9HAk8dCaNcHaEAls1RyjiRKSpKw7Dno
8XjJlgozgaWupUskU45PXbs9/vGH4zZzyB/ZnwsMLxiVIMx0ApYwnNcQS6x5CG4xkWXBGDrrTLCi
a+2dYmUlwhe3v7zXd6UIGOL6+HLe7YZ3JI4qwjz0ZPU0M2atpHiDfhSZE6TfPmmGysUmtsVs7/t2
ZEToBB1ZvhfRQGE0ldBLpVEha42BVwzav3AnsfB9yZKhbmX1Z/DZKfRmwpEVAVh8gD3QidQ6udv6
rkRaUnFh7w8AMAKBdKkWxP+exBdf5bPeT0IYKhfH30L1UYjazGhojQ1qGRyydPDQt7lmfNbZUq6A
czHDUpm1YjMLFr4XrTK+004CDl+fDgBy8TH3bYn1D5xsS3VYoq2sWtslXQfJUKtp190d670Yu3Md
p3cP68LxZNBlFcVw9c+Zpt8KliXr+g5dZMD/+fCqpJ/hRmbogXYy+yZgr7DWPwC17tOmalQ5Bo32
eFeE5ET+WrpqPL9jt9m2sjY9KpqgiM1P2NWF8Q6F1OGbAFjjlLXxC0SgyEk+M2S2ymsQVIS7AxpW
QXjn97QlPtTEDszMrQTUWz9GGvCuHDILjX4x1AG8uVdc0NBu3shMcovzgKIA8eeQxgmqYdHsbniD
p+7xTmC4QrJOThbxVRlFfk99y/miFKXWx7BlcANqJ5+NSih7W0mSHveY8641s8ZuUiyZY1EZQ3DE
pDQNzoEB5npoeSMnbY8QzNDnZfHts1ZimGI/33/3gFwzXI58N8qeRml8og5RINflpGwQOKLZ83Uh
yAfe112kqOA28FULRa8rdGGtt0r9lXDXfxWaH8suw56v2L0+5U+jP24B56HQyfRNfNI6nU/5WfP8
UjagqovLb6QI1p7fgRzwRal8cJsfw0ECOvNjm+7Jcu9hhcCnlvqlG6fEnfgCumuIeojH+T8WQIws
LllnBFnFp0Zvd/ohDSb7I+mtJgwCUuU2TKsalgc5PeRmwa0VZykInuDY7wQerCvIIOVcAF1kiXu1
IndLoqCTcBHhaQSP5DFJIQi3DTuWw9XByFc8helUFsXRsBjWPFW83azNM+Ddrb88AcHbZD/n3FEq
oT9FJvSM2vZ24IjAYnObQWoGi/B3xh1SSi7UPXI6yyTm1DIVy/qoFyvKts/mmdW/omlwKzTWvE2T
mJ3vfUUzOnTcC7wc3WxjAZv9NPGBxOtrVpmCbDqxizsSUzH/fZN8Zs2ikXQala7V5NOt04enloFJ
uuQumBsP/H5Y+EPBzXjvMwbQNJaEwJ4dHqS8IHecvB9o2iOjwGVWyGmNp1kBdnxicMsC4G1bXlhC
lmxyHwK2W9o8lTGuOkgHbpCM1ZSMf123HR8jxjuK4a9Xz8xj3T7Iqn/6ZlKtONypd/weSve+r+YY
qkCeg45VEdWCQvLZGlMrCH813vGG6nttnUz/vn+4jZyk/z3Ud+3KILwQ+jC7mQEc6q665+Js6Vg4
CZTta1UgjNxKMWeSVOWoJEsgfDH40ouzEoKX0+F8aq0JjyqkG1cHqlcGlvL9//aHxmSNX1jm2LdO
cCCW0VLbtVch4H2AWZ/1T9VV5NVIihgpGYCG2Aj53UzxMT3iU6UrJt+oEdT3ZWbPxSs7oJr1IE+x
myZCZeiM7PNV0+k1iliFuPcjEcLvuXDm0sBEKzOxDe5VNBrCDngHmxAeg3BD1g8Nut6MTCUYvuDf
Yvog1MVUAgdhHdTQUvCgALq5tfF1FiMNviQ4fRHzxmska/CE8gpoXYsoaxMNeHek8iQQshyxwAjE
PK3GmPWUp4PJ+KN4sZ8ZCrIRX1PTP83aUe1Tko6lzv8hJuNk0YZQLQGZxEtKwI27cYmDpIXgHMr9
h23KEYnK+QfEXyTx213wnAyBczx1PfXsQAbCHG0+EzWyLe8q/ZBnhpjTuELmzJ+2Ovk3/nD/mwny
31qA8GCfxR6jW7+pDZoMNPEJRRMSPTNYUNhPMtw2i2N52lG3S1C9ZJsl9PM3Rv4U3ds1Ju+v/u2X
kW8lkwenh9Pb1mg8kkuEPZY+Z0tEf/6oZv6PqyuykpJPzvC/xVbqMOMf3a61Z9pjNubZdYSSkylD
QhGQlcRFsIxm+SLfM+T1NHxho9BysUEhycXJPBReuhyNjNdtZ+awohtZqSuqrGkAsVUwp9etq8nb
WUS+L6QFHkwhK8CyPEOAF5BQdDnWMqjASU3GATT8VJscO76tqBiEVQ8ESv77SF7cLcZaWGU3cXlX
KgccgcVfmiLTtjATIbpixYpeThi9kVf5ZEwdFWrr8LujVQu8BulCXyQ4KLSTalZ1dRXLTZIPLO1A
HjwatCnCvNMSS0E9RKPtBww+no4a2rkZNw8dHewvlBUYgmeCiK1tCTDO5vRn9ujmYFJqJOnhf+kE
rNRC6okziVfr4kgM2GIMTLPLkU8CfPna5299O27zwmARRm01IXqPh+izoxvcvM5g7utCfQxeU9ae
xrYRLnEogFnYM/G9BMRnNvc4y5pM7YL5wBlpmZGVDW9HgrIsLWMgoKKEDkHofclSAMVEH+61IwQ1
BUS80DMMZEjx4lmbAGbGLcEC1Oj0vlPMqJ4nn8jHyeNIbPt219wmWSvtvW1EnSEOOiQwucNgcneL
QprH3ix5HPQz0kpfMMMY82RExNRwb3sCb7UvDHsnSwqsQE0ENTp1GimAqH5aEc4FS8rcDdXzzvGK
9ZyPYjQ1Habzpn5QWoaMhRG73cQ7J5VgsLm5nxmA1fj+MSpCneCkieZgwy+TNy3cKtGltwX53U59
JhP12+bv/czvaXmG5d0CnCzkGhQipoFD6xMTbz3jczov5LlCbArF9NrA3Cw5QaY4COPFStv6QYCS
scHsr9Pgueu6hOk91iOPtbo9pG8wtRjnFh6S0ydAB7+6zVzw/Nzm1aWkKdYqjgMReW+wSFaE0DUm
nRD0uKy/b+ZuuZ+/XxB2HwiVWgNYCGu4nQGHoI7gOv8LhLMu5mQOvi+gx3pM+xMiceSUcsXObC57
idVKLXgODu4RTE2f/I/It/5YRQsWGgpV5iMlM8sq7xvwl72QMp2rlb5fp2XWoiG9jh+MiUj2ddAX
EkNsa36SsOMHzbY3Se6gZo+2+kfMJTFvvJk7OVDJS0oTosDBvgWbHwzto5QHh/2M6Qz6ShkePjdL
aD+S6aJGGvq6gPX7dOtCV2ucGJRRdBcfhGw1NKavDl+ggnyCvhh4Q8OpK7lHT2ktyhuoEt/aFH2Y
J66Scm4Od0ZZNo5i55DwsYKeMFUNFdVmEyPo/BZRdyGNesgn7fdNu5RvrBSkO7kZngpn0Oh4vAYY
meNU9T7XaEUu19IDdNUiqtJYakg5F0C9FHBSKNf4SyD72crEB3yBKOUZAyar4FFBJCStaFCnuueP
0l0TUWsZCjqndm6adnvptr8fwaxed669v3BqxTX1iDw59IMe3YCswgBJCbmtrxdicSJxNXv4oYFV
a64m6ERCNT7UirU2G1OANHHBy+kxUPp4/Ekimjdd7qwQImP+xcGihpitoBEqBvE29fU74jhIa5Mu
w5G2G7z/o0auKvwRGcInTKJjP7JMoVKgua4wEeNU3h6A5hjJj5SV2P/qn0UtzG8pjCmIKemRUO59
yEyR7TXp5lUHkwTwqefPlLlMk3UY/xJVrd0hyubW6Xb4URk68v589IqVSzYykNuzVfRGAgpsJYMJ
WW+2y/5JGkYo9qkvloNZouTFYFLLo60uQz4Igc4NsjxXTRJVDKGUljE2qaAxKh5Aw9uCo+8LPpjv
k3YBGGyn5yemJ6ISVk7P0Xohg0gTig43FzBi8GvKCKtI2H9qNQ31qqvsH8YmiLR8IJwjJ0tXYNbb
djI6lhauhGT7ZnIZtlgf9zs6lbsfiTV9F4ti0ssIMv2TQmPlCnbn8RYuhn854Dw88xNPGrReUZ1I
APCmuW/7PmNkr1laCPgVFSKk5uPFdVvif0Z7ETfr34lbkd3PHNYmQ+1U7lY74D9tVySSfosTZBpk
IJ5maWU6oSyJjZ9gRXDu2nVGpFlmq/5sYQ7ybYeYa7ORxLXJa/xFtC3oj2P+eoNS7XrIcb/f30dG
4TmrOn0SnvFCWd8wjHhHWtFja8pNuzaoyY1+dNY120+NUUDptGWphLg87xfUtcg0jWURSbP5bBkQ
mGNDH9w6B6g8ehIlfQaeq0efjPVDMbWdt05uzoOxjGY6t+vl2wjba0RxO+08JZ/BarUtC6vaz+52
dKNwp5jW4MrOZ6gmFDKpRRBlugdIC6ixc+8c4OaDyaSn3NGlRhMZVhLiDpiDk1SZMMDyxgZyv20t
WVz4P9UTe9GdqnZizpg2ofx+Z+u8/HLLzRSx6BdRpFHGSsmQ7Y8b5qCtAqqcLAYBHabEacH1580U
B8lx0qc8xgBfOV00UKXTOv8PjCzp7T0BCPz6QtZAZxfUOmMf7iiZXihg7Pa1jYfn8cZQd/+xiBs1
ZPLR7KnzShRYXxwjzyAXA2+Uq8PeSSAn7+RxOPIfvFyJ9n6E+TPrKrNwwSkhYwl4Zz5JqJLFyv2p
sR+dHQ+13gwpMP28UT/TItHt9QfgKvODHe+7Rafs2SRiPhY+BFuhZEw5eHy+HOW4m7Vz6E6ziZuA
aCcpoHtQ99YnqsqMn1zfIYneb5OHD3bWTU3uqUAhpZoGGlWSU11z5bJZuzslq0tjzBBEAcn8fgY+
xisWwyHH10xu8U2MZGT3y9XWfeiwjwsciw4ZRFImF9yHAltyKVf8hxCS4YhbxVKOowUZ1fFuySth
84oxMwrELDAV+GdXY6htebZvZdDjjaYRKcO/Ud4RzMEigMQwKNq9GCEvFql5mOSW8/NS1SzkNj4u
2oDcANjkkUFSSF4KU6EKnbnxxbND8kEjRQr3Gxv5251OLD/d7uszB/a8Q38NVy4lmog3wtTxgvZ6
s2LAZqg51pE8sMODdYH/IGu38iSY/bvUfDpSv+MptkZjm3PPwUbzm7Kq31Xey/qeeyS1WlmVBsXk
eTMYzH+q1KNPUm4R25GVJ3airTS44X1Ss93nVKTtc/139qfmLfYL/boNe76FSqEMW8spyKPH0e9D
qBK+GFYg2HitADH5+ATg9Wt7TbukkT7fcJgXdBvfDKu+TK2OYo/The1ZEmA2GAMC9Pm/BGNExbCC
cEdVbJOtwOxuy/Sfs5c34Mp5wg5cvQeDnUGmmtl+g8OlczCDUNItd6UpSfRTwE6f7l9rRpnAUGOg
fDSezwAq3QX1mac7AsA2QamW1FBDUr/tfD4jb+r+wI4GRPfq4JGgY1Tr0g8wToqPsGafvj2xsgSs
lmiS6f0hdF+CAafEyTI03Jzem3iwYjZIY7yFWA18sFBRl+rtkwPp+qRMbHjwRuagVqT3OQ3GO9vd
YvQf9uBtSKFoMraHYIX7QD7Ib5w+tYeAZUR7Y0cLHsiPxvAtmmW9/zpYl8BIR9ujQ01zc/h7iWYd
oXPjFH9oTkaT/WFzpHbz3ejuPLQXtZNqt+nhDtQ+0MQqpEE0jQVf8hyZI+bc0f3qCtZ/4VK/qIrY
EZbJAbx4yZwmnZjq8dm4UXqfMWMuK8j0q93yh4zQlGOT094Ks6g/0rCLyJuNKnFroV6uv7v3wbvK
/JDOkFo75WEnX0gLAJ6zLIir8aX05SsbjJrcode4xrme2Pn+k+2eoObTNoU1CSzyxtPlSPuaN61w
o00Uy8Gmr6MoaU17EYdEVuZKpQ1/TzDkGKNqfAx8BoRnUzgyQkMSoiY7QMzI8ySwqc0VEfjtx8DK
OdtemSspYCcJ4iLW3/YFDP3bE6B0ykpYWmM1yp5PB/YC5zWD+vNiE3eSkW8mbpFRhsR+61X78qJr
PgC6mpNzPmgjtYmtSo+YcayjDcX7G+JC7qrXM5BfymYLN/wcX2RmlxKaGRwxSS9iDfcl3P3tgQCj
Z4p/7Dw5mw20UYWFx4HS5DiUi3R9H19miPz/vzEiDC1JliRHPO3+BORQT3hAWuJgV/id/cimm5TH
Vk+QuaYp4enx2hYqbAi/oxn4aOhfhiRZRkb16DHWV4CTydgbgJwE4RtfL9CuQYd4qkjI8LslIw9e
4i1oeOcTfi9zaIMPp0F9YaIy4VIA8fB5hvbPHUdN3w1xV6I+j4+mtmjpYyuJcufsIx9xnUjDo0mN
R1NUfST4nSWbMoshbhQyoM0apUm65gS3Lui7oFqi5U0iDUugy5BQ8cSSWtMC5ZqceQrFDdPSOfXK
sG8AE54RQAZ0KTp0v3dIhpM/vncoikdVkQaNofbfsOpqxZIyj9F6UjNB/ZukRx6QJtaycR6oPcJU
y3V81CRHcVjO5A6L6//6evMd2jOLykFS5Zii8/dYx5Qc9ZisGPndVL9k0DEWapaq/AxTfCDC1e1c
2PxLEu3LzGvtiT71JmWsH2iNxr0acbHYy00ekuelRo/kEM1mkjHgLG2u0OJIWMoUo1TgXJK0xVmf
BC2GLLX1Nb1GGYeh78myDcBdgw2A70ZZpWofazok1QbJbwmGihrRHkZ6Kn2zYbxIe1vXXXwP9NCG
01QNHeq9aUIiFoliyrXFFGqeUF5kXsSFYvUtpddtXUlkJBX3YCuhxifFHUMLlReaA7CuuR+/pkIe
c6dsaYTrEU9ISuDleLeLQJoUkgvr4e9HPHPbyoiY0TfPCzJVGZ2S4/7d2ZVK8ZvrdPuZbEaLv0+N
z9ChhB8XrV6XYjwkrmcZ94djt1oJ8USxLoys0rpBTS4cJt17JryAZBy5NQ2d/FvChPvXFY6SI1Dy
7JM+vvMQhmTjZH6dk6aHPGrkAX1b80pXunqezbZAK0d7lz8ZT9ls+TV2ky2J4qU6vK+WPEow6wdg
WZSFxuZGmmSfghcalryr9xseiywf8UKxhuj00EJBkO5+lmR53bWIA4Kvft4J7+O5gB9crXsE0Ndn
LYuuJAnXeFHvJL3Z3PQHE/nV6Ixa8sNPVaCaDohoK8yvHHlWaITVNBJ5y7Gb9CFmi/Je0EW6uqpM
BvC0YAieWVowD/Og/JIj60uH9ZJvFDwaxz8KNaSYM2oRL7hxWPNH+3cGkChd2CVafSrB6sCavfa4
Lmo8JdLPZ5W3xQbwpxs2XpaxhrgnxlwtOaJ6W4JpwLaGLMCOp7LmAzGSCq5rlZkIU9zEaUflvajW
PyqiT7ppAkwxf6bbQqQtzHZh72nsSU5CMsjt8AyPr/IPHWrMbg38E2V0Q2VuncGy8/yYuV3N1pgI
Bn4ftrdgc05HDoXvSfntDa8DVVoBdo/9PJuyuJLeQLJA5Goon5O6gxh5JpkWkbSH3Y3td8zrypW+
HM/QAfcycmhVDCfJQNwkX5AGbyE51Dq/SiHExIqDpkpctzUr0U1wygzw0wIYkTONOocfDPFD7f9p
0V+qYjAFOC36OlDNUAltnKdNAPJMTO5YknAqanSmrPTIi+UXactOb/Y/Grj8aPdO92J4GsqLP+jc
9jEaCr6F9CUbvoIkerV6atRdqgCVysMdccufgWxcyo+knVcGNfMpYt+DyXtubLTNCt8dUPjjLkkR
COUJzIAReJXgKp/MNlSSXsebB2kxQshQpMuyITwLUdDASsb51AGU8EHcaL34LNn994F9Vrqrmt1V
y9A4B43J4kbDFOxxPqJWdCE7ES7W9TklWZIrBg5VOhRPeiZ24jLlLFJlh7buDH22eMXAb5By9Tes
ujFS9fJtP60GXj82Em/AHCEPfa2rQQuYhjwl8bzakbnViX6DgSvFnKKBmAM+k9c/u5z+X4i4Nm+H
U54JWhsl0GPmjBp7rYitzfcVAcxaElLIX602SDEw4SjrtfcTKoXMKokzfDw435VZFzrkx7Rl2D8r
pQi/fV+C/6wffUXrPnKVceTomYSY/xmk/KpN5oKqPz2PksL3io/uyhrnt9z66b+/X2VOL9rllafa
QU3p+Hkvn3amX89hsVBEGgaZGxybieATwHyIaJeJ1m5tFjsnN5/nHpwEUlOjjq1ZDJSnnd+gCuDB
xGXk+b6ab+rhGFrvp4u+TiBv859D3HZ15CtMLeIhhdTb8Q4y3T3IcbY+FaPGrORsyUyZkQrnOn10
ZUIZJMm0BMI3ubo8Hw7WxiyvMsKyFOlJragsuorAajh7oOo43SlFhriRDFt8SuPBoQji8sPc5kof
xtsgF6utjFJfilIARw2Dv52WbnBj0GiDV6XZ8mkLDWFrolazJiEvr/mb/TrZjzpI4773mqg/JZCq
D4vG9vvPtTyzGjKuaQEgh6c9kQiSTG54b6O8ynpnV3GdVyzLn+sKDsHLsd5jRL7j5gN+GepNqp7b
S8EG0A16fNg2zuIefAjH7Hk5C1i8Zc7U06y5dccE1ufSzqVdZyJqhGyclhZz1+Q1//tGS0p1ICv6
l/BAEAm8PFO/ebVTTlLFCoauXra8fMHpl/LwPnQAAh44Jnj63DkhxhZDUO1Xw8gpZ3ZnJbmlCDMm
Nl2RFvK7pkPshtzIQ5MF2ilsHp5jIL+hjg8SUyvh85WMnBNOpuNTfs43lRZ7BExtFIhMj4xl9pDk
qcAcVNEDoQ20eVc8FjtBHw9yzcsaUoNhIVQWaTgHyAp0yTCbiQwyVX9XVL+nqM8ck5gKT7+fWc1S
dGY/vm8JQ0UVdrnWf7WY/h1FAA1sLfGR4XjSkSsWuOS6RO/3E2S7FjQ/iqqw8FWx54ro9FRZU8LR
0RMpcf5sDFTTz0y5AG/NHXWzPeNgs1PDwqJukN7TMZ+N8Qz3zKlu32xr333cDACmyoxzq5RJpTKQ
tjbHXaQym6dL8FIVtla23U03i6/Is+l7an2fiNVa/0IDDyQwpq5DT7b3doBVIlDIP/Li//9YHbNs
tZuVQRvfZ4cNEVDz9kiBWklTLkrSSU2WV7yZ4a+Y6IDMV4HvMwgZH8kbL2OHV+3dBeXHq4nzUF28
nBlsZpqe32jYjvoTTS2geLVYj1P5bAGSVDLtsm7tbbVv4eSGInneA+GW9Yruen4IKKEPrUyTUPEW
73A0uSdtW3Xm5kHd61bFfToyWZLPtlH0B4nYdBeungo5TM8AhzkL9KYxmRUr8nCptkiyMevrEG3o
ABT6RbUgn8xHjgtU05DHNr8wo0KZaigxk6JpWIxhTv02ZSqRET/N9CA8PSb7CtsOIKXFdfMTCu/J
OwvBbEsxRjJ+/SGYXRs4w34z0SkfuI2UCxptKaGdUexkCYURSbhUGYOZn+bS1Ypkvri+JOu40lyD
VzB5TnjEXe8r6IwK2+8QhChnNCWHVnVrKQ9ScZ+5RYYXWAYmCqgj0Yx50d82aqetm99kW7/6vozH
2K+S/BLJ8P5zWgO+aHtpwLmYQCYFsE4aIJyKm2vVpVn68UYdYzDDt798lzHOkpBxo7AEKnUMSJ0W
XD4G24N3F7KcfkLBhC0+sYrBVscwgZ6QghL4d9NWl6ngUzlZKNZV52syVlzhTdI4NeecqDmaZcHM
/stp5pCgxHffCajzzVEZUtfaiNiYPcg2VJIk0HMXOS/K467hZBQN4Bm13O9mbEfx6bxyRARQNPrz
j3zAK0iU7RI4CkgTj4NOZzuUhX/f19FhLXbAj1a0AWEosB11McCqAMOUlDDySXFxR00mwT5SpXGP
QVUF3Vo4tn5VDYmApZAwL+ncaH318iU3yGh5+XM9xCXqV2Q+O49J+phKwHhgIQwEXkVpWli17+6X
lUY4z0TQ7vpPdqsX3NJudL3lG8+rdxx7t0G3vFsZe4NMyWd9OrzPSVu9o/Bfh/czNDmIbRHFDJy/
h6Dh6LIVa2subTgsmMCq/GFZ5LWcZOSMchIkyBWVy+Qxl2pSl+45SnAaNhdGFEOpnmDSPEx+1K3p
h1vfWq6zxE+vV8kwo0sZcfIL9z5o09sGp3KxURvBg91LxkvP93sLPTW4/eTrldkqWD3CMQxPZ86I
ieAppKqjFcPQ3HH5ext5rmOsPRWnFiJbqIt/AEG2Ow0s/k/S6Wbh8HKM3y+yEKFBkJN1hl7YuM45
fVWQfVB7bxzCzig/wM3jaZH2D6qw7MIMtheAMVyzRvBJDdYDIcVu7+qqcRUUzqyt5324JRX48Vbc
4JfdHqJGeoG5NKFia2bWABgcNGE4esJUl0rMV2K8WKvSTywa3X3ZgQ+1BpNIcCA27pSHvCc5LUn1
6ovUjuwcIypipa9soFkTTnr7AHq9ApIboYeYQPN5RSjBCvyRKbdjlNy3tkYnXzPh562Hx/DD8fHj
I3FyWNMl2OL/sp8l5TmTXbJUvZDKYGmLy4DJvxdBMHr/LEBQQa6YylSoK8K7e0or3zfB6Sd27QNN
IB54LPcslnSmmSo+FcdpjOh7//bPI6/b0EoPPvyMPKZjuPPuYRAHnKIZeW1y3WZ3+VnjwWggA9LA
OgVOjeCvCasKl74KiQmpT+Ogwo8pFeoZawgSrDJaWRHb1qDTxUbjomMImiu5nn7zY2+Z7xdEK6Tk
8C1w3Fi2hA+M0ILo51gUO5vUJ4bq3ncBHnOcQRaHF3myGO2lR1JZ5EcMRAoXDBuJy3FrqyGkttcb
hw5oSIIdu2vSex8O65MldqKgPAJ+bnCI0OyJlQtSv+PC9CTZI95hP+xpR/nknr1Qjtk3SCGVh7pH
mwcB1NGsElO1xXarh49d+CwvGg0Yjnr68cDi9nO9j62r3xWIkmnsPyEXdGXqnGkZC1SqKQUGLDrU
/hp4ssEkr/glieRFqBfEjbJsA5DnTsCjMb4bHx0BRqZpMwPYA7AI31KQMDnjookW2d3/f+AP4DTx
9OhfK50Fs2XmF16/3CKAFGRix0GAhc3zE7AavbSYRrSVVhVhhWqIBj2bcnQcU+H1krL/+H1QDnyu
Ej7ctwGxeOpGX4WKlDrJM2b5tBTGQUrhFVPOAMEam1Pq84qcZ7LRK4zA/hb0ByZlWOLoYvgV0wS/
X8gzm6X82UCex5BCGGzW4835XMz86PogQn4AX/oopl7XUczE0kpi47U5yZCABGTWy69T2YgQJtna
8WzTnwUdJUs14V5MLtKlQ3VNlrem4fQSf7aeDLBiTy/poMTo+QR0gQMbeLlz/QV/ZFg6hySEmHF9
82s9AQjS6M7kThg2zs3Z7/E+qnCOAOMriI6PWcDxhOBpiF/gWCSHUe6G4IEr0m/nViL7Vz/N8nnD
7V0PT9r9pjYZXBttVYbz4rHdzER+7yL0iLobh3OIfJho4Q0t1t+Lo34dYDolm3H4Rn/0KqV9CoxP
Ewsg0DqUE1xEuCMiv8C098zRNUmXGXXNSjiCHLawzqSZn2016x2azMovzhCg7vKaK98FMuqTJwff
1IP65A0y+ZdFFOpBircUvOGTyoitjUcZ+QNEH5IxymLwJFuXRXDuOMlyuzpDAFhl9J5B6YZO4AyX
DL4oiKHhFwhSVR51WkxcQxXsaVrJn6mjbTC5MOvi+WIiM0A1ZFnVN9XIs5zE7FwIuMkkrTKtNhpy
wPUUOydE3mMU6jDwlhEegtcXJpuUEW7FjKHUzJC2GX1VKp+FhIRsvyoUqDtwtPs6dLNpWPsCDGS6
MvnfoYujg3lZcpfPk//w5bc9NFyRmC2wX4TJQglhDQwIjYH9sH+9w7raNrqPWjJUunBlKdzk6bVQ
K1Fj3ixi9TIZIODDhoSYJD3sKfLNc/yPfEV1Gocl4KUX4bJci9aRm3PMAAfWUXhG27rxxiIc8Cz5
GofqZweu14hw4/KIq7MNCvkRFdrNXyA9wk1/+ew4ixB14Jzqh0mMxbpiJumAClWqiRyayDWX4lXw
KI00ZUJo8Y5l8LCyrK0zmzqFZ2QxKhHT/4VkPTlDMA/f6xEQ8XCyDRJsx+k6segru0fL01VhlxWW
Ty9RU+3iYQpQJoCKYUbNCY9v/1tvGe30w5nxlh17fzMJJyhG33jYG4vSgldaa4OIJMMKvMGJJ6w3
sFlquhYt0N7Os97G2+PyAH2oz4QypBylPGCychNqI204jSgWH8FLIrdbx8uaOygGAXtpG2BU3s57
F1uqF9/RuneeWCgsJrI2ZE5UCNsJUP1cGpDcpznWjQ/FZEMCQTpET+WdAGr9duP45rDNfvCimEL/
iIuCcW1Ghp5TY5SwvAXFZQV5XpSHddp9etIvR+Vfmolg9CPWYg5lYBILD049cmLxrW0CnQieyATQ
PeBhzsJ1hOKa1I3WhE/BmyZX2EDSqF2eS/5Y5Kux6bbnJKJYUyVghiYgXzcbiPX9jjnkF85LDvVB
fPMrrYkjqbB1DFIubhP6zfT0it3Enrc0GttKdU7X6KY+B47+uivtQp3f6CNManC4tqvHxc6mNZ+V
Suc4x3XvszyXkHjOKKMQRn1GWXC1O3Hg72UQGYEPryF++UPteO1CVfkeW4BnCBuCz8d+hbvIojd2
2w15SwMiiHNT+qZgQP+QXtgrP7nHy0nrOhmfG1NBLm7vb9C3D69frJx8IKNTKZXlh+h9xlX22NAa
f0tKaSzXssQXAFLn98trOBlnPa9SDybWi2jyQnoigz17jAsxl+yv7MZqWYdagH7nxpN00xZPin1Q
N5lZT/LNcgsXvUTS1YNSGk+QkfxwPdWODooATm2priBYFNImyzRJpL7ZX2zAsmCNh1oVXOJFD8hu
fW/p/UtXls3Ra3IkPRIq68Gy9Sqx6Sny54KjFiOEqoaHxiSpObhg7ujXO4iMTmiw+wAeQGB0tefO
ZrqthtHKGKMAGtnxK97sLdSWzzDKFcBM82j8a4Oi/LfiOhn3Odqff1k0tHdiThDSsUZLmQsDCDwt
FvYpW6hyJZOVKk+HFspJWmAPkIEL7dHe6bJSVotfaRLYdUwJXUmrZcfesQqdzMnI7MA8jfzTc4Ys
8vDi+s/9nU0g12O3pjUecQJmMUbO2oCKUUsniSlrBxuTmhBe7bSK1jlLxAlHrQbEkfYdRyisIewE
WwdHJf1m1toK58Q+Ff70sKxaeiaKTuKKIvH8IhFglEHCla8g+ksyH6d0n0ZSxm/feRYgJlv0z0zC
K5PPYVgNivdt1T8ipC5FCIe8rZCnuLAZCPSwcZefjZx3+XCSWlJd6oMwc1Rq09ONRFBpECqLpXiL
cTtsHNmQsz1TrjAr94i0Lae+uP/3t7Y/Eyq/Qskae4MZKSInHmqs86v8YRbaBIxkCv5ovQL89MWC
A9tKw5VWso32LRpuU3ZbagZgL63qXEJgmgMbjtsMFo9EA1caH+TuqSVipJwRAWtrCXBNDiJ7z9xE
YhWGAO2ayjC4cibPwIwywHOVUNFjtF6mnWpzsiBnm7MstGQdVGEbdKWZYC5HCvs7HuOXo7b8CFhz
ICbRnzdUnaSYq4n1ffNXzEKv0kVfHkQ4TXgfYIT8cVX0qscd+gOqP96RW0mVrYgBPttmeEgIBuxP
bIluYX+TVzwRz4Fdt5hYjoKH/xdDuKoi/MtjNNo+W3q4AIYjoBdu6FDLfVbffFo0HziMsnk+5Sff
yhSPEhQ8Rc7vUCIfhk9qW7tZ3ZjRKKRpzuYHO4yR0O1GalhVLxBgTGvxLK7BYgNRCbuLAA5D01AN
QNF3mrG/PKCHbYljk+bCRAtm/nkW087hzfroGitm5Tja72MSa5mCDHkuanHuY5X2wCkp5izi4CvG
1iqUnXJ68dwiI9BdLTNQonT1Uw23SM5W+/8WpGklbS6fvBFcoEsudt07rW0WA3gt65Yh+h9O17hN
JhES8BJz0WUJZFKjLbK8zIZUihsRgXEO8mmZB6fImlniWXpDq6pwKSSkv//wpqleZ2c8ipKBA99I
0W3rp7ndu0vRKE5Rq/r4qYzYR3UoxwuUxjlEqIwFm0bkuzQkF/Dfic9iqeHNlKGp+astXkJ0bzdl
JjdzV0P8hKOCemlwtJ3Tu6MK7jvlApqyS7GogfQ2BEzwFzm4vp4XRGvHIb4Upcr+DDbF5GDFuT+u
e/iioK07IC8YQL3ZFWXFY89r7Uq7HHrTfRn4sRxWe+RoxsZr/olIzY5iD5PJDDouKq0gCizhJpaR
THs6nggiFKUc8a9wDz2bM7zfTsae7SvzINJaHvq+5DbhMRad/4q7Dg7zjRvgoHOjIjPUcXyV5JxH
Z1g2CCfTrkXTneEeBs5wQF/OGMOgKPx9gf3l3eIzFVtt9ou4ReSshzd4E9W9McC0MKRU2sgSBllu
eUakYSrJqFPEeLs+NIXLumeJnoYs+CYUy6gnQNYvPSIOghLsvM+fOISyTYoWn8KkM0Kdj4SicfgV
pjxY6GcUz4tmiL/IM02uxrKuVyEhEljALPX+oS3C3MJ2XXiSkV7XsauQb00vj3sNDbgA7SNYI71K
VTcZhHj0EPAFWmph3cMkYHko1CYerwvklEP6F4LzcR0dEKyGphxGuJ1mRyZi9m7oFrflVNVoz9iD
YtVeTXw867YLwRqhwKNMZU7bY4+qAvd9RTYWhZLL7LRuNplZwr6hZB5I0dvxKwHt0tE32P3pAnMs
73XIgSqp49LngO1Y8qbsvkoK/aPqkV7Y5QS3BnIhDbXOOE+F7NVyubs0YjYONZDwAJ1KzdSI7XFn
0Mjb9oUesWKy1m/p45tnyYZ47jmugJ4dqMb7C/glSuc4YSvHD0e4ZGO7cjaz6+Z1WBDqY4/tM/kE
V+GmEUl6DsvTXNp1I3YsyE8RDqiYeCBxg8bslTLSUyd72Ie/s7U2p33tPBe+2RrnB8DLdhgpWgGN
jWSGGQhHtOBh16tdS83qp/cu0lLhNC/X5NFKlJAhT/UAU37l/9Ob3TMh5/ioJU4dDNAOCOm+wOTd
7yadPpbPzDOc8vCQ3uXiNEpWNPF/F3qdDUu5LSMjTtSVKaaVES1sKJRdJ37P16U3RbKiuIqP4fov
xk08SCLxJ5tzJVJy6/4u3J55q4JhirSGpq+fNZfpaWVY+yprzrjaw/WdfsHCegD3RPWW9lYMRN3z
rXJZKENyWK1bdUU7hW0a23KAqr0u7e1Hx4e4gjy8KwpBJmCtR/oxi0ZI5WU3Nls7l2vmm6dPdZg0
/XRXX0lxc7Kjnz94mQxgWNojBj5nFb+KMo4mZNeOscjF+sUQHstoPgfw9MtzPJrRJ23KAE1Hp9JT
NdQiW8nqPMvNnPBc2kNGCMbnOUpdeONDapTfd7UBon45rXabhdoVLuP83TvWMJ4lcEeCR5shuLk8
KIZNM4pCd6prkxkIdvM3OeQqtLtX7hgwZsQXubBCCaW0a711E1kn0E221rJgUkgYySGQcbEV86Yy
5fZRzvtiIcs4pVKyuoFNl75esrhBKafKPWoyz5NerJATY8GNWA+qTJkM6gi143wunvpGMNDZTr+k
1wP6E/zidw5Doc6fKdUr9yWdhAbMMKu3dx05FvTrZT/29tE2NP/FNfLGwwONJkJD4bci6rbbT+Mj
z7un0SbX3DOp/ka5pX9Ir19UQxGhzxD6ApQ7pEajpcB3EPjGKgqJHm92awC9gkQeaiN0cVqstlQv
Nw2PdaS4Rpf995naRgJ6qDpm/fCUL/NcB9qMJeLojPCKvLjVehfMDRCfrcs7LAV31jzNLOT6Fpht
WFRsXS5pGDsZqpXr6P25Z7qkRSWXEondrwEbSOxAxK+hgzHNqQ//YpzQLFIjJUE8EcCg3PIrtuou
09YouWyagB08Krp9kaWjoMhggSPxT+Op75K0babBeFVOXkCirwLpzXFK5Jv7auEwN6ZAKfkywnHf
ObGCZwbCbztoedshCmBh2C4FxErEPv0cXLs5V9nyqAU94+fk7WJ8NK+7EcBph9UH278Kp2J3fhhZ
HHlCybN15JgfgH/uhrqe6DzMNY/zWaoTumzAFSZBUiWe9+6RwAL8w3O9FAZ0d8wSS+vbwe4chgyk
jqw6ViW1fQyqGWQEqs3a4JeKBzVSnF6nIQRs+03yQZvm5muagBfsQZ89AhFxUll2u1wxVjJb5OdC
CIxBQiIFHxZG46R78FLLmue4egiT5ZDVkdrNmLhS8p8nTzkNY07csvLrlUHc5H8wUk9KDSic50wM
s9Dt55xtWhdrzdj6SGRTdPIvdrzjU8wTjVX0bhPyav6//zdwMUFOSBNnEHEhqJj7IdZ+s4l1PWfs
3sHgzpjyPm/bx3zsU+9XQyn3LGANPiCl5/eBWfx6KJFE92bXbZGp59JK3wcTuQjoyIbrJnt27sa7
EeGp8E8hI/Jk8VHpBN93CgPV5H5LYOIjV2XyvNJXRpOkhRLVXORhcU5F3vNQ8EG8Oz5FHtx38zxS
alx8G3H8aQe6ikVSyUMD5ZDa74Fn5EV78P7ET5fzyfU6hAJ5iIZTcl38Dznbp2Hfx6m5JjimsDFu
N7oTE8t2wkXH09cSn/v8nRhagK9EYf+pcyDc6/zQO5sTpXBe3UnuRxXWp8/3bppSHaeIENdK/n5n
p63f5MqcKFfFVo9vgLjlMp1J7kLniFcCNrWXkEqqgVTVempio6rLHpEz5lj2I9xR3M/DGn/aGXp7
PMzUaa7YlvZpYQTcflrnNo37vvSzCtBoTufxRB4NkOe/mRB3vPlnarOZcs09s3qMjX6sFMTbKR3K
q5XnG1e3KyM2jFf88Mg4v3Yqpvg0w7nHAllnoYKcY7pTlB5V2pJHey05tsEmNKHmaNI9Vc22h5Lj
dWfODEnqJTCwx11/HjC6++8d1CnKWRNPfWEoeXP8PZ/b2RFrNk0itN199xqdvbGA/o9ZrVZ3DLTM
kt8MUHSknd16It0JjwCZk1lB7sOeucD3HwBannWEWDMWiEwQPGye9vo6VYe/u7aBz23MQH7wkLos
Ta9HLpJKs6FcjFzl8oJUf6xLSMGv/B1Zos5Ucc13zr4U+vxoYOurU1z3ZT+1SHbDGZzqvR1UFUwg
kk9+6YITLzvrldix3/nK3YtWiWqsMMekH3mAIv3Izf5Zaay1pyRoO4sJY3NvzeJtAkdjX6XEn2xI
GMVle6SsQjTG0Bz9eQpAA2C0WhmGwfhT2GHcnuMEB1q6qktggaXiY11aXJcg9T/ixBQilU2RHA6s
YwSVnIaCOXC5Vio8viLMDk3DQCq0TG4KS9bM9oUOjSCwHH9WPbQntt7maYkEV7P2B7fynm2MzHOk
3wtnYDDyZw4iCyVT421iaqBwaeSH+iG37G73yvisUlsD0qlOAXy4sGBb42+7K5HRHAMLrE6wC3m9
oRlnTxetAD3edCb21A5z1ujageCmsgSoutsQPJl4GF3gtMrHLhXTOGNKv3MxAx9EJISJf5FsbakY
JoZ5CL2c8HoOKrW5ePebRGn3DAH/3YUnwXOka+EJT1iK9WtWcT+ApiZ6OZ840+isZoxu6ESD4VIb
M8F3Sj68ultuewj7DY14asOC6Eiav3T2/ipawCbzR+W3kFxoAxIx/fwQbutfSVRNAg/UnAc8eeFL
WDrVh0+HmBWLKK9lnhP5G2TQPBBCr+ASY8YpGdXsDFylStfEK1fp/5Qsoxi6JRfRQIOZ7mMQwBx6
Dv4vj0kngR5oErxZGUKCfUGzzpAo/CodjCGFMq6U78DerApBv2ck3U3a3T58GwqNc2Mxl2Bcys2A
vpL3F5f+ZXW7axSjCwR2YwDhswrH0YjWQSXGMXpWhIYiOoXfYU3+Rs+xD5ruR6bE01+N1nauDRPo
cYyHBxGlKwb2MRm9FBoLkAg2FxBJF4iYw6C3AmeWyoD7XXZ+c+eKYrMa4TdtDQGog8IGUIPEE4AI
uJ1YKbPydGGATKtS0213XZaMv5morqjuTO3DDh6dcG88TgPH6wav0CFVyDvCvPICiyelW2bBPZG9
0tAuk7maA6tp9yRRq9s1IwVs0aBDGVHn9oOMgKOa4tqL7y5XeyzNB5N3+77fezvVtJk07VicSDoK
MdGb/UlZ2TX1J6e54UcjHHVFLg+gNBM6hEF+eCNPC/o8o+ACcVA+2Oq9MpW1XMv9/yeuTVlDK2gf
CM9+XgWQ01excGdupSmJFT4G2ZpswKvlpL3Dje9jm4Lkkh8Aoi469VuhcoODpr2BP1FzoM7hTgc1
mbn4x5IyvKNjfzmlN8YnmsAvtHUSTIBff6ax0ErO5hOfnmkogHAN//1tcOZOrxXaZ6tyESWjIKjh
JOkUDXg6hMG+OlRQZPYAhaQLLF5satgNZkaAC6XUXmUEVD6Mo+OSKxi2SYhqN3cCIuWxefDEAZD0
3tFI1AV6N5D7F9zgpjqn4GYTENyO8PZTK77U8ZbjM6CjBemvUEPGHIZ8n62F3XSBnI55956KtCLG
bLzIFG4Y7VIxUSvPFku2eeSMV+7f109vaBtLD/TT/a45lIlseXnaTDOU891vKATyHnnwo4vTZWJ8
XQqbWU8d1B1ir+cBfGgxD7L/+PlnxeoXgNVuJScfTDcyghYAWCFKyLxXNi9ozXfM9ynMyalPpQoz
W9nEpOKwoeWvzLHsNfn8D71ziZhDaqkVRRuGDGKjKqn2E+KaFP/fNifXNYfyBlMxu1W7EAL/GGKR
WpvofWChjbZVh5GklXmI4b8uV0esmZQHR2TD3lDT6Ki/q+iRqyA491ebyun/9xwaVNY5sg3erHH7
q6/gNu76vv3PNQ6EIoV5pmk6QAURkdAEQoIJGmg5GiLjzC2EdJ+OxKEEWeAm7CA1KWWBgNaAOZh4
yf/MMoO/griCYSvl6x6r8tdKOxMMHkF8jnYZgDudm4y3DnVzPLpgMEGpDMuKXS9YN4Vpa5gwDG0E
hg75nLoMD+mRoN7A5L0KQEHhcK3EPmgpwEWJlMEr3WD6LfMvx/nxu9yx3ShP9/ZpyuEWGGlR4HnW
IcV/sM3JPmNrmJgmSNv5QFOgGiDl1Zia0FbsFQu0CE5AACfpedSSnQTeWp+RuEdYJX80FUALVYXA
RVBP0aC0czestsyPeYY/cpxAtJtfuxd0a0cxuPck2YW/8dgUcmYF7L5qFRk8yfj08L2XH2YIvtBL
8w5nkid1Etcf4RtctBYG4ICSvEL14prgB+duKGsdopcVc9lBOXPYjEGAR4Ng6YoxdgW33+aCtrBV
jZAZbClvhRfpdIKtAs4r3GPo0l3utGxpgs1iPJOE9Aaqnc19zA3harquKSqevbv30oHwVNHOXUZP
VaKYCvsg4SwAOdHoOS636YljFN/QADB0DxzpnwVLvZkb4fCz0wv+kcH1sjbsW+zFeP85jA8gMvw6
m6SHV4WfxrzAuP+9Lu9oqbIe0eX4w/rMBpPpCSftTnoVepz5aAq5qaMkk+Kbk1mkdiyM/zDktln4
2gW8h2bnxbBOjET69cuEALbw1fW9x+ztGNS7cjw/0AMxzN6hrgfLs9LjGXzCo50p+fJ2rs764mT6
gZoIs9lwQZ7/ASw6j3Nou/8TCYxEOYtVYntVPQD2EfwyQWhtP2RWJjmpt6eY75+HwmXC9Js/ZRIw
fMWcDU6yXjMQzyb1Ex/AxO9XokyAq+9RKnr8jFu1ibrYnlnJdNM9D4piZSCsfW0MPPAinWyyN+Dy
84DbDOLeXaZtjN5Lhub6OlUkCcsk9AEG4Dv/o4Qff4lBsrgfNTWi1E5cilxuPCvbNx/2LASzzxSO
pIGG7R0jCiTW9DXCbM4OxtLGieK58w3CjP4DiC6RQSEa56pUzHMro14Uc67J4PtAwmOHA4US/XF8
uwLE3k3Tt79bd+m8AxXdzYiSpIlj/etuLueQSFwfS/DZwBQmbJOOD+jscYobs4M41vBJmWnsWmii
suphZaj3HJrhZDT5FtU2sq/MV5D2yHSzjP+hKIlMoQePlUx61x8GsMFBQnGphO6pEWrkbVX4tnZ0
q/NuzuqxooXIwpiJtpRN7EcMiI+RpuzS1aYl+LD5Rk0WRtUUV1SRugLP4kZGrtzUKwqadNVrOeHf
WAqKosfZXTXrpRk/9szsBu0BZTzihMupG0P4lYuecvG8mF6LBeur+Fk/gxeOyU2m/4EJmGFpxvDN
0Ad1V8p+HILo2r3T8IrPLlmqF0GDvrR/qRnJzlwaPVBhu5B10BrUzGP1CURmqm/z24CwemfBHHO3
Fcp5wzCGMUrlTa34jsvITwJt2CaKG+NXJFCgmXc+sQzwBBFl8Sv5A3gLs1jyqN6AJuyPPsUR6dK5
x0+i8ZeWdNsJFkqD9NmRh7nPHvmoc9KDvz490+CAdOgQVtV9hD/WptbnATkrTPycUzTbpmWjnlwE
zaHryVFeHtek7upulfaVuhqz8DLWxx1Vrxdk10It+6gFcIiwHmdhnWnO5K+9MRF8y6REF0Uj2X82
7QL8EJwxm55D48fSomv6QVKzIrE8tEDYdTDeZypP61p93ZdgZ4QXhGvZJnx9IIK6b0eQ/jKhMPY8
jLaqslFDX1A+y7xvc9G0linEmX6yEfFUSrd2qh0JsD2oPhnZI6027umqNpvZpp4lEa77YjYpqdXp
uxazIqY9HsC2heTqf9t6Hk/FQLxGCPv9p5Trg3jHgoafJRD9OiUoTmK+ufC+BuoG8OSL/HowOLZa
xAApgdYf5+flUPCZ6Up5CXFcTv0YJR8FbFXUm4T7ut/hibe3ZoxX4ok9+t6jP4QBzrvL4PMyrZij
pS9tBaJHyOQZGq6hj7+qpUNd1K0DrKfU6ImB0koM+bC7QqDXFa1m19uULhvKR5HwrxNramvCTpT4
/P4Dj2D9hF2h+66zzXTU6/mYNOAcKnMUlXtNsdNpcBRAoGquBB0fdvdxuNJyzwve4Pf9GeExHvpn
Fpvmv1BPShXCjSswdNdvcQq8CdfzraD4tRp2CrIh7mRP+HZAyDeFWIN8olrxK7kFctGkYCWy/+kl
YJqwyzMerdhtrMSk1bDgkCGoKh+1ijLQ3Cndw6dN9amJEzxudTVYScRQkxyBOW1hfvxJyIm4QED1
uGU581tKLuP+WB4ZXCEfY1AhYyo9DajnN2PDwnOtEH1Q0IoCYuqP1VRtiTo8XY96ggP0rO78mvkN
qA0QODQUPOeEuZzJxmBnef6D2RdWbVldP/id5WpxajCf8hXUUQAWFcdIHPlS+ptBGMXCbi6oSH6z
rH7Cwf4vwIvi5BLZjG/OV5CasPsFqrwRhx/tQbNHWnhtQ6Fa9oF7uNvvxE24bTdexx5N6x7QkXRl
ooWijF0+tpu6f7jgZkBzaf9pJEP619PvrZpB27FJRL0WLRpFjcGyIlyZkkVj/tH7+CPw1D4bMV33
B0sWB6maRK6lIf01NFaxZT4Zb5ElTyLoLRHDTk3QgoBRd/1t8YePD2wD44LtYEs4m7NSc+qkSzk/
ns/BdZ/zDUHDxYQdxHWXoDXwwpMwlAgW0eAHJfdyFiJsu1s9IdCmuy/vCcoKdE/N7bLE/pygU1sy
DxgWZAY4XiqkLeumfymXw8yLL7joUlzbcTg1iEX++Rfg66QjnRn8JtGuFP4kKvPiawoGHcla5PKq
Yr8K/0zmVIZ11O9/LI/Ys2RLrcH9ste68+3DQsMBOXCyf72LO5/+dbnmLU0zmdmUC0DRN0OssLhV
h1dSfmzAJwA80w1/yLA2DQGmbJ0iYy9gKC9iQqI2QBsidEUWHyx1+heKXmYLD6x5Lddjike4ZcTS
FGP87+YQlDTSuoFYEh9FHGIxwzP8sVeoTfdKJkZAxUT8BFBzZJ/dQWG13kTYj/JVdVdD3aetZXuO
evWBD9fDnN61OeDy30xEBGMXLHiZ8xscIlL2dBScF7bESAyOC/o/0rpdC4mfl7Jqcv0TEPG2Tdy0
4jeXTwuwqpMC1zj1WUiv+TMayJ62nBL2sfmvAMmiPlg6V2oFvKl5P239sIEWt8DTAnJOQugezrND
whE/Yii5hzRSeNIQJXeXCOeZRKiPfNggcPi7A/5aaZgnAtMD9HhRxcDAicj3S4yfVHCIRHTF84RA
rXqiJeedgD3tL7oYl0AVUGNRR/aj3NTTu7eXUPMT6+abiR78NYFjJeaxuck9ZQBDDaaGsWaeS66K
zfO+qsbixxTeWRpW5I6zRKT3wx6O0IOifrKEKTJEnyzJA8t3H07u8Qm5/RKqY1IHtSN45b1axKD4
kHv0m4s0mBrHlJR578gIYOLlLTAc68VIJ+p4r/Ji0CCFzlxPBd6dQllB/r0+6CwGqsXkhoChaXd0
6tGf/MJi6q11LdVe4+dUOtZDmSbzKKFApsG1uZ5DUZ7Tc7HiiV8tcfdiC249DPYpSFRTkUyZ167d
J2b3yDE6v+BJnRvXhHFEhIl5axh0Dilj8FnMmkmIrI8xzw8UV1iRn3BpizNjBYm6kF0b9tSEFl24
sSFSQMHLp23Lipg15+NfGDCqmGUbGUZ2C7d9GECtF2Qbw1zwvzmOHs4W2n+SgLLpgCirWyQgy8Js
fkP1L1VxwvSWwMXq8qjq0az2/aXnjG5CPOL7ObIqktRH8TEcyIJJWDCnVcxVRcUIGL7wODi9FPUF
LcqKBG4Qd9BLQ/Fn3zhd0Q3YhyLesnGklrO7JwyeWo7G0+Th3plt+/PTC4wCoCfWYdMVDlgDqq+x
qNbaHDXuERRv1QmfRThtJ7H0KQxz9R5BCuoevG4JTSUiP6EGwralDtpFyUoovQp/5bzNVahE3Vrw
Ojv6Yfx8MzcoCMWdzW6NwQrq9nsxTgDDWwtppr9h2bBLz5ilwW37ZrHhn7Z8xhV2eR2uNQ2vOXCe
5gcDXCaf77G79Zetj+SDiDZfJXuavckMocJVj/UpzVZ2KrKSyAvBIoiE9cA7p+UxihQb3c4P3axy
1k82SlG6CnnHDxSIqyh+I5pWF5gQQr7P/frPUmdSZDI/fvtwIeGn6OLNldTuVhE3aEl1Jj06hnnH
M1E7EJoXYi6dRz7Crpwfhwj6hjEA+xtLTJjTwLyFN13MVxzrcIoy9iikpX+bHTeGrAS9/oQ+7pQT
2oeRSaUmyRuweJkNFOTM6mu6qhvxGVJIagWjk4LABGYWYXyzqaueDCsJ0VhgBxGDnydue+l008zC
efg0AbqJSI0xD/xj/zklg06e8otUSIB3EfW0hFzf6OXpttoa9d4G6eFa1rSVEfJ5VdT+TZDTQ/K0
14OvlY8Jng6vFkfAZaL0VadcXy4b3ZghVV1IofyL8uTYh8ukNfVupBQhB6ZuCzN9xmgYK78Okg+S
/Plw3Sx1PRk/o7K2aK1CKdY8BFIiirw+9biQ10CPZnSZtZnDigT6D4szYy1MM3d/kx1DPowW1E7p
RtrMbrLiofca7vgGp4ZMXtwTNf7terJJ/lU3TCb+FJOl5dOu+Qw+/SxtIrhXOlcnJ7/yZfXEss9U
/GMMIZuc2CNk6rhc6RwoKXjI2M+NzPQxkdNObmuoz3TsZ4GZScJNMD6aW3KfMAIl3qOylCfvAwik
rYoFP4Gucgkz7Cip6nevHbT7JbZW8pvhovFthUQptSOThDtQFeha0K6HzaYpx1rcc3AnVSRXTvUK
+NpNq04IYMczOzIxk3+DyG6Sva6NTPAm2l/p/PzmoNhl/FIhgfgBdOAgHfmz2PVxJv6H6PGMong5
ka4OGc6eIzVmUU15J+ovF/DEgjRlfC5Rr1QxPxtNK5/dJdagtY2zNSaRGCZYd9m/LBVuMcap2JiU
qxBU1bzF9wZWOsgbI+4m6qnr7sRZc+wu0LT5C6qiqzYTvBtLYUAJK8BlJXJXQisQO5wp54oqIweb
lwoIFarGflfsroq9kEHuHxmmcVUZdzgOLknVYEhMURP9tIViXShErZ3q3x6UrqyoTAw7Yydb07SA
4kqIak6/ULyvWDDDFX0vXmS3jOArZXl8+eLFnscDBh18eMBz/wC8ja08yAOYxHx993Ni6knLD7Xq
L3mIUMbfBD3+jX0DPuKCW2FN9KaZhbOgLW2suC99wMFlVc5zXaZWfYJYAYinZAh5UR3fAmV3nNxG
q4mvg1HryinUPqDrT7ugLBl9MznvYF0FFIZ3LJdiKj0VBi7jvmRkf2oMKAhdtRpNcV2bNtlfLtr7
FV8BJ12YBRf8s56r1ImFyYGU5klDjRJAMo6/IU+dZzSf+nnXwZlATHmMGmI5Wisi0D0C+5EcW4nX
vVw1tUtI0z3v/3mUISr+1fHa7JxS95J9XrEDXOfAoH5M9F9F4x+MJNvwgiLd61sI+DU0E+5Cx2Ca
cjNYwV4b2ts4e5SwPQ/hdz05pZ7C2B5Dv4znZ/016VEQaBpq+JYGNHO4TivJKtjsRAXsqpsDAa2Y
mV5L2mHhR7AHAnoTjWY1uPp1y/9IJJQUwIyN56EwQ18VRht8HaLd+vz3nuSEEp1bZajFnXip1d1R
05JHj1tIFAV3NgCrH57nVw6vghj6jBWZyJUwyoMqK7eldN6vZnJCBVSIVeU/N6drYqsz0srAF06d
x2k2KYQwiArv8W8eJmbMVsrQoCNYY8apA/I5XjEUewW4fF2vCOSlxKVhGMiEJzeihH7fzoXMQYG1
rZJa77LPs65msQhs/CqLlc4K8FkY+1pquzN9ti3Qm7soomTFa5WIGVObJauyE0yWu15ugb6gsYN7
uJmEM28MkYWdNSwg918+u7eXrHcgNjTUI6g+EYxf35EfhPwvmaG1XO7fDFstPCXNDqs3poHSX4eT
JJ/NWpQjQhtnG044oNZpvD+REEeHn+PIWK3Uva/jrInqclwkErYxv0Xo4ycO5hfY07oCKC0RLDY4
rZ/RVAfR78YG6lTOAQMMBaatCQ0KUvA4z+aonrwanuX0VdK6I3ciADYyMlrPfigfCIHSxKd2CVgv
YllGhuQmyg+lXdiUSXb26qMj8e58eXSJSS5jB1qokUoTSs8K4wzQELHFcCLt0a3sY3mTn0dB3fW3
QMEioIpwMRoWg2AY+kDT3h1MAQvStnu4BP/NPvS7q1KuKTfOcayMAQyTf1T80KtXfdW4yU90skys
fVn9OBQfe7xSsrfHBnSyjgx/si/FFwznNCvh0fwy2i/hO7pSJsyc+R/ymGK0JDjzoNPuzaaZWnb1
gCAb9KLunovgO+ab83t17sD2SD20VNNbdUoNn6OY+iP5NPbjMvQHXIaTH4h/KkMfl/9Ie+a7GiPA
Lbn4QZXWGbic9HbKHxyt+lyQN9+AascgB9QNhsk6z5ZLZg9u8f80OUG0MvBnEJ5uZ3pxVlQkZudc
2MQHjbgfrE2iH2umhWS9aBlFFxqJSGz7KXQGLTUQv1uw6KW/WIlzc5QfTMkoNfveQyelGQjN/0mi
oDfGQU9cDRBhgkZgluURSgBvyUHTo0K3nYcwroehhh/8EsWoYQg/elTfd0plxuhmW5WafZktZSq6
LnHZ7iwTOe07RlKENdF62VE8YhrDAzN0gLgn7HplywxmtOB+1cUNRAe6zHqzQLL/KVE103GaKz4z
PkLV5yObSdHHsvU3PW33cyIaeYKavaw78xp2EZ2aGWWdZaH/8QyArSwvqjaPx6aLYNWsDllYFWps
9CgIKaJJLbvmtASYNauAjU+WnIDZ6qxdKvF96FPbHF42aj9HiUT+fWZoxmJRsJD32J+3HIm3rz9r
nMkZMcN2wvyNyJqJZvVckcqfPfQqSAJ99PTrZiDuePrV8xtTLYxM1m6bDtenGppxHLS0L6m80TGs
c1SKk1/fog4S+yaL9Y/ExtnSg2BKyodlfBPI54jjrvkLD0NtSY25UU0PlmUjpZgMXjvxIgudfhMY
qVH/8eVMumh1L65zMpiisXNrTl44RWffm8M3O+oCm9+ZhhGCXFkPpDF8Tbzi+W2HbI9yXp4nUY7J
CPoVgzAKmPaK40rWM/GsQzvforSYtk+WQE/uO7ubq02kh4Aq5+hy8g1Z+2fMwdZZVsIYt2HoyQoS
mJs5e/p/SBtfSTI4GtspeCnZRtUAee9/Nz7/Af4Gt//t7te95o6fy0bkjuEKwlOu5iCZQX/a02PQ
0ZF5YPS2Fd0FT2YKZbqdmxsQqZM+FYD3uE35MRhPJtTt/m5jkQX7HfKPNfwZivew0vYADtLlN86+
qPhSU9VftE84jkr4JkQSkwGFm5UHBa0Y3NnqdJqfYB8VXRgwC0JobBuEJpT2VZvTl/L8nyz+HSWS
Mvwv9435ajfb9pePcNFOto1qfqdrK/+iXVcz8PJD3+be09MLEk3vA1MBeZD8a9fKP+5sww6OhjBu
9aH/p1wM3bTJykZdUccVPvS5u3KqS7mUuNtTy+YBgNSZ5Ss1V2Cu2e0wZDjzMsVuciR8T92PqoBH
/hptp1IDJMJaV464FA1i71+kcNq/uXf7+liTQnOA7LgMtOJQ7tCCjY644Z2LCpG8Ce1kdE88+yFk
uaZ7w4p+t8CWUh0GPo1vJOdaLdUDYW5JfcwJZbKirZs64OcqzZv0a1sV3TjZNASpHBxevU0HUu7o
vQ8nkWbq4bahWJWnR/LkawXm1p+WGNFOZXD9vv2XjzO3d07mq5V5A8+KGRE7T0t+e1K1is4jFxQ5
eqKLuaC83NFncks/hcv4LKSLrPzqJAavzViuAAmS7ldeRzcS9Zr4sDUtmVx0eqinC9zStWCYk/zw
9ekr38VHxyoEsNhc3TlSOB1CumVPkK+iNzTU04cf7qLG2Yv/te7fQebTHZ/L0yf7wHCps82qavtH
s2oQ2flgjyn4324Vzbxznh/03WfUPKoetzrQTXFssM6j0gMcBG2B/mxhPDcrXmV6BiHcNCgCi7Hq
hdlXNMa550uoiD2HzSrhBaT+//V3j2Oo8vGT4fQS3qgZ9oh9XKk9HKhlClVZZMB4e95zJAyJL2si
/7tkRhnfDoPdlbsF4koNQqOQMXfoX0Ng+rluChJv0mrNbeY2GKIX81ks1ZjFUHZ/IyrMvWXmxaL/
iE+6sO9JTZ6pmmPVqXKZ9HMHjp3PUA1roXTLPOeD3hmCb1yv0L7oCsd6KufkTVnVZ2f0AEg9teC6
DlFwJUgv29Ov+Xj+L4I0qWWEETine6m+V44WbmYJfcBLZO5IPXTBfR2Vp51g0dSra7pRJzmZq63y
azqMNKzcEA1cQdPGvriKWpDnK9KhadIyNYIJzNyW57KzSUNMzfIYFlFZ3FxLZRWj8WyAhfnL6PWk
QcaRDAzEJEj1CggWWblSTS4HpN0VaASoLVztV60nkuX0j8pVn1PvMKKcsO/r1w1g66mrMISNdtTO
1RjH8TqXnFvRT2OtA971Tspi7voyaUw1V46Y7ZxKUdIcgDsfF/heZVS+iNd0VXUudeTYfvTz/NbF
iUpnBHIel2lhRo1y+IuCNy+Ble/W+1OPSmf9ADWEi4W6rY1k1R0SdvrVB4m4iGE1jjfh0LY2GFa2
vnZq5JMuCMR3IW24fzQZSzJIagTvJETH2GIqYn5S45VTAyKMO6hC0W1bk/GmbCqlckHKc+272ogn
Ac38w/nGGSJUU6qW7PYge6ftWtYA7lRb+BaCqSyKoO2hzUXow3DsIUmn0rchykqWzYUwo1oTZ8JD
ZRdIGNGRKsR1JaR4b5m875xJNY3dK1gXek9ZCyWT6YNMqSmsz2FlGkncjRdoNaNmbKriC8X40IVv
C9hiiLfAYbDPxRDQQXJrbZdKrYyDrefV8Cr5VZCWbfyskYV/pEb8t/sAAV4wVfRSfEMei4S3N3/8
Cvt7ogkYB8oBT5B7cXcSvCzLBFf9yaluT+vzce1pBUXv16beXG4pi1ekHgVoV+EWiQBFULb/bx3o
fPA+Z3yOrg6KOkVlj4dECMsUFBmSEBLjiz/4SBsdap6/X3icEtqhLUTxtclCpzUz+i/DHPfdBwK8
R9C+7uR4Q8O97XjHkVDa2kujmInW8AspIpdZPP0zpujsgZl3fdElskRfHm2Xx5LTrZOeEmiGk5EC
qMFUlC2/2UWhQ7U5DLlMiBQIeNB4GjA0NRWmLATsDynKmZMsrIbnBNg1r7G4liNHf/UAhN9U5v/S
DjUJXYFInMKjDd0qQZD+gW91+pCGKgNQdePXp3dDrvHuG67Lw/wh7T1s1n0KJrxCTXXs6R14ATt1
CudlF/i1h6VhKnrDi2Q/JKOl1jb847R+LkeMsQC3Zi4+Dfm2x40+uc041EKrR/Pa9g6fqKe2Hd3p
JPpNZudAk87JBZbCkqMsC6ocMzcscThOdY4VYSbE+ocbJ0B2xnlI41B+ohxplIy0OoFr9hw17aIB
uMhqzgcYdRqhXTHDXXGMXj3CU26/1Dkn8hD4g6UWa6uSZlt9XLLPK7FwgWmHePaH796hGBUrff3s
enKkBcG2M13jx5ve21hnZWvJHoiDdluflXYFn5xA7LAAKmeVpIRTjSakvqeKdcfXi29TiyTDuCSi
A/zOFUByw1fHML0TrW5FZrN0zzEEYilmdslUgXEVsMS3C6jBl8sQaXgkwdxTtM4Bn0Uigrl05sPZ
XD0UKW0p9EuYtRih5J28BD/tw6bTBWttugyi8ttWgp3P32780mu6CAYUNkcePu9yPNVVTbruuAps
1d139VnqSCjTCxdjbQ7XqGDTY9p1p+a5bf4jYUcX+Kn6+JNc269uokKmzSyjABtaB1XNZiqd+9Ng
nyDlCCFLEmTX8xrPkEsbOOFdc1Tfzlo9cZrHI2S9t+4EouN2FelrK/gqDMM6IYbUY9CtTTz0rs3a
17R4jdtIfgmKQRf8PmT0rzDgwbwEBk3P1ioYpHDUOiuP70vmXoSJ93mGru3GphzOpTRlIRS3N7ZG
4oppLtSUU2WuFhFxMI9m6X1lduDQ8Gv3RTz4AcDlST9XOgiwQ2waF7jnFJb0m7QbhV+YhirDzdVD
Pn3+rl1Irry1zgtp+rmlIqQX/8QH9v6ucbxMeUx4tWk4soNb6UwGGYIx0+oKWdhQ9VMUhFUGd+es
quvf/xE3BHPnDZbTt49SvXVJ8dhw/pQyjKD47Np1oAcW5lGXFEcbz9kmLQHNcFZ1sl9BIKtEH9B/
XFnnqbOrRDbDyITnXKn40QinXEU5a/FEHWQotWqtBhcmWZ/qti4H506KMGufxNZk6P0uO0WJyL06
ktw7fUEqHp1gYzsz4w5S1JIoRBo0k73oCfQtUtLGFBffPoN18tXzVd4cm/fahNk0sp6/ehF5rPPd
slyoBTI2oYDvYlwfhaW5KZVC1xlt7Pl16lqPKCjp++kVaHJUFcWHLcyrBjFzr2XNx98Ran5lT8Lu
bVA22Ylj8eYQVTpiff2ZSF2vJaa7QNanIfImW57XKLncHtQPQ2hc0tmAbWiYRzxQaNTZqFug68kJ
myfoUSAGug9J+svzPvAoIZj6VMSLYa9y0opEutrdwXpQF5sgHpNMoCKH8Tl1dAh4JuhshydoRvOz
UaRxJ5p03SZ4bRCGK9aBpct8fD/+QRE4+7qr+tV7e6wFOKH32Nq0jCcEAhyBspJovAswEEEp8Dry
7Cxj6Zi7kmAUAZqSK5Agx+LCwsnupHMKeD48xmU3wzohytbrGw6UocDv0AMIdUqQygyNQ5fkyKNt
qs34G5x3QCEIYsN8AUpBcGNfDCiVgYYpiaIwEcowE3X1AxVbT3KllDkQ40QHu1qvpT53Ojq67Ggr
F0bsJjf/2Ueytp5TbPb0U8fdkpWSmQb8IzRsdr8AYTu3TGyZit2AiaAjW4vqOyIksBWoUmcRQ0An
+M4bLR3dF1n+RbPifak2hQTfkheKUDFkjCOejH8BxAfMwoAfPUElolAFFM47s/i2yB9C0xu6cRdn
xYg8YOC95H1YrWAMI/Js6tBbnT20q4S4QCRYN/idugtH4keAMqbygWw6mJAoIlluTIXPMcCK3HCH
qOINX8hJCR8KE+m1EKER9zVIPio/YPPcdlpcCbm5buJ65/7Hl9XzBrC+0pqy+2/jNDBN8p9VxZzP
S/DVgMjckRlFIhnZYoOq1Y0kQeA/VaTHkZ3scHq6m2RQfvVvusz1jnlD/kcxepeH06JLhBCLla3b
o0uyiQPem/K0vk9HQS7d4VXEnG8jeTLBu1ou37DcQD+fvYlGnsslL/r1sXFmjb2Zm02IFjyd3XaG
BQOq3/UHOp7EZfwbjIwk9K06lZuqcZ7r0v5YYQRprPDDCYgoXqy8KAw1Jugt6rKyBOQTm57iH3aD
nbO34XhCAR2SWJjmcGL4gyS+7YXOn7aoOFklH5rBa8Wf2e5rEcWal21a8GK76C6hy0ydtKiKq6j/
wu1T1lD2oMTdouWkhi1+XyLWGJPvHLXURpJR6S+wHt3vaqbrWi5DGzJkQFjX87/pLO9UUcu6q6lM
Y47mOPWbcor49Fs3Ker1JmGbDuRdawJxo4V9mMzOPaJK3kn026zAwSdkd7VkBtFJmNhSkZKHrl+X
sKO2fCmew+JXUTlX2tuyFG+G61/4uiPCdyMy1Mda7XMI/GsD/BLl6+HLClpA8OvX56Vtxw24qujz
f8+5tedwmsYQ4BGgtPlPjux9h8pYxBWMyoPGHEDxzUqlu2ZiLFR3I34WPAU8sR9hWm6xyzNJQFzI
wpNLS2gS9Db7SghRYOP8y7pw6xlQHHJwVd2jQ6edl4h6Qgb1yyd9BCa7MPRmkWFBv7tbA3f8lzlc
uUewyhM/UElm1QS54dGx9LbiXUiQy6AYBJHkwUUPtbXENd1mh/0UI9kuAYLY82jW279x2BqhvW6l
YahQBFpX6bH4PfIrc1ss7mlLrVedDldmlXup512cowN9CH+16jzhoQR80udPDMYpPK+4zOG+PkZ5
A2No6mhrP+Kk9lUuJCLibcdsLfmNZ8J1YVcX+R4O2a59l6fK9aMN44t4VEj7/qduhV7IRAvoYFgl
CsJe2xpnb/dCXDFVw+hU1Ohn4S6B1Jimg00UPCKWe/Xu4e/o8gCwXc9RQeACTVj8HP3Fa1IFLXjR
1x7XGb7F3vdXNYJGRHPDXoDDoE8xyL/0nn8J389ARZpnp4pMrdJds/iCw/RS/xuMJlFpmU0K9qGi
3WWWuTGW3t8+im9WnYNQNKjYeXiaNRBcS6KDwUXM6pEDnkvxSAcRKFzLUmzmkwxp1X0BoIM+VIYl
zFsMy24IRKAMYWqeihbrk8h5Z/WwqrOPTXySZbNx7KLFxPXXKMtn/seXB8C1at5I1JzzGBAOF+8L
kiGGq/KbMZMQsXcHwFEkmx2IIWty0mYyRNFgqwhrTlSomu+oNGrhEbdwR15C/1Cdk6c51oUEaCnw
ny3dUJaZ33VulEd+co9nc5Rm6FKX7TW7PNQmoLYGJWJONw9kdJd8Pp7IX5dn5uyL8bTIBgdGinaR
mTUarAjBx77uDX8Uc5SMltdMlpzqo1dIivBHwvtuPCNlrImShN8mlNhP/STA37fvbM0v5LLRLhNv
uLY+RrX3P9w7bNauTzVqzR7h9VJSTUPGEq0q2r/Qc16HVAhU/EgjgZ9zqD6nDkSoMg4YNeUu568u
uaepiH/26HnJs+GcfQ/5OYYQLfyhU5jQ8SP5Xeig27+ek6/L4SWS8vq61Od4J8JQkUHl8x+U4jy/
mloGDF0JT5qepFUJly+cl2BB1y+l01j0phF2JlBdfXEQoTxCKL0lHVDMW728AK0qUY1FDBK1s3n6
JdcQrL7cJ4VzemDCkDqEYD6rjS0IRF1E54mmgUGNIa16nFNNd0//ilJGXnW/aypLxcs6/q9/mrzd
m0Rx4Ky867A6w09tckwQOLjfzcTspbQtxa+xfqHBtvfn0gef8M4G9DVCkoJM/u9zG7+l98WaasFQ
m+Nj6mSYIZ3JrkAZVhgONsdcI5VHu//nYO7i4O2bd4yu3XSlRPAboULxPIh9oXzwlh1qjTGJqVCV
XpyNTe3XqhqYweCQR8Sz8UTrjRXZ0DI89l6aaa00IaF84Ngz2rD97Djhbt9Sc4/E9CJo1lpnrCDG
aJE5iFRIzmGTcW8svWkAb7Ws8OJqn+ObmnBuLVbg7NPwFHwASmYPu9a7vQNoZzz9D+ODbSQj9wkt
xlCFP6v9fgCLXWxUUFjI5eoeI+Y3Ll5MDejjbTmsZK3b96y+k2Mz6GzWdobpUlPVcqRrrDw9yrct
ZOZVwDpvj6h+fslNF2bp1FScQfZuMtUonPUx1RgUA1S0XEkenVjja2rKcyqowkE8/LHH23GA47a8
YvX/SvSyfebKpyUwA2xDKV2DHBbxzS8aUz8OHH9pBAh+SFIYKvWTOrv5jpreuW5vpg21uhz3pDde
zNnn9/z8aSDeHrkp4S9GYhsxMhJ/dPHd30dcVtr5P5KnEf9zWIhXtS4KowDmUYQWoSWAqjhxJ5Jy
CABK89d32J4t9Lw9capov6NleUnnad9Q07qwLK81BuI510ZNBajPd73HCw7/63uAZcjnwghLjYcN
UzZhOLzv5VxX+gPKaGwGhsPoF23ZwKzq1OS5qdfFZKFEUZIrronDPdKKrLu/K170hX5rcAUISlXx
4qnh4qm/DVVgH2zhP/I+WsaU9+aKFFyJ2Ycp5RK49OTK14kMWPhKwHzjZkxCcfYyMs4chKPiR/4k
D9e9rWMY7o4lEXHWAauguoMqosQB5ltNBOadKBR3WbhZkyAE7o45KIYSG2XxPO+OtbMqPHZiYfoF
IjQZzGpux0yJwqxjnTAVGEU6kP9CyPxP2Vxybgx2X8oV5/nHZ6lN+5IvvnUK6QrtT+wmsufjTQXr
GrBl4LnlqW3sdZPc4ivKqfqYY1UjtFUYuJBlCFa/E6DxuV0nPVgOB7nBMDZKb775ZUZXlDu+ntxX
gu0+szlMS4r2vW870J5uCmT0/jxmN+loTAG0yqJoPPHnlCMsaptwWoOyguCLwG6AcBal0s1N6W1u
bdNaxqsv5Xc86eX6grfHGb/IlNH6J0el+sryvUNgW4//51+Pmoe/tD6fsZLFycqs4+Qnfv29YIir
GNwB3Ut4Lx4T/hPgvAF5nCROHbLoxo5B32+Nc/SZBaEmZh3XBXC58OuZ6GvFlB7/mLy5OkBWUNLB
Xr5RlTIS/5mX8syPBvSj4Y63ova8yzZ6pW3cEPSMD4M8V7g1OpY9PfP5ybhcA53y9FN6w0olfz/y
WTonXznKjdVeWjGUsLVdx/hFbiwW7IzjYvaitLSbxijvwR3T7D3Vhj+EG1V+9IfqKMhFk0SRvoKD
6F0Gw0ROHbkiCx/Td52+iwyglEFEMJ/oM+0rF7v/a6RRD4cSXHvCWYPfPCHrv3hMk9k290wAvLy2
SDKQwLWl3m+uRSHXoni+tEVI7fpMhJjx8fAKHMlzrO7aQ1jz1t80PcffVjQxeelR5wAYUtdEOp46
qDTuy3SxGual9TpkiOvpn40ZchHeVDUVz8UPt/CG6k34ReDgtN4IQRrAvLEwK0u6YCRGh6vI4GkZ
VfV+xmqfUSZPZEaracjTgy9AF6Fst/ktdRIqJqXn7pwpzGajdowT1HXkDgPiykvwAeunLPeE79rG
SUs6WY8PqVgYdVXyKnLBZsiEGQPZN2TXU/17noKNCkoL2hURDAL9pSCPw1qZAt8NNs4lehvV4Af6
AhXOAeengVMStYI7V1R/RLcucD5pwHB/lrhLt81RPUEM8OOjOsbbPWBk2LZY4j72WLmpUGaha729
mm4rjRAQmMMkVqevWJbLA6QbyUnNq4cnKUbRN/QcBEf1VYpmPcVpCU6OX9WJcSi+IeU3ba9t9er+
TtAyKU3/O96e1PQG6akj84mdUlDQZGUC1Jit1IU1Jn1/cfMv8+zetH2xrmzPHKnQ33Wu4TwhSkUO
LEbrkC/8LdZB35f0M85SaoUzHTuSa2S95gk4Laxv4iwP4NXxFwYiDXiONwTCN3oHUHC5+3KHt13E
D9YT0+9O9XYJduDmGgWitBxpowTkBLHFXI2XfeLw8GtV6qKJTVJzqBpThaUNyYRA4PRCuh5P6sAi
sFg7WJy7xwU9Yv55FftUR51f08HL5wQ4o+NTRRVPZPGLZ3q6YmrgEel9xcx6rFNXloD4hcB2Q1GP
CCdz3ieCqXfIrDnpbLu2g1WR8aZKzY+YiuK+ObScCyU2OogjlnjWljI/WCfs3060P/LjeW/pZoNb
7Q6ZzpFUWsAFXcaMqoeFYm1b5Re3LrZDFlJqpZ8upnH1N+RRS84JQPR9NshknOUYMUTXaNYz01Jq
6hi2jLCd6sMLg3uhm/VmIulXZds/ZaYz5UIqMqvGzLyF8B01rFzLHt6AHt6g6i4WzBvE0DW0gBIP
lDOk85zKoi3o9HW0iqi2gh34/xYxK/sXbIUJ1ISzA1lBIjvTtnfJL0ZS5DintdGwJAjFBA0FpWGN
bkpsGW/lXUGm+opx0a4nJFspRrW86ifuSahtAcb2mgHaWlSz5/S59krJm2AcLD4r4fY1FBRBbuFf
uF+CjtdpdcBzRGaGRXuHR+wHAKQpL7pTS1EkypMObs7E/U9jvF+EOhy6Dy8d8W2ta8E/s60iWCzC
iHSOZIPOSlOAyT5wnd6COMYZhQDwVGpGZfY1ahOqC5gW00ejkcwnt4d1BLTQC80aZA71IxS3zo/l
PjKZb7dKs9AQHAIe9nJQLcV474LdGa1/k8WJFjTt+TivGyPi4/S9dZV/ZCyCNpPN4d2ZXTGNLlYm
ymX5e8ObKP1NsKBCmJVtNjLziyFspd0fyOF+J9fCWOZbv9Y55nqSwueLWhmjdwPXAoe60YqFi0+/
MMeJCmmEDlZ6M/zXomZvQk3N03YePFQIHTKGfzHmyoU0fXBBAnufWokf3Wl26QrclzitbMBCB+2p
kyawI51ELmym7GZm42M6DX87bLOxz6ZMIjWxTP5G3lbau17bnsT1pJUzOJsL3Bam2ZnFPyjf07WU
OApd36CH79g2DRSNUzJQm0hlH8+TD9/hOKwPfy0RaWNdprALnj4+/ZVivFnECjmQ0HC1tRy9jvkc
nKOsnCUWsSoRMN+t1sZhowGSFHkjF3cKP+UvQeFQaQ47A0+WcXAXC6Ji/XF2+Oilcg2rJzsa/mP2
4wN86NzmNfTu2scyQcJTW74I9Fb7yEaWmLH6JQgAb/u/Lilemgq1fpl6v/TU9WmVZRy9FwUmJ/P3
BeJ0nvpANjoPaoKtWuji3Hlllwo/6YaGD9ZpzpygHSFHeXYBviK7ZYZNA4o283pcFeeAH2gC/2AD
VBTks7oPM1t/K1T1/eBffJrqdI7NNCKsiBuUyWfAmvye5PqUzvmKIe2+3THSblZjDqIRIFF1vPfl
HVCxPIQhYVhbbl7n8Cikpbc/6rV9td26mv6X10gtBUX/NEPJtEIjkxzRlEfpya1COoSKQYAVWF25
AHMDz6kwb2krekgJTgf+ulIOvUsCKN6th0o0r4vUhbWs9FH4h+fzebnZCY40k+5TehFwgDv79fMg
9TceorpF78faXtEo3BosReKMC0eDu7N/xUQlAFSs+G6qloQH8lh8cq5h2bj3J7wW2KqZBpEPncop
K2ZxY06E94vFP/OA0cvHG6RCUTuD7IdJuOkhuYosu90mec/UdNYPIQtXO/meZM3ZZ9aT3ylRid4z
yJf34tT+VdsmBPWzi/x1IyfpO8rbHgXQFPQMqaA7ZT3i+7RDn9Y+oDkDxDYgpVKMvKg2M95d3XM3
ESUsqzBuxExBELJyn66XVdQeRFsv6dWh30FFlEVLqw/gmEkeR0NgIuzEGTYmNx74XbiQrtzIRhpi
p3oP1/GtaepDuI0/+CSTmrcD74O0lQDqE7IvWl0cyaj4IKMtniPEeWT6+f2CaLDMIiVVFBuh595h
6OFTiuB/x5ZDO24ginijBlxGLOZkVxiEkov8ih85oWCddU6yfVainW1YSV43rFcEqTE0QWauOVW+
O/YdvbJkU8jy5wFRh8ZomhJTl3+Q5k+96sxe7ADl8JBiMadjGR9QncQhh63oOivVmE0Q17odDvL2
gQWvcos2WajuNpPLT3hSbqV4OsQnjZWy3GmRb+qfh8pJZlTDiKueEfryJUKx/A2es8K6fSCzRkZx
wP1tS0JlJrQinYAadcVmQp+Lzc+1RxXibM37XFgxWE9/+Ko3ya2+c4YXfmFfkTguQ0qhzZffo8AI
W8VBCr2PWoaQ+UXCJa0VNUkFmz6TOTPD8rXucatTqub1FTmRVn4G4fNaF/NNn1jUcZyJG4auGjuo
+yK7cCQgHwKWWJ5ja+ROcy6q+PAHCjymOkA/f/l6f7ssgxuxJRqjP6etkwAeCzQn16eUjbB/gUnz
uRc52kTEay/R0aR19tsOOo1tUiLPz3LD+ZyFC2rPP915TJvAjDzLli95JElJOM514CUrC1jtRv0+
nmw6XefSC79xIcMk8NnF5gxoy/Gc+Mczwb5poRfro6uA8I0P9YDFQyMARJbYX5YTqR98gcryukc1
kF0iwKwSOD9rHqstyt83RIDi6+0MlirLgPZ+DAABHkCjuXLiA0hYwAYbCnK017Q27/vClPDwCorX
zdhSg2RWFiEac/ktQibANpbuGDT+vZsOoYSHiOCvP6gZ5tvc55SWtxhxSFI0gyrxeD7+EUef+yzr
enBjHryAZ/sJOHLHU+nprkMu9ZbXnJMOboSTXm+P1S0F0foa0MzE+s1q/egw0EboQXiliE4A6Q73
s1TpTG9okXZIz9tM2F86hldfWAVi6wEnWJNgLJQbP/9Qdmsy9w+5usgHBX9CWkY7xxm6b5TyWwIc
RdT7kHVlkWkeYdCPz7u99w8lljl2Nc7DzjSn56ht/nwmew2xDyyaYoQbzEKieo9NcqFvESm7DXzY
YJz9Y7mawttQE7ItADDIt91ddf7cE5K4aUSL15mceaPzdyvYXyhq19/WOtYhRf8UREzjOaYv1IjI
XTMO+48tphqo69KtjsWC7mb24/U1+h0Wo8OlzQFTc+g6vkQmzPiSU81V8ulRGpkQuX8pYXUWe7m8
c/5hCZQgHGMFnetMCRN6w5aYip51G1dv+kRifJXoOPpI5n0ZLOcRkdRjyLMFJLij8sFbSk1f24eo
Yn3ICntM099R+WkJ3/xMJ+epDwqKVCYzvMdh8+pw+TkWtzufcEcsadWz2KhH2U0LQkl8eKdfZLP7
s50ttlvrV9dzStbuUvUeVp38+jfXsydRQFq7TUKMu9rLS74qPw/HBS6AKmbvCwYaSh9GJUU/PE3s
eV8RpWHugjC26XYF8djUul/aM6tji0fFwLsVOzRQdh2MPHACJ+s+ywiExRiIDlBYGdL1yNriTbUl
WD6y6FYzhI/vr+QT8+7Xfm1wA+xolfmwlfwSeexNzaydiTwr1Tmdt6wf/xEknO+g3PzKIrBAfwiE
4BPBW2EcHxfbv5obk4RPL8Ou2qwZYysOxK9RDljvJ0EhmMscKcQyZY50sULsudp32Wm6Zlfv3z3q
ifD/mi1602rGVIGTF3GmJGS8Oj04Zb/n15z48ophqvLXgImGUNBQLTBkc9poDDSfBMIegix78fr3
iDvCRjGdxrgXRmrfY9AXPRejznsYyWmOGoTxffs1q0tXvqaipc4Kn+lKoYw44TvViN30XlwDBLzy
ElGA68H/40hidMZpzdnMfL2N3jxUX+dwksQ3wP+w6Nvsud7xKjoJVq+sJuILfVcUdSLKzJOs75mo
jzcLSw+Im5CfoW/N/6wR3PLufbtzmA8r8jutWD+Pk+Y+KksrXGDxTYUkGLRjAi93SqJPBRdEDicC
cUWkbGJiACwX3aWhVbMf3PC+OqtfTN5HZ/Z4Zc1wE0+SuIMN4kTLaKg+aiKF9NarcGebETERXPQj
c9MKXGbrNKJMpKri2ciMiGKL43llUMrSTFw2ypYlIGPDcflSs1yIDdqcgbrdI4Qbs1u0D5j0NTFV
b8bIRnd5B5sXF6uy4IoTEBPqL9xAFcFI/IYRrkck+senRPCgrWiFJhG8f4vwuSSF5bPxwIIZ3AC/
7hmc1cbZQW0JbuUjPJNUIazgEse54atsyvB23ULiSnd/eZfnRg0C/y2aPTYRGEEQH3/5VDXBAoho
qAL7sG9rgscV5F0MmUTyZYC4NgMlNLKUzHtowwUrDhViERInd9Tn/mY8Q/xdTwIorcSk/9u3bleL
t5fhCMXOJtDyvBJUG8dkS6S8+Tn1zneY6jpQN2lzz408hLhEWNWST1lRo+7A+28HeHg1vdlR5e4t
RpKj8+xPJcC6kGT9i1X/enuSEgGabkNo/PU8iKIsZ/bcfMx1WG8qi0uVs3rSz6ocFnEkw7rDH+TU
UHWxGxIjsGQL8IGWgr3SEbrqBIPP+Gq5RKObab4bbKPEVXXM0p/kjskIsW/19vrIIkEeEb/A4bka
R4mbB4worVh57F2CusnIVm1jglnoaEj5PENPw4M7AiJ9mnYj157aAAL/4xEs4nqAYR2NhFuEtGVG
DmkMt3fXfjs0LcGt/OyFm/9loLbbmXlshyS5LzHi6Ki9j+3eYy5Cww5GWWgyayp7qc4xEj4AxCqk
xGJY1Dt7iZCEjarg8RvD7xJoOWLaE4XlHaFQjKxpNdBYfgB0W3pojVuyeg5Vgw+1dInTAqcOMMcF
DL7qmLaV7TGIPDWx+E0j4T3BNwmidQIbUotBUvtrVAwD90dm2MG0SIRF2Fz5ynslgH/iUL0uRtsF
r1I1Tp6mfpLW8WS99bSa3MytPQKbiEIrSdxB8qyBZ982Zckcypk0m9GcseSwgvmOPkGkAR0kUIdS
N+0k0i2x86rXkKGF6EMAm3QSrYCY34HN867DgRenCJjDPF1KsTovlOSFdY+OYF24WxuTC7sJ/2PL
5fLLfTJz2Yx8zZGdRpg2YEOi1od6HOy23/NNY6o0yOt/b/I+J3at+cS4fe2xcZssiCr/Gt4RmmAH
FvY806l5qhUo7QRDCU+J7H9arVUpVNnP+rvy7X3QVSHuMpX/dFuQjoIrFA1qwp/Cj89hIt1sILXV
s7iVYKAb2gQWZdZLUphVRydvHNrq1/BDLFpMwBSyDi08dG0ULzCZuHkI0VYuNV6EpgVTytOV0bYp
TQ+5aKwcR3S1KnqHLoAHw57aNklp82XvlY7g2+oqOZE+YrCNX+rGfse3PFfxFXm35TCKZc6aHsEg
FRLgY3ckvuu9S9YPRdj5MwzEBEN5poqnsJ5gB1Tz6rfBCFGkLx5iVofnt2BR/+jBKB7KinfGgW0+
Vxvc8Q8NCMPgpslLi12ArwXzijTgi23Wi5KoHqfhWB3UNtzgPF7/mZhkaKr/FGnRjLKumWPUC69/
uLN9MnFj1TEFZJeEsvQ+WQOU+JfMhV1Jx7kGmjLB1e7LqKxUfWgoYzidnBnPx5tyjtVxtrx/dCuz
r78T0EpTTDtvoM1pkkAcFooF4AbnXiXfry4Nn3+0OPiwyuaEpzwHhJRw7YkBapqddaMmVB8tERoP
eCTaUyln3YuQfTS2WW7g0MkXSMzAZZVV+C3zt/5nlkTNk1Hy1hkaiwuosqBSSxlzagMDdKj3HkrR
W4CIfMybozVVdXaIjht48dqr9v3WWZBvrlsXaCbOibWVRP1YNf5JjV1YtuMGe1NOwOsgf25CztEk
8TqE0M1b3H3S8fIzB4SQ9f56qZQaqon8eQPzBVK1Td1bs2Is2uZePhf6LYCu8vRlyyBBfnftdps3
dZVlzEwUNQqQY7bPpj6eBMjuSjI5wgdBKCutAZ2kWTc6Qnfd6cn+SejQ7ecWwmuMLIKIPj6/KUhi
8ZhLq0vu6J2B51rN+il1BKfzoAMS27jwzBYGFAy+YFQjxbGQIQ932bd2w6KZlH8IkK9X/NavzoP2
wYJf1fx348KUlqNJYzWOzxlAE5Fz7Gkq4GDuIOGR6K3andkobIE/PwL9TlaThb1tlsvlTFaX/Gko
H5IW+2jpp8RLW/+bxUAMON/Vs+WbaBpLD0npROI0ECYtWYecvSENLDgvNaomGL5+U0X+/pslJ5if
QybywGBA9R/Dyt3dPKbb/s3eC2xAowOzf2bohjfutrdsmLwikRIvGl65jti6OSKzrRyzFMyvJcfJ
ait0Dn2U/AKjrqr+bnzCVq/Nov+t49aAVk4Ht5Q+EvpffAoDzIqG3YdUVxmo2O39U7LXOMRxow1M
N0m7tngXDKZ/+y3X7CpkV2Xxfl3UnWWg+o+NkophmLjn36nrbEBJONGfB+dV//QbHJ1kDSkaRBEP
xnPc+pAltV1V2r1ZV1cKVN1OwbUc/jvhuu/ce5b7gESSUlLR/frS4ya4gkF+Hqoee/MJq5HwcKGw
FO9T4TNRRmMMAeVcVx0xe6SvOIEGZv8EQfcqYSnW8gWJVFFGeVdMIZQNmfWETJpL1X05x8XXy5P1
2wJiRs1RZ9pvlgVmEGZYzdgewM35x8vpOD4ly/kiYAPLpk4ufwX7ewPH8SrsvK/JUF2/iKU5mdmD
dr2auR7+eYjOSOyEDPunhOwA4ngicFXQvT6/iW4sszgJTU7mRL5C+2QTlp3jldjNyRvz9VszYgVX
R4C8imDRRBpNqDZc0fg5uqTKe55t25RUxmnRPfUlwZGKYeNBMGT1htLox8YdEwqWj6P3aHFrit1H
j3vnYJMcUUdIZvEPzghHu0pQerfotfoMp4jdaTBITdLZW35rgHk4eVGTfcLuiF6k+m+VqKvH7t45
D2BzdftTHqQ242VG+SGpBGrMUtrxtsaJ+wli3/iCIYdO6bTZRAXaYKRFobeWYRJZh4qd9lS8VU6e
Yk8Y/Yqqcs9EyJKI6zxhR7t8wM2Cpdokc0sC8OqmTmqPeuFEXvQcYDpLxsjkVRKW8fxkcoVF+2qm
gedT5GCfWrfr7DZRndEEFx5zqLc5TXhgVJmIoBcRyt52uAp7GbhzysUS37xZj2LZTTIeU0UKClC/
fVwBQyR1q8/A4wxm7poQypPAcDJtmK9/+1GMKSN5d3WEO/SkvS0gul0dp+v4OMBAA7j9bcXWcW0r
SJ2kUGLfUbOZdB1TLj/pn5UcLAx+kCNERFYo0T6dRGRs0L1at4hVDQcpsIywqFuuCzmCkgBES9tR
MSiQfQcdnaCyGevQ2Tp8B8SK5ZtgFGo6yEJ5gKbFTNdFgSWmb/RXBkC1YLnctbCLL/95C6UPw9wB
u98lRb4jDKkFMGoIDQAm0k7vJ0Z7Pn1GYiFZ/vnc2YCTHIP8RK8VsoKOwSPe2vGsvCwsuLugOOyT
s5YaoHPnxH2LpA312gJLmcxzG2knxsXyq5O0vw0p5OVjdMy0H9m6mdD+yKU04CCDVwgPsWLSvOqg
Ol2dCWCW/4Ee0LXVxI9NZYqQ+DeVaj27WIzRJEFcxFSpAeOTb2xHmt8sRsrrH1THdOjN5fLWLgLV
QlEu/D16tZEw1y3yj2+eqs8QbgPl/XggU22bFZLgqVG4bf+TmmLb4dqvLPNv+Rg5XGAL+juN0EY8
VzKQCeAtbz+oR981/IZl8QK+2ClxpACbcXL7LjUhVXSMwD9B5Rf7xWYR/qN43N7xKPFliH6yXJXW
cXF8X9FpdAKdBR+LbYj4fbA65RWIgopdZqkTWuj5gvEprL26JmHP33mk9fEAnz+0qiSJicXpMWPo
R/xNRvuzIRuWwFv9vHD5dt15vCFJ3EGCAHQjMgYv26Q+yOmiBTg2vndHCgGv/mq2wRJIugquAFH+
6xT2FPSDkh1KJsgrP7Th/m48CIO83dR91Q5iVu5twSzbOj/4ESd15ScXudVl9ReUgvkvEpVCbUpH
K2GBbT5i8qzuGzWktqZsAY+aB7yJHPUQevNmnHqTcexUJIsbWDgUD5zFZ6kUuYPeqDl9qbqWZdg5
ro9UR8EY9NMYY0r93qGtE0KGymx2KxUZR/PTw0jflLPlC2ntXe7MZnFLnoUTIgjc4A6Sf6E/LwM4
CUYTIOygOMOxLLd7UBkmIIh98oRk0ydimMANtxGksqgaog5uQunKTmjVO7r8KvrkBX+IXJokhAco
hL3wxkit31vN/pIPYXwKY+j1nS4/+dWm0PUy398S3rWtqwsdKXp9w0vEqDUc3qLxtdkHBfsUubsE
P0IGWfr4x2KnxqPyiMoNLJC/MswzZXkoZa4EXY1KwAmsCJvx3UBYWbRqcZZjgcIa5/lCF+9wWLia
TaTfjdbgu0p1Y9P881xl0dbHIIWxZqnL6TEiihgsumLz14r8mar4W5wjcT/8sORI+2yY2ddfy3yr
Y+tsoej8fdN3BMYb+fCq4Wc0ue5KEIL82jkrMJtFyQ2RW0UeRFJ6jWdpqL9X/eFYVdhRwRypbY1n
BFpBdWrzpfq6T/tevsttLoxXbUQ0uXj3aAMTtftFfxCtBWWchOdn/Q8TlLUoeGoGjUD0gfi21P0y
EQLUaPiSKdiSQ8KQv7hLV8rnH6WIKaG/pAB+x7S/u19IJg87uep6zjGegpSjdhkTpVdzjy4GjByg
P3ulS1xEqPRl9/L13jY7z9gIK/pTNd0zylpmWgZY5XNz4yx9CheklaLxW+RupkZqGGOAUwM5fy4a
LBx/r3YcGutjxXogyHd1TVW2sgvVtVDfT3Mlamt2df2iWmVuTiE8QxpGfyxsKKpY20VdAUHNua9K
niHkry2EZHBM8mRFrhl7gzsLyD15LqgrDaG1FwdyDgCELqyRXbeSUx0vPtDIwpdFy/eIVb4nAcz/
+7O17hN0TUL28j97UvWBkBjR0+ArUaNwWZ8e0jGWBsc2/YXU5o4/VmnlgHbPxK8gUoHeaPfl/DZ9
GJ22FSJZpIp2U5fUQIMYal8hABJvfZLxYbTjl2KT26Onc2C6kj+703868sErJZs8QGLjmN37RJZS
EmFMuRy2z2o2PUgW/0jexfjRpKvdT+GrHP0IKglaT4Vti/fbwAqZH7Cq7wTYTcn46i1uuPCgBRoE
KZBf1EOYIRy1ruIIJJaf+9Hb1banE752kc3EMOb770E2LJ1BuhIqdNyl3DrlqgMLBpI/HiUuqW/E
EgRR0KU5C0wa9czJcJAaLolzbcfenoPKdYT0J+P2uYd6epC8klCHatJ8eXTZXY2bUoczJj/QXLP4
wENdBRty07hrKDczX2bbaKYI+yPmYqyDDoGlmuhkiuFZ+/W6X2Nd/HEePS6zN1gUbP3qXsNhT+kx
W06KAwNAWkQTv8hoYVcDE8X66fTLCPxRRALzBVZg3xf9LurFn6qcDwXF9aTFQ2fweqd6CblO9Ud5
5p4vaygA3gglKemIYB+tDGsYyUKKt2fBVUGn679ngoDPkJ860OVSm+7YJQpjHCNYfRV2fOd+mePl
CTaKKZ4sPZalrTY1aSV1mCSlReqcZ4feu3WPwamwU9R9RnYc7l21aEZ9uXYm+VkC+qwMWrvmF0a9
uwOAgy6df4IVQeNIMO/KVmd7BlYLsyJQYb5OJwKUOIn66oFKoTrSIhTiNbOugvbWbpHroA3rVWIK
hnCmkMnlJ1f4krbrKl8ihtprbro6+I3hykiXWRKflwA3Nmdgj/VvemD09xwKoEPl92iEjFZAamIi
uXqsXLWzzYLyLLAaFURs7g9BMxXwz5pBE2fyamBPOqceB8Su+2MFRa3efohRBcu+W5QljerJgvQe
/AD4Iyuj9c5cLRJ7LYHUOKC0I2av8I1Nns4XWYwmWNkUOt48+rCjaq3S48jlkdb7Mx9Q1roDn42J
buz9cHVf1RRGO5NqEVsyfQFHyMLwxyGa8Nph9wE6wiHC0rGdwUHsqL6g1d295/P7iw8OVihepTiU
I/uX+4cAu3f/6MeER+47xgI5mlMwWgGMgrRL/lO7tDpzmGh2voU7w80Rulz7CdH6OCVYKGmBd0SH
kPnJgtuyhFrL3S8euOE5foqRqdDzfNwP4KBLGCexWHn+tfGhU/kIu39bdNA47uggeZaDtou7lFq6
BWdQ7cDPGQ9Ts8nxuPJVNKmfNzZ9CZdTdPaTmPM5LyJoMUUB2gyZ1dRa97IHtELTPh5n3+b//hho
7QKVHEk7hb1o6GF9dYvns2iqO585Som1Hv8rr71fUA+86OwOvgpIERvXA2PaQBgbHvMztDcFNtao
dxgFrPhwe6IjnRIAKknKXQaI5oRFoeP0KxPLd0Uxbc/Yu5Vpa1TDvgZy6V2zgkp7TsscfuFMtH1Y
AkQicdsswe9jn1ndYy+DOIAkB8MJJ6jqVfBkH9/kRuN/lS/M0reShEGrNa31H4U6E0bVxYEXTK8O
2Zq5O9OzoBp0/Qfy1URFXrw+/wHDL+mnfwXzlX+h+xldmiL0qSOprqzijhH9laeynE14WkSYn3kV
4OKNqbwJg4wfdWrdXIdIDNMNdVRy8ri3DY7GzE+xWs7k1qgGlM4SGZl16I4mOcXa40XE2BZCbCAz
JQ+duN9by86nncSauZ6zidJoLtuwNWGe3BQUXp6XfW3ZvfmDejRt7dV5l8RTscxYOKvmOu2zf77u
NjvNdmxuS5pp9LdP6Xe5D4yPXxDboo9onrFDRf6Dn2VqcVIXSvE0x1pkZbDVclpaWK6Oflq8SDlC
cijSuI6vS1ec/0U07H/ZS0YvETK+nytGTYDc4pqH0fTBT5zcRdLTejRu0EN52Qqip9hTPl8pTMvm
tebEvL/XYPmWRd9W3gHBIFyBxlpKcKF1ay62CGtsy4ku7bNqWZ6mMlSFfuO+fu7zuG1dtwiL1x/g
15YbYu5viwJdn2Oq+SiudJK4ueCx4mtRpkIvSgCYuzQM2rCQWYL8hdcWTSgPzz2+hByZbb74eFCx
qSVLBYqq+i/wwQlOBHi+xJGQnzD0QRyp6aMNyN+DKv+LitnVnJOmyMmh09nDG0G5G6fIGTGuGyfs
NW9bcl8Gguke+Z/RBUM7poBZZQqflqtfwG7ZNPsCkQqoPyfIjqCi1vCJbr52Cr9YODvOM7A1GEFF
Nab4BDcZ6TWuzcS7DDHs7TgglQ3I3jQ8pvwOjGenAL67upGzJaGI/mdoFlhntuFnA8y277c7fHxa
pbkRTJBXmDK4+H7i8mu4qriVdfbR/9OyDfr2LZItJEFLznR/0kwEdj4t0IN9zlEva/ZBw9Kmp5HK
d3hs/4HT0OIwrSYT7tjanjD6h1qxFD7i4eQ1oDxVsoB4G5L+1ZPUGr1UzB8jro7A0TYvUUXFNQyl
r8kSRn9iufHw5JhCPktokFyu6cHN39XTGm8BML4FHiSftxUgJ2bXG2nBoFbaMwf31gKPEiXM523a
RZHDOLRnk9dBXDo2ei/qCttrjDWbJI1oDfOzUqdAV/11yamgAYy9S3DUsgcM+Wv6PPGHHhtkocWq
mbfCoZ51Q8KeRwpMD7am0vmyR7FWH79y+E2I/cyodNLk59mpah9Tezwl2qphlFoSys2UV96EpCWB
45sGl1uaLA5cyoqgKa3S9T8/VxjcdyCb5UOgYPzunzvwYJYYwHG+KpvDGJeh8gnWpjDb/6CTIFk4
mFxD19lZflYlGbmq0VHz9LUMa6VY9p23Q0JfE0n/1uBEp1bACAy/pLmbitBuhkOIoV11j8cdr6sP
EkDl3bhoIn8uYKm7y0LfHqEEzbVC7CoGxjLc6fWlZgJFRJUA588NbG8SrUI9Xk4aSPgf+KJJ1GuD
c11xeygCyAwRbm8DSb7ZOT0wdSCMVGcgVBQBGh6ssRhzzUUVCLTr85nT6xaLPCN1e9iXpT9qjgPE
ZS5Cv0+1aI6iPGU0LPA3dPbfUzPvRe+BV7ItNf5v8CEdrS7fO3BBauG7HiybwCmNbSN+5ckNaIT6
PTwhMAQC7drfGEZ55kUk7WbRWEuMSc2LfGESet58sxGk2Gmxg05lwG8lz9M3gCZOEkAnQ233btqg
AGdQ21zE3SuGWeyanKwirgus73MMUb/HXA9YmQVYnh3plkgDqMWEBINRnoAm0u5OJeA1YWg6FF7G
9YKK4hJ/cN9GWaCcQfNukv6vS+kVPbpL6PjcBOZiTBxVoN+Z5qhDCZpdvb5pwqAj/P2QM4+S/2Q1
QUoDm1Lu35I//0Bb6xPQ5cLybKKbUAx5FQGWLOcjAsgjzDWcKgRa4aykN0dnHibnrgGhFHFmHhd0
Xi+sSA0D1JuZlFrTGDIBHEdzJW0AaDhigB2rWmdh4uYLjjAFsSMiioHhE9sZezYQSS4dgzFCh9VL
ejM4o/YyqBx5xxUz61WB+lfy7QEDh0cNbkk+WuifWqcrUWHSpFueohzzJ6QG9jTdaH/8c3dkbdbA
WNnR9zAS0kUqG26/esb1sp/bgtdUEE2CJHcHXDkIf8MMhI7CizWPYE9OzY3fle6P2U3+Qo4SWRVy
kmkp3GDqxa2ZSiepsC16PL0MeEZEn6tITLyRd8MEVHTwK3rV0lK9r/xoYycsmilV+etf2/q6GM7Y
SARVgT+siIWzurI2DfIVR+ZvaTyMDU2cba7646NoDuT83xdQfxAxdg6VYKttbvFE74IB5XskVx84
11lLHwvYcfTnNPUUVoZPB6n5zjxbJRGeYIp6qsVzCZZ2y9y7/sDmtPp14nACY37zOyryptxOY3Yp
dQztTy9lCKSqvWf4yv3vh/BDU2vssgRs3mUux+KniDd+aV1dBI0ZiMmcS6WIKzft0JNYGVYNopLe
lGffAft9NUeab0rTwJpGKIfJPVtquDX9NDOtk03eC0G/pibAYCEhaS4kOcmjnsvp43pSfMnT8Me/
FrVMoeZ5V+ZqGBdQSIJ6qiEPMGw1VG5UDaZWk4zrwDCeTyjJsZU9mmppr7azPDUc/eCDSherEP/w
Nu4K6ZuJGiU8d5kCqozuY6XsPWPUPQ7076rmpqfMkB4017k+LjgGmOuyL87XF2pMml/VQaIveqx6
xcAkEB7f1ZTv3uajSAdQkFcqJCTsMBr5Xx6c8WicXizw0R5QGvEdktrtiNyoEw2yd+OW6II3PzOp
rMgD72RUwSz/nqgYrslai2t8wGic9S/oFXLQX9iYR/MfNhJX2iU2X8qZy9OQE27g4ekfGAy9AhZr
su+T3bFfAE70iqcUyE4Izf8HaX1lIpGJhoSq7xNXjdgzd29HIUCXjQchSrFHrrs4magaXspo0mtG
ViwsLro5CEgVNWQp6fbOL+2MigQ/3tAD8Uupe9MKJZwfMk14ygWxBHBBr/c7Hjs0xsVr7BPn/cRd
Y2IsUWWU0YjCciH0I0dmX2XvAH+/EnG9moCUYkxB530EnmQ37fV64xe+VZM4h+ycSeHy/zBQnotT
txPvhgV0BX4swdjrfvKgWz3z73rrZO+4GlWatDVHPJT6vaEpl5Dx3xUliVFMr1NGKDW3vbMZbRw2
xSNEj1rZYqUosp138i3pjmD9WwJCYKDQbDmo3VJZuej7/z4C5GTSNuZIDIJwNnuNf8gK1st86cTs
oAWOOI8wvmEd8WPezysUvUFwc7nf7KMpY1XdC0WZ8LAxx6n9Wcj4lgTVjSzrCvBan3h6DOLDeeGY
EVt23iTRKxlmuRvQm8RwKYtno+VuGaziAjen6vfaUdJiI/yzCj5+oSlxkTcSVY2neibpA+AeHTXR
ouuETqA45g6Px9NIpa1xoEFKC94vhGgVd9Gej/mtet9mKgLcIAaB8yXVTDtGza3VOpufuUR77GmO
n6ZSrNxZCBkY3jbX8pdIq5F/Mvh3DRAGPEMmpPLeSiKR8c9E64/FEEXMSDZdYqMGf2+NMineOMjv
VtpVWmzkGZSTILJC4ID/YACEGqTE0NXPnjvwqH1bmxa+xJwg+aO+C/J3odvN4jJBnCjbCTk5NrXY
vcIqp4Q7EwHR5LHRGzDMbIqtn/lZwcmJi/X/75lF4gDoI078Nty6deaQ4WUnYzI6Gd1fdRq/m9S6
yDmCnVBLWBinLGrhfOEvic0rw/5wL8RbxF/N5c5Pe8U6sCB/1nIAwWPSlJwL7wEzRMfyFURXifGI
jsnjvIbxzETEsHr91NP2NCoN061y3E43ga04ZnqojI5Yr3kTc66JoIbVMueRe7YWVpgENNvupWi5
QRa79qRKFA5nnd0WBw30ETOe4dBDYiDMWd+Nn2oabZhZUm/BBtulKLJYAt0kXaLnSMTbUTyo4vCE
QmPL+NUKoakPMK+IHJXfU4+rri2+eWuzXBr/2/oGQJp/tEqHNM32UmAl1wM/9lhTiSs8rOsoYbqq
s3UV6m3Ms0NbriW+WqP545ya8HQkij/r3qY5XqPMRhm6wrWJNvt6vodVllTZT9TDd4ba2Qu7fsUX
PDnSH0IYZoqQu43ZK3NaUVrRpHi0/x13y/5z5V2scrf4O+Zpn+d5by78o+ZlYeUQPEBpj9fzM63U
QP1NHtRM6v2BuMfCwWI69yZ7WQpMs5sZp4nrQ02OHSLqhJ8TmmI0pMIFhTmx9NFuVc4UkKc6TRkt
tZSP6TgfX9BK6C1G/vMDl8xibBhNaAAaswHFLLzJ/q+orwr2p51XvNq5FvQm8JKUNOrRVXg4v/Pk
ei8foATMW8M4bPag9++vNIvY+MTyUILJDaMqhLdMGLBGa248f8LhpRHiDUo+P7uIlFtJQrGoAQmV
9TkHzUaoemuvxrYtYq3a5I/XTvhk1Sq5bj2bqVDj7FQrzlER/RpRS2UwPfVbVVRs5Q+EPl4UieNz
fB+Z5jQM5/NQzE8qvFDlR0KZKgZVP7Bgg9G9NBGPx9d+8vlnGdL2zFSm501jjngMREmlruhJon66
9Y/Gp7tduBlYfKcO1mdnxHVBQ8W5msOLwaFuHIEYq90D8c7mAHKAT/ZwF61rJWOuhOiqPwhFeoDv
5yzb7kaRKjLHNge3jY8cRG/GaUA2B4Qh7CToAxwgF9PVkA9RG1jmn4H+pZKDFKZ8/MNW0F+H4xrn
jHZsAaSQA1LNaaOf2geOquaC7mp2FvtJLQw3meelwe65BpAbwpNLA6sV6U/Q1neRwxCC9qAtgZCS
IxX9Tz89j4GKP2JRvpHH+PCFZt36suwsmgczWa54bhA9Qxg4BEVEVWBNGFYV97jvi0Cqzgof+Cuz
nzTZugi/JgebITOcVYaj2o/arnZTltB3qA+eNBPCHK+cC5o603gL9Wc8zMbEuOpsxKBeP0N8Q7qJ
e2rMKKMg1XJiHRPjRdYs8NWUCZXooHddiFW+hCc339SUu+/jqdz7/5Kk1FPzNe6pZ+H4nsf2DUTG
mcn0t9WJteZhZA0DGRM6vFIUXQv82WLiRRWk8vIgg21sLFefaw7/Fi9u4RHKd50IUUj02FNWX194
Z+9uCwXjABQ9/W4wCt1kL2nj7/BwCxGV57ygzqnrouxuKujpHQMLSTGR7BHfA9d1KXWK2JmXQR92
rj5FKNc01NJmFCDSZaus7+aDHJ9QvmFGMa8jKrKl3ao8NBhdlKTnS5Avebz6xQUvIIpNWa4gIAh6
WZdP2dNkwYVAP9h9NkuL0f4WL+Yn4l3Fs/e7pFjqAPQplj62cpd1jGr023u3CKHzg0Jtqdlt+Ex6
4jiLQ2578KXNntJqvEyHNY9YXTcx7cx8RZhfiy+b+HH/s7COQnYf4sNoeRn94yCIhNIpHkn7rhed
/Ome9PxEfbpUSdh6JFcqpGnav3iYVl7Yabzas92VSyVpWysPQMbYwa9uvV02ahZy0njYPzivIVqY
cmzLXiWDm+tDaSJaOjE4sPFpwilP73s5fk7w1E84ENabCQPxA2ccFGZVjDP/W468wmndmMhlSVHF
bUKf1bDff+7zWhiNoV0YvmW99IimFvDzJ32uymuOu280fXw4CO6Ris72g15ukMWbT5vGdGST55YO
6mL3JA1SNAh8Gc36WC4mNQhAEutVhwkfteOU0Gftq/l5bjbpTYBpohFEAn7gT5/LBFFPmP+kRD57
eIKvrZmJIFc604e5SsyRl7QzyD2ldWjxYt6EIzFmTce/kAeVwsQoyL/1di1ZBYQEiMfbWYi1dKj9
5u/vb//Jzhn18xwG8pX8lApYbwjBQhGD3B4X0Txb45RaAZZbFKEXpqHEoR5ceZVhtQI9S3tOKMXH
c6lSbpcxuG4ENFmHo/tWA28wMiNX2LasgqL2db85ppWZ7ixHt9EU7bV6TGa4K141QvX4b0h6BWoY
ji7EHyo7rmv8ZZgyh1s9DVLvTSQU9+JjDPZOUOytcRXarPNroSSOvCGt3u0WXl58IWS/P0LIhq7c
6jtT70acay6azgL6y7gMu+dQqY/Qa2zwv/lvimAqo3obj7KfSz2fqSGFPwaxIi2jF/T9QWQGgibi
+mYT4Tzn0N+MoakZTLi16Lsh7SvkgwPsVjZcZpuNPvDQXyqXsD5pOez0V/jdGuSdxfeCXb64kqOb
L27NzduvR72F8kx0DpBvSc90W30ZuQXuVRuA1xQisv8q/ibiq/t6eV1gvL1l8MKbVAoHUgdsJn/y
VsIlFTuYYcLAKk4g4+Lq+y8VnuXQhIC6dh02OY5Yb0cSnvRmrPQVv0l9F3JZrqNp7dCXYnhquGjs
eF+525Z/+pP/kLm8ugBP4x97q3uleRnePofFczc4FLK2hVsqhqSK18kJF93wKg7IuIUbV/+BBMFd
fsY7DWH32iXXauSg74CrPjbXyn0PVVipbpRXpvcJXqY0LFt60lHg8I6/yhm1gw+/tzt0S0AUk1eQ
vfeFblv5oTF95NO3gVXrniytBFoS11NlsfMe1GcUqz2sblWwYDHzsSc6bqRCgEPhUSMDq76pgx/J
Rx6d7xM36aiIyIJh4PRAIJs0pMO1jTNQdrzTgo9OZr6DtB/WpwPXPXXur+f4y/yor2euxNsVz4zh
ZQylzZYC4xjcPZJWzA8izOKDgh5ILnKfXjvdSrlYHGNjd16sAHCtvXdtURDWVySIJ+T7BIcDjw53
RRbjD+iPIzfTBdsA/sQa81TAI5UF8leauNctkiBFhziCDapgSIYLnLKU5bCDRnkmdeXW53u6ikZI
l8jbJcQLXCw2kTeArlTIwsfZ93uCGvfejtyU0vkPTbWXxGbPpnK3l/WuZV6s+89UvXdUZUIU6438
FfBdvI1CFTxl1u9Eap0n3GfeToOi7K/rt7QiJRUrELTfA/EB0KGv6IIgBckKWHr56ubhR4tVVdL9
ATuv21Z6S0PEf7UrqVnBAZ5uAxYPCDcq8O/3ikc7bgogIqrfWAZwDM6s3VEnHSh46iUSCPwr1gDw
mdtpoM5ujif0GkBXwbemMIBbLT93mavEk4A7nRfnNMix9nefEcUFqIKmkg38nkQaAazk74oCreWf
k2Ds1gL+DOWSgd5gz0+KKJQ2CdhHvx/7VeIZwFL4ZFsUCeOB3cBuxLyBzZc1nnF39+BbS7oENOxQ
2I3AiC+etQtaBXaRm4HpIPU9p5CeuNnarh0Wn5/trVqZZ9YeKj6ZCeWrQVZDQGDDC9gjkigc/lsd
1a2e/LJYL32Spphk/LxMNiuEAILNOzDN686lmPcgsE5c7mEhsbKg9hJzdVDgI5nH7nGtZdAEV3GB
gISOsndwM06eiQibs0datY13GkQhmRyRv5pgLitEnMErCaJ62XwVJgDpzhImsE6/u/0YwMIeQqn1
JFzee5V9rtx8LvYA/n/3SsKcAIS+doEAUhTmUVqnbp+eL7i0Rb6iqzd3zmla4rD7/IMrHjA1ut0e
PCSEU3dx6tspdNpHlMEB5ts1B/pAGrZxn/NWikzvqWG5MyyLhPHNNRWYzEsZA0idVQIvOvCYYLzn
75N5O4fQZX+Q3FK2s+mFewivRXY0jZL+Yj/Nbw/elm6+zhpF28o7NONRO2QRQ6n6AaKyYig0whX2
ijjXKIfWSdDmB9SoTdi2g0GJ58sQNqlPqB+vfuuXKg2ssEHxU8KfF+qVWAWxHQ36+qPO77gTbsho
AUSOBmVxpld66ezJU1wV2TMiBu7oGX0R2uXrYLLdDR1LJ3+8/DMY00ZQ+Z5aGot9s3jasVEQ9JZv
vF8mNnh2OZiDFI/XYz8BM+GXIuEQdAtB0B8QOD+BnoiR8vB0HMweJsM0z1g11kf7z+F+TALg1+75
CSZ/Gtf1/ajyQuB8A2zHnQQARjpeYyddME9G7B4cYecB/mCA9ian1RCQCYFd3sIwomc3zHvFeLcN
uFhSB4m+VVQU7ZV9OrWNEB+2Xl2M01oVU+lx6damG7SboHEEbhOxc1khdL5lM2Ho0isw15onnQgy
wE/4M+Z6nAJl3gycX7j2XGlcPQEn9ImrNoObNqzhu3KivsSGiCxR1BqBfMydOlxm9lrG6ztA4Jh1
AMFvusnKOJHG1DShERDjwDSDdd2AB3byZICXNatLUAu7DRJZhE7/I1fUZJsUmJHF0k/sxb49dK4p
G/Ht6K56dJKBBufCb7vsYV3THhGvA5DUwfrBdNqS0p23R1OoBGr3bZt1qRbVaDT/BRhhVOojLISb
2wnu3NCIz3Tr4cmO8GfYX5nKy/vqiO3mzF/Jf2X2iuu4jbPbkOrNqNsFPlPJ0xavJPejZplcm0bu
bsF+S32hZAQNr3Vs8p1vGpkg4pKdR7ribgKwsCownGd1kZVqlK9KTm4DZs/B+nCnbDjCOvLbirq8
UfapXZbxVfL0A61KpbJXwXzzQGQ+maZSQToEkZnla6GwPGsDS0gxXKnvwkPxQsSxF3Evn1gwpUrY
qtBO+zTWuHta1VVvsm0GFKv26E2bv0+zIfvrr+c8Z9LenfGNpUAswpWihYRoM6vZYiDfarOvAqmU
kCZ6hGWt85TmHuuy0Qg/GVNrG8FjOZgnuCRdCW52ZYj0XmByJSqjwPw+IJYwAZ8Q1uS2GHrTG4E0
MlhM2ch9SeUJFpaCVhvBz8NaxjXDD8XnHmQ/XryWoeFfbckqLHwX348vVuzaBS4FcHuZTBIJ6CnE
pSylaNgkeqeeEQdeD0nN1uMD4IkWAtBd6uk8KRB9Kipoqab9WSrWBUaV+DDHtSfXqtYqwcZv3oL2
3j/KcoNjs2gGxyrUeqor7WhhF9pkPh9sHhNquWDjL77tL7gvBkCpnqa3FtGTta3TQlGDxlvHgguR
eUMp8wNMvg2TNkNgx7Ome9l3RJHPTB5f5lORUqSTnHvOBkiy5o5hU0PxAML8uedVWgHCylyv4K1o
arhBoauA10k3rofrBX0J01G5nIqGAlfLfVTCLlYydRILcUBfoorbSqUuOsb+uyMb8+aVaxkTJXYk
SU5mlE+OGMX+iiETs7ny4sBH+bC2BRW8uVM5D5xt1JsItI64kNIntuF+l592kmlzjlVrprly++zb
k7/8iEsguhwuhH5MyW8LwB++65yTZ6yKFpDFbqw7UOhvwRLu8Ns9r4BbLLTpmw6Xk7llSRyr+rR1
3qeZHuNA14BLRegg/I9qfD7v2lkSB0nvsV+CQEJaNqZnenfBetauRK23+dKczr8G80zvowqYZ6nd
vhdlMUi6ut4ckPwzNI8XHVeC58yBna3FTcNM0f1m0BRrM/97cjqnXaI8iULUeL1jJB3jpusg6cEZ
G0KOQfs6Jac4EcDGAlKqdlSkKrHmNKhXD4gJ8E/Nc5aNK+eVsEC0B2eSb4qhKipwW3VDmxOXaZen
N8FpiiBjo9w3r9pF1eIVnlsgeIr9TFkmzTgocZuD0uQE4CNCz840NcEI7L+TYWtlLYt2raAmU9UO
kVgDqw4y6QJK1bok8kpVy3HEnMF1Al5lIPY+R2dBcq+Fd5ZADh0PUr1u0UoEl0tw61nRzcrpjmCM
QBsUQ6RyElzSjxNH7NuRT+j8gtkcBQLB6gq7/TGCJosLok4VhGL4Uj5s9B75CV8kRAV++c39IVA4
+yUW5h04qGWMP/CSdIqyQsYM+PR/3i4LZPvGEXALdpj1jtypLGoN6CN6IxhRLnZN29hxh5l+ooed
Gt+j+zibDutFs+E2n3yIrwWetGw3a/N7RN4R6NaO5I/2Z7fAHm2wsKFqo1IK9SACxaTqgvevNRKQ
dnRq62wQXBJNbADBCHNGgZ1afbmAAi7KaI1L87nVoBhneBEeDb97pvRznW3xyj4R7nKbfCMtyPI2
Hx7bNq3/ebrbXii0m+uLPVX2FjXxT5ARwc30a+mvPuX81yStVoyv+xbopM6poEeAdiGcDWq3xgN1
NgrsK9VTXUyKG7dEptPw83yIvIq5kXbek7ckRjthx/tH4P/jlZ1KNfxVQ9p46U6J4P1+VJxdoVaT
GSpWTIGDKFCRRgoSveoC8JRh+WUvlKrlAAQVKvVQcmzER17W+dfrdsvD7+tZgF1P2WLE+IHlLBVj
J10cU8SHs2uDNWVU7roWwLaWk5Q/k/E6YyGih/T4Xgzt8y56MWSsOdv0HB/kwmBwx96f3YzF5umC
UBW9XoxkiuJPTYzBQJbPB78WQachfP2VHsLEJ5fKTFOCJyYepVQfEdb/O4R1rLPDuIOTAlYiZbv7
GJ6ZVc7//parinKaCy0fEu+/DiVzGG8SZ7YKHpA5+q9E6qpSe/t8WhdzIspjY01EHdmOcoin2aYI
xtJsuVVO6NU6GlUAMedyKP9G6FDmiEGG8O6/MN3tr+wR3SnddZE/Kn6ihd6+zZptMlJ466yt2tYw
5JiNyIQymqT4hOAjYAgBpfltWanS6iDVjcsFFztGeomXEfNVpP6W2EIBP8T8SeIputVnwT0jUWhf
bQjtIGm77HgDh7noaD0sF7CiJ0RsAlEzXAOm4hjk90AfoX7l9Y08fOLtoE2ou40iqRuhgWQTVNfm
0YObR+aVHWaH0+zY6VToczk+cZ6m8nuH3gBMo/y6Dv1D3usxWFDbiUO3TN36UIBofpDKVdr8tluT
w+IVTqaKegoAzKwgvycdjz1h1yt2YT5TFtmKtCidgBd8fRpPbbPrW45oZOPixRH6FpK0bsWmgnqc
5Ne4ftFLbq95JecI2+2JJ9tjMo5g+QzJB+MYSBTq0JTYsW4G3nPD9Oo9vfsgg0vwHGag4Jhp/QMK
1xfNEjBGujDqc6j6Q3gxw+Vzdrp+8hY/f8pTrA/Erxb9w1uRusIJUOYMDx/9QX+qat0drv/vNQMy
Smt/g0QuLlAoNXCLXT+tb8eduvAzDagwUjarQJF8a/r7e7jZcZsmLaAULDgV/6oV9FFvFyNaQDgG
pnGb5IbqxT31L3Wgw+AxKdd6ZwfM4Xr8JdCtO/01WOKeZZukc3hil7VaQGDqdiHA81yu8mlSrOPv
LPLzcwHeI57xC/FxccXtOwFRKYNMq/UpBgf+UUYwDxXZYzEPHEdUg0wl1Zt//RHRWfQKW9/44YAn
1eeLirlAL//uVPL0NkjAbQWJTs4u4VHZ90jOIyxqIAh5VfddcECix7YZqFHN+cEzObvVf7rWqtoz
eEWEckU7bD0jrAVZAPfQUW9LcDr5EVXUqyXE1gcjV2Olo91PHvjWHb9gj7pJYNBKfWr3n4avf+Qg
5HiiWsIpAjf8+jEob/+NJCkaadV5aENQ3W83MmnjgYyzMhtPqZJtWKmZ6MfXVQpGYk/b5PubWKjT
4RkaZhYAd7LxuSplHP6osvw9xQGdFJsLdyy1y0KMvHa2H41zg/UZvQENHYrgbWj4XrO0mmPjE0y8
WUG13wJz1gs0hjkJvrtQBJ1gBxZu9O8n05pQU2lCdytYaZbyed4M/V0MmXPxQTv8ip1hj6/hVM6B
/9BNly81SVHQMSTqcp3BjxxNG6cjyxazIndk/+9W0yWNY1W3JGqYSVR60QOlGI5PNguMoldVZwTr
ek4r23gUl7u9pipF1OTToxvxANLrdHoOVnst/VDH2QaHJ1gI1DMuTCwUOyThHkn1tyC8Cq9yVnso
Or+pSSHO5aRH0rD97osnVNwLYLA0NY7gP8OWCxnHDtZPhlTX/4n8Lr6GTrrerG5O2rvSqSmN4xH4
BeoFWkl87G1NJRo5HnAzcqqZ5uVufcYlXg6nHTFm2AmbVdamehWL1F4Kl34fjNm7qbs3YYqokGh4
yhIBlQddzT7UtzQn16tgxjpPe5wKGiK7AMJFwMAMF/80jJ1cM1KBfxGm51IwPwRmN+sRxjbkytb7
MfGA9Za9u48e1NfOe+U0RpU0NgZ5Pt+WvQl7tzh7NFUwhdQDZw9537KPjCePKurcNBWxqHeHu0aX
D0YBTUjpI8rOz/GChvtBQ8f2zunom7wmDKUKoDjRdtTfBtNdA8W69XUgKOqqtXsdecIZBlBtSlXs
xskgAU6te55Rr/wKZU7nvhOk2IpcTka2SP/ntzDj1SzClKMnwHNeuyqx6APUHr3Fx93na7pyJXEY
AZhxFtr7w9fSd9Awq+Kiu5tFeS+MO5MyAaPae6QHqyP1N7NqSPnP35Lbu/NJqZJ/FlPzOHZRmLlb
4agdKtNFsUFqQq0Y26zNjYVoLJSfBOccU+V1XfhsHREjZdjPR9q22k+2F3lv44t1qm4+8EaeynDa
binlO4d1Dpj4OvjP4FfpcyCXbogpO1e24rSQ9dzMqd6LFzdU+o8tMkRWU1OLX1DIxFM1OJgPBn3U
op2BYp76eVZGjgs+jJp86Zq/m3Q1bGzIOUUNTW1p+6LWJJchqYS3AEqKQMY3my/25ERKBnKvXkRy
J053CfZASHQxwRJCOE5y+6kdlhkUImI5oT7ho+Fv3vP4HVl1AgHRALmRM5DZyoQZK9Ct+FfMEObe
gtqapETlR//gqW6iISM7WBQAPwcX9Dw+b3PdffGJNvTXv5k/zy7bpVv2DeJ63bAC6mJWrAsxC+V5
KP4kFtKYoBFV0z2RIPnEB+cwo/iWoDAHcXfOYoClQ4Eqh46msHQFJ8qyLfN0VuDRQlnlCpaaYevO
OrHxUNRVjX4FAD6lsGJ6SU64XgjHE2PTrRFzMVsSNTaKcoawseGt9QS9U1Oe3ot4rzqHJOzJUjE8
C5zA9S9WnG3MvIg0T81M2yRuMcLpA/yVpD3q0waFLI08Fx3d9JLd6DbXvEazPEWt8ACD1/BQ6MT8
CeulZctCjanG6YgxfcVzN0F6Qsd6OuB4YKWbktrJWVjDEWm1BGmcAywA/dSv0OXPdl+SBOUdsU8p
GOiMufefCNVNu9oYpuxv5FeFi2evet98kaqmQnPwwh8Eyk3dHEAh2cO2mdNtyam5D/Rakb77FdFP
jgczbIQzEqySpZp0h2s2WrYGgYqCjcHj+nUmaqiAusFMFfkEwCdcIRIoVsCOIykfYtL1D/iLV5jr
ILHwhK61EBQwZpBhr8x+D10A4JS894J/CfVTk/Tg88YfDKNMvjMcyYDRJFZXwTLaJsgBnF7fnYjs
0qnHyHg2Tu4ogICMFGCQ8+qwV4HTx3UJ9SIlp16HFEinHDEwfsCK986bPkImqvvVBkPGhfXL1M5n
SigaTbLEeXk5GSio/HQTSama/F6ZJEoH7/IEXRkjN3QMDHcydu2SoC2E7HTCkREZbvytKZ/V332C
PwztqCz0MiDUrU4NYVB8HLWN49nBNk4wvt9tP6U62Hj9lpd5YXgqpS5rPw7QexjvDU/St0dN2Hmi
xI2zqcx5tiMnsM2FrjIhXX1AEl2uGJqN54hediP4TUPrY9drpniuCCz7uQ+HbmsTEIQ6SH/vH21V
mzB4UafQUS2Sl2DJXqxbDJEdMVmEXvTGsSgEPv5sNtILIzlENfc42Ez+1UYCxJkx6wbvDLHYrodc
GR5z8M+J+Aj1EzNPfZobUwQGl+1FyAlvg4OOPc5lo11D5bRRTMcln7Owvon8RSvOu8dVvv9rY+OQ
JKv+N90u3RoH36DY1W/W1t3NJ/nut6acQJcDrrL6Q9hUqtGPdfWyys+Q7Q6IBk+rzGVGhBdSWKm+
zNNjUMqkMphZ7X9akW/1RGPE+lKusW+t+7P3ZkaKfs13R74HYLSi0G+uevuo8VIT1LHnRgcmZN4a
fM/cLe6G76qVH1clvCnq99KG/i+bROmDFEqloq2GoBYrNQ2jYepPgy5JUGWo0sLzQQUrKvE7qbz8
mvoYKrnEr8ct0ydcmJ3oCb+1YaaD8LzVViBYJ+ltM2htG4KALtUpMpJWxbefu95c2eavP/QOjfig
j3gyU7L3hBCpblWa2cK+uar3BTeY1freSbH4qWJX+RqOFDAc0R68N90VR3lqYOI5iwqyod39riQk
hXEeJW5dNaxxkG+3HgpO+jRCPmLNpqy/xf5yrBzmJ7SCodCGpH+mn4SdA72kA2Ib1ezHqEXHTSPr
L+jqKLMdjc8Mkvpe5din8homTbDRhRYJQ2kSlrpe7b3UOc055ksCU7eIrs/ds5JG7Gayl5UQefkP
qAyFZCZhuSEVbZHYzMxyp0EHz5uovo+Llu2+C4QZt90EOsD4svC7BLjaVKxi/vE7AIQYdzBOudZY
T1RaZ54+GM0O0f4YNaDujWdUN0BE2blG/mQvp5qsGuAFa4qTdpUfQTqJ5X5x6fUTBKSoNJnbZ9SV
RMRAob7HJRXWLhqBkP6MSYby6SPILyRvG5oFY4xny4LjO84gvqYa/iJ6I0eisSx+fPwpn4LZ4hhG
NidLz/DXKftUCKnO4J31KytuX9MdkXAynOsWNZb/16RFeB6S8/4m6l1+tvQBbuZ8inZ/ie7qWa8+
NOS4EF0cKy/+4calwXRBy6dlzN/IW/lO/wSWVWdcH6XRf4TK9AwJk9ueW6r+h6UYxuLUzGoe2npc
MW8b7e5XgAVhvxAqAYlsJIQGboJByO3A2poRIkRreQgVUyJ5SC+0EkldUqeyJvH0BuQ9ooLZpYhD
/NvtZmF8NFsb2wZegN1Srp4ANV+SzEjlbi6aDIaHtZt0F4vl7abt61yOYnWgk3cxPqoUPsuDzK5a
hwTAWwy/A5gNIVadVO5pzQhEesOSTTa8rOX155OLn259f79lDTdDLv8WIUQEMIg61IC9GScFMN4T
leepZ/FNLPa3FNoQczz4UuowcInrfjiliPFYnraX1J0VYsWHKcenW5KJChpSJ21XSNH/8BsAFzYu
/5mrwiDAf6sQYrQEIC/usKyWmUUuULvVZ9xGXNb/WXdRwpyCXpUrmjFzwRPHabyJW5CI64xV34gG
dIrErI+oTQIvS0Et/Loj+cwORUw0u4bfHHEhwzyERSnx4QB5ZoEmFzNun2KCRt6x7DA8wkKhGsn+
MSgIyFRaOrG/IsGA7qb0hSZdsLgUSFb+BkgQy4YhASv8zthOVKfySi1fa9Vj+a2NgZuvCaTdZDWJ
Pj+VvhP0QYQEPFpcF4EIC1IaZQZVEEo/kjt5sUmV8Txxmwd2a3FT2It9bzWgkZO+7T4tH5M0XSYU
smrOZTmZ0yjzEn4OPvrv1M1vm2HB55p4VTNSe+anyPHLakDAt2SbBdXG7fz/H1fKaHSK/VlkNMrw
tKU9QQMOMRnCrucZumRVyidnPf/rS0dZCUbEb+2xI0d8bF9TLtW3sKxtow8sIZ2/eJaABmjdgLQ/
3pOEi1eEudVJdvHLIwqGvz0RL3ASVHq80wS2h6GGBINyhXGCxcv57iMixOD0aYa7xBmCZmmzBN2V
GWvAWP+Wn7PvJXzKoHpIXOd33KaRTxOvaeIsY9wMYdyquqmfnVM/rwXnF1X03cfdQvFFV/U506I/
28Crh8isN/69ir1V/E2WF8ds2N7F6dcOkRzvKWq5krnroJ82ruCucmBLbBwBpoHD+sC/kAQfpnNL
cp2k5YXvJ104TKyj+dqV25AE2O9X3E1lM9eE3dRK5jasGFtmglACMqo0mdquTcMBUj60t3sHBvuW
8vYYYq9jYJWx8r2W4lI8zXgFYqc4NCqlWtOXM8QNYu1mK5wOj3ZMpQmJJ2I+xiKw1hk18OAtK6z3
cPD9t8eEt0ClPyrXeVUrECrp6Cvnrew8KUiTZOvbWczQl2MAg+vKFzOj3JOjEJrHIK9zmnziLSM0
Zgm5GZ8iefWGcSUEWFbwTpY0EhUiDd0D7BYdd58CuhGPoR69k4X9FCJVL4B9toxIGT2lLbJRGFuC
g/0dPMQmGSn8vMpkR61OJ3TQ3yLiVJjJANWm3TRIMgscukBYYjZf+41fpV6rUdclcyQG9/OF7Du1
V10uYxDZa6ldPFftmxpN6c7Jyj7/+07AMqKExkwFU0TfDUdeIa2NmmrPkF5sTGMONWIK55wFn5Fe
bkw9rDA6EqtF1jUjuAnk8R+DeRYzHwfSKvnppv6DkKFnkDQoeOoBS1MKL63zIHG3phwqtS33NLn9
CMHRTPeOkzBgTfKIJLUB+O8u9LX+8ElKFltEfAVmtLK3G0sROiGFjLUvspuaS4veeJUesSoDOc5x
T8OCuD18dIJ6dwZg5qcIb6d0griUQI4Zn14jeLqQa6zLR5vVmNDgC/trROlka8UTJxgTjTZP/6LX
JE9yIvKEuu47hG2CoGLI6AdORTgAbQY/FdLRrv5dVPDA015mZqD5jk57QWUujCpkrvrjoDpk3+qu
afk/j2clJ9+9ZAr/wNWmi+PVrKbQwf4r1z7wJAAm7/6JYHEEGOJ//rdGh8/Kd/F8GIInSLPtbH8f
LGcvEtnVCesTB/lVa8o14yr5UEd8K3IgA9f7rLeUTexAaJFys3KvBVL0neu8w4kMxNxuxm9CTfoc
r/hJIIrxXOUgaXUXA1AsjY7/8t0jxoHpkeTf47VTLWGYlbK8VaNz5WIqGa/E1Hv5lvJftADTyUIq
3gZozFfltWvixWa/6UkdWY9+TTBcQ4eTiBZq9cDx3wAi/nHf6JHiJ6fFwdzHivaMuoE6Kc9SOWCh
znHuM/aaKNwLvqBH87i/pT3nYB65+BdEVDGhfcycZxXQuZrG+OxnxoMao96yDe25I8i4yOrYtsbY
UkQg++Qi3Q1/hNf49Dk3D73knq1FQiFiUlvwY5N7s4Q8PxpKWrlLRTxkRERh5LRX5R4b2MQGipN9
7I+J9tHFMsEOR/xPyB0We5d7XECOKsYUcYtrch3PIGhNfw5ft1qMj6Pz7PYzCs8fzVlAJrypOcBA
RDq4K9bvRZ8qPVBEZunwLxg8MFxkgji2WE9137ifCVXE0q7xGoDpgvm0L26FS6IXypBb8oEhXiFO
tTsnu78tC4QDUF/twXo+2msN04x08u7lonbcqMMbxpYBVvrN5FPh4vIfajDhQNUETjr9HqhTY/Rx
6R5LAOkCyCt0lcrmIOGYt93vRh7JOjAcby94CJ78OGgrFzhmupiLfqfEecAWD5+62G8/+Mp5ba08
8OcFZbwgJ1WdAjbeX4K1XpsDsnDcep8/ViI037KLbOwKjRNJcvDubEviEdWMkMHJfXXLhl3Cabir
az8RVQ6Urt/yq6m26mf7EhKueDDSiiT0En44t+IiKykGKdBOTEfakSabGPWrCZJqxtfdqfk9pACp
p/nPnsIRfWlGwCGx7gP4kBrhbk2I2s+xmyMQc2qQEMnAaUfhaWYHRjV1CbFxnIyh7smfDwaAEAug
J25X3zD+N2Z1IkiiriBgvy2G2lmL2J/fz2JAIRed4cF8pMSZtrHmu8i1sUJlVd3g02Ij+TeyTMqU
sc75h0qQ4IMYDYftMS1PW0oR0acaYKEwfVTo47f7Q3N9dK6l0C0htHichNRpA3B4QRXs3P4kx4B9
jcDU7wfhpw/6TG19DRrovWsqS3FyiACYJ17kL90ZPBDQEboUhY2iAokFgdZmI6M1tcMNWn2HpAEB
LYGkfVL+PARVRXsKDhNxWLBwPgqFMIiGVDBnwQ/ps+Ni8ddy5PiBWyN2VyScF71sw66PHT+Go1rT
6qCaVvkeJkvIyhCbmp76Hi1ywr1eSkaPSdLbNcqohX1+3lod0FEnAno3BgXklSTFR/J7OeJ/BtDk
PjPkGBiezH1lovbK4cwF16FM9UmOgbWxIXM5Wspl4xnqdbODCCTEI0TUvddwzb2koejcsfKzb3NI
G4cpTv5UlwZONkGgWR7zOMOUhO+dPBSxRBejz1E2S4LMKSXLl71s4bOQe83po2FhiFtBEV4XO12z
o7Cg3LnagRJsuhsgOy3RAJF+nqdOkMpNW7MHAbcLIvsR8U29HsBSjd1MBWe5APweaB7BdiIXRluT
yu7fwdNVO6hJyViA/BTPIIZ6n/72zvPuQZ/xUszIF+Gkn3h4hKNNN5lYTOBKF6+XNnij9cBmLH+t
6otc0cNp1+wLv9mioj4EjuddxlPwmJDhW6J7hYs7LiSKdmurx6FyTc6C4kZosoSjpmbAK8DlOQh8
h/kTxLO6djGQG75fZnyWkbxPFW/GaDJp8d5QypFkb/pnrijlu2UA4km0DGaPXLyTy+QxPDp6YMGt
x/O8TO7qcFiaPSg/QAStybM+8sHFXvtcw8Id/KuY9/axiubaoZzT3fQ0MWkucNYmw+oVuiI4FBvb
iNe33qRAK8pF0R8JgpmBPCkRRAjLOaGZZC2THIkT26BPmxc9tRUYE1qQD+WceEGw6cfbiAEUGD79
tn9rN97F0OXYQuVt8L5igU4z3l/mywHUTHBPSLPRkOiidchDH9phjkcZEdwZa0lFr8wiUej7j4jP
RiPl7j7fzlGvHxL1yJaHLcFIP6qbsrs8gUI/q45FTWT0f9p6bmLuPVlw+DqD8FAEC5353d1ECpMl
xbBuEvJ47XmNSvTg8JE4kTW5XoioT9ySoLSgE1+pjBDuVWljRp27Brcb5OLPE99oiLv+4/29836r
rQEd02iHj8N6L78BHy/eR5N4DzjXEeDuHuoJwon5OJjUcc9zKIBCUFYdehfziXzJ2qqN/f3vewzI
e4sxjrF7myFUnHJSB8/asDC+eLFahXvvTSeu/rxAgnJUq0XYzaZVr0+KSgN6kdjacReqC2C2I3PN
B59S/PK80C38VTUbBGf2GDwF5cheZiQUVtDg7tflDMCajGqOMA2M8c4Efk9VD6v5px4sYxai0w2t
dUHMkbNMjIqAZtabUuScjimD4M2hkBiy8+VNJAE8qDFgePSlHSnKM2fan9ZzHLDa8lwWFFrgLqbC
QXsZqL6s9Fn3jKxMu866IYidrm1fTfZLRZpDDQXcVR8WPaWAA7vtzuxmrax427X8EuhLZE0ig4xU
3v1r5uI+KKL31b9IQ0nLfFeyamnrNzJKfCCDkHKPvKo/3QKm0suOWU+Tbdmz/NtlxB431X6ARFeZ
afykgXsPZWit6CHXYfyPlywBop/3s2N5ayhyfJFk9luSO5x2Ejx7Blq0XiHtzciP4lQMLogxA9Cq
sA50TpXcSE5Lkr2ITF5t08+idI4lZW56rthuTT//+Se7Eaf8XFNBT3wqE+Fc6paoNcRsz9ss22lS
j0QL9NSyMjUSqmvZ2U05CDNq+psGr2+gybWnQGttB/AgQrswCEAw2VChKdaxSfQ4PZAPmKOF7zWM
nLF+sD9vjUffI4I6RbFEeMT9Yf1sXNZMUr+KCAh69RlArpuIHXstjDlNo5yZ1Mi2vEkXoNTOCJP4
utyw42TFUGIVTPTgbjW07Gch+WwV2UO7oiEqKNYBvAMQ/s0f8ioGz+bj0eHR+Lw9scsOMU5vGa61
6KK+u3QRk+Bf1CoAHJ+mjtNh/asqmj5OHoSPH8Rl0YG0LC8NfRMmYQZuul7Xfss/InMtkG5JlmK/
6Kh8FjEl035gjcwQCXxquLNbBu5mO0KJRFAUvh8FOu7H1VSshBGNq45x6w/TGTKVY0QoAL1L5vAd
/rNRUwFktBAI+c7svaNjSd2/MxrVFjHjjIzv1gFRFbouxQwkvx7YimjXOP4sfzdgbarAIlgtx+82
AF5TGqbB1Ixbuwj+4olQxzjLlfHJNu2+fuw0fIU57sWQTVZg8Y3eaDcjd+Wp/Fby/EYmAbrHJxys
T14BOdJYviwZOnDdzO9Wr5raKFh142jhsiw+BfbT8NAvQMV1+uAOJ1wKuVKAbJoNLOd8d8XikSdX
QCqUKUO6cEYazyfR9BRVwg3Etl9gLw6+Rf/qwkyhJYJ9szepQt48CHmr9oIaT2/4QY5x3oW32sxb
MSOdaVvyDxZSrMn2CpVKvWH/SoQpnxOrdRCE9iFCwofF4BqeWHQIyriUdgpowZVuv23IB2tMo0j5
4P2jVbsjlUO7zqMdSzXRPygddk7lgU4SBsvhC1ejgJ+XHbZgp85fxKaQT2o7B5z0pnSFfFUJCO9S
e4L6ms9gOS0cUyziaEgEDgoB3e6Lme35O7d40CbRH+EV8OicQHoslBjhpiWNh/HIGtDZl3y9q1oc
NWWWxWkMcnidcFlpW+PIbB2e2W0Fd6oqcAxAIBBnEcZNNNw1JmXoIoSkycrEspwsogIEu3pWgEHm
SkoZFc//C3UDCEIYBD2DDwcoY9JqKjzbwyWIjZt9cFNzs0LTNjzV2NVnbG2vs2cd9a0c2d+VzwA2
8RxgceSnO8q/g611u8ofEdNfS4XjY8Enj4xwublZv4WemAe3wAa8viPkPqAzG4xp2dMnvLvVI8rI
V0pKxvCFymA7GCOdOOi8Hq19HL6r4OVv3qbQe0P1L+fSlMMazCWq000dhnY2p2NMug3dZmrrXfIc
S/T4U+3L02llcitp4E+vry+wQPmexaZQn7UcsNl0HbhSenMx7jVceUkl2x4YZgFx6kfdHF7pa07e
nxdAQbHkZGhzqDbOWZiI375stTsyY67YUa6UOUIO9sXscASCnrWzx6Eq9tT19MTgkr0r9xdBje5K
YRZZfzGALEq3aibFOAdJJgcb8L2BJFo312CWD6UTRt0SOgJvlmUn9NwN86C42LR8wV/avSpExBI7
KK/PIqc1CiHf6cPA9irtb2bpRW6V1uj+ko/LXrol63NVuD6sxxGUJau6sJ5gEkO1y254DKRJK2sp
9mAyGrDvTpkqBmvEuggRPDbc9l9DKB6pGh+Fyn3OJq4DWV/FqrMwEp6WNZoAk6BY9t1yXzs+xxzE
hbTHx3WCjwqsSUBKjABPueZ6KV5E8LzJ4aJfL8oITAvk1KPAVsoHe+UdjYaaSJYwJMIHQlU1dg8c
Y4nrDXrPmoFAWDjpkrOA2Er7I1LvXqfQeq8kGEofVRm3mKN83mZjaokoFr5FGSFCAA2thMpVPveP
n14qhx63JSaRjcn+vpXtPWiSO5D0q6Nakjgi5QE2mpD5VqoHRzuMkKey8zP6v3PZL3BhMTyGYSaC
PVGoW0BbiW+NmaFlcEECqGITdnuBw4V30FKnjfpGzbkWv35BJs64XK79IZQNv91CSEDZvmMc2e6v
28kue23bt1Hjsocd63cvAnxy9xlrdKdwqFYmdiBYxx+BxeVVCJ4xKQuSo3HiBxZz6F31yi5qNv1d
c0zHycvKTh4qSK4KIfot7SkTiMfKfscIM93LmPfTqAE1ESmn0s23cemPeK+gju/tuwXc3rVv2Jcz
tKTQ3IMslIi+GuvbyBfsidaIxbaUPqZhYgzTJomxBrZkklXu0qSbPkzlkqDWWxV3Ly7vmy5yAr1M
6IK4NrCKJXiOI91MZTTeSbp0okfjzwRXGgAR8YKr2K7Gjm/w7eiTwd02b6/wwfx9FFDfXh6hLu4I
6KFpa5yXpZl3KiVrnm6paOW2328iVcexhXke79XV3ja5oBEijoTfNF2S7XntY/btKhsI9KN3R4FZ
ww07P9NTIyjuGKbtw1S841cJdAmqCjP072hcjrqW+5FvAdpP7l7YppvlHcOojxkFqFaMzPFCZVkk
/K0QUA7duj8+6hNVWDU9vAyjzWhE/oeY82yUvXltrU42gmCtxt8Cn9S/2KUeJeBJQbF25HnV7oqD
+hit6CLgre9ipFyjh69z+lIdVwA64IVr31q7PGUrQoYNdA0qgA3Oq7axo6OimXqjHokDVeIfMi4A
f+SSWfL2CVnyyXqr6UoAbaPCHjLz6hp4UeA/HJszfQZfZp0PlEhudXjk9XRxaGDRDdJG7MPnM4Gv
eE5AoXglWiu8g3eLssYM360fzdrkFvfMDCToaTOpwzy+BiBo6Ws3RUbQjvai3MwEGOtapcIpCjk/
7uEyXUXwexjncg+MFPVwrBVGT5SNmteI4R+ZpxHS0n6Z5b8rAmqQ4ypu3nxASjvwF65L7RXOXz3i
HNlk301pmHLzzEnlMrqgOCD5S1cqY/cMx4k93tnEXTHd6hRhLRptYparo0+GnsLlATDZyZW+3opl
HH1MnntdAd6iCjYmd/3ybUwCuIyofafPd2VnbhFVYB5FF7j1/doqHOhH051NVHGQdBg6juMrdKDS
+H6bH800ZONCOShAVtscolEArUBIdao+g/JtR9oL1dycZidNWPa9qtMZIsB0rYqfFzbQNlALwpVB
upACTTkXlZ6tuqepzmsdsvlSkVTdz6YBXZhENl0eMsa4g0jKnTmyM4Yc9XW0lOOBnl1iFnOOXr+C
+e/drMluGr0KZI+mduwq2HoACYueoeCXTvxpiQt8impfWOQQSB07HtGj7fdft39TyxDY1zfsWySg
vaXb1lVgREwKphke/hKFEupfa4sd2SbqdrKDwAaUXP9XQLlJ2wzCgShexx3OfrKZmt576T+Dgkvh
wfc19o3H1/xWZuQCN8Zu5qVwV0Jk77DOKeOzvNlXteFYftBoDHbgMEVunk2K4LVqp7wPQx3lPif0
Szu/Whnq/ypjk4SnuDESHo0r4RUHYz9zEnhIinMV2jT08QmsA/j2Sri7MAFDfaF9TLZnlS29+z9T
AHCpcGI2tabtv2I6VSKgWUs88VPdOVhk8sVNWCF4n9AopqMf3HBVI9Ee1++aVoZ4eHtSGHFW7d7z
YhdVcJc6lBZLzn8H8e6NUVDlbIdp7MwC0kLhhKcxPhdTRjI5xNnSebXEs+ogq5qWfSnvLqRm7xQF
OULUOagoZGA3TtvmalyLFCr70ZnldFSSN+w2pNgON8Kit2g8COw/wEaL6BFImQzVyFJoS8Mrk3j5
fqTfeyDeiMqZ97A9nLlI/6ee6eifrYeVKcRyI3mMeR71J1yfs560SaxXR0/Zbipbt1BEXzftFeFT
kRYqbS2vD/Nvk3m1XHrMSc+AqJktuzl18Lh4sUZ9n0mw1FpmmCWwd5DFlB1uMWo6w/RtW7uiRQro
lhkrrSdADhfEqMRZwpjCxGn39NyKDbdiZXzMlWb2p+t+/boFHVJPQC+IM92FhtQDUJSYe81epdGU
5HxNcUJlncPYgNvLpuYZRuOUDjaf9Lur16bOHrvQp1ZXeDJ1HjgRa6B70j3l8BRgk1DR3pXb4fXB
//eTTUxiMFI+w27QDvGSAaMydSnqzyMl6rkAhHBQ/lVsy9vGtmDaNh0PYOw+GbFUYYx3oqmd1/MV
lpdh9CJo/7YQl88yOuFajPvylJfxw7XCfi1oIG9WPkaejzUf3bwE2IUnRZdsFSYX9adJOCoVyFh0
WPgN5TAEfnuBOy8dfax3cQ4+cJ70w3POlTJw+abL8/BxEr4ZQwCBLHl+diVotpyuV0pVKSzyBDeV
3+2Jl3AaP0xxYUaVCOzPf28ccsCcqOHHqyNnvK/pwrc7BFgo4/e7jtyII7lp/1KICM8mjN+Xhmxj
7LG+ZuXeaioHatD4HSa5Do6ZerYnhoWtSGauUPRHiqSkUIHMSilOY3/+28Mkar9J0py0pLayd95s
zno9fHscaVoKWbKlzjq+koXCINHGvZMjSBhHsaS649pekgyWjmral+PUA4iL/Gd8x3kAYQ1LiJgm
T3tDImUJarLG+OYJJa+VdzSGkMW7ariPCjVI28UGbMYrt4MJAh7RewDe7W1paOWmAos/uDxIY5b+
zAMGVKZjhIe+kWpM3zM727v7Na+sWTeEmZGS9zV/kXaVoVs0wP9Umbyk0WDKZNFnqwGWIXY/5j8q
um8axHM5f3x+WLa4vi0Pox8eT11AjRfRGcXJaNH0iVPsY0SHaZY4NTJkAHM8lOTpGw23unV19Cw5
E0qTzMcZjLNbnJf6pZImFUgdM9qp5UwmCCvVzfUyTrWQMaMNsiwpQ1byQAWGbmtrJEGntgc1eGl9
O8MNlVMHFBmvPF7Z2erBzmCc+TugswjUpYL3nBJjGZjP+aEt2yYVBtK5Qa5FxExPka8/t/NIcyl+
bN/Z9ZfCM9NsYFhTOMRUuf63EGlARoYpTh8q5ErvBmpLyhgyRW8LZXUEpcSKoLkPpaSixcPgg1wT
czTWYDDE2Q3cedzegRVGUYHUX1sQW29ahsThydByH0zx9XweNiKxPRJdABf4MGvafTSoMM8X3vAf
L3uVixRv2uR1R38wc9imaja6hk0ExHRGvyDbjYAahsjFi1FBty9yhqIwEt6+WBtMJX+I0gDfCVkW
aHZJwMzSF+1XMwqhf3aOurGAa4FYs3VIzTh9ZPoNEZ1+CzeEB8Vh4kqO2Ub0+8llMaQ2+DoyZwuJ
DI8WRrDvNY/YEv3f8afQuI78du4QvijoQ7WOS8zCy/T33xPrhyzsyC74dyYs0m2VXAHTl77xCDr/
UvoUJmIFV/cfri1zcnct6nPAwbn7cTxmdv4wb6m+sXrH1bwzCrHcmfUAROKuneCldm6ZNktFPVA7
O34aumuEgDpQSVMq+imT5Eiaz95Edu8vQ5zssJbiaDMqFEZlKvHe/K8FsaecYBdvrl4SKKtN118N
RP79f2Z0QjHAy53DQLf8AuVPdI8ulVZVytH8Ithc6lwW8upYZmGrCTlzIZJ1AnGdz/D8It+d2oMJ
N2kysujXAhUa6dNbCxjBG0y3YFq+onUW+2pe3HxOYRe1qPh5IaODlrzeUMK+MLban0b2NeaA/SEB
YqJYnVgu6Np+fRVRnSUax/2EYBVM0yCX8Hy+mHbmmBgJJo8NSsB0KJDDoF+Vt5T9Oxb0WtYT0NFj
f5jbTFguIAgo9hWJhMbM3kTF4L/V9Y96blMjloDNjz1DH7vv790dfxEMB8nxI/zEeDpDGcr7u2a1
d8Pe4u+aaceGQdvjxv8IeWciA6eAgUKv9LvWBjg0hUm3Uvb94hA8tQCXvfRFt3+uPuitsmbgpddX
i2lwC740Sud5NlWpeeErUhPb5Xo7akPd5LbUVtfLysvV7EpBNhGsbcaCDWExYmdV9V5XsRIzqPcH
wTUlTnXv818pCtzfdtYGbby3EtLzxfLvKtFC6gFpcbS9vdFV+0HF690wPIJWwXB28ydJ6PYw/lhk
19Y4beM/9PoFNaJ6o/u204VO7EQXcsXqVHWa2J32QSGlEuBBPa6HrE9FUcWPnLkXrSLCMLAB/nvC
0RIpBZDd7fgGr4dOi9z88bgFzOjB4UfMnw4TJpMBxGYzXl9Xl/FmuQBNwViNySmzd+ESihrD0m+i
gfTgVedKwd69IkvaTaO0A7Q0WZ9nyebeD6YpWgikegum2v/UKfPpRulrLd3lMr1VOd2raqxlodVf
j2eQEhIiWwsRM+jmJJPn7YQtwKpoAtE4CotkzvaEjS9TI3AxqaHHI9gzrk9dGiSUjwjsxeyb9eHa
Wwt9DoTBoEsATXnzN1ajf/qzfJ+eXFLko/BGVGNdkfrwCL4Z61a0lnBBHKfC6mSSsWnMCBUvyUi6
djAFxsBesPJl3Lw2ICS/ap8fN6oyqg4UfA9nQk9CN9FFKXTY6m4qZbBfKIZ2r8fqRw4j9uMvV7PS
c7O2YHztgVXmLmWtKv1wG5NXjqgOmmTAaYW5XreicXgR2F6Rb3BqypfEqB3NMrLFipQq/28HO+Ga
DbF5AWfdashp3hcvLihRyjmoFv4hSvDDF/WD6eJiIF/riUWRVP+0kNhszRLjC0t96/uwnhqdM5eG
lCuNKeMS3C0KRjzdGYl72fkRi69+C5SqInSx3SvIP0v2OZoiBEqiYR8BOzqNo2HrBDQWTuEiaASN
enPLvaGcZiisryoF0+hzoM8XWodaqVPj94U/YlUMgjDn52B6Pd64Ip/5AMz/KEGeP8+YMgDNP0jO
9wLICRuw2lU6jcJ7x9RBcvXz/FBnH4XRz/1PNqFpAHvA/VjkGGIOJRHCxXMZ9yadnfb+iHTlEwUP
1rI7Lm2ASaQ5UDDtzFCuGu+EdAM6eQVubkz8Adsh8cb/nKceJAbHC5NmQZznfmUhOFn05MqTo5wL
DalF7u7K4WAt5ulQCiDUoM4H9k6h++Zbr3Rv7mA4gwsc0QH35l3TbVJzGrp/Wodj0QO6X7JpCiOd
P6k2DE0AHWzXYSgdTeL/ly7JN3XzTNvlezI6CM9yXuGpzqAXkDA1ZjByriQQOtFC1s/TQz2Nm2aB
p/zfGeEqW3hWlVC2p6qB1OwQVDAoJ4MoyQ74lTpIycz2UsvPcfllQfhSCZ2AEONJIKLlHSCmNivX
IH8edzTzraJEdtMUTPobylFW8CnkmggzkcWJ5M6vjZCoLHL3QEEryGz1umlmsXucYWNwnqcJZvrP
ufHN0u7SesdxPmCZ5+D0sw3ED66NBu+aq6BYaNqiSdNLv0TKWnAW8OrFItaIDBkAHVBsrY5cmT3Z
uNXrMzyy4J/Kqm1gSEFzL94scQkkQsB5xm8FgzmtMbfV4YE0sCoR9yC8Mf7iUTla664L0XbQlXHB
ocYloOYk6VGMbbDO+4itNBdaeW4ARhchTMpHoOhAc8aVvqYHX2pNDIpPjIJJ85ksqURuCTkoXdL8
pr7iS2IEY9Qfpct/r1qeq5CGOV3pfHsSupWh17nfhx6W78CLDVP5jaSKaM2VVXQ3elu0nm1f2Y0e
MTrkfVWRiHGWP2GBHhXPk43rnpIZad0sLLMmCv9ud+ZusuHwBg/l0xe7PWYaYZLDk5ud8lIp1U2J
cjWXboO96BJaUC5ZLxalnRPPmwz6y1HuE/62EgLjgmSrgH64z919XSBdPN8aKA0wmIBOh/+gZzj9
9JCwDZJJCdU6KsHARAA3nKdcCRCz2Q5tK0Gs/dfxCBSbwGvFy7iO1hPJBG+pmEBWyyKCoPc2Hidn
QFz/EnJMsxAt4I+NywBZR5eTIVw0u1smvfQRnHwj3S5ZL22dysKhSkQkqA2af9b8qVLfwjJltT4z
52k4OzO2G2t0r91zUWrCJQmvv88vvAU8ub+gQ8uUo0pEllRWgYJaD+geGf4698XbjRrckk2/BRc/
UFvp1mnG8WRR5WG8SEPN+x/vuJc/zAYwbr5JtrjbVgEqCYb8vlr+IyLJdCOMlmS7jq++5MrOeq6X
jh5xpHGyG1vCB/Rau26c7yfz7i6MNs8p33rYgZx2r/iNnt7EQRqm1Xxr9u0y0tT4sKeAnFbx1wLt
OtAHa6efunVJKzQDgPdpTPzyzd/eSzfPmw96a9Gq9a+FB03fgViglQqo2YgO1R0HS2GXnRewXmzb
61+9NcInPD9TB89bt2zecfbOvcfvcAIHCIwDNl20BLIGdKfcnw2sBbOhH75XuOZJqWYWI4qbc7rF
NLG1FgiBIGRbwfFiV5LmLdxpnBYL+TsgKmyUGfHFaao7Va7sqIfHslJV2JPYRMOSxWXWVKzlUSMl
or72ZOYoHLFNk3ELSbDwniEv95iSf6sW0AP0ANJPZD4rkWmM7yriif42U5RVURZSy+JSzOuqX+uR
NxdRowv6LRHTWJy9ytzdT3S+uj9PHT6oKBrIEncnEaewBKX9Ei3zDy0hryMTt5iKfUxl0O8PTr47
5DmRTcNqGyHtSrrj5MZ/hP2JjLCnggu8tpjF2MOiluQspico0AMitnYu2KDPQXGpk0ch8O/BE7wG
ME/t0yn4Nz+MqCExtcLDFpcAV52MzZnq65/LMAi8qdDuSbs41eu06fFUDDfo7yszxh8BrYpZTDee
FjEbPrXjQV66JK8NWwSWMIAJ5mtYexu4zA9WtNRSoU7uy/j2QJo08zbBO1mG+7DuuKjJ1F6Mf4eL
/KjhMzeC5Obi1Vqayh8dkyRDAS+aytkKujDXWsvDffpUF+hsSKgT1P2Gu6P2kkPQ1rRLDAhjKygN
b+kCAM5vfGI2QWb1OTzfeVE+fQd4DHXxVbuwTJjky7He0EoYpaiWMvj+8aZ7osThVJU7EZTTPNqe
z3JUoqkVeK58zj+czwwfnHBvM9RtdAg+h3JnDWgEucSLNrOWmsoz2lv4eHfGkneCP/rhr3GHbx0o
e1ERXKeyI0yWeyfAYhDHLi7+NNeDobbllzYHMs7fxZ3yOeHWgTndYHfpTnVnRXNU05qZofAy+TGP
CdI10GwmKRk7EpumIBNBNX2BixsjUxZEbanMIveZsiAI7SNkLY3FXDgyz6y0OWh3njS2eLQtZ1D4
WmvfjaFw1KoX5y5KpPlzVKN4Tjz3jc2ycY90L/v2rbZ31yMSrUG/NTnGPChGO6tsQviBfBrx6wcM
sVrGNxMUFpdf49p80BMnDrjWLEgMJHKSTI8PQ+Y4LmQHNBwByNbFQAUO3nQBJosb42CeEMpAxub9
nb8J7CjlAdtRJxxTdkIYMOogBQGhXtel7uEsi0CLJB3bUgV+5Do24RJ2QVN8emWA3azjHhqi3lbB
9bczGenP/Td+IxKETYktbtznuqA2MHV9yA+DiS4EXiDVGl56Pd5HaQGcd6YQ/sCXA/kUm6KJulIW
Ekg2pJvSo9y4RxQ9QKKZeQslfzpb9yHRldMZfCvLQtCMDK/2rA/sCAYKSgQ4PDXFAzW3a7J/YkcR
eCzeo35AP7i2BV9GnlTFDCZJFFNmQl7eB2/ETgjx9mPKQO/cGwYNPUp9dpn/mGpSTt0I6k8kr5sB
aqs9GhJ/W6z5sHSYbR58U05czZabIDRLKQm+CZh22+Y50ghrusygjRJuujWjXan0Kn7/pVcf70x5
D9f7YWkF8tqxH5/T9PhY9ihdACAGfPTVzTClanzHnigH3CBEHVld8BnJIx+99fntIDwpw4Uhd8Bj
PngoVi4Iw46Qwp8/aZZzypaW4IBqcOfPTpAuAJBw5iH8AIMu+KU8dAD5hddV3INZRIrJwnqkvjVO
RWAvnT5K30v5462pZNQc8Wgix8Eu8V9oKW/OIVTkh491gSKqMFLvohZ7kg01hd84BpdprK1dSpNi
+nTs6/Nr3UZ+fnUerOwKUkwY0C1TqZ/aOq+TzRQcHLx+B+N5ed/Y3dhiw5Idt2J2bRkCBbxUzjiu
SorNH1NBw4NZKIRO5ImnOs+sV4KkWDH1+UpdupYZEF5HEw0GnsFmJqWkmD72x3x9byldWGFVXbPb
ACag8OLuGEkPAdiNgwOPp46WEzxdov68js9x8i03HgwcZW4NvjHydbt0yvp8nGlFF3Jbk/EHk3Wb
gxVNPFwjty8ySz2mMT6BsoDXdhtHPJc6g/j3A7b1ItRv/K0cKKYoS3wDUDbKn2I+chRsmL9yj2/Y
BV3rJciAT/fZSH449zT4QAIDrluE38JI5/rDu9vhxcwHq6XAhqZnxgnq6e2uKTFVKGuec6JKVtCC
4z8nW6NDPNkxv9Lgqux2jaZodFZKgHXObWDmyboWlow5e4PGYDnR7INyEzPoOiiI+Xqc/FJTAaZJ
KyMF2d70ZRmz9bDZf6tVB7j2Pwg+RCtAtK07HphbrLzSMRlWK5nvvqVRjHtiJzuUWxqcqAI//1ef
EyIBxv/8xXfhXpdb4W3wh1H0ClK8WIUeIMWeXuY4vrMNZqf3QD2TfNNEnC1CqVTFNGbTplXiyLvN
5lKqjwcTDINozeloeq8zv97AhW0p8x4k02mnEJsPa2hPTB2Be8CnomqvZ60nSJik5ScGZlVSSgR4
pwSu8ugQpvNfDppM5QsLnuC35ByrKb6J/glpMXAZMunND7nWz2MJ1J+seKhyOsNshV4aQJnBdcHu
/W/IDQ0uIFA9afplko76Kbfvsgk+ivQrSw407aXFM4Xv9Q1L/E9ZfBCB4GGwc2Mfhnrj6byu9n+n
xMOXsuFFVXixSC5fmvbzmEbQLhKA/LKCdvD7tiGbSJEzQz/c/jke9beK7GfjcyUWEut9bqpUUc5s
j/7pmsusX/zolDIBNwDiMjKlGJcb4VeX0u016GGy1fX8oWAyBW3cCqgwxlImqzH59FAjQ0OQBS7t
tPKW1lMo6+TOo373wBC4PijYdiMsHjV60kEass9MNhTlxKBs+or/atBFRlRYJmj4yOJm6ADV26rS
2nZASzaOiRvvkYVkvpil1+73pgQRTpJpnSCEbHcrumu5S0mC6DpYUKEA3egeOAPg8FSawdgQ7Ws7
k57fAtZvYi+No5TN9qUPsbjTUdjH031c0selcW49Ro2OPNEZPa13ruEAgtGG/pZNW4yEoGcUHHbr
JuyBNJPfa1kyFPp4hiyQUiG9xkLTUlzKoZFpQTCyrT3jpb+Zia6cZROijqxyfV1KsoysGFB5+xc5
8eGk9LSKmnZ/+iLG9/Ab/Df6DYxdUij1AepMEXbtri/GbE6BK5nXChYUkFFimy/YtylqIEk2ylCC
k9EM6Iqo++jSaTnoc2TkIted9HbhnmzbLbb3TCOQ3axL37hro7fTY71dlTTkrZk3Ob3v6Fzfen98
wi3uzmCzzoilm95ZZ0rDDL2ouynMkOgFR3PlSZciwi72sQS6rLuSB0rxJfi30iMKMv91UHCY5lyn
zuXsmJzisg+ylodUmSX1LLTujBsQrleh1GSoMziElw6stXD0huMVUDMn33ulCgoF66Z77NHuTsVf
UwgpVPf+GKM7cwwkBH8LV5Fi+pViFCrl4pA/wBC0pkiqVgMnpOcVAycz10e6zF2Cwc5NVAMm9V4e
4qKER12wpjntYsuBZbyHI93ijUVapAjMkpXZY2/NFeUCXJeeUbtHFessyId11Jzaw1Sqk2FXVlCf
3OXx39BUnQigA7BRIy1MfgTNKMt1ouX3rg2QrrPi8xAwGR7cSytXR8sHv7bYj56kedDHZFTpqpSs
2LXWl8yLdGxkNn7jCSljcxI2T2Rv2OwcXPZPxE2wQ2tiXASbIv7viSf4seZbRWEs3NixfbDQ2aNB
jT/Nco6gAxHGoKYRBF2WRrDPpNKK4xHf7pP+sItaHkTTGyQpRHp4diP1UXE7JJ1Oul+B5x5wr30Y
k41WIm1O9FLIE/3GKw4TIM348kokqc1kp6ppH93gTAINfwPX3eZH9GEDV7gADn2QREY4hH+A8aaX
EaLVouo4/fu1Wq0kpsUC2hEf+jSq2bBq6nznMC725K7za4bSydx9iirfArY5phZ982C6SbANv3oS
e6yb52R+AbZXUX8cLSUEqKjBRqJ6zGR2tLv5foRpBInbocXV3b0C0NDAdIoXMGSdsZc8+OUatZLk
/rIpWX0LnhESE02xt8nQ//y2Vu9SveVgSdyoc2LiXQXLfpj6fSeoMTP7MzuG6Lq29CRFZ1z6CinP
VkE3AuWJCajwcmfWQQthrSa2bpyC6mL+7podxsXoZIGQbcQErRGztFm242T+WRvfsx9NC95BGqeJ
n02ToQ+chEl1t6wseGnXzdWxoCQSxvpU23KDZmCaFcmWNVJmQe+CpTkazXDrtj0mz84Xcyh7vGlC
h92jwMbUZZSkoqaqkm3Q5cjGnUejyKQfwCFnfni1/+u0lyU6Jiq6f+h4xryYSAkwwD/EQCJ1p3wd
dqHy1s3sdqIl0K6puaonj8Rmby+Ndm7PWZmCVM1HPvN00JQSAyGNelNKTyzmxhKj2Di2r0t9zAgP
pY9bz3cYacJjQsoMocQZ1ZPRofMBLz7x9/7z2bqqgv7wi8TNJHswVD/9sR6alfdZAoDHTkeQxOHg
QWybj2rDXaCbdQbwYqtVQIErvgMOTxGQGIC6k+F05le2dut7HO0RvJ4Q1UyFL6pTel8xYAKphXHY
W6vPY3C+ztgT21L4IzDsa7CMKuhUg49xjqHxE5naoL+mCDyweprZYeSc4ySMWzJrIrvp7K3Vm0+d
pKUCIzFM7t/u3PgSgqxUboqjM27jYWJzbVGePdA11+KlN8SkXP6Lt58GV1H7NP30b1F62ddSFbPR
tYe+8d5pYBqCwwSXCzsxBBT5klrEFpYmqkbJonX5YeLpWMBd+M1pMiADlMxpMuMqRKExkKGvY6Wn
2i+m6ysY4wfqNdxOW3lw8pMrzchCTaO3HwvWyi59VsuS75vapU122sr7pkVArIkDYiXqM6PdpLuu
CFbEW1ezRViB/OUqBK8792+rJmhOIMQffObtf0iVyKdWAoO4zCm1Y6eeepJLGbGjmU0z1Yggp7CZ
0H1EZIWPzVZJ2DcTyxTLWq+AGw37dx+ofBLi5PW9H6tF/0IXQhJTMwQMxSczkXUaw3hZhMomdgSZ
jigySl3c24igWA1CmIW7tB0XRgCV2pvjvrPxmFN0mhIIL4BxVmR8pZYmBFSsNhxowsK057jNlOIt
TXzmOT1Bg/0lUmuoBobJ5pa9vGoT4ytygVnRKSHsdCz0TVTEHYm+ozdcwM6P2jIC0hFLMWBsAXeK
1SbXzEQgxF0OSdxygXv/SzOcf4Oio2DqKrfnnUrrWtDkJKTPrKnURRL1OlEE4s1VzKEBV6mGjgx2
/Dy9RVtRQCJOse+MEe/WUtUDtvs2QtY+wAUSa5wtJyyha7V6W1vxtmkaCYreUA9evZ/X971joSSJ
viAk8TGgrqK1k7PMOBgLpLSW+MXxaRv6AqDt9MkNv8AMP0vkIQ4KUb9fEAfsy1vy8NcdpvZrnfpr
vZELQbdA/AVKc3wwJjpEeR2ghW46FgqEDdukXJbL8od/U4mJTVBnShj/0BF9ooNuFOPAqI3C5One
BryuOizDvY0CyjWxR7cHo1berVV9Dwh+xGkOqNAotzFwAueVPPAx/uAWWvbGkFEXpcTjoXDYxXse
gqJwsg5/hJK5wiBdZw9NDVE3D8gN+r3hp2njbVdjkgXpPZzIYTbyUc0kSu5zcVFzQ53rqHTA10Rx
NAx/bnO2d+++YUxhJC4HN0RzfCcfYbbj6DRBUP4DiCzKCjmszaPjnLfxGjGjC/vuq31uIpzDXovz
sTuQR9SOzmmw/o/Kk5Tp6mHksQesRNZOpPKpwZgcOAimup/POm0mTBu/jQGmn9mLG/ZIa8R5DnBl
17R1V14vp9un89rH5bRePazW9qwnENOk2chS6Jctz0TY1sjKQWCj9yJ3DrA8b5ZhX0iX3DUnNzUU
wOImf/XE4qIFvxtHqXnz9LkTLJvgdynh4KGwGtAee0EQWUJeGTFD0I9mPM6tuDbLkAwmSV0WljYO
BdT1V5sg/cTDuTeFCX1OSM8P+4YMkbFjuqZRarA6lVsTnuSGgbaX2Xk3U6eTG7J7RX0hYhPzglFy
TTpiJ/aN3e6qDzKu5julm40jRuLsZ+fZOVPwMWAJibzx7qGBvNJGLprHJro8fQ1Z+0JI08zOLPbU
sRkhG5AOTJqgVLR3N03kpe9tmHFfLv2/f+uPhAUgmMA+4UlgXjOF/8DeML8wx5sOMOHuzXm1GPzO
eRAPCo+7UwnkhNKam6GrrwBiN3D8u8l7R5c0CSqjE/GrER+76UKBuLthjX5ZPnAnk8zYucjuurGy
/Zw0dDf6R28QiQpfRe7dg+XeBBEskX/S1MDhW6hxxkk2qUe2izFLYw+jcSCDZ9tncav9/dRVFA2i
aRxk9D6D2BL2gNi3FXOE9804Odl2KzGThExhLCejFvviaAb35dhpRX2QL/n6+j42tWYHOTTFe4He
LEgtoBZh11uQDSGCLRGaePAMHOq2zZp7FLXvnkxQjRAdKEe+Owcwb1Erg8Vy4Js3RwngwZM66O2Q
T500b+eG4QlUSNq3oFSHGrYwRkyMdF2VKOwuGeEuSsSn3bbr8uIuyN0TO7m+Oif5IzpoD6f6UrDk
Ww1cnYF3w4E8P+L1zOTgMEhvex+uYfmOTiNKtwz6SRRiSJ1r9FMohURbSNlpGUbS3YqCJe6/dmxi
u4uAvy7NqXYDVqlQOtV0Js++irazHjNK0uJtRIrRzlW5ClnFCxcxKTZXFlr7Emvoqq8s7iKHt/Xu
DZCSinYUr0x7P1Z29zwXaFREEFpsMWcCR30JJU5aBtX9j9uVu0CohCKOfbJvb2YRuTjvx1WyqIsR
C4JGAYtnvoqP6Y6fn1qKK9Gr9tVnE9oKFkM/Fl/a5WHUNP1v09LGNbG9lnhRWzftf1bBaK9/EfDv
dtXy0MbIJ3/8jobwxeLwZ/4vHwdVcc/0Wfv9VL6B/lQcgHBXcggjHXteVff98IeN8U1DxQNwT6Cg
HGz6iZzGVoOogK+EaKtkUtIHeRRAjGxORUzsgQTFtAjQDeYjzb91+8JcIzYrODKXDcjhmdJi/y0m
Y1RmzjSAQWyCTDyhOmSFzwMSkauVADCSLhMAoWcMNI8+0EtCOkAAXAiw9n+JbaeqSxyv5GpEfVgn
cTW2nDfbpJ+Fz/7IOncHkNo6/z9ymn9rgd80WP2/k3asD512FDWqjRmfEuvtVyiYyio+FZE0F7e9
qFN8a3Rbtwl1f7QuQDF/VBGmJBzcYQijaJdKs8/90zGSfRc1z2c/AI4rz29TQ3x5QT5uNrHji4Iv
8IjjRLyXAbLfF2YdVFWqGvluauCaN2xUzbLXEaaVE8kALRZDFHys12vQ22qEvuOhiEOYM0SAZ18J
FXeOWTk2U2Gfv9AnlGx0QKqDKa6ovBfyOu+vDTgp/UIM1ps4mf43BmUNjRCuAT0LcAZ1YyeRPcIq
ygP8mIH5kQEcuZJ6SyeStoFbJtDJf78rC7ultVMgNEs/MegARMCAHq8SGZ0cyomj85hVRNzk3Vlq
alpNQah0rmp5pZM/dL7Q+1nKQAd21vfprjgUf9TLyv4HE/kWQ5GJfB+gZndcZKcmbLVOt+VhXKoa
svTEw4LoInmo3+EI0zJp5n/VzTCOyXwoqjHRIvxUGiIREcpAVAASpGTaWUg466IaFuNg2kLhtUKg
gVck05NQ9QlhjpI9C5xvAnuXKy9gMLzxXPctkygfapwkIJm/5LQ2MYE6EMDU4IlImQeORJsg5SH6
66XcNnN+fRI7zyibGE28pmdFvAfQW5QEKxFmx4QLXl6wZNI32yPTgm66F0kcF+kQbLxdVRKiQaTP
OcH9IThoWSYsxL8EjB3495V1y2HfepRHebJISHaHhzAJkZjNzOcF+gdwz342OD1m1KhIWG397f/E
4RXsrhVlaiDpI8EOtxGUACcBQKfn+E/DWfaiR3sOIVZP+QjoBP/wn7fCr/gg0bWcrwoq5laeLawW
JVcZXiir9IhGHgB8nrKG+bzf54u+EQ0kQoiBiasCKahEeEnnaBSC7sMGwicMjPQPT3+UUav1luhV
e/BLZZYZQ1F3+Potsoynlg1wT3U6Knb8BkPJ1R3F5idCzQPzrWkJPJRAy3TLfi2Le4TBuj6Ggx99
bAgJ7K3yuA+PTO+Vt23OmYftn5Ry3l4XKYQ6oSRkpyR20pNbrAHGNNYr80OmwGa06xeleQo7DPRd
kva3Q4dbUBZPMfV+szBSSlSr7b4hgeaeYNa0QHlQSlIigWaJ+Brzei146gJ7iwaxiJD41B5OYdde
fHwSQqtoAD5qDthpz7P7S5OYso6FcSBdvU7isqSqrsgFzbnCQqTCwPTm6DnyCioodaAYkfLj10Li
0XkusA8pm3GbuKO9/gmF4rXMIFZxLoFMDAgQJTF38g7qwGubugeTl3fFisr+onzX3BvBz0/LDFDP
gSgeqou5gl0JHBy3Jv6PFo93xWnU7HVAiIfgCDHK6y8GdEL/kSYhLnr7P6SM9/hp3w11QcYvjQFK
a6IgNZbUuNdMW5Tz6kzX69L7KXo2cSM7OB5+y0Y0UGO5dukag8XC+532/lbOUoAqRP1AZ7/PYyPN
394a+KeUDFmvjgZrxHPS3fztXpBWSc6/mLdpEP3RoT3CnsCFs5ggAmvrUAl2epJ5dYDz98DeXJzb
XcvlsEMieSdZE1LLgvKLgx6o1X0+sKb1J5uF00cHAuTsnE1GIF6AQ9aP+24jNDvCQDAl2ze7lRxv
Btw/rOlFcXGsVnS2PprqEb147D2eROeT3gQJyYYXaDJ5gFd7Y/bVdn3iEwu0LPi/IWAQtOJqfFTp
Oo9rDanQCRqavlRr50hq00T3pnsxH/H7nuf7bVLWiSWNdbrh0EQBjUQT5Y+fhi3eD6/7MVGi/7lV
atFqUtabFYJxsdYMu/6N5V3Kh38CFNAzVnfr58Wkstz9bjWHwXG/8JJElZGcoHp/AlY5vMslVFTP
xnAGI3+y0IkbcCIVMSlvVnv579xwC8FeBBv7giJKRuiVp2LelHRRt5ynX/DqRH+Mlakrb4Ko1ILG
M08rNYG0QCyRAbOA7oY9sYZJNXh1qQql0WzJ6slFmyDcHdUhdZewfY2EdlEUor2iuxE5h7vsJm5j
0t7Ob/pE6jw1X1K5pT5Yc4k89NQooJwpfd1WWG9TtrkSGzm3/E0w/3vMLvYhei9kUtVGLBj2CSko
KTEL0We4oMa1mDjZjPeAdHrUJEYcZmjFxF+i5v3ru9OBUVjAImi944aOWWjlPvkYB0Oyi2BaBvWZ
MGLxUy4JO7kjCg+pHfi0iH5V2+Uj7iGMcXfVt4mnfBihgG8S6vEfSg+WHRRPRJfTN0cDW/BbTLJD
1QGcnMR++Ob/85og+HJTaPSIW52hU1OAtgPW4uR4UbAya7ORPXZyz9roAHFw9x2JZ5SUqY8W/HXg
6pmJoXPtZ+RaNMo+VOeDY+A3aOSw8jjurEQrE6xKR/dLpmCWB55C4x0iIPVh3tfS/BzygFTpNUNz
B/R27whH54xk5PmnrNFHmSddaJnOLq9RzSpvhRuHcHBJQ/w8nH0POaGdwaX+9095GUlScd4DQD/+
wuuZFgP4gviz3QMmVqAJUSS9X2FHQmGocMBYREJM402wrLvtPAEOrE5+zQe/Zo6QozJomwnDNqjK
EIqqyWVWSp/rRKKNzhTkcmyPD2rDoT5FdvSkVepdpHSbpB6VKX5aYR5sac4Fd/hNj8Codofj1mas
FiUniLsgmf2CRXtTMOOdP2ZXS9R9m1p7px1rWAze4gwZDHRj2a59nsodUWFbL9MwUS41Ee8Ep7JA
9Q/t0VBd0jrxi487VSdi8NxHY5T43V9BtyTK9XL7XyUSyGc9vyMCoBWnuQvoEkQrUCy5MXxoTSIr
3typQ/mrA30F3MIDscPBUN7J5M1GJc2U86MiwGzInRetBATVtGjJlbbdHulDgp9+c3CajPlAGkrL
fm0uygwoR2c336ZpPClw/gipyyd5kOzz/H2iCdmjViQgreHt9YzgfX0e6GJvd7yayx9uX/e4saKp
D/5LUyRhzAz4slpZBbzeHyNM4mTTdl1Lh7BRHKTzJyPruVfe0EBb55L9owsSBBOPuB8+zKnOZnwd
FHAoFKCr0WOopnZqWBL2NlUsnAaxjcp6XWpemxK+Qlav77FfBeNVWXJa87gdqMUnvM4RU4BmwkpH
aVNytW8sPoLbl3uq3crYIYhUYgg2G0zvKMEihPLAMSmlhmPLkoSFEE/s48GXftBcIADhqQd8rfHZ
/zb8z5rCn6nfXRXTi89RVt6CxPli40BeJ7I3CNIbfnx6E6UflkaLbeyGGwsEq2mWorYSf0Yopa2J
yDwBzXts+BOzPctU6B+GhjX9iLWUD70wZKp+eqH9CM9gqgI3CCnk/BePz56MM1ZskR0XfNxTzdhO
IyIDObaqcZLcYrsZzVqkj9A7QyHERpaV5La9eDqsmdACVQhH+OOaEKCsg9ik+AxJrmmYeN6kUZk0
NrTbfWm/38v+7OZWEJAcWBNYFGmlm/i+lvDZzWIKHwLvaqV80BAaALa4nNqXofzxAK4wm2/F1E0Z
GD0qmO2F9r9fkaLFPMPNwXGz6xeSXN2svf/Sae5C1WLV3fOLNoIr50PQc3MpoSkcJd6wkt2NVR6a
ZZRWBNWySUXtJu61AXArvmrRj9y75aC2dxz8CZHHVB67u8/Khov/d1brTiDtyJQccOuWeWjTqQBu
GdTlldkfLGXRBrPgIb3wdmL98JW7b1vYmiYA1UAYs6fRN7J9YMRkaXpiNqjmM2KtfZ7poRQd3Io5
9sQ2Jh+ZVx8wZZBb609VwNAWOFK8fb8GZOQgGWJ6KWkvyK2JpOYF26YJDXncYcz5HJovegraImDH
SGZnagaW9gLS5+DoGRz1iCJ4J/UfK1UDCmwKJMY2Z8PTg+7PQHWJ3F6MO8D3FkpSMJgXDszAzIIA
wv8FxTxbeNVuH6LxqU4y3DTAO4y+Of21HrrPZYUS6fxYvConM1eM/JuM+KnfvomOP/sJuQIuwdNp
EoI0fptLucElNS/MNo5dR/zacoIbYR4wLFMrFxl2CFxu5HB30K2voobWMF7hOSHoVMf36hBnS5nf
uo4h0W7oCuvwzpqW+OYq1DELj6sGUm1Jw+abjE1u8KYFHFLqr0UnGjCgqIkX0kOQrl3KofHuszZo
OZBu9qvS3hIWlO0w++QYl7F5Uq7Ef8blySQEzo7LhoiNJIWjB24hQLGO4WXQwztyBREqff4qZnZf
qug7nWsETX6TGFanM9UZykTBb1fSGsTh3CUoOFZ+gHSx/N05hYkVd6vr0pA2eTw1bvxtzfXbBRxe
LRhXy9aOV87JcG10MfPIzcIBTARrbEd4s+TQBI6qYemJfIf+YfafDhIPaJmSN76Bh4DwtjoDUXI/
X4cvCZ7HYGzrF0n3SwXpMqRH2a0eL3Z4v8ukwGo0e2fqXCMJIQNF7wY+bov2SqlDML8DF5zWaT2M
X0QN/HN5yQx12s7G+D1g0T7/ye6JdicgMKpJBLYcl0nw4gr9plkx6dA1JuquBw6Q6qRboWVrYY0g
sUVnUDaAHB2StWVef82zC0y8HHEmWqr2PyrE+gi+7I8TX7DfsifpPY46qYfkReVgSudwuw7NqV/6
Xk1FaRgZefOpaR6z3eamQYf2UohSqsL/qR+AuwgBV3WlStDQRwFY4aTPBMnuFGokS8RXfTMX5kga
+gBUX3q+F1ZAzo6RlddxoGIvnWxSDwIumzRS3t4hj6/myNSahjOaiccWzAQxZOMszthqIqYOqWaj
R3DcCLxYM3mLR3EF7btnKfMRuP2XT388C5coMbleeLF44bYFxcWyKmfRdQXqCaXuh77VrkC4WeDH
Kw9HnAfwE7lo10vAK4cxUX2ZwNZXn88YcEtGRSmI3B1X6lOpKZsE/047YU6sIL/qWaNcDkHx52IW
MY7MC/KiytFMFmUQMiiCPZLt0oq8+BHG9ZqUdc1HQp6sACdyKs3kEN35SWcqZ3Q569x9duVQtgs9
0xHLAyDrZS0Itn/0zXblLNW5JC8WpWcpDXiQy+YR3alV5Etv1NVe3DSm6IEqwSb2RCteNGxESOaQ
VgQyRsvM/TLRwggDhkLroSv5bSZJbfrHYk519kip8xy+OP9MUah+WeL3KvsoRCP72duHnbMxH3XJ
wG8wqoxGmRJOQU5+8pf3QyvuZ7rQ5w7hEXdgVkfgGd04m2rJqUy/Y2J+9mK4PgHStsH2vIPhueFB
Pg5UM4fTqLi+RtKQkKSsm5dq6qg6reQtO7a+zSgrZdhWxeLIII7c67xLhpFQafyzHFDivhIkM07i
yQFdx1xlLeysHMhKPB7v+3YRDse/Iplp71g+KeJAQh3k5c7vKfnpjCOlwlpm6ssSS+i0FWmAs9SU
jFM0u5buce8htU545LkuULAIl1hMgZJj/TSwv6A7+4sJaLA+xTmJp9s9u/tlaZCTeq0C2GOeS96h
tcCWoguJY8ROU31+L7PbKpy7Cu9mPtYoCBxN0IRX4SMHW/XJZp95yLXHfXeC2G1NIpafgrCjsdDA
U00LwjmORoQiOTRr+LvK48jlfARtzGh69kYQ3L2DD3T6YsWEhINq/9LGnLWwYhFFtxMbGjJrrmCR
V6i0Czj8++AgEwJBTTZwV/Wow9pcKm14QYQidYhOVXUKYsxQ/gEbmWvxPOOhz2GEe4J9IT1TD2Ce
7Hv2MsPZ7CO4o/gYQNZM4+hTUZln80ZrMdundN5eTjEUZgc3T8DdEXtTelDEDzEgkjPsyersJqQL
aYGkgUEDvryyaidysKrJK1M6gbKdoEeIk/lHPpDwNdP+CncolDnJQ76MzK0oZonLZpM7m8CyIqga
4zAwc59OusdY7+cPn5Fjrxesfma+gAxNwy/sSALYz8l78kErSSjEq+/wKqZlsAFHajqpeQOOX8/a
Xp+T+HHZXtKe1H9iOmkg1qsUYZTmwRoA+bXtj6eNqGlEkRIxaUYtUqLSs/kiHad0kqu9V0j/GXN+
eH098CyRFIVbB24FDs5GGpgnJNszfJCfQW+zQpwWlDO/vXMEV21FodD3Lcs57X2PdgVwe8ksvqrR
mv3TOE8vns994DGcio/mRhNrEWbbnvF6rEikiLaGwxXygROeVlR7fvAkboJVmb9Pwi1OxgbFIUJQ
SB6tU7jjOk7KB0YRJvLY04zSJ969DP09dORrWRwVe8ldebS4lTURX5j9RbJv7zd8ESJbCfN7LUtY
KX5gfQL/rjUvB8p6B4tGqncyLWN56m1Ne+vHWfBHKe3lRI7RG7crvGIDUJCaJqfG0oHk1DcCWLaz
TYig128RWpZCpvzy3iv82v5fSPSXf0NVu19A7qG4NKXLJuZlZaBvkmq7vGV40jcJ1q2o9XMgoMR6
qw+dTxbel2h1jfnBbzgLbNMq0t5eKNQCPGA7Rw28y1UHI+0hTOB3to2fqmMmScGhsmjzpetF3kdP
hhnyPV6AUxaX3U4KdGFJebObISPIb52BS+mSrF8Gx0qb/bEA/A5eW56OgDWan0CzF6sMqflc4zIY
KxXpcHvRBj8hFHns4Mn6EVqUe+hrzHI3wklqhIcI+VjDMQEu9PIOg/+Nr/ZrE7JTEChObxCejnEp
b79l9TeeBXEYATJhlP2scO83edLTykiriHutyrYGQU3WkkqtFziRvzAu0LSL9HZIKpHWy2OhDDkd
nkK4azc7z/b16sZmwrdl4DIVlsU5ywWun4pvX6BqYWS/u6aXvlN0Q/p6MYNkqhDcvPC5A83f/T3S
vqZPgu23I5QJHTPSlGIgcmKaxYZ2562E9X1YTAeIyN/eOCYwOxq9OMnGzCeRx5d7+g0re2Ch/nYx
jPb5KZSqVBsRZTE6gNuOHR2DkPyGilaO40EmLX4lfjRXnTviw5mzbwgwvsyhWjCyMfp7TjBpKhAl
MWhA1MHyLPrGgx2soOJz/8bFHTyMnc50YhgkTHgh+papTWgXhXAqvPXhDOKBLkx+On8UyVRoB343
y9xuUIQk3ipmguoxQvx6/iBsQxC8FoQVQHIT7qpku1bF1v5Zf6rZOqm3PZM9sTMKMKTaZUfKsZqX
M2CoTuluW525P/HSrEEDZmXeIgSu4I5cbVqnTLfzeHkEDykWu+8oQZ9HkgHf6JzPhGn7w4eZukG8
ixK6t6Zz/XEjB+eakZ0DqzWjV2ImNwMCvwwci/kxdpdjszT0APXSYd5EEhN1RLeKoR1EZSqFFWX1
hL2e6d9aHbAMQazXaG0FjSftS1qQGqDeTQLdJKAPjG6BNglyxkvv8HCzkCZkYuAyt6UGuTUzvAsu
eXoQ74zzI1lqCfPnh+Xd10sf5/6SwQyerMUSzDE23cshSDKwS+pEcIERSF46xtLKkNY29l8vabvt
1KQFHrsj3+Eg5LPjkS4w4Z1t0HCDNk7OW7AgYnGTHDz+gWEF6JnniunzjrFYxrx/MbB690Y9IVue
sQCvXPbfTCje/zwd4eL+fOEsKDRuYfybSkf75SJFv9rGEe1JjL3FWtxnEEQq3up3nzOxObicQ2FW
2VeqDttXct0znZQcxbC9idj9n3dFVt1EzmhAPSihRg0e6V5hw7hYOWk5aSKi1vsrmMklimlwFL7d
pTLYi3pTGZcIcU+xwWHecdB724mkm/Tq7P8o8gZNOlsuc9C9afi2oGkb/MubFZnx5oeYrxsd8wZg
vOGOYMFu4uW1Ph65RS67zslgYjHgFGMzjihZvTexCXeEXrr+wXVqSaiH2szQ8NIFKLRo+B0MOzLu
AsAiFUY8z2I+v1CzUYYVIrw1pfLQGpzsrUjD9GWDTFdIltQbj6zm1gxBYPb8u0dMHj9rERg6v/QH
nVVERB7e1Y565ZbOA/pq5mP4IxVsMg0wUeQA0GSRUJ6xTi8jJ0RiDx0yRZE93o9ogqQ2+vT3KpBx
0lQ79qXtC/XDgyPeTAfJ9ZP/mMQF+zGSkGT8Ld2jAQjXBG2+kdXeC6oPqZUDFN+4hhQbnPU6b2uv
JNz5k1gBCH6d6rc3jqr5ic2ahPkkPE2coXWQ7EebHrzj6aVv109OQEmqz1wRbtS5tSOC9KX6RU+7
rrDDMiXPEOyeJ74dExP4Dq6h1ozsrTVVH69aDVA/ZkaFDDHSaDf7QeUIkqJ3LHR+7Eiw17nEAhL1
6sbcQ8qu64nrC+sqkfxcywMd5ZEpw07N1ioQBpdNoE6ZKL/qUnYFnL6+JNuJwkKi/0NMMJp24UDx
eDW/wa9KzGXkI5Aqucz7WJEbZ1jIY7CpTZ0JGUeqKu9Ym+djxIq9GTsDWBHWZ/lLIaK+lgJi4Dvi
Z6v1W7H1yWmn2WJRqAG2NqnhzdpNBHCtTUfJs0EkTsmDtbxgz0bM13XzGBz794aUe+w7qYJ/tnDa
29bO+CxseGyPD9h8t/JgLvZh9nnSbqT9E7mPw46of2W8cM/c1WoqEPBb6Z9c6Sx+Qlr8JW/jCjI+
Cn2hVJstVCg0OTzzmhJU1uH1JcHP4OZs4OjSrKuYFJ80FPY2cwlwE0V5GN813LcZfTG3W5+NvKeZ
zuDHq/vo6zdTF2WzYgQoaE8puYey6zSK7YgyJCoRTwNUSeebkNwu6LngaeMXUsnSb5OrA9AaHAd8
QgEDzlGFurLYV8cZ4G2xgeJcNiAXSW+LjT4x3/NcPoEbfgKs6e9hWyq1uXOgOtGqJfBt0GUX3vVB
vHIUDBplV3niAJaaEfGPl9lgNbWoon0OdnbimaBUdyewYKHtIfUXD6Zz4CilNUSjhjH0dsI3R0ag
voIA4/1CwP7FHOdJlhZrc+xFz2/2OIEWI92RqmruP1hFZKLdemQ1JLQAFiAwMJ4QqXotQ72Y6Pb3
CmkHgjXnWDasdGyLfTL6HLy0qnoZsooOC3djC3NcshTBwn6vA6LeX7QeDHRlzBXTW9gC1HIEGNmo
Ts+52R3neCFe1KEGZyRjU76Zht6/R354yhn/FohnUpXFrNAlZGSQ1kSalLa4R3za+V/oS4YOd2co
SFwELgBZRcKgxzyvKXO3Bh4oH8csAGCp7Fz7alrx85BxTnw6pWZPG52dOMHLp6Gz9sqBen6GzmYg
l3U83X7xck3SmIxgr1V/Z/L+t8hwL+t9tCL63gHT/d4x0AKgw+vSYe1+jdX254iT604xeY4JM3dZ
5FdDvAoed/tluZLHe6PIPkAGlWr+Dd1pTc+KoYlX+zTtUswMQXRxfoMOt0zYLGevm/fblN3rIp5j
PPodJQLi4lIscsahyX6LZglKLefO1qYZJWI2U1dYg64uHkuHHMPcFm6rMrD6NsaZK08TX5HlxgZR
QmkUy8ywfd/1RVyRbNQJdjVGBHudhpfXP2Z/5XhWtVy4mhtwXNGTfhfRtD9Jh8X6g9WQF43ZZoWQ
fFanOC1OWJi4cWPI/FBAu/4pvysErQqrUqgZurvjzH0EMjpV0MZwz26oWNGpyNHeJxA9tmUyg81T
oi9X3FJVS1B/J5LBQNITTeDjvlTRiGXTLdt+qULqRbOkgzxuCYRgltUtG6cng1OSyCcu+A1y14J9
HF3H/uC0xYVoFlbZXD2s1dUkg8oc4ptgAWCMd6SUB0NLrYuebcw5bLwJBvuQJjzOnyCZmrSAKOmY
t/U65HYuIezFYK/x2D2ndfN70gADFY2sg7yfmrkPhfal/UQ9cy55NNbaPgCc2LNGEBNDgnCECJXQ
ASXGJSLtShcrnHJ1OmODCb3yHeW1p+OsoPSF8nFgql57FsZSWFDlLLdhbFWQIIP2V1v+uojAFCiw
O9PnxqdFa4ysdV5/r/l9NBz48JA4ep7WjK7mQcM5aWmp7r0ZRSVZhJIM0tMOpj+/T5HdUjoxXMXE
Yrk6jRk1E1tBPmA2OKzRQ6ylpIzngvJFhtSq3JfcTS9XafkR7147P47w2nxlv8EF/f0udyJsl7m/
JKSlk3N2AAzDTUhB+6CfM8H2aes4SdRogTN/fnMERhoQyQ7YU9kGexjgD/9P092aX4fl3LXLwACe
FO6EAGXy1TSbyiWRp7GLbHxnzyG6FZZvTKYoryBcTMABXQ3Q2xUOHOJPmzAfA8RPTz6ruaixZWOW
2MZENE390UPMVS/SMwV83PBIcJYRZVBMAoLEkx400iv7ggvC0V2bVrCmj7WXtJRiTZweAQijDNTe
qP8GhGDmcOe7myoo7iv7TWL8thZkjUHJ6lIeCgbtJiNwhGEhPmivkOrTc0/QogFpaa8aUv2B1eXB
K3EgJ97gqbIWq9JCz0qKZ3zytAZifarU4bEi9eSEP8Mbo0UQWq2lx8RXJC41T20Uq//XoqUSjJQF
+UA9ELMjdfcyowKChYQjsFBGNxLReStTQOa4j1xn6eUmsSrMcvGoxx286bUYBf+8ecYVyjLr8erV
reuVCRp369zVoeB2mXWIj3bpYHXLDnOqE59wDKiQzs8HXyF47i45eAqlDsAMy9ajAWjqpLc/fPsV
d8usddB2PruB2wDhbuFxdI9++q3v+d8YvCGEu3K1EgDbpJjNS2ZlU5wA3Gpzqun9GkcYBsPTu/TW
C261AR979f4B6dUDvRQyF0nJQ8cz1himQQaReC4X67woLvXDd+2CftCmtqlMvfumdtXg2fvtDrQT
sd+jPmg3WqhIXsppbD9Q/DOQ7tthB4mh1xoFTJhjFpoc5Cvrd4D23OoopnM7qn8gFs0zvNRmoBDe
klqucqQaOgSxDsZTQt3g/JDCWDj7FWYB3fZQOv8NQsik+v+Iqeckcwa50rOgaYAbA+GDu3Kno+Uo
CxYgp4/T0DV2Gf3rREN2nB7I3pvCapsmKaYx7q0YdRztQaiKXA64E3DUK/yPEJPSMwphazeSCe0t
17ECW5ZzWu6KqmRknwtGBwfhIBBZXNE1I8EAcV0I4OHw4f2fqBINRKOsm3krcamgrM0fEeu5i7vm
Gdmdk5IgXjzYb3h9ObcIFyKjFrHLoBml54NkKFUVT25OdgE5ZesFQwtjwqc8gm7x3Mx6IIhuY7bc
Hj4vU6Pau9ilbWE2MgeIVfUFqB7RmNqFEbKQm4mXMWOo+/U3UrlTVuNCiLrAKyg90KLSBcKR0Xdn
HsjIRcXE6mGks+8lRoZK0ndj0zyJtRiFlgr7z+wxtEOrZG763jFQt+lsjjtvamgLkmb21v6iHO1H
byPL4++yRP+b1y4Phu8qwqc/A51iCxCbPLCISNGrF8/j5NevMAW1TrLN7Dpd6K2ZhyruRR50uSkS
XfXv3/XSdaYzOsla9emhtmHfriq0r14A7GHh4a8Pp7/ZDgQbboYgt3sxYTu/tiSEfTd/tBqNhLdF
6vLYhvq7CkhnSlL3hLPWi5R0LfOf8jGmMKI30M//Hw9IxqwgEYLocn688kaylSVxhjpfbAOTJirA
BtOTEkOSt6rWenQubO24QqZ01zwtGUVuXFhLP2SxvGuAk4zf090xzlm9pSlL5bLeJfyYANopG24z
f9+BThZ6MunE+v/aNqH+6I3V6HG9QOXM2PvSzd2KZ71Ze9GfkHe8rafcikxrUcZ5IeZgPXCK6FSh
IrRcZbbQguuSqrqf/PGptCRjwPvCxf3xFd1Ke73m/dHdv43M6JyfIL5veHyt+6gJRvA6EfDbZKXn
GKwPEeh5HpBTwkhPLPGD+o0aJ4lEC5V9PaNgD5pZijHxj2KGeKBLKjrs0WPFKwLHdMMGKARCQR/U
AN53kem07qi54LEInk3cf/SGoqDUdpWYrJ+B2FsM4xAg7N/03Q9EpmKUfDjp7n/Q0K5mlYzAwdxt
h6SELWGmHSIGRv1nBhz384xe5V1UuRzk3nrT8KjsXNJfNjydrIzq4ldmJ2LB0omfyeovWS71KSFp
63+tsnPUkSw4hzjzMB5IJB5f9xUgCrTwOtD2go0GzvuJSw34Y5unaP7o6ybSxx8IaC9Uz23m/TXF
kV+1lkylyp5392zwqLKZ8m09Zfl7gOdc/cxa1mthaZBg01uNr08h4JINMLgk1DZTB+Jk/2DlnLbx
ACI9Pife6XYda/PAa+wJmcY/Lqi9lTpeCFkrkvuW8KpcR55uHGQrKnmw8aUW7cCpk8t2jd/oHdKh
OeIM3J8cTK8ewtzosq3ExFpCNFmwHmqO1hVnoesVUo9AwlSYT7FaMU8BhxbH8wEvUAuatwCGfBsQ
vii8UVkIOARHXudzDwRC5IUTDbxnAjpSr808J+2qk6brNHR55ociCN0/N32I/6XL2NbQVOMhQHDO
/DnFWs9uzBjzYwMUtVmSRhmcCyJEURzf79TQukDWGni78bMsaWn5lKB8OwVbJpSJRP/f0vdu82oR
9PdiE7IZIrcu29901NVGbAJH2nPe/5lRUhMzrqItN3zZCNmgvLytM0/oFflWdFlZpZbjIQ3rUnYn
GQazePD2c/PENL6Nb3kPF7mCYEwVTYSunglsjyJYzD+M0GBcU/74x+ryBR34wm2BMDBVSj1C0lUH
/HSm1LxnpQRjOiIK9iEAeimO0pZH8iKWwtjerwa/+VvDooABC9UwiMxv61uC/WQQnfUA78PYUBd4
sNk8URaNRPhtwa3dmN2oc55J2WHX3k6CvrfUdUlsH1HTqHVYfRaybJ0Namv+LtkPgG/PZDl1lgdc
ZSi/M519m2L/OcH9RRPcPqK1N3Tg50W0vNTEkU7hRZ1jMVZJ4FN7eIfKw0iXlbp7krmvsP3Q8/x2
OXP6ECTfgZRrF8afuHdrIt20wGmVApT/NiWuom+rJZFOH4l95mTPVDHKSDXHIMF9OuZjPHaJaf/j
cj6wX9vAzoGt2HBc0AzcoQOiH6qgEwwO5BPLi0Lwdn5FNK1WG108FZZDSHAXzneJMtu8se/h5mz9
F6VQjXzl9v4S3A5L10Pe21RBl6qkkEw+OM/b1o4EDkjqTp07zjEwxnzv08MMbCWnNvWWbAesB4jj
scag4UgSvQ3mhIdB5UkI57SO83xVneDU4kwN8pWYXCl3x6p3DIG8mekFfOSoSIq9NTMkiNNt1wzF
G+15AMBfr5j6mgTNgcQgtqQQ9tY51ZJshpyMGLWbyTHzi9iFPVjJ3z0Mav++Set0derC9aELjJqB
araSmcKI9EdWfzCjb4gVH/mlf5ZBruxorlKsn3PBelOIhp+Dpqkr9hRhOaUUF1cHahA8nnIxqhW8
DIBB/bijyP+kpnU9MkqtMFEdBCA4mLfRYB3YThvfwD6+MLfx2e4UGevfepBEwJQsrkDijzY/aoLD
KUNq8vaE2c0hMcoVMyA1mCgk2uRT6EPlamNLuJwz763VQY1Um8zQgK36kAYCsHUNhQzKJHr3MskY
8lT5wTn5N7lhbj6J2WJR7bC6cTMF6OvIF6Bp4EAlzDggcMg3SmFXbbzhSQz8x3HeIY981Ua011Y1
lswF/F8qoGkD5esJ4SW+Lxrs0GDaDtgB+oXOMGxl/Cw/WpsXrhVPZLBrxTIMzdZ9NM1+EEHnbcEE
YEwV5uLl820u5usE9+cbyQIxTUrWUm9FuxSrE/CMShSDXYTwWKWc3tMilnosgj85RTaZC4Dr0qPY
hY/fe45WQX3gU1GmoVP06CLWIz5DizR5mBmnpeLLqe15SEUb8XfCAns53F69X2oXHBFekDAjbR+0
7EyruPsMLBovQmNp6GZoejCS4nuo0EsT6EFGLklpFa+KumfJUX6NIf8CFbgWq6iSN/+DoPLuz6Q4
CQiwOuXEqGahTvpt9VD848fclRBii1it6NWqlK5PWZbez1hORpVrO5Fc9eAn5aq/BQ//qGCBGDTV
ciyZnNFt4dNQyV2hCL0uxmvK8rxbEGKQJAz7RXlMrY37Fm+vwmKY21c1PU08+mMTrj1dWVs+FtFj
MMvKDfwiFER20WXS2DbrEQICyuCHQZDizLSN58cRX6puidDoOZAiJEJXeXgaZRYeKoo71Gk4444R
eaoM9LBdJKoXkfp7VGVr7YaMBNGrOW97QBokXf3swFlYd3XWOUtZ5igqIVPSRQ17fQml6+ake0g7
Ix7RYZn8T2mgZYOuZd7aBgU2Lqn7Jh2A+mL1wU/oQKQ5U8u4beCWg0waTjL2r67LOnELyPLFfIs5
vlK+MXdrhOd1wPQM8k972lEALSRBcxZNIr3dMfCtBrHwFQOe0JQxjWrSX7ArWp0/hWulyGJTBw+o
awoAqckb+fOn03utNW+MUoLuciagkVLcZ/nkINaGbUlDPDTF/b7mwb92hjW/Drq9vBigyni1UcmO
XhTkth3WdklHijeIMTLv3AA95Hvl/mOTvnRIU3vAH3em6KoVZHj9I0ebIp3EplESd//esdR0Nk4t
oAqoNg9exDpiydNYStWxz0izTw0QKSd9DeiHFbPz9Rfmho79vCK5rH08iGFEA84hM5FTS8aGpcL8
cttmdjWd1BhruviDX77R95u6fUhhBxvobpNYnXMAGuy2UrgzW/9fa3d+bEH4dBZyPuVqHNkrEw2x
PNyERaRplslFqMQYKFDMFteYqzkcfwqcQtDLkYLIZIkwYk5DcOrwiy2J8serEOTQGDK72wEmF+6H
rQpS7oTCeSoVJh+czITAeYxc80FN1/1N9EcO8XPtP5O2OgWVhsLj/UuxFhTxQu6nrWnZwrH6R7th
5NSCloLSItOzq1cw5EWoVwAZySGTKjc9uLp6JKDQtjcFbxoLNP2EuMDCAHBK8lvAtN5cc7EbB88B
l20nFRZfnSDYSDyVdYcMR+/vtdi+4aCWToyCLbq54WGWJMjZJBt8l/yh2pxp8v4ubSjjTGl5ZeRY
KPdxlUJ2+EWxY8bm2R4TjWvNg3TToQfkE+4GjBoVpaOOshjHIgy9/FvIW2C3HS+lkwkgTGhraCIs
PfvidciQad9CkCrs6iMqQ1spEBfEbTUuOsWYmY4lKMWEBoStlUaXgduIKRut7vQoYArroY9PfgzH
gOIndeaA4iIF/LS2oj6W9Obr4T/UqvZlrnUIHy8mV+H+zt6wqVmcgo20VjfgAlrIC6ngUAwZhwph
qfoUfOOiYWyItbEPKwec2k0HPF5uDJE+9gttYYJDkTixQALs12KwIE94IOgxkUVzO+CCImeW/Tcc
YErogp4VB8rCOYD2FMStBV/NjoiUqDgwve3/yVaNdYv+dDgL3F+1q8QblBSnANjNMjG18C8RaxDE
8XiklGAZSos7xBK1A81oMcWZLbV0HUm52iyeY4w1/lPvVSJQWhxz9LHUDZNxyqkM2KME9BRp2Qs6
BwrbuDbsVnmArj4SpKY6rh5FtfTp47S02o9gucILNN4TcbSjGSqObX1Q8SJBBbdBg3o56mmBR/oz
mqMkoL4OKUwCJal6pVo9r/n8roBdxfp750/5eL4ZTnAh9HMXcFCDEjq/y6iua/R+B6xRu60Y7wo5
/4yqPufgYwBXBz1jg2qbAdLCRc8bTe9PFTmf6qtg/AEDL+iXUkPHWrH2YYIH0jG0zI5sWIUoKjzT
GStA6NkS9XqCzZSoQvHhRkIQiIN9dQ+zjeWielfPjHGDux2+nJYoKpwQM84unSATxpzlz9ODdJtp
8G4SxMqzN3AyWigYh56RCu5mxnlOXo/V2dmcF8JWHT14zJxdvzW0LwGBLOdPTQasQa4WrOFmi2RX
DAR1MPaJ75RGvHxPUw0o6p36ev9k5CG0iN1X2u5zA4bEfDEaz0LL8a0cnUQCcQS100pauQCyiIIP
Xen09PgQyY7j2IGc4sDRZOJS7KPiQFCh0BKOsYUXFkmTigfgQPFOBE8tTtzaG4CIm9FZboSiC8we
37w6yMRnxBep4251kS1GCMldtHd0kHulMeua/I/3Ds8BzW3a5N10Da7Nc3GvJAFb4nHjG5BPA/V6
A1dSELVO1JiMIeyscYbTGxlNFFgqtkvj8dVIyCD7NzL4zF452GS4xHx5KQBQo71nGaigz8yejpWM
zYgRwtf/x1BUz6g/gobCHKe4sWo6AyZmJabTr5rhBqjY8WtEMy+JeZk7GXa9t5rqJjrKGHq2+ijm
t+NKWSmgMntgUEcLGM9E5un3nC/cjSCkZR1uOap/JQdpx+3fiW+r0v/dRcif+8Tmb3yC1oNY0p/8
WR57ytOUF2wqAdnUlBm8Z3rJa05bRxIMP7o/8pkPoXk7vdK8dgWVapKzkUPo8CrRDiDMXjNp8wEi
aKHpmJ8LqjP0+nyHvyr9XeCwoiJmj18FBfBy4aTvJ/EgrmLqWCQrhhydwrkbhtTgmsznh+OilrOV
Nf89WkPxdezbgh4k1BfU9a2ADc6LwW38skx34oTA3sptVzqG9Fxwi0q9TXq2LrLHerJHZ0P1LJvq
i582b+WJBxOJa01sZnj8Ul3CtYmlqwsCdloyYx7/LoULjsLdLORVM2ZVxZFmi0JUYnuokT2pRvEs
mUGud9BjtkMOpjOjc5Nru1MZXiwlkkEmHTjg4Dbr6qHZ1fLnfmOC25qKivGLqHC4jY26OKUWh8CJ
yd6I8tFmLK+GgLGnLZjf963GV7QRK9R0c0HTF0HLICXVxG3DAC35SIXntwtGUxIFmR9UwYWhNorz
LyeyA6rfNFYh77N09aNKBBut43lI2lTiuWoxbvGskbVDvSYL0MQ6tcpbZyhq0GfGP0p+3FQ5X0BN
3MGwEpWaRtRzZ3rKg3ygb73g4UltKj4C2yRk+kWv5PkG2lotYMXpim8Ay3Ov4jT/mZdwCEtD2yMH
2PBFG5wm5KYEnaHmzG0KkDn7AQSLN1q6or47ym3bT0lDf4cFmuHUS1vbYA2OQS4dyjEajNBN5Njw
0cRjMd00rkKf0ItejYMXaj5ft1kiQgJkVmhJ1KlNdF4jeMLcAFBu+SB9X7tqVxQn/sxx0KleDMW5
w2O8jel2gGxrRNl3uSTDeXM8rz4ELNtkLD6IRi8MqL5xO6yJFaDjORvgVEIJLjBmlo+mC3+jVGaS
dNGTAvVamzvjwYxDJATsLQG44sXlf9ZaO+1H8weelsXcjtLXu0+gDntT1BBrkz3XiSXHACK9AF1b
tkxsYWmeDdAyZ8jGMbF+xiKLO8bpb+yH2yWvydqNmYTz/Gd9kxQjLkJMCs5gucNqLfF4xI/CucuA
usF+9x4obVE/JRIpxCpeUVuZGYba5RPon0WMi1tXBVd4EpvgrC1rhExoz9SIKulxKrfOI09f7z45
akGs5SOt5hCZvRNBVBoMv7sUsWtt6Xhdk1jjgRjqRSRrJOZIUqPgdwcd+ZbxVOUf0Dl+dni48zIG
VzBSZ43QmrrSpER01+VD9m4Z65xfin+QVBzQFKg5deY0m+pEMJNHFB1krMaXb5Gne6FzAGjMqxJY
Tt8YiulE7O0msi5BUeQDESH2O0EsjXaPhHAosPaHMCNcMaFkHNwjG3l4UOfsVUUxs6FF2ZG5SI+x
RbcZOfoHpYZsj4lDiZncbzaTZDKEtS3MgRlm95cWjLze4fquEe06cjBcYKDzVBsQvvcbAvKDTKIF
EsMi7jvfRIf+H4I3/vL8rWWB2F1fxbomNZlPk86S7u8ZkuaxxnUWfMgtfsxDMm/EeggGhY++o0dy
NHHJM3ldpWcfWAJaKS1bWAwI9vCaYzpYjAT2CWKN9gYX2JbsRbcsZXgLlB2Eo4An6iRX8lDlukPC
g75BLjIA2roxIXB4GYe4PKfJX6UdMvgwLiHAhhQQ4tT0vQPwCxeJ7O4FPr/snmpF49RntSm8V2N4
GCoIva0E4qj1p+2XLuv+d0LjTLXoLY5zaamZKe3Au97V24DTbVz1Cwl909CZJJzwCv3J7/On9IRi
A0RqFfvQSPLtLRs12oA38Oo5xmGE1kadOsbLWDM/Iww12pQp5dbVuhmwy8XQglWHSimi2jipYFbk
DNO2lCObLJRKGuDhyC4Nxk35WWqhRg/lrnUedBKgs6DClEPPawl7fUuMoyV0bbrDt5DANb+io0L8
/QSPEn9kizfeRmz94F1HRUGw9C0tSzmRmcyZ7EWi6sIfAi8A22bD76928YC4wZ0nTbwGmPwvzFCR
2NTFa7TN0ejSCKb1Kgyj1J+MnHAbgEAOiWy/An6GDGKvYmj8DhHvxrg0FLkIZ2zp/pvTNCsCdyle
8jhYFEi/4sXPC+2PxwFNjGiG2DbHRTHKh0bO2tKDVvUL+tHUHcqVNPXbDP5GqcCDqYO/Ug4vVecs
kASFuhQGbK4cw7ZqP9Qxyrb5LArlj+fVxAdHD6dFD5nCYiftpfV/L8xv82vaVAG6f+pbjKKsoCLg
gH1tmjD0SJAshE2Z1dsg8vRCZ1TH3OVnzh5yoj/UQZpI5WEDhAbPM9WGPx8daGmQA1aOY2IvzBSg
SWh0o9rr9M+7z0kZAxEUfIg267XfpuCFuGFPk8/7wkQHnOmNuPJTwUZ5YMBtgEN3spC9DhErnLYo
3SKXM+GMMfoMdMuxE9eh2YQYGr+6qCx4HWOn2z40GoVNTc/UMyC30tb2q0DbXrk2eBcZy72yyTPf
sbAto+S8XSN1C+XSYdVMQvzJDw+XFDvARj2QJcQ9blemZrpb3JVsR7DWZUZGzpRynnP3kBZ4ZJFm
vr007EwhJgVXxR9br8KXE9Jw2JE7tzzpXEPQVHU6GuxFSev9vVWEsCOfHbj6/gzBUF9YeiFP7ha6
Gnyu1kS1P6nrY0nTjTbRgnmjnWhr57vvu9CqFKuGhLxPi1rcOvt3iPLtpfukK610v6XqRrHQyWCI
oEW0baS01fY6CqwFH+u53GJG5yEVqRrOAiwfp40c6CnXWJL/zp7J5njGS5DkkrwFAaJGS3wQkEti
HzxX6eeR5oISi6DyOMHXEBwzSEgoaSyvLUKme6MJ8MO62PDOOiltKePdKj4qs1j62ld2B9F4f7u/
CRz06lg84CeuCOnPrtEKzFk//G+Hf3Bqybba5+Vhmismx3jyBbeouQxWdbIe0/RZFTa0F1R1BwIM
R5OSciEmyxWDu9P43IU99iXwxof3rCLuWEx9RNT/uAQclFRxXYp9eTovkmZ7x66lXZaHe0sPDFY+
CVzW4v/TKFMCSR3jjbxuxjXvL9GwB3rq4quVwdCXHpC1fvsgClJnyGYPULMb76eMYYRwk+5pADye
A0UP53kI31v6PVRKzhhvNY0EADRfK/SOiv76cOQ0tojyR6x213E86zXBxcLkirl9+LNHny0LBkwr
xgu7OojCwpvMcxtF5HW2e4feqmafGsodirr4ox7XCh672YtCGof/pWrObPLkgfjubsjvfeemrVSI
C5LsGPTW2iGLynBtspP6lM9OikXC956NuTTM4d1w998TRuoQCT+iGcHGySB6EPIhF8JXI+EDArNy
2FfY4Kks6BjgFhfD9YC+k3iXS2HB0XGTAe/suOCQNhHoh2qX60TuKN2uAswtLN8X09MbwcAlwovx
0BedmeiacM9wf+l4hgotEy2POIgl33AJHfdfCLzQH7IzKkCepc0CXn9KIg5hlT6fqfp9hK9bwE0n
4NkV3xd3wTfKyr9azA+IL/umc/YAipmMkzzrNfsHDfE6EFeqvorSl4PjPQ5LuTZ9z4DJW6nUrtNL
4N+thdb6j4MarplnJyJU3SsLOfbgiQRPnMZo9pO3fP44/fng4MUpLHIdfOpI0Jnzmxixd3ZbaC1e
1D6EsgprRm+RMkYnrzXLlnqE+VJKEGH5Q03TIG8OhwOSXz0octgzeNRMenJ1iNR55JB/Ltu1cy9u
b4MeD9VCAUaw9n/bnml3Qn6OftsVYSFOy9qlZUX15uD0EkFfwgH/1HJv+uyUVAa75AIMgpgttbA4
mdcRReWkUsuCLe8IsAvcv2r/UbC/Vw4V+awLPmRMDz2EA6mLJ7qfpm97YlM2x7bvvWhy4WyUOvf0
awrWuFEChGVh29QUWVMmo4qumHQ9bX649Zo0LdZB8FDPvdO/Bz2r+Ril0NpvmSCMVofL8245ezf0
+gu+E9tieLDwmAc9ovD4b+gFnqWr5n2hXYS0gF5wejEkMx2WFIYmxAD/No4pD1chw0DqmpkYqbOp
nbPE2npp5SG1r5JDGNLPA4tMaEGqhQd7YqzgOdMIJkJPlgx31zOS1z8+IM/reaRzupQpM9/R/eGb
nH+aw8I7I5VALi2wHPDc+GZCp1FdNqibu6mNMpiLSFw3ajRb+m4Pgue7kUzNeqXH9CNQp2qiW2CN
DVnNaYnSYdnErP8PIpEI28prz+wXYA94z67VVv86TupTNZA0r2seV/w5ABN3J1+kIMFquJtPEMhl
V4Ec9fbKVY/p/rUm8vcIrXQyCfjUVPEJY6/AADzjzecq+NwrWGkdx+1B8Jt+X99x97SiuvQCJhkb
KiaP7klKVTMHGF8a3m3I0EwA7TQ0qiXQlNrhgryiHnXHJ5fJmAs0kFCyDCXhPMntMBmY78hq+cF4
undX4rQ2imopfis0ScxSEcuGOgS5V8p6JQas4Oxxdn1sOt6UQuewnTWhRp3jsX4SPCN9M8NeAq2E
iaTgy/ZUHfDZrNZqBnxt1CMu4I4NnJFu8ld0nPVbgSqj2f4wUMWWANtzRwHdGXZj+5UvDuEWuUHl
PhjcZlUAfvGdDSxfFhqDRKG8+WI2bIGQJKmIp6NcGPBkW3MNBubmA4ldLHmmNhQj4iJ6heWoEgJ2
yC2aCV2hdB0T37OkRf4QB15wEAwTqs0UOujUxRwlOL8zeZYB4oaJZb0haneqC+y42ht7WPkrYC5j
7+4t804MkwIdnbQiJPhYaaJC8bl3xy2MNeexMSkp6Gpa3hNFjon1ep20U5A1IueCyMtF93hemyo+
+q+aJOL44PDGEtBpG2KwVRTBaf85QGsGH1WRg1bUSQDqjYXZiRmMDhZJ4OR4tiZqtvbWKOwNZVUN
tXOgds3iCZB+Hw0QiJIfQ55OjOZkvdFFQFqBlpwW8WVHECXCk0LuUsymgaw5oL2oK8bmUN8aYqjc
GOK7Q+MzMhZ3BGK/5dpwFoYIV1OR0W6THZJCstA3yJqwBY16owkdbv7gzZoqT48S7cgVC66Zcdip
vQYvDga/mvWgCW49/t2HpCshdO1O7/XnT2FRakBFHGA997tDrSewOzLNvyvXheB5IRD4T+DPL9zl
bYdUBLM5Zw+wNzH7NfzmrKCzV70xcI52EUk2BSg2R5TtrJGYKaL998a2a0S/cALs3htUpVI21ggT
T+DAyl5J6mfLNz/JcWFQNAbHdYTqBYwDr5STlSu9a0PNhZBGiUVzc+aZ0ktvhas+4LIYr59uqGGs
YMnbRK1ToMnQsaPbSASEUlXIWEtjvDqS3OhK+Kd+lLVrz0srF0zR0Q4z8sJKicKonrESFeIUnYXD
DW1yvMq8/I0rMH5FUOGh3bZVHfa4KF8r83inltZ6G77PRAnafM0s642dc9UXBo7m/hGwxJi/1ZFW
1OsXCduRMF9xDrcOvPim1wHfFne7V5zstxV1jjeWdOutHFGdyg/oW+7Z47bqkq7pBfsSy5D1x4MJ
xkkSe9upO09NFwtrYNNli9DlQlKPZ5+gK/PmqfuPL9CD6p6dByqNJqGqKMq5We+6ti6yZnIKncUI
if+eWsoyl1eJVo5fNNtsPXQB8Q8Nlb74cGe+Kwj50VRT4uquouiK/YWy8PvkVAO0ixMHA3k5pfFD
/1/noKCn+/IQkLxpuDGXWttq/oMoog9ywagh/w+FsSj+HuOTgsK9drseea2NB1eZkI0JS0PoluMt
4/X59hYLlVomK18edSrJvebrhuYULy1Y8Y+xmGm8IQW4Fhk6f5aNpjLUssIEKu+lLmiafNAhw6tq
9Khfyct7iPZAHD9hQSdbdIApZhc4xeJANqOctGNLN+UFn/AV6qfWki1sdtEeXw/Gq4Wfeu1ND4i5
Hb1Hl3tAZajWxvJOqyHxoX+uB3q77SiBQiF/4whoUBhSP6sfmRMfVQo3mEH/PYJg76kZPKCpKZ+Q
N/LIGPQGBtKn6FcxXaKNqEGsaDlosMQ8OIo3iBxOjmbKkhH8aTaodMyC8lW407KhlTcUPdiaZUPG
21/zHL//88PTAYOJynG/BEfyYz5rq8oPyX88VbGgudJFHOe38IXj2kZrmIE3UqzD0qvTw9EeSA3t
JKNcFv6lGC3hNNx3nAvwfD1/hwAuRT+JtVqcS3t9wH8f2Tz7MgrhWgW6uYlpN+SIwJv/BysAo0I7
CYhJv13uvi7YDkUaX/A6D1zK6wg738JrRNa2hOP944B+KVP2CoEOTia4t1REEe1VQFO+2nI1+nI5
zs1WzQd3tGrDFyPiGSforHM09FnimBOnBAOTyJFJ+W1FJ+tXH1LumquMCN6ubzCSQlZIaMQx6bMO
ErzfQh//OhAMuXjd4/FEaQTxr8W1WN1+CECNdv9aKx5Jof0Qxp50saqNPfedT4rmHihcng4ppo6A
pmeWsn/D7cKP9A9kk9pnIUi5xCBwPcLLZYYZD275BriXqNIWkYvDALLW7OGtLxQPEJwEOWoqwVzA
rzuHRMa9gAVZVpyYaVt0DvyIoQvPGsOn1JXNNPDUHLRIw5YujvlwG+mUgVxF+AR491wagFZuIQdB
87qm68WRtPP5ImeRlVrE+PCNFJBgLGVEmnSm/jU5bOEKrpBlfsvbZ1h7vC4mrLJUKeiFPZ9fdb//
ClQ4Qp0dTKbVbotF0Si25CpEbQy92xmPsvdIAWBti1+Qs37szT+SO44tedYGOkZH0vc0fyeywSro
v3T1ecRcmtjkVZ5UVn/FrkyCbJO7AXmlpPTi3o+joY+uDVlgyc/qm6JMYrTqHpoxSD3Cm3cUfWg7
AMeHVO5t84XddvfyDL/42XfZnwdXyLuG0dXPlVHLkodRP2Mx0lVr28RrhP4HEJPcqtljOm2jqmKB
dbAHEcGvpr4VTATyCeFB19KwPTdFzChFLltk1nlOaPUuJxHlBhTmxNePi+0u+2yfAmE1qH/2tXrS
KvBepNnJAmXkpheKZqwM3XoiW5hWEBfPEG+HWe0UGasmBztDC6vKZOCtMGKPPEAE/bY1xlNgO3N4
ZnM659CIH1eps/wk99Ifw9xB7hQdnlEeevlWcE04zsuzaCWC2cKKu2IMnv9Vk0EeYDQivmV4Zkw1
1jOoynkf43vGF/DPlJ2xrrxwEpn5c8AVtbD704UO+00tnJvgm4s7Zgb/OUz0tZWjA47vNwcNoSCv
g4bts5qZpsUZE+IBzt/7Z8EcH/7aqrvQY+f25O1dblhZ88QYOjQpK6Nvntq8Zg113gNNEcWTs8gG
F12Vwc67KPR9lFj6IC6ObJyrFGPT2Pvi07DssisMBHAP8q+x505jgwNv0qWNUdzX0JS1L/f03PLw
NeBbUwzK1dyHSBZ4Vk5AJ/7+r3bLwdXemSdoXxtNI43WWe2d+yrjAPiazffo5iS4Riwd8NlczP0K
pvkRV6fujLrXHtMnG1vnAQGa9kFMTxyepkN/E7Odt2dYZ/1yASoREsbDN4JcfoGP+v70i0cI0uEh
RHN1pUVVQTrbk8tRi+x1FyEifbleI8daBO8jzir23qaoQ9UBK9zfd9LwjzkJWyTjTClDEEzAYeHN
TgFeCys2G+A2wX4ER2rYkWMYz8oLKEDJAz0kJLyoVAgWheqdbo89rLSPUgI+R/1BLV+H1kkQ+9y9
oOau0zldJmZgfPieogRNp7C+pU/RPKL+xLxUYjEdi8ZupEdl96fmn0bbAxkhyy3MMLQiyMVj6xml
nvBTHHsVlNiEFIW5xU+ufd1z91Lul41w45kny3V96fsuzb5O+XeXY2F0AyGHiiZX6Wx8rY9C1EvJ
4AUKEUkCZR0ccUmL2/C/Q8Hu86cHdRloO35gEy4uy6m1ZrQo+t9bf74ObhtIiuQRZRQ8P9rZm2kI
pouSjUEh1plg/O+mcoZ4+FcJ7KvS1MqpUJ2uZXaURof9SZ97ZxhFf2LS22O6bQ7nXV4KN6vi5cRy
2RP03VX62ZwyU68xa0gsFq5KOLuVKzG1LTiXwWMkkJ1VpPoMfZHkeutaeZozA2Q23SeFCqFGTMDE
ja9HOEBdO2Kx0UvGHUkQiFGU6JoTlNCLShTalo9TioaeSfMYtYHACEMPNi9yAzqHDghP48/6oxEk
ZeKmwq6vxeg3kPQMshT1jHefxvYg+SfFUmh2/9ssYnZBqKefkS3jAOYMvdxC+yrU2ugsJaFnVb+i
w2wMInMjvEexJthxuErncUuzzbM83BW0XjENmdm0YHDL3l2mD5SjPmlK7Yr5KP38YMQV8TeZA1r/
H2G6vlVHEYg/mZArD2O0D/uhxN71sa4zltDzQXXYa/E+UasPFwuvwNsTqjQjGvthvNFVO7EXpEr+
FVVwCvX1whmTEpGYfPR3EYHoOKvgluRnwlIfGfLXXTM0L3MSwVowjaRtBv6VVoe69i+en0WLz/p/
O+MzMr9rka2JTRuK0I0S3W6+NRxTe0jzECibggtNPOUEbCdQFCWbcK0KwlzJZU2X5iTNUDkOVwLP
rWOOUdkPefsRBUjoIjQyhNpgBL4ki4WzEU0tUOjf5QhdlVlqktrz4TvTCD1Ldi81GoLQOtfTi370
y7U7ArGE6Hc57s24lajMaaT+GtCzatAsuacRGiSIBp/6j/4d7Vi8fDrPHiRkQeOPjU3jlxnqHtPS
bdWi0vI1iGKuvqz9JawtVKbcEM+IzcTpKVWQNt1RrI3LsNYJyoxKdBSLTA5n2T9GYDXAF3e8Cvd6
SGNaZylZwpNY/C0uerR8RpS4VMHrQTDxEQ6GRvYGKJ+8gYeD73slb7uu0ZcefncRSyaU6Pf2HHWC
RNQByykexyTd1ZhsWtSz3nH3Zx4dvyZG/YaJk3YSJ7az8bL5PO11aj6ZEUAx1cN9jf3ZgjG0ADef
MCO1UZBlrL6FliF2V+QC92HXLyhXzGdV+G9choDp6zbx7xa3nzeJ4UMDF+3PhZJDG4/aWJkTxemQ
XUYZE6X9M6Uuj5SaR34KTOeF90XsFqKh8FpZmpz3lPYVdRBuc0aZ2iqHPeaUhXRu6ZKeOnrdJg+N
2NmhU6gfMPoNHepCCjqRiMp+t261xjCn9evvU4ouGakSTxlJhMyOT3ysujBcZadsmcsPqGH5X2BS
n3gMA/Valo1PmHXGSMHpm+uMvnI+6J5s7GeT2cGPF3nU8gfGxtYHsZ70xjc7/2VXWP0XUOfFSU9X
pwij3rwE8cLcwGUoTeM0HW0/ZmA7sCVnxVsXNl1zGxx00J42IiDrSyZ/K2iySJvSEW+qypcqzcBt
jzqAg20v1rhEn0dq8fQaZKooQpXTpNfECaUF763bfT1JIFunngjLt2FMmUwFFMDTGFNl2d4pFC09
Pgd39N2wraOFszULmX591e411fB7OIsAP27F1T0CdaNa1k0thCT5NW+7yQNLGh49yLYL1ZeRguos
FEf18RBXFutXGhCZKb/QzGAgdQVElhtVYT5Eqe5Mk9sWYUSUG80pIiEQuzUeiewTviL7TZsdTupi
VAzTW9epKupLR4gnpmUdDPR39l50PN1LAeHGSHdnmJ6FYGFu2bUnw9Qbaqj27UZQx/gP2HBMLjRS
iINzWQJSUkz1XpiSJD1fN+mJVmtpWoM6kdlW8HmPkoT9lVlFrxHJ0jbQR4RrRsYhbp/1+06hwqn8
L6rCsYMrlLRgSzw+LM4RshnFe9RNDbochexi4pGIbAX4HJKPyNYIFGKaT1UAVx/Lhr2z2JWNEs9Y
9EN+Kjx0CjgZaLd+p4hjiqHu/pf7rAxySjLkditgiG8qS2F4/+Sy2sJ22YLAxZx14emqjBS2mmgv
1LQAWnbAqvvO9BsvjvOY1owBrv0SYt8JPZawEBusKBKNj3aooLP1QxIbzzm0YptBmBWnXoN0mIYp
6s5aLgc/KEo+FY8EljcJ1xCEYygx3IPqaXSPbSZKv1n0zRlqYd3I7nRebUksuQnlgKkGTF3H4lqI
F8TyxBoXEMjplik4Fa4SF9+7BTGq2yOck9TYKLRcVGgdPHu0FCxCP7v7M5/PTMzEIhUKiGH4iFRI
7zbFCwpyXnwb3OxIJ7UJxAhZSoGXG3mZajuxIZYx2epGFAD4aFAnuVxP8zXUFUwSdTWciuCT6+Ri
BAkp0J4n5oQAWomc99iajMCet3QxTQL9nxH/Qr0HuSMeOH0IcCHW3HhItW36VVpbjBQUIpt6hGg5
MbTWfYpnV/X3bduDNAEWrkScMRiYY4McOYHIeN6EmSnqovJQyf41FKHMiroCluWglSFYsIJndu3n
2TGxOJlP88QpHfVILeWx39egRcpXemknC2YQEXxazsLgHslWDkRpxFWAlP8Uacn5722MttOyQyAa
vTtc+TzJoC1/1jMQwh015MEHt/zczGEjvbPPdfH1Y0VdjpIR3O7UBeDvzmGkVgHeuh31hX7Jp3Ut
CpwqRjni1iRZ2a74opABlVvz1sNFHczTf6107LxI2+7xMqnFDIeaqsam9+/8mmaFG7GjIASJyOEj
l4zkqlHeGkaOOIAXCW4wSgaFul6KGmMlkEaZ72/qTt1+3rGykzCq7xDXcE2hsgTLWv1xlKBr4HaW
DLOQ/NJGjkUitpxu3liteCerVCm8SxEmWXNAn0OWxqWDaJNIv+WCKMcElV9ZitAQhYP5E6IufCcK
v4gHh59WSHBlAjGgyYdtQkHgerqKPk2hDzZZvayrC0tIYLy+XC/JeUU0m/At+dLbDHzW8i53aEVr
ttxqN42dFftjpjiEYlLCTaxIyqmNB+OFFMhKtgcwq3f4wLHTeE93DdMeVjshefnHy9AwhZjwSIm1
Fz8XJrIhQ88Hz44yr19TVzQEobKnKcq4Ebz/DnBehi1eERgCmTZLbfP3qRuZb3z3nu59dy3LXxrS
A8fWjoL/jnqwctrB88prGwtEYzfEU/Xh87srk9XA5SHMTWPIvwCZ/9E++GgO7MI5EUR2DErUTyjM
bC9kW2p9LeSEyuZuPTCCWbTxiBFcXyvgAoSiiZxeUOMeVVqoKjpbTrhASHjO0tGAQJRPRhPbRkd+
t9xc0bXj/ToWids1JMbZVTlKbTgXl5xgwJ5ED0n3grOtuYtoroOP6gUPtTh6ED5C/ML+MoyCLreV
SDo4Jx4IRturg3weHPu0nYY10tnnZyykeRlfKVRVQPB0tSFejjRW2i92DHnIuLGUsh8uJsPv6GBZ
S+k4H17CYliyoJOCl3ljrWvyznoNh28JQsu5hpQrMssg/6wNLC3wIGEiSS4HLmP9vj8k3xc15532
/pfe+vWzrRyIXStwf4RZfCASb32ZMRASojjBva+TkJdgvjXa5F3tp3KTUKmzwcKeb2MLa5JexX/g
KBAtCBondC9RmOLSfeKiOrCkY6md1BH1CzOwPwqbjhuTfghKPtIdYHrD3deEL4UaRZDm1+R0PtNg
Xvg8yq5qgkbOapF8uRWxKS04kdATZihwpMhDJOSLzZ5vO6tQbCTul+0q1hKeRD5M9qSwzfxcPByS
Il9sWrxIrogP75MH+q8DycM7RQVSvxVdKNBXIEGZOskGaDiW3qwlifCFtEAYtx51CK8uohhX7bUh
VupIRlHkcleZnjW5z0EwS5nQnn0imks4floEQq0+GyaXoJWOmndqfhDEEQJgmYZNlvGGgSRDBFci
lHVKGYjvJhCio53KMomCjsyDKmXgUzzvs+PCyV+BZGzrnz/0s7xI4hQW7q+1Pv2yoHPel2hBQv2J
g6/MuIMIf99VqfuMPy9C0+MiGFqhY8JHzkHjLPlRthtvJ40mkm1Ait54eUB4Abr86UOcTXKtrhJm
xvUQqVf9iw+fDLFJi4+c83lj86fZuGSYDEJirIgMCED2MCMXUScsXyQO6hOMNeB2yA5elEmb8Zks
g06B5DTUtkhbWZjOpDiJeYCEMgpl/mnG6d2OvWFHPQ+e+0Uwm8GJWeMGOqtqlCQ9IWV1YHcu/B/j
nEsXSlQrX54XJprAQZkVqR6YadCvmwxUBmovc+XCkuJmC9LH25pf1a1txaoOZEa9lXlZeibIuleI
xwxo/aiCYP49TArN1mWFRIpkbwpidWxCXGAk3o++VzfY+WJDtFv9SortDxTiKHLlcw+I9g4zvsAb
PJG71iv0NmEViSZ/nprUiDONryXlgiT6NFWPWE+Ot9uoH2viPhRm8WmF4+6TD8Nh7//ag5qtKx4/
njR+gJZ1Hx4QG1B58gDm90a/WS5dlJs9GbVNg64evHF9Ba2fxEIlKkNaSdR/O02CbjpUzCWxsaiD
EATdBjBqI4XBEm8dbRho2pBbFagVye0AHmQWOony3Q/fNjyS5sj5xAZdRNqudYeBkm99uTa4eGL4
NavklKqAnvtfmHGWBcSBfei+c4qnZdYlzFOcVBQYYuhOLgNDqmBH1qeK1yafVLe9LzSsUQN4+3Je
SrZplPVEXZsLmR8sxA+eUASkLU35m0wCtLweJedog4xHp7a8+LfPTd1wlTHQdiP6W5b/grW1xkjZ
g4AVpzLmnrAFusCCluDrxkos9ZhZxSNbLdAPfVZVmrXaRLkkaX7vXdZK+20+T8VwCh5G5XRLffn3
bxEi5GQ7YUVmmD/+Msdo5zSOpEADSuBjSa/iml2gFyAv7E47VY2NpdBfz+zVWzfFGUOLSQX6z4Dw
4yMX9lRPFNFhNTsSU2BydZavDBAiL3eSmL0uZDIK41Qm+7Q23UBEB9/28ogidqatszu0e5w4fE0d
H1cvDNFzd1gtxWVru+xRp/TnDRPBdO4/369CSpVBef2uUIauYbrXg9DpBlLTEibkUnqi0sVy4I0w
FXUUy+1xDe2fWKEXEo5VFcglr2rfTnycR9HwNvCt6VTtexvf/7cvaFdq4/KQ6XwPiaGbEi1bBU7H
xHvxJfzJVItfZTUergFE4GxbZdzALa0iEsXL6XLPqAy26LUfRS2BLB0D/Pm5vpPfw8Rh+M+cg/L3
C1RIhqAezl14vX+7/fqLqjsOFleCGDnwZUdVdR3iUYBN/Ke/dyoLNRU6ms6QNleX73EYfSF9Epg0
gDL0J0K3MAdlqudriKqd8plBl1qmHuHFBie9P9Web/OUmO+CdtaNZH0u/4DpT8B93BfhxEKkpRF6
mWkAIdqa2tas891C+uGfFEzXomnUUb2VF5nY7tMVK/GeQOMdNRqjMsyJgj6jHs83eDs1WQU7rFZU
B3JIy8qoFtJ0VptcnSZN0EW3sLhym/eJ1ZfP5vu/E3oLaXghYd1qToRhy0ch93raEr+ETFWi7JCF
zR+iOZCGFLelE5Ewvlggvr6udvngmqDNPtdZIvv5RrzvqLOYjGA67Ax9DtM9OhKCSSPq8NFKMBWv
jXBz8K3kzt14vwciBR/8Hjxev6vFnX94WF7He/XqvVAQbUTCQedjCFzsmWjXighcKfpmefu0p9ME
Yrj3bENDDnlWA4lG4oq60Er39GM5gQvW6Ty8zOjAtlfR9jGLJxgwZPH1uFRfC8jWyXj/2ctKn4Tr
QwBkNxczret+TwzQcjtnhKEdGdd3RSLClxqUIZiRraAVBjTZ9pjkzrBZsrp33Uvs/9qWCDNxEmsv
fwSW9ZJ+FSUXsZUbnl5DXyiMrEIyroKxJKdM9VJ8iLi6frM62IIJpB1wMogeYkHYoaoPOPhmBbXt
BSaypkPinxPEMSxqU26tem5qsKbUHHdFioi/3fzk9oQE9U4VSauAG2ePUFnL2d6Q1T1S2RKHTPLT
sb4xAGRE1m/qVNJOAulhrPzD7TYaEDPKhmAyt7fI7tk+L9r+5/HT+HGHLbGK1AM20+a3W1WfN3xN
1gxEV74Mzm3RIk9KKwpusIH5e2de1Sa1UvxnT6ksJgy3HTqJPlKvXT1dHCNCfaTXqd57y13h7J7M
P9VoZ/o/uc6O6aaB2tsI9U8xjt1Aclp7dkXsG9Qma5fefA8Znwm93LAt97uxX2L/M3WmSV8wtiuk
gIKP5zTVjRi04bn+HmNr4H+qybSJuoXgeeS98eB+8Wh2b462H8btD7GLPYqSfzseJPvIkHQCtmBj
zHdJws12fPqaq6cg2m7BR5Xp4Ty+8spkOGj9Z2+jzvJ6b6qvXGMKKFoPylVnl11L+35NV1rS4sb8
HtadidhEaQ0G+f1MYw1Sc/aP+wu6f1F2U/O/jpWt2dpomudx2ZXLLY0W5no9L2CpxXiI2LF/QgRv
9S//UoYXKg4Orz/QFLWDDHFB7cmA9d8rfjGy6XBJO1aiTxPW1uuZwW1pHtLKFXth2/TGUphl0t44
v4O5Qom5WjOHCdb02Mhm6PiEtPjuE5g8X29C5gL7LoDcIxzrVKpi1QQIMFj77x9WEu6zRiYpdxTg
PHRdR6HDjPjQgck9N6/mhhTvGh/H41XnjkicVSKA4J8AfGearyhBtLKqtNtHGMjuIMRFaeTGVK9i
0ovCe+axkKca0D34qYAQAqa7mOHqqc/VlfQX0f8jKksUYt+UyWSttM1dGZX83Ravp3Hsi5/ps6Ko
D2ls0dhd0UuXMzkPtIvmYih+mQ9SvOFsrMI1W8nWkQk8rvoUOq1taj7ikGE3MQ78V1DIn6xRQMfd
cr1CmYzF1UM9jPB6MvJYEtqw5udnWJHrG+s6zWYpSUDSReeznaRJi9rYJYPkFIhUJvlhxmum53dH
OtYRbbRHPfPwA1Q3Bl2HZa+yQxNbZIkubvf+9WXIX7bvwNQ6Fq8Mje1Kh36yIR7snxpUJnztexYY
o0YP5vxX9zsG632v5DIIGv9mRW3mFrbBlpyzTOje5dLc7PDLd8BjeV2m6wZCUU/0Orx+/a3cURyL
AcBuYCyT6Uwyvgy9HY3q4Zh2s8sShPtealS7xbMnMmSuAoha+x+3aiJW7HCGTl3e5+8jNgm4zYVv
4IaWpW1Z8njc0aKVA15iYtNzpfYJf93kw2FU5iV5Esl4ssF/RUJa7QgR3M6lYG28DGcXHNWGNzb0
rEMU5k6IGberP2OeNNwOwciETJ6TtniPBBIn0w077cuCYIAoLHi6viATHzkIndsJZV9dQ3nFhm5q
OzKauUxoGETfObv7oG+lxENzeENAEnhEQIz5FxbB0r/iM04O+q59b0iojk4ltsuHIfS6MACzTs92
cbr7f3MnG5l9o/noT8JbjnqwypJhVnRVESXcGpadJI/HwW6vNsFg7XQfm+nx09v2wIAhEn4t7LHP
vFlfIrIiTq0EgyDNdCAKrq4YAKKwpCsWyUJ+NWSErrc4eQt/rP0Ua/jig801LZMo4hFH4pZBzXyk
oGcGBA5vaG6lUPp7AeTqPITzk6g9T+IGmFa37VuZXZrJMk4gsk2UMI1GzjPxUwHbw7C7huwyIENt
+fSUWFG/VvTVFMfpSJIvg5kBjTlC5m7O6/LoijvwHGgakXcvD7aIkR6abV5eIGip86S6yID8Ddr1
fzm41U+e8BfiPO/DUiLNPIx3XDEKP3zwprCEKEhoDOWgrXa8ZQrdLzx3rfJElTsZBiGqYxBFYJ0C
GuNIbS3TvpbHkdn8Io9kP9Zf6lZkDe5KWhSOhE8NOKhavPFtv9ZcHJdwC84cE2z1bUtPqJrSeY9X
Cr2Jr8TjwVIFQQnK1b1PGuAHitNoxxlDEJRb8IzBZrWyRSwZrnGpihW2qifx6KFV+h6zAnefFEcE
yVMkI/JhzP4hjp6ZA6GGmO1mT1+7goNmTQ61jw3NwfQOqjeMNsE5fPiFIisQCZNrpZ9oUwZyUGpS
tcnCFRvWAi6PtX8JEnDn4bo+Xcd4vbVwVlWEdd5d4Nb+RscpEfr0cKHmHBmZXst+rew6Ld9r3oMN
LVlOFAeewTkpmHBM4K+TJ57oFWMV+UgmWPEeKfU7x1rhiq/I4geJaWuF2dTMyB09gMeJxkicWFD6
Xh1xhsRIyWlBj3jAZox9k73P51MSvxnyI9aavdzAeS5excilP4zXCAT48nuy41pzZaXR1N0mNyrI
nIBz4kvxP7palvZSwdG+ELLRHRGMkzcuSD4/5vsFEQZcezBcbPluOf6YwCjNjXEP6W3+Rr30ATtp
ptW8iJ9dhx9faTWbysSzh7Z+ZPVYyCQ9VSuaWCOO/04koUUMWjZ6Vhqcspw0nL4RMxa0PkJKwQhF
AwvK/Ig27WIKpCrEgpNyhJYiCab1yMtHOLius10qXBgQOI+x1i8DRHx00HNU+OIi6oCoFyGF3XQ6
45qKWOQj3lXhS5pOfgOrTO5MJohhreQOA/dobZrunDrWc3LGAeI1vmq3H0p98CxjfDxWoP5dPYd4
tw5OLs1fSXZxZIJJ0CTe8996z4VNdvooxCJnuF74Ckg/hCr9LTXVScrJQZS2nguGOLFwlM/SY1hC
XrxiJQ/TpAiuLHm7FRxFIQb5N7CaSqZMauJ0KN0Htm++69smZTlI1QfExR6+z+nQ1Z5AuJ1MiGWX
Cq07+17z55Oj6bFAOnTyHT9NcnIN6ZgBI4mvbL3Wpy2WA35eX4t0EayBn2y1dR/5D2SEldPtESyq
G6TNFWq73dl7WhcZi6IrIjNDY/cN01sUCFIYloI7EHqUeqdAxVZO+FH1I3JxLTGfusT2HbHB6uZ+
fU33oVZNnnc9EiNRodcdjXz4wHek30dtL5o+QLQd8oCdU/GLpBBH38tjTl8r16pgMAbiOkwSr07Y
arAKcT5K0LwCCVSuV0Ur8ej10nv1fwhHQCHWumORb+cMfMVb7OEOVLg5pNuD/0rkr31IwGjrTuxt
gcHsgobFT/REMTPmCv0CTp/nOAcH4MozhJjF8u15K9CF4115EIDuhPGOYIY6U41yNHflnxzmsgvl
4XAlPYDZfxE1VscC0X0pUMi6TcS/qbSLH63YPYRqW1hr6WupazWJb2o/S3eb6uhrMrr9w6XunsVn
73lLdCnNeKcH47jD7Dzu7924a45x2pjob9lDLNQsoIJlsO1dXNjYNXb9bdCg0djDOKF0BLJ2uw39
sUKBRLNsWSYSWqwVJi2gGFEMl5/fGMzrxvS8OCuvtEAfCZk+u2H3ZH+n3tim7woyLG/dbd1LndIU
ItZ5miCafcNdjjgo8ArkRFpb2hVed8JCkTEmKOkRKtPqPs2uWLaKSJlD/TgR3EcBxzN8WEihpAEo
SWrp9mtSkBuIRJGgM+m3sRsDi8+a3v1MTxt6ZMhXSn0IVOGA4Z5oJVYGCjJ4HSXTqiBaSz3KywwD
NZvdEwt/gqXqZK6J4hYZXKp4d4GQ2Upemto4ZjyaS4U/6fdh6Wa8E+rZVXWXre6hfXmK828YuMek
BwpDThYZdU0lIXZzh2yB4MCqahDggBWnFonPQAJhv2LvFX51SuhyF0RHTAnJPzoNC6xKgcJy6jvb
VezgLkKHioSSy5SrMvNkbqWx8S0GLkEXIYqxdL3pFehLhk3uHmLuRJ0rpDuHv+9X/mcnrUzN26nz
Lw9tyzP5nzMefA+ByzDoppNU0h2poKFfeQc+4stv/owSe4ega4CiiZx2pBNbTTC++yShG2IE6ra6
CFbMYPr6K2M3kiuabwz8r3G1MRUOV4JLRDMYHPIreETF060jtoCXNEgdpCW74ykpK3enWb8tA4IT
NQZwpxQ/a0bB7jmdT4KuJwhIsK9rJ7x+jTy91zD/TqQ4pGgnft1vaBP9zcUBtRsuzL1k/zayY5H2
VCnyLoA1WvhPfI1oPbB0r/ogy/1O283QwMN6byMMSKJ5GvetsCM0ps3PaMHoZK5RZbgc+btQGdZe
HzDj2HYl5MqObsKAI/FWABQtp78cypQPejCnGuxCyaJLstFBGJrYXBsn/rWavMi8U2g7tarJsRSb
fVku3X3iJ9xgN2jbGf9siADIGontVNVH81bxLtPghKivrshVHP3+vQ3wViqeLbo8TArvEt2JYdfR
BhGfwnllfIZj2zPGOD02/Tf6gBUTQPsWaPPWdeDiYVrC0VjV2kIci5LXMbPNXstxDAqXTjukTzEm
nwegm/5zG09a3yqfh4sUqULkE3S1t1nER9A181TgIKE6asMFp3+ftv8LZ9v26FXhdbrv2K8QZKG5
69aKjXVSJ1Gd6+Mfio2QsBlSCth54BeTQayUW88Ik89NJBth7CCriuDU1UczvZzgCvJR0Rh9PALj
Zt0OVg8bCF8qT8IPThDPqwNvLPptSF2UJ9L0Pc6DgWza1w+BJfS9tmQOvEqk7szMlIRf5Uu1C6li
yr+B/kZSFqR6euYIhKx5pnhCRUsLBoSufU405WUNv7E8MHbD2Lf4beHyhoueLCIE4QQzyTKMUguw
FCMyIh3CXqEVt9bwCkHr6PhyPxnIE+R5qPZoQQ3VwfihxWKX/gF0bhqmAOsAgGgbzUSeAE8PxZTZ
FbeaQATcq7dn9qd51+o24gYg2JjZLjnGG3gUtwgspqDJfXs/fqeUGwhjNxWwN18fI38y0I5NbyQ1
vaVHA5c2orHXflHJILvhsZgfoB5qhbY5Ri9wdNWyqLxUnkg9Ab5eIeU3yEUAUTozbbj0az+BvqE/
v1G9xJLw511yXXDH4GfIwSLUwfOpiJNSaB9o3sTRvb6SO3zZl0WHvLUo0y2/FjiBxLlrOkwcUdC+
FQi8avDrWJrFGDGK3ph6E4REvDDQt1hE0Weu/aOCZb3vspErNlyDJzPT+YFd2WBmg932GB8U6qQb
jf+lzhe4CH89jNWgF53bOqHVUJM73koBxWY/vy8MY9H9PYx27+EXl3tx0lJFi6MR6fG3caiOUC/+
jyYhrt+1iK7u0eR2xpCCFPrSzvqe1WgFIOJ9sUmrIYjMWlPMnzmFI/QBPaM81/R6Eglk2LqvQMxW
w0KcqEAXBJEIZixtlUmi71PhUnh8s6QgSUHJ9N7x/LDCUfaDSLoodt3pBMPEaXh4yoWClUFdBtVX
eWIJhNMh1x159DvL811Z65d9CPZRr7SnVbamSDwnQiNEwM7UjA0RxWEcSye7h6np5MX0DN7fJkiv
vanIcFLEWRfDKr87DAYUqWDzDUimoYL8t6ok0ZUKGxz+jOsFRrSZkYCUFuDgXjT2n9SvwFVnhHPU
XsGqwaYxOU8AGvNy8MF5qt7uwLpbqMwiSDhw9pMehSUgMPSOMoLd/8eGP9gMfDCQe9uYtWsr10Fx
GO07S3fvEKiI7EKTZ9UqL5XWd4XRv0K180eXdmrrX6rOuUi/TyDaRgVNRomSLjg7gVlveDT5Jzo4
WxxazVIKR4+XQgYhxEZx6R2llZwhNxcooAV9lBbTgba03Z5QbuJgpoimw5ZWby6J/fUb6esSHiQn
q/m/ahEv0e4EhRD/oLfZ4s+XkNWm7eDARsj7Lz8Hdx3ZSr3pz1MEaZWB4eD+31pSC8IKmpKVywBp
7cpwnljzuyJKAm6AObBjDYaIwSSRb1j9n5OF4jXTympZSUMQePCpeJWs+EjjcvSxdnKjXM7QWzo3
3oc/jYBaQO9haYEGLB1lJoJSHgFcUH9VRLiaCO+oGOnNxsuIHeFWuQsNN+Rxud4z05MNLbO3cs4j
5WG0m/s4D2jxOgZ275zuiWku0r001CllB9yOFCyMIOkNS72jHRXeIp8tqijwnWvmD7DIJMaGGEqr
lGGrCcGCaoExxKmc6bMGLwCjKlwg8C3tBGX92qn3M7ogPsIH7s+frc7YV6uVVVkuFNuMBUSNjmSm
dMPy0RoIjN/gKN+eqfmqIYS0nqyxvvkWAcQR9K01BZDXpCGBT45H4GZCSLEy4Dl1x+Y1yIqbOMs6
uY5A/YC8VkZky/HFF8oVeLrsZYgc9iIWA5+plt33XNSj7hUoygqYap/a5dkHVwco7UfjHC8wHZRV
VURZrGumPPaW21/NCugB/D0Mg131045SBjm1MX9VP3QMSbidH6C5AIxGu9QkpOESFLj/GfgIvw/q
++5+qDpU6QNmydObLmhLHKQeD1r7Hdc+9TIJSvYGS+fso3u075jUKDkoMRJnYDZM3jBBjv/Xyksk
mJ+4fQJr7uhL7f9kI1sdTRs3EO0bB5COqu0jRze3C86uVJBoVO/nOGqR0hS2kKhnP+T3u2UJYeMD
94Hr958oWyW/4MGbLmrtv9f/dOwXRDmIKyd3TVoaVy+mGEeNxNRyNtKpu17vbCReS0Gb4KdO+vLy
ghQkp4+CBx/25EcthNqBryzdLC5hagJha2w5m9Cv9WE41gNg0zbE1i1MX0wAaMN/52Mm6O1Nf4mt
0rbU3KDN/ySiVsEzgNsf8BTFFNVj6kCZAimWwOXXr6r2vveJCfZ8x50jLB/9QF0T8VTKrz8sJiEV
1aErlTpdQLeGdf+tH+CytBHQkBmjYY5rwWHxiDNQLKrcyCZxCLv8rucHjFX8AoXoKzv0aFOZIAzm
EWmC6ACRVLrSoaxfkc7/JNkjNbywVoo072DHwwFAXLyd6keC/0QvFLq2cy5KmVTjzlyS0kioQuCF
Jt63d/TperoU4uLJ1QxT3+3Z4byQqbT7/EbLkFz6ZwiyCMDA+YvAvPd4mEsRo4bPYc5g54b6gQRZ
PTe1tspjcTSDRgtHXnoBhQI2gHWOx0OC9fLGZXj98ABdgihmUeQi5UTW2Xb7KnAMy2CqsGSVBy1E
O4dFB+imlM4Uh+NgOrmlHkC0FNtQ679NqLRa93iijkGLO3FlfywUQtQJPfwMlpxGzl6rraxJJFbW
73Sf5OuBa9uRnjaPlUpdCN+vBNYAEa1xqLR9E0HV8yiYCu6ZQglKmVyUisBiFz9KVOlQf3B2JH7t
qNNt1G3fnoKVFZe+nSl6T8JQyPRY4oYosI69HnXqvU3vxAotuAcO4DYww3JPtmTQBVBQnbYBm1sO
qXEmbXEhpgYm7zdFiJK9kP8NX24ejT5sq6czmkJbyu8BvN20q89/H2yATsYAfK2SfM/9HJe0x9kg
gGX3+5qUCDQYyN0kvAw9EieMkzubJPXNLcMXPUVXt8LGFUueMJOyRefKgT51GlW1yxd6n2MCyDEG
iEni1uFMBv6N0JJ8gUfVsvK/5LfoRZSamgB2xf+cpJ8PJlfICwjD54rveTtOdiwQPQbsjEKa8QHf
C0c57I1UJ4IvyB0Tcmfh2gl5t1eP8JHxvRuwirZbRLJhWhet+XVUBKaXMYiSCAkahXrxRcjZj/Ou
J0VAgkGxYhgGwH1/DHduNbRT47y1B1L9q5iWNHO6YYtQWB1k1ze8PKjgSAT2hRLWDZv4WeyFJDkJ
BYxvSAhSQ5r+hjk21nqWjfU09qi1yVxCWFiuJ3fipz+lcST2GjiNkdABqsesnZxQWLwPfkgoZUNq
LNN4AtNgJnF5GUoz28GNSEsoHmy+jFZ5hp0Y0KaFLMqQQztIOpfRP0sFRu8x0+NBFpOiuopc0hOA
eBPI1bjCNI29YPksff0Zp/WiEbBuhJXykA6dQ+lGo4uS4um3R7u5/BjBEwR1XWgxfXBkun3mYLsX
++Z0EoCUhNp2jPgWLPC4CNsYOgK+Zzw7gfAe/9peqCSplusnnxFh33g8rOZBuTj330JCwUPvQrmF
NgnamwnhsfoVZ0I3n6Ab++/Cq56nxI9t4I0OdZ3bWgVtRLX2SnBbC/VMIhbYZ3jxXu3k27f1ArqH
WFAxt9n6z47AWL973t/0/3UNej/SnD30XbX6D5T1ocr1jEF/9BIVKcSduUiLVz+DTowCkp0MAwco
uLlQQ41N7nJltQr83wO/pPyntKKwII/JdLw39TsaPQLsmzBhXVEZwSkWiW29uQmDqLcM3agUwoP0
bHe6UqLYyRugITxi4aeE20LjYa6qEJwoynAttBsgWdRnSQSFoHTdDZq3MGGXJns4c3TrBde7KtTw
t0gFK+qUBTlvAjqSWBYEQt4WniKccjCiq4n825rl3xSdVrbB8JOkyS3N5EXiuWPGPc0LxYivaeD4
I41beZIwVkuqnitFZMoRySogqES4THUNGEUbq3uCel+n9HwBtO0ktyQ+tGUIxxHRg+3r6VOybw1u
WG7WJxOEOtYSQO+k9mJ7EwaxF494TIHyDg/RtW2ojp9xVHFvRx1FL6t89abSqudzJzM9BhhgPnp6
1D/xRwr3fiwKZ+pchaBztThFodsR3+fhQk2XEsjNDuYwMpI2HawWi8fxelCLprtc8k0CX0S3yZKD
HuphMGExPF/b1x8CKlbsIi9qsEic3fGRSgC9P7/tAOtnhIxCiRLd4kFZ9n0ICXsW4jyj9wrkzpmp
uEm0gkWh2lxVJVhOe0lL/cyZ/S9VzCM4xBzcl3ciORr53zkbvl8Be33b/edug/3C+oHtA5PPticd
6PxBVXwXU7QpPWR7HvnKFt2HrDjD3QM5mnZicqW4yrMpfdwxDCP45LIVEOELC3jn5eDrHlNnJ6L0
5tkUDDIQe9jOjcE19ANrXWpKZKV/3r+mpM67ncgTRoSOM+vofyCN3Ez5njfkESwZhhrWhWNdCd7b
WnqCD1KU5f7ThPIA5msbJxXEQjM1SimP9ZfpZ/g8DN5vbNyP9KoJ8rXLldFZe8At9Eji3bHqeq8T
7lYJs6W8qQ8UBrwOelJiGRxmwxXL1TVoxBM3vvHuDliWxNfxq5PN0WIz4guBhLnmuAQT+WFQx2Lw
J/HNp0yZ0ltNRF1RUDSsFjHwmTfrdgg7VTTmjUgy+LWptleLbHaN1m1FCSByZoEF0h7pnSxgI3Ef
sHIG3BfH5tXo0Bg9g0QbFggZKd/mLXZaT6qSlHo6DeXDG0UtjgjqMrtjxxP5zR052EvdRYpRv61C
go0gOLnfpucrEovz4kDIprF2lypqbQG9AIe9rlHq5GbaXII8KIS3XuFFRzZOVSzpc9vGsOumutKf
a3qw5HykmW4UBsABmXTo6incALsXgDdhGVA5t7JAW0vNhhqLX63BCysOFgSdCN062LDNKc4vhXLP
t+nRfRXI4s2MqBy4+BOwaVsl1XAchz4OMft8xnJsT7aA6R2RCcR7rdzxnYG2o/v+irztBn6ah8CR
x41//wMYaLlh1I36Akzi/aov6KZIPYLuh1UdVWlL6Z8O9NCwjZPVd3GKGj425fEYCzFXSdznXdr5
5YFXQQJWl476VwIxKi8AfOUb8foHGIKecwLcFX3Ka6WUhz3wI/vY+3eDLgUpNf6YHGp4GdM4RYWs
hO8M5HdsImeCGshHJuOWIcclaWhEdhFEsaHUtsUHLLdCOnSojovpd+2JnxCGc/MjZhERrG5mWVWy
uKeK5qVXYmNg/dsDChDC0YMPNPlCNwKVDE2kvsyMdKIRtjWkKBVtaKGNFhw8PsLkZ32ljVqGUf8T
n6Px1iq55WJ9i4T1zBKy6VT9t6r45xrKGkRtiXDzqV/IoczfgkbJxtLHn1y/aLbRbvea/5OlU4/w
x3P86K8fj7hdNV67mqeuqjn0ME4IllAbVZEZjeGRTplW8bVlBRUEzmw0eoh3eyFNUpR+S9S4Ce+A
z8pJqDmjPY18LVhAhtHk3d4W8GCOLmwtIOI48mx1YYEmq6IbOqD0TRIDsVHctCWhONP09czMjOY+
hfaCn7uKkHFoDo88xKBSS8nyV6ymEHd2knDnhgSpKMW3DdTaRZUdjdS7ublkFxMk1Re33WUKd/om
MaIhj316ePM/F8ccsuG8OXN7WgP2/Hoit3755g0fei/MFun1aSWXmqkCt2VGyOW258f3hY5TBi7s
I+Lc7NjxootmKVSPoG+wPYujLrtSRtYdRhbJyht1XhoQ+f/N5a97oHhj9h6+u1E6xiIaW9HiBvyG
62ck8UbqUWxdBbVdiuHgTYbkc8M/VkA6bKbGaJ+f+yYtIRSKRlxeinhvQF3tB2GTBCqoFHFZks/r
n2PTwIlP6bW5QGWPnK1nKZY0RqGUH5zSHHbDqpJrJHHjkIxgL0jbtD+xx1FJ9hmC1UPgagD6T4+K
fTYfHVBu5NvAnrR6UNAmz7+63PIQXEREQ0HKv6RN09puOUZHfuaVVBVOz9UqiG3+A2/yX4Y2gWLN
nquexZVF+T57fYlj1h5EFvF+817vz+e4Jb+uOWQ2wxm4dVqf/fvQbesQL57MXT18vhZeP67rlS3T
nByPKPSYNQOzGnn6X1wkVtUmH9ZAhy4RWx7rGM+a3qfANNMfrAq6p/dsd5b4IYPVefdEun83KJoq
Df/SiZdXsf7rseK/iQ3AQz26MNuf3euWgN4jhVLWTQd0J1RyX+R8oQhbo8KjyQPFuHf3wv+5FP6N
DkqPXigWOZcYdjlx5kn/HZWLmWTFskP1o6jL7eSX2sz9ad9ftH60Rmwg2cvHAt4LX7zrIqEMcYmI
qGaM/EDPLDeVSPPTlEuhFcAD3oNyUug5Dp5atEDNWzncHgff9Mi3JXr477RXGq/M9+z03YyBpZWo
Dx5yvDY8OfHF2MU+d4yanpWiFxfpva3SYta86J7eP7LyWtdE8PnH7KFa7BlzvNLPTCPcH8auQVtG
SDlP826bvFMG3c/ld04OKtu3pf8FXoI40KR3KzeCCBTXpOYmQ8jfFT+JLbzMHPQhnnTAIwCix7vk
e7k1HivxvtOM/ot4BoC8YZEHTTmTywP9cwap403Q/xCZA4U6UO0yhrJ5agr7a451PFPSc6LS7CGn
6x1WhQ0LXIGFgH3JExlQyZ+z+L2UJ+aISCpWMPbBrlneCHSBM6P19fsCGjtEWIEVD40i5HkpZVyM
ggqYW1uUqNJjD4VO4dzPWkNDIl2zepps9l2SZF/3WjSosiL9qQH0e7LexJKtGTemTYv8Ojb0RWLj
39VGWvATIcQL0fPFYJ7Bw8MQoMNrDZNwCyoKPcawtK6Ai5b9eoPHy8fYfbEUqM/W/DdWnlZhVock
1Zq/brBqvf2WbP4uogP69V0BrmiyqhMWcTW483LIIRl3HBZSIKTu4o85Q7OwQIKev4X3w5j7oPUS
Sb1B7IhQhK1dZ47L38Rb3KlObCwBW4TeD6KYZkIPHkxuYRpo6ROsmibW7DTgLRDggogM9Yl3uzUI
/ddpsKlHIjOzC8Y/JDDoWBHAKIVqwwFXIoS+yeN5+6E40n+wbD2FUhhUApzkaLMapxJukLoi5JXV
vcEFxm/eQorLtgOL1UXLPE72lI71l/JdN1lWoBgcl4dS81ui3Za6TiRnCf8ChqIdewIdrU7u65PP
Fb7Nv1/+9f+kyCCy+NsS1E9whhfcaaB0rnP1qTBciQEX0hH4cJB0R5gLbOwP8O2nZClXzYDMp8Ao
yd2G206HrdKJ/QKHKOmbpfeQuJ4T6o0X7bxjUsgDq8uuZ2pSXp9HvrxBRaFQab6r20P2BMB6smU6
U4s+X51SKOYoRpYCurh2G/wA3FvI7d+Bn5ZHecO4iQ8A1wvh7Bl325CIM/J0ygyQG6Fjp32qZNEx
zNoQBKyq5sVG0yEP4UPjY8o4Djv89HGbV+3lkJlyFwE98PoN0j6OVS8bZDhbZbjztOXHR6+xG/l8
1Hsww25GSHLmP17q5kRZae4stQkyfqgCZ4yF8zuBgTpjzlFEO3PaTvcW1/3jzIcnzNeXx8J6SKP6
FmCxAbKqXVJ7UVHV/hJSkF3IQGrOWxUr076H7onebriAwpOkr29uQ4lWt37GxDq8ZdCISavKscdD
lCWxTaz27puwCHpIyA2t77sDwjfdh8iGQD/qbi3Rz18kX2IToToRaqT8z3Ie5EnPw6O54Or52T7m
IdXzLlkq/82NU2kUOMB8Xuze0TS9M0xPaPuJ9qpB1Da+OecTcynyR5GvsRpenYtvLteCiYTK1gH7
2h5oUZLF/WXZyqmCMpEwwNBE696yRDeXQg11CV8hWw7MoD0gn3ynVrJZnOLI1HYjTmMHL5mn01xQ
IsLXkVSzQP+uIDLWGMtSvU+IgxHEaPhDBENU3JcfZOqnKTxUfvG5lF6b7OJaqu8lYCGKv7MunQqN
l3yg2sZvP2SG3VbD9o5vsIo5iLxAa443tW40sjZHqiLEXaF25DA5CjazO1Ndhr0s4GuxFKaMbcGS
5DiuLVNSDOpJ7ICeaSAITDfi+8RpIEfFFHI2F+hgEMYuJbUnJvOrR/sLO0hFEQef1FNgAUH390G2
JRPSMwiuZ74+prdJu5pmuxTHb9R5EAcDvruMbWD+Ir9vUPukohm4r15XF2QrBbEqhtDxKNiX++rW
FC7rtYyt9PAHktW9TVxaE9bZ3+drv0qjkwnf+sUUPaq4RQwEZ+iKR9BHInYJ7Qdql/ctobxbWbfS
idpnHhzaPScmmJK/RK7JEdIw3pDrKTFXVV/So97kLUu8uHgpAavvPPAXY+IuAQdF/PLuqxvLKeEj
GrXbIJIkaifMVGxt7Y105BEfCvOItWSAPZpWb9T6N03FPNR7Wt/xrV/pvBXUjXTKaeIkRpLBvI+J
Ly4dmIJY8VB7ql3bM8RCzDz08aWWsgdogOuVSpCv/XLQ+LQ1PNtTA1wFr1lEmCmKR0TkFtI6CMea
BK2UXec4FaS2o/xbGlFf464FSbQBT6Dhvk2ClLj+UbofUTi9uD4HkU27KdQZH+AySnFUuvnumHEL
4ImwEm/v77x7HRhrbZWU5WIRlGT4y6zeBdtuJdrXt6BJVAFCn4SBUdaCROQH7YRep41N5Kc/cECz
AkoYYLSmixs39YhkPgrGWfNZfDqSs55foqZW+eOspDEbj1I4L5Up8Y5AapoyLiBw8QD3CevOFG7w
+jJqUaGdfp6H7ZiUj+qOxB3/76OeltX3vFekrXGGDids/ZR5WUb+lqsHa0E0z97o9FLjNKE3lc4C
Co4LvkccmU52CKxQ5JPns2pexebMzKf69C+CPmmibUZ0cGeGu5uZ6Nrzj16Z679Y72SPsIKjWoPf
/KNKp3Vna0KXRXDvvoIFubXmh3hSVg9J2x3nxnENoLOJU5gW4EuwX4mETJsl2Qwve0H8wILRnCIf
y59sQAP2MHHXha1fCD58YAg21dR7n4e6CrtaidJ7odRQe4Xlk5uureT8ZRqPuHGnS7XNpyCjonfl
npWmUprXCet7q+PLLDo+0XrvPpFr61nG+qNfs77ZSSGoAQA9vCDBZQyRWh4sC/ZfMNUk5A342+3c
S/mxl2vPxAI8+X5syNljFluL3IdD25i5V9jFfPiUbw9+iXdQJoZ+ShP534Q6nCcokUCKG1NLKmaB
83weQW/00XPTMDIdG1qTqs0dNv3xU9HtGpO7hSxC9wJJAMPiuVcxgcksJTGog+3s6JqgWIeg/vI7
5FMFr/tbQ6TazA9PXheS9T7fNFyci9xRVCRfufieJdPKulEM4B0Qb+haX1sVz1oWlt2CRz5E2seg
Cydj5RqU/OLO8Ltc/gZCNDvMMPIE3Ke4tOuupv3tPGiQi5wcTKpl0C7sa7jWCIVcie12G6CDbQBB
K655iohP0BvyT4jDJ17RFy3Tkq6ljXBdD1NGxTTS1h5fda3jvLV06ZYrXXS4MThIQyYHKmn8lwmN
Bn/U+mOsK7PB1lJdGytpJcf51HGZYBoRAFIPH7w7wcUgzm/+RB6AbGXVburJesk9eQ7yji5ffQ6Z
xVeV4Booy8l/8cMM12BBkteZuuFj3BaYkNLhX/gSA2aT5zi0S0FMPbq86w4+CPpQq9AdXwAgUqLe
sQUCDctCCbPIGn2kkS9eQDwAaQRuSmMC1gjzD8ry7XW26cDY5TxzcoghA2ycyXGp/InFHISKJPAU
PlLi7o1dFIVDe89tTdsXfwZ+/IfKHYsB/bHEtEcVslkagNYvhBoNlLduR81qIjupSev9h1DtmYdc
RWFTBesnvqizJHre6e+FngJxivsNA5UX9dkgX0E+Kc+WgrisVAYconXBTtqBnZqlfVpzrtWj/Gk1
H6IEp/NjB0ijtykRxm4/Z04pRZXmordcoCOMEmDAfdmEzNJVnI1NvdDYgfoR2RZx10CcKOZuuHfN
NCKQRy63zfuZBRKyiM2aGU0VVbZ+oYtyGttEUJfzv33vyJCCZECOOrlLaVqr/JzGbqLYiXvAjThj
k6YObwO7FhQDxAZnubqiixrbSTQ3Ruv6pbLmZk7OgHFpJbpj1p8W5rvYYbnnapxsJZA3HqhZJed6
LQdsoGg240yWagSoeQz6En6+sc90D0ToDm3UvzIP8B/svtyTmKb1d14xrH/5Y2UwDmG9vkqikp88
Nm9+ZreyUwRVnNWrcGO0LjK6CDlKjfMcT/OKe0/jGKThF1ccHwCcsAKsXpO5JoROa/rJmSXxI2LE
Ij5pIKWMHYwPwuNI6XXqhs3jBz3CMy5cFnpgyf1n3NR4MxbYG6dzweiR0Jx0wTJCqAVj7Aj/ZqCb
N6wPtKD//yLvgU/sAEtcHVcLN4KYyN58wF9Rnbp5ijkryMTlZ/kSEkQkVH9a16RE3yBeFSWFbT7s
D3WNTDRI2vgZHPyDkVfnvmqzp7l47RST5Fwouyg3l4/u2xpkxx6KUKv6ckVkhUX+Qm6m009iclyV
4kv8I+5SlJftNMvzb83Iow650EAn3rIZuKxanGiKI6Gu1nS9LzKebP3ba/5PLXj132jyDcBtC0a6
ub2si3CMzfXE5PT0wygQsARByjnWcm8JmO8hLLDeyY/TUQq6/1BxFFljMN4Cq6K7uuWDeb2Z6/SI
JFSBmw5TZc84VlWW2HlVFy7WqVRDbXCQ0TPSJCBpYvxg09MSwDu7AzatsYZb/I3UpsLVE3gRBi0V
xFOhKcPpoJMrAZaG+okDgMA0hUiAFBvtVUUwHoWU+WfMRBeH9EeYPILFC2bznc7+/nARO6VsWoMB
7nBUNIAFBQEFDObgydIa0Uor+VToDX9WFvj4ApObA191tCDouV57gpD8JF0OXchvQp6+hTX3fo8o
0nLA/b1ORxPgz8SF4wZPW37JPPUeV8UA11nOtw566hcbZzILMP9J2v6tFAaqC1q/0YP7Me0CY90z
ryjZegPIPoqsHSvJjuA4Fv99YLqDTIxUXisziOM5lKoXhOV3mLTaekFJUsICSCMYY+GodTcHokh7
+D92isn4Rn82Zrc5GqZK9M9GbLv0lNC67t0fcuCX1XixPnjVOIiFcE+oHIv6dTwHt0k2byejWG5J
N5TbOPDhC8pCwK/LYjoBa1f769VDR9rT8iIIerbvfZS/gn+5HY952A8+FGMl54ZA9GbJ/UkeKEdd
AFUVrDxh7r6M5B1LKkOyyXHONavnTsq8IwRkaGrN/ffsZ4RLo/+ox2oQeZqEtXCRsVAUPwBetTir
SqeYiEur5uNjaaVzh1MTg8q2o9IBlWyZG1EgrfmQ+aj3NBt9JuSE6XPILg1tgU4fcpRrwQyWmRIf
F4IfnC2GSv+uxX0xRK7R4wf9rY6PUs1avx49s2A+sFze5vzvXfEfa/FPb5iv1uolyxqoaF72iizv
KNE+64G7TkW4dMkzjYjhaOlD4/G40Hu14Ys7sLiwY1fZvDs10y9Anmou/OXPa2yZd45Uh4KFZPgc
SBm+lOsdngJ6Lo11xvr4z+f8gtHTIWRnv1fKT0lBB6BggHFkg0BlGGX9icckKhxMV7YbvgRAejB4
W39XJaOX5edbjKKhy2D7vQWMzjFgZhc6j+MsbzyLJ1gwpZvn/9PA4ZS7dNRImQkfFT/oiFEeP+Jr
VVc7KyZHIp9WCeUWP6+FVwdPwNs/7qrKu8CCliTeFzFEvZuOU+2pro05eodyY+euZDrRL32roYaJ
NpqErmxphwy0b7G1yeYreDAUDyyFngIXghMkePu2aEMf+HCNH3GdTPxmHW/URRRwrGEn8X7Uhk1J
Pm6pVN1BTiTsW/lEzJ8BFBR7MZ2mo5Cll2b+qWkhMK0EkkmUuJw4GgVV5AIc6V7u/0xNxvT2euDr
g0+fsr80dYVnz9zf++NvpBuVPrDoc/e8J//EpkYdLOIB3H5xqbYajgcVyOvXt+UcGDtdeHvV4m98
FBfT2X17FeEv6FL53UBVZkxZsIIwGtW+yq1KnngRoqd1i6m8jdwkb3Qw0IXOD1UJVyaJ1XE5LOpx
nDkspc5mUDwz5nc0JlxpoqwtCiBnNn9DSMDkFsudIAYDcAViP/OpGPksH7re/3OghSj29MfmGa6s
DB4JAATuRfCpTsmjrs/nnMvfrFiQBlxMJvMxCWs6Cxm8k8asRzPwgGBBDYyIC8wrRGmX9+UprJOP
OvVVWiM1s6mxdxOUwyrbq8IbsjVmJl0I295Z7JdYQ29yHDvnngCyjcw1oU9ivpZy26C2YrptdDmu
yyimDO6EsISFjHIcuShgmhCLO41Mo3t1qkdclRcFXTSBk3BmRNk3o733IyPtHhbA2CLbfy9FUfnq
w+lWsa/OG6EBEFWz/X8ga1Y+s+gBzHaxwfZZ2DuiXcmctgBD6kNneBF+yXhuiwFxIoGwWOwfIyuB
ztUv+vgwYwbiYFb8oQwy2NvXApbh/OP2wiw/rJ0KR9TybjOW051LhRj1nTBqQT5tBCp91fyeVApn
Li4t2wVWnuoKKpVnoF3apMgrD0c2lGSk/a+QJ4PfiVYxQfXuW9Qeb9PvFr6Onau+CCPTg71yBwNs
FrRCTNxmeyw9/HMc6nvQcTq/E/V/9/lN3MVPlbPu+ofIJqr5LBbY/NNsYYNQZ+3KG89QoGRbVdhS
zfepn5GjoYTagsTYL+12LRRQa+fuICZlDuke9tHtIYNFJ4pgnYmylCxVYjA55a+1uXzYXXKTSFxn
K8Fm4Evp6BUxmssnKcmzvtaWAP8lO22neqkzYmFV7jW7BVcQ5U+tf5zZFuVvFYNeS8bVj0Ll91jv
Bdg9C4gYS28Et3we4O49HlXzJ98h71DTKQbEq5b6fAXRSqzySndLfZoiUHABNmbNtMUxoVmwzJXR
RgiwSVfU/l8a8Nihg088vyu5ui57qGK5fRuxY3F2T79iAAvsf1brRiRri/CtIqqyPyyNlPHThnNx
M36dL8jP1jHLjaFsSbzZxOtr7fJCX63PMI/qDHIwuypdwqJfaaYouYyUKyqfJof4z0TP3k5d3kZ2
3gAOnGldHiYCEEwS818prxAWI9FM/R+ZVRZiepW/GQeJXZ6m+0fkBIBAzx+KBef7ATxtPhyw0DbG
qFRipkLNG7PtFoLJXQek2QYfPLlGSkCYqsYO+Rs/k6Q7c7rsI3XusYF7Z9FkdpWP8XGrOh9fXD5F
H9rf3wiX0gHu5lOyZbLAZ1G+CLg9xExpuhmNAzcgZsTecuv05wfyFBJpqXcDUFPudultMwExSVKE
KiZHe0SCPFQzoGgQPhgkYXVtPsn5RMQSipGPFScrjH+cK8TR0Bh8iT0f0pg3DBdKkeSufk7xnKo/
dvZoPHrfHXqfxMYXgK0SqAwbCNUX0erYe1IBWz1uJu6M+V8tDBdmb0OmyXAtF1FlckQgTt+jP/Li
9Pb5wKSZPX2HJlLpCypB/rD4Kf4dDS5q78aYgLpdVAiC90RoTfZek/7CTeJfeL0MBzWEJzv9CKvh
oGfR0iBQuQITwob17DKyGQb7cFwNp5DFRototNELmOCCJI7NW20G7QHpja7T1vKEyoAJ7tGWXx9Q
Cjujzo/VrSvvTQpI3q332oVHll36Bq6qKexiyrBzumZPT0mKJFwGoG+4c+dwKaJbO/BPSz2Ch/4B
tOIk8q1+pTLPbadydJgL1OC54T3EvC4LNU1zJUndeIdSWHOn3NNCD7zasF6TV34U4DvLmBO7uWly
NgraqC29YyNHBODb5bSTEiM9o7CGhzWIyuupSNi16taHwF6I41M4RL+zwI18zmSz4R5XPJQITX2H
cn6rEhwikSJbEXHMEAwCTzd0nbTkYYuRJiifiOYGA7mMy6uKU1MIX1O4Fgg3hBTSzi06L1T2GMbq
7W5OrCZAQVuXPk8NwXNAcO+1h4WBIbLewNwPfoPQgCxKttTvXIYVXWqzdgXaGiY+5neFU5G8wZ0H
ODwlnHbbfwVC8nk31gCCqSMKgsnS3/nfnU2UNix1lHcvPLRew/ERwXz4SIDY8vv+ZdWXCCyMQtrB
xk0nY5wtW396KcNz+5zmDIL0j/voP48+Fut+YrKxVdGLVvsbAfadnPeKrah2hn8CpzS5c/V5YBbq
FcNHlcYYt5JEiZFJ7dj6WYzpiZX589NMZTwvANM/KL6cvw45QkTXdcGWBDzQSMSXeoKHIT7itKYD
C5i0f9bCq+FCwD+YCkm9osCGx9FousFvS2s32kB+nxBSXCXc9QXIKG0JtwkwHmwEYQDeFLpe6vIv
EQRpvJvdmwOFcPs9lM64gjpOPyiKUEOHgt1NogC4////u5ZaX+5hWgKASZXhGK3Yin+1eU2zS33j
fxFMKfjIWA5GOI9uWT/byLRkCy8/ZiwGdXLKh++9rbqe6y/NuvgM7Ut3YCxwSjA8D5BQ1fRbLv6+
9mzBJYqHfvO+yqC9G7+DsVW89HGQcgdZLWvUx+mfCKsU12vH3LCIWDIGhO7EOHU3h3LKlRRMv0uC
dlZj2EUK4onwMLvmJsmwC84tnuyNgP4E7VOR4Zal55IXSDH7jjEQbxwgs+AQVf6ND30jr77wRU48
wjJwALeRpCX6W/o873M1FNN1I1ovnEJanhch6D2kskxN8Kh/VZZt7fx04oFxUHLzrLFe1uqzOfl7
EoXpnHAMQnRvI+6ErJeLoyucajG8b1QOkcYKfbR0/vRUOKJCAAvqASCCh49yiRPCUEu62HuPJRjg
p5ey/g4143k+Bj5KTp5ho7tMhE3dFNWmiSEkIocGGe70zILPM2a3287XszTjEIrZwbjkq2tiuTaw
bTYLjOMHWMqPkYH9/PjlxC96tDO+4Rh67NbjjRkRsKBasBEH4ju8DB7tTd3kPwE3LysMILlEuGmb
RziyqueOWZD+hJ7f4VvD3h3Y3m/amkDgyf9Eegma0QJLFLlKrX3Ltg8KF6c2oCL2xx3bmAehtZRz
Hs09Tpdj8oGvB1IWZHk5Ic+VcINnCyZ4+nvKoBg6wcIn/I2K2+izVv5Ng8iCMSgAfIUU2jud8CsT
o/12wIJHa1zHbCrizQxlXkHPsEw5mVHCwlzhrfheYHMmodNeUS79ieoAavd9rgl5K2UvgrJ/pajp
PtfsNG2WmyjB9BAE7e6P9qpYU+wnfPfOxFEKunuA+Ic8bkR+6FgtJ8Xk8qlzGJnc6qMkis7LdwmB
8RD0B/VywTFoYj44FJOgEa8SFGOEguzSTOCQzEfNXT/GJFDBaw+vJlsnQ4xPjcJVnuMheNjhwmMh
kEs98I3f6EXdKHmC4qEIbPE8iIHidYCbASfblQblrZfA8KkQoaeOUa6fsLisfkDNWyTL2pjTYMtK
sOk+YdVyVc9FVbvREhLHM68uSTQTisS6p5YiOUB62+bZa8t/H8jlut3lGVZfRWll6l6yPu2EzG6v
0ECbi9B7NgsHv8kcEfUi+xyRDC80NYlBCvQ3IkN2YxgZbTZ5OcEBdzgQ3/hxRtCq1Os4SdJWEYQb
f9tAOJYLav7EKnMzo9Kuk7GZwUrtyjYhfALS55GPV6tc84lE/iBUVFX5bdQg8/H9/EGg+zlfQSGC
qHbkAUQJN4sH7jP3FsRDKq0a0uH+BSK0QM/5JE0EwHCh5GwcxWmGnnG1g05wEUVmHruBKA52CN3U
jWYzX7LssTzqeHCgr62tifWGD3Wt5/XEjlSAdEjTjXzhXb5S2gVlWNbTO9ALUA2BpYOWi9wJA693
FGvTnZqYpsWhar5cl9dOF80oPx54KiWLlGJVJCDMsLfBVhEQAUe6CqaWfSO3apq71xV/fkG2LZZr
TqtMvS7ftVYKqDbMBVwnPNW5JDdTiZ9jOfg73kJ/UlTmdaWHg+JA4bBirFzPjnvfVs/83zZh5Rky
f6EQ1dvlD5SblvCXQ3KTRVG5T7vS2GFBF180pWxJN2YjTmBJId4MsjpdNFUwCoFOVHicdZQ53gix
8KwO3mCXarUnds4vtDVAJ21Dnx3KjlwoE8mVVGjOU8X9dOri1ynytMwvlGpEf9G8KSpZANCtP1z7
gIgUw5gKNzviV4amYTdl+i5bKbg4Su93+eZ6zSqcrZZVscNBlGaUv49mT9M4LlzxoEG0HoT3dEfC
sXC3FLsxvKWGdv9eMByxVc0ScPOWb3mKDWRCA3v9tlHwON/0c7+Emq7ycNPSylFrQMsv+6E9Tuer
m2m+lClB4Ar63L7yP1rraQW9HF4qb+ScnJs/tdgO8vmIxEWb3NX2t2U60H8dSqaJxdCRbrLQT5+C
ZwzOr7qVccqlDyyUWi3dGF1Vm+VqEBqMN1ILjekL+ueafcBews9DOQzm1BKxSbaxBaaFDyhFxgx6
5vk3Wtcq/Z9eERO1/sJg/pJkkV2TxOPfsWqE0XRxuOqyPjRUfvS44VqYzsXjCtYQ/JYk0TidMHOv
I6DsgWnJ5JBrNeW+ldeKizgUukLRUyLt2ClvaB3CB1O9t/ZrV34hrNpV1aTfl7lBT2/c0ggNwQde
vm8ozMTzFBqyyxRMbnbPvyv1r0C5vcS7D3DICeYq8s95a28ScG3X3JjAKcatT34NKAiuL0aYrDq6
je9XcTmQoqncqcSXfM0KYoNL+CvrVI8UJGcBJzk/puGkipnIrlslbEHnZxdN11Wl//HJLZF3tsDV
Rdy9l21u+v88pNFqbXZqmOXo7+0YjCghHhSpRJyfl+VxhuJPvGT+WRfyC6l15Msd/4Kfvv6YY3c9
k0IRNN/5L8odHhoRh10GiD6NPTUwHxZy8MdEbMPEN6snVsOS8NnVnj26PIiXCBp2v6PTTtlmKzgK
n/bALvvs7i96I92gQdT7CiCyUXWJwRhWbB3dMXEEF9QzQsyBD6f8jBr65PLcWMCqHubaKwE1Zsrt
NUECp/G90bJCjO2d43ysvbsB4z3gzZxMEHA3/THwzMPnPGwoRNaFhPDPg7ba81VzAXqpk/YS4FER
xi69/Kr3ipfehogAw8Q8b6XLSipIO0wNVmTiXXa7zItBqYs5Y1t/nJp1MVuajUf8ymqmglomcVmp
mTsHWFVsXPun3NCl/YhAaUPgqqyTs19JBDTkWoPN0EVb6eUQNDSveJkypoHiSyOJz3KAF2zTeWAp
2bQMV1HxVwFZWNTxeLFpBjfE7jYeg43hu/hFQWXsrtxFCYMfjrfp6LUxbny1bu/nlqvnrdyFi+eq
hHZGN817xOPVR4IrXJOumxgR8I/NV9wOpuYgmCXdvPX0KhynC7T2aDq9OG4Kb3k7lgZgrnc8M/Gm
+NANR/ZhIrq120Fx/6vAaW+QPEkh6M1xNjQMxY7ksn3gvhsIHEu9r/doAuANj7TAkuzmbTqsjat6
H9JSEkfZ8HWuKsY8lP/Tfc5cIX6n99RxVv3zLYxk5+PJNZNdohBfPSuuzTe7A5htm8ppI83jPLhM
PMVHkvLxNZM0XrEMAGOT1Or8mBLDiYuLT5DBUJO1aIAOaSypOGBv0Zy8h7wjfcIx5q96EzyjzSEc
cwCD/gbxOiTpo3IS0WNc1xzpMaqkQsf0HdTR9+SB94/AWjOz//FDpoFeovHQKDzPZ5nPJ8ZPK3nh
z6ioJ7iSRs+y09oyR+UywQfgKnBaiGowPVFoJ/pDUk8gzYL40pjzvfIAWsckN1Zllmfx5YbxfhuX
Al5fZJyjsi/pKo90Nltj5KMNqKIaduONsL7eIwNA1Z9xwT+pdQ4nT8ZpVj44AiUi75G8UoetNy8+
catqLcWMycAF6n2DfrH7GRxTfsy4n+wZZ/QMM6n2O5LStjFeB2dXTMmhbrVyTRr/lDKQY24MOFay
54OH2LrYBHewRWfb5VTxL/r0rFSx0kfTbIAK9hdpKQzLBbiELa8BNz0KMP9huyQw9o0jLFcmOuFA
FLskrVJaY7k6ZEQ4nqIkBAqcpfUnIOikK1kWnmxfla660aJHmghmqyuXMYt0eEFjyY9/12FNdsTk
JoEZQJjOA2hlT1KNM+ED2UX88JzFgimsFPoWNDABK8u+PqKaHRqAT3BQ/BUxsy0Z8kdef075UYXc
2RJ0/ka5GBX5wp93apn1NXyARIpiH+nWacqFIgABBPVQSPnCQJI2j/mQXMIr0JZCXI5kC+7CUKZQ
Lf83wk6i38OTDI1Gzdn/hBXLKczAuj2gIK/3EinKaxooDrNh66LycyB371veWvKcAmEaMJAb+r5i
+8q/mXdl/wYEMqGQWG6yO5deas2iagRnbNS+YGRvsHPXJIIBS931+fBBCTeCOneu2pyrDUzwB4dn
UTeS9c84tRzzIlX5DCb2kbYeAOGihvjPFe9Ip+NphUrYQa9XSRjALd2+pXguNAmYWc7MNIefAX5o
CMuDnRmMYuhkQYTOebSsT/JF3sttsSY72Dh5zagL6nHrDp4qOQypUHaSVWdVWkbxQkR9cfgibXBp
hwDoOc2R1NeU5fu4vd1vxpmq+tai2DzMdTSCOSlPIjrOw8NNFHS7Sxq9QTgwRRFIk4appdWnEsfo
ee0OyCggKoGCfiWjhw84yPE87fJbmJRElzWFvke8kKinvfWuF96HHpAuiW1hRRC1jdzOnDw0/STw
eViUmR35gaM/NHiTOqlVjgm5YT4LM1vOITjH/ZiP0X0zcULxnRwD9CNdbR0VmOh/u1zQhilMWTX8
/AzaviFQ3IsZeKYmTUJNw6FEGbZCKbng9mPYxfy1LoXWOzD07SXzekF3aXsQC4T86vDB4PMwQvt4
pPpDpn3wFUdIj/OHqc90IiVVkc5e/5FwRYZi1UdJJZvEf5vwK8s6atVjD2BU43cr5UlSbsg7aeDV
/t0rLs6DeoscXFlQ4ICZxkuKwgPpEKz3qMb/qeMlZ3uZhlfHLoudvshNXxA6rcFZtagiHYiy8LM+
eoHgPw7N3cvBOsiIfrPbbBZqI3z14L1VULtYLjSk9HgY/dgrpF/0xbzJ389BW64/d9uGbllvTYvV
6XBtOwB7TH3Hw/teyrE48oWPk9X5SyZUYqZMI5ZWkol0MEId3cuq2tr0rF9WwXanKw0PkBuH9fiN
Nk5BrfOHp+BSiP7JJyF8cZSvX1WCOXAiJ48y4Yvv0fPIjncA5ViWReFoiV7dOmDDxdcqi1KhL0Ve
fL63Lt3WFxUVL6uC1mxq66qx/AgoLB7txvQlnKaqc4cjQskNOqJSg8LHjrQBupweL6/3cftQGlwW
GXnxAjAmk2M4NtUkyaxzbQfv9/M3eisUdP0GfRGg0ADn/TVFGhCakMOlp+4v9/2z/dhNmbQQ4C8c
ZTcsjcLFDEmgaGzWNSEl5BIRRpP1IjBTs4vTsOptOpEoH/icev9YKT/L5PoJKKxrAhutPWetciGg
f5ExcyZyCW85oHAvAmv/xLkGmi8lSuYQHi55GNgWXW+QxV9Z1TJ5vJD+QxWVEsRq40ueUV9rx1Qq
cnihpz517x8I+EBbMeP527+uXOidRYlSMe5KGbkZDXDjATozR3e0EPZ8uhlpkZcib2UT6rB2xem9
DWkVaLAYMEK2sajoyWa5HzqpUbYExJmlNUG/UdGmfJw14rplXgVIXQD3HsNQQAOOFy0ElPyluSk6
0ZiGgIqC7g7lNO4znpO7xX7uIPUIiHM+xHoy61fmpEF7itgWaI6g9w3tbuJ85+NoXL6f/ihRN6bE
X/r6COldu3P3nwLUNkT18V7Q1v3Gj3FmioZc2G30HK49XYgAM8mmGmYLbBTU0ykJxjrOFp9Ae4IT
qcpLbm/NUtYj4VKadIvhrDbtQgwHHAQUf9zpNJ+de90dAu1fyH1QHg+W6WxarHsR9tYTVxXoPogJ
Gyd135K+qBYrja4vHhSrWPvJTxZJ2B0b7+3rvSdfijYrWqy6Xu8rUHIzC7C+GycIz3OKHX1LM721
Vv8UtK8W2osf7wj5zVrYW8g4jBVW+gcI/WSLkJrDpvNqUD74FU4SemCvcQdaw+c80xNH+ChEyxSI
PZczmXvYWRWoI2iMR8CjlCjuxMIyPoN4SUZTDNP1F5qgwdOS+Me11IXl5fL/uk9bNTdBQH3fa/nS
uNOm6r7oubkLx+bkeNkgsYs7gTKbbyYl1eJ//6+1xAbxaU61MHrKnW0hV4JjNNnKVwoAL7hf0q6z
rH3XIaMuGWyf8XEUmpeqDq6GA+VHcueUFcnfRNrCSE4XBq7x2sxHWEcrGg8iwTKRViABq1GU3oGb
XGk/Jb0J2NjSsQBmF2hnco39C9Gs2OZDWboBYKEpZl+b/gkdNjL2gkYrN4f0wnLhS/P0q8Y87MGe
3AqP3cfEsx1gx+2ZHuqiByPk7D1HR4dJxp368w2bzJCLhAd0ERG36kkN7Gv37jdIlCtuGB3q4DIw
8iw4CVaghqdh6VlIFde04n4O+5FYkOXCTDV31rOOrmkvCQW9E9TcdDmA2i7Ijj/GIQ4TOzW+9thd
gOMkNedGzg7JmPpnw2jSnoMAKOjfraHBr8n38SR1+3zAxXLAGdayXyaQgpnR4XmFfMoKN14KysZK
4wegKW89SUvoMeMHy3EuMrh4niGvE27GEQPAWR7mnJO34bmbDnjTjlRXqgXTKbYTJ3CXRkMMX2Bj
3ow/LF9krGDn1uNMUmh2FFe6mHLEzU+pxRfN/omVmfi9ZUWfJaGXpryyS8U7Xn1G3G99K+ROouY3
Ol8pLOWDKArO7OTrO6pfkOrtoF3QCxv9tYcpEE74thEGYjwXy2NsIIco0204YqAL1bzf+WwfXyZ8
U1heTUWYIcRgwGRhjotc56L/J+BZVcTRwm/0g1XzWFRB/eHD0YfnTEZpo4ANvpxtFEGO4GQ+FWx2
arhOfoO/UyqMNU1V/FRTW4xzEUydj1NloGvze47ciEPqiH3IErSblkFy98/v3+GiIPcBCeBeIIGD
Qa5ik0rnpXkhDA4movhoMQxALKw5buf/cYqo4NJQDg9GjN/GifxQF4sLC4+Ob3EZYV9qXHoS1AMr
rdaQVPya7A+065hS77J9XyDJ7bsideNaIe6oj+FUL13n/yExBsTCHNTICN37G0nv4sLR11FFg490
BShO4EUGsYaDQAwZ+IxtYsULFGnxTOZyFr29uluqxJ0YUZD2ZKrJJ/wPqqL/5bOr5TMdav4OCAYa
SRVuibYnLvj+mDk1XYJreQZGu4RqvZimlhpvqOkK/oySrB71wQ76473fGZ3CTrWUE8tOpM72HKFK
nx8so8odROC+Ivw/oCoMRwVZbmSFG61M231t7mkpU9vumAY4+hcA6sAfx1fsBvv+mtVgmKFopWm9
lWD2plr/IXVNtMrLRc8spnuDSFIcjKwyxlEDaiIlwPdrwZUp6oFSs0rBjADwGVqMHRU4Fw8Gj4P0
EJz9BpZqwk+MkGUJDsE7GK5uORPU/GGEeLWXYXknS+3vLYUpOmoEIXPJAuQIQYo3ukIy+cJPWaGx
f1EMTaYCrdvByeP+P9g0nGXLnTuVqNl7X5pA9ApcJY2tnAuqtlxdCfHEGH9R6BGhcSlTrqSWlR18
rzK+Zga4kWnzSY1jkVyxONHx+s0yEjHCAu4ggO73jYBr9MEeHzl4pMtV9NX1N29w2glow6EOOleA
JKvRxL3m4M/O0WocZJ5ZY3S2Gjl2tJS7Hx63ZJm7nMQbX68ru/Az9tuKP5WAUYaRWKzOJ/gyFXX1
7kBoXwN2882gP4DsW/aDXl6a4Yx9E1u6KyDPkC65EvmGyLMuyssrAVQFz0urUFlVXwqnejw3yrKk
L/hQ26yNieBMiucB7QSQyAYOUAy6dTv26utxKBevSeiwJkGxvUf8V1JTu6Mx6AmVmYJqTXui9ncH
mqm1fmPdfl55fNiCP+XN/txycyqT4OawKCnhSLUqymc0V3GJ+0vSgulo52KMYQBvtZBFDTBNS/g5
GE4ui2xa9mV+i5s/YUp7S/LjV4iEqnO+iIpv6pknL/s7rhp1Ux1hga3X8EOppVfjoLBvv+WPDnQZ
oCsoqpm4uoH7b+9nw5vEU24LPU1UT6ApX2QzgJ6mO2hy5nVPHTkoCxXGF2j5zxY/onpCBBBfLndL
Aa1UqxgBQfYQifbCBLFI/pFvac1wS3zEd5i+pNxXTHqlNdl66muY/yAjH00Rf2KNVrEMJP/SUqZ8
HpnhpwsqGdWNr8v9i8uUkMQwkq9TC3e8fbC+VLWQIuD6U6yy36EED4Do4PAbPdDv0+xnjMk51ZzW
btgOY5Y5+kqRQKxrwWgwO7gGY+DCOn+XKMdjG+OuXPnaoi/g/yzY4h558WC0BvLApqf+PGSesKNX
brKMz8vxmUMKXpH4zA3wprD6kZbn8ozln3klIDwnlQS0DcCtwG6QItJaDee3WAC7jZ3TJgs8Uanh
FO2VHy5reGj6xg4KjvQ604PTaj4uD5qlJHu6cj7iZM9xDG86eooP6Kam8Qp6FSn9NFaPUMGoLsz6
fLCMsY2dax1w0HMfhX5ueovqZuN24K8PEFeExUIk34FqQqR8H8yIu6F6bOW4DRvXPbl81cp9rTmA
6uFkyfsbtjXI5o9ePMlulIx5xx8dhtFk5/vDTWh27aBNEaQ1WRe8TdoiDroSSxIcSF1fcJltQ1NL
23kXtkJ+ZOm+aQf96yrT8nP+NOgRVvAIWZvIAtpBq/FhvFp3b78ZtJw8rp7zOoNrLem1zk8BzGtb
/VcD8b1co4+1Dtr6QBlXOzoEWhOVWJEQJUftaEx9AfoCF7591tWDgY3zarzHep3QjVwKXrEbDofS
2Tprj9XQU1rvvkJRHxXvqK5sZMlcFFBi/7LjLphBCXOuKf1oG5EtNUWjNPPgTT7kzKhCeb1ZQ8OH
txdnnIxvxpM8DtD4z9cbhtITIMqH/lKUg/GIjnmLq+fiTzKJm3QXzt9XAZR30LVxKjXVCMRBqcYA
dbLpjNdW9Yze8r/G+E7AYITZTQFSQ8C28SXT9aMgrees40QA89wTq6I57iRFV9B7eMO+Q/tnRj3T
eTp4/UdECXkZn9M2ncp3vH5UbEMNMPz+8q88QsLaGq4SnERwSzusAaE02c03F2bhaVhy7OLFinda
z5de45CNJZJnz0iTliH0rOyoFR/8Qovum5wqLfTaQUo/r/21O8KlTDPzXL7S3e5bWiRrZx2FYmFJ
JtDBbXRHbUeMK00MIZRFZJ4jnJ+EKk4pt7U+PbaOVB7huJI8jYHlWG6Uf2gqVsGdugavZR4p68Lq
aFB6yWQJAkwrtJGE6+AWszdOnnF/TmCMiCvlxunZVdGDdlnr0LnuPFj5TcvkSc58d4iLH2R9xHpJ
M+pjNiXAw6TC2AjYjCkg2/2wz86mtE6K0O42yop7iekFIC0RwQ0X4K1slwiZpGMhbscp2aLwsYjb
lA3dZPC8B8RFU/liLrGWd6oo2paNWsSJ3WVYVUkzYvtEFOXeFvL7MgHyPzTMLVC3+esOFJ5hmxXz
vbjORKD8T1az9m8ScuARbD7tUIvMCMGzb6ZjrVKhYID6VixasKsJMYjy0ruTB7yr2ozH5yV84Ggi
tKgtEc9xFjDiyrJWv+1YqqdJ2NWAZCu4BKyaS5fGIiop1dfdUrdndYVxtucPSXJj72StL2OKcxXj
u9SxIp2ZR4tSMQi5kWnbYnRuGw9KYI3kTkfn0Pcen9hBRt0RPwFd5Sg03T+FLwzono2yxSGPxsG3
jUKHjOx7B/FFJ2WvHoPMHSH1y2Z24Otf+vK8ZoPWA9Bec7o1RjB8fGx8M+LXyLQNB+z8QKkXiWoX
L7Afp9Bd7wxpuLHlb6FwYFhjsLLzJplX+PXjSFuQviG5dxWjZVbsAwCFUh2tUD1fZHjvWG4DP2Xo
YEWT55uE2nUQzFI7RUQvrobHa0tRZ32fBrubo62mtVwmUzQWCWc+P0vv3Pji/SKE7c6H8isnpE0Z
fWRiDcf0R1wr1nkU0zdkcWHc+lXkYCIJvFjMdEw4UY8w1MUyX4Mj2fI19SWpy5k64q40vmDQ4rSs
6SdFP1uIWWJsd7axB6lSKwZUsqX08hueOlvrm8TeqNDAATiAvWlqnoxCF5Nak3eyQRdK6I+s9hQa
0FR3Dad8naLBshzQYy22JPUixQQ5Ec33nMJ6x3fl8bcdjQWJbRz0RkTICj9W1AlwrOX6/4qkmM0g
/d5YxCwPx4x5YSvKS30U1HZPanOuJrARIwRE28fkbeoQLtCwmwfdLdCSi6+AF7Dm8Sz6F4dyZrKu
tR5HEknZNMBGW/c1r5kfd436i18219O4bG75YXypJ0dNnBHHLcUvUyA+ITRWo2z3x4FLjuYQ2iSM
5PQyegFwD0B/BbEcOTGY5YunubTbsjJYjK4QlirvAdICyNHi1dpqIPwqCwRSo2oWYef+YqNyF3aS
JPvE3ov01oGJUbcpj4JfQOV+Lwj3jZ8P419GFsoEJqZ01Pq5T6PZPn8iYP9RXgCCxhDc4cuuHib0
N+gxfIV506eyjM4CpudSvRZmng2KEUS1J/ogFh3kTrLYHEAGJ2UK+oRKr/0UBJuH5ZhRM55oJ1xy
26A0YBfqbjmLpnX8yxCTvap5L9Gid03hXg0fAaJohD8Bm2IoTC6I8bf8i/kJkZanmyY9VUI9hb+t
nnLs4BOWu0SHT+Aa22D05/XHPax+kJymbfglvsAYxjpNBOE3Sr2xT6dIyzc4dkv9iX8SuQRYL77Z
a48HeahfCv3dmWu3bu7P1OFuooV/oUkKvdfpgK8WoM4jTKzC0HDWrceBw6JaYlQ0eP693B1o5mup
yrGGNQcd2lrke0fogAgyRp2f4Ho4GZwhA6KSU/YRaTZndp7+LnqoZlOufixn/rV/kxxBZBW74RSk
OwyJHLyhRmkvvFOBeAo9hOtJqcwkdG4tmQt+eC1wqVsieebLZQyTUtBth7uAArk/Gq9EUKU0laI9
42y9hWsgnZH2mNlmEduUUqDEfbO/qr8kV+AOpEEm/VgIYR7CfoMy/sQ5KETRcxEoQdbdABWeAEmM
pSqrYAUyYhfWrAp9aAgxqWMJqmpk9O7K4a3fDGKvQV2lPrkWg7Vm63hFF7r9gZrXziyh0Qo4PPrz
oZyfGzZCHVDhXXPjNRv0wkb9xL8O4KwbHkAqbpgjH1OBamztYN5nepixVR7tPN1eRutSQoi6Yg22
iGIT9JPPvRYKpNmN9QpkG0/gDfGfG3dfOuU+D5mktEh57SF8D10uTAQuIRwtfa2LU9n8nN64NmtH
aED0Z63mIjfwlxcsKvWnAdMqkfAFTHWwurz97jDOydWfbFlHQ5i580MdeAAWVC0aARcnGxX2W/Sc
WxQ/FFpDidJL1XHsWjF8rp2VHI5T/nQClvVOwWrnJrZjdlcd1y+BLoXliKZFbBYkB/NR/SAa9E+F
Viavn4OkK2z00rycFlcoHq7qybM7cRwsgvXDPyLFhLBPXDge601egonjJSz6POHhoSc95/6+bNq4
1p/Lyr8VFzee90Clb7IhwS0JVwlYU2Wd7HZ3XEMWaqtHp5lGJj42LZ3bLbprSLSVlY17iUDRcESR
EqPHHmHSbf3wPQCI9j0I9xTp5hA7heWuTmwmg7jEa7SgJhNSKFw+FvAJaMnkfuDVd+bzyIZrxJHe
j6pCD+WPPhi5biyRTWIgLMX1ETb5aQVdWAvhA1J7R5/MvQlWtzApbD32KplJNJ0thbf9lcg3Sgu1
7aRlHbSNsxRSiNO2KeoPC9LaYS+po/c3k+r8QSGHlqr0oer7gjmKYQy7oWNJoMN1B0x85c2SQP/b
M0jvrhZFjEoQ6C+oFHP1BZloifJHnOmhyPuIx4WYVholG/MLZdQrRxwqzuUT3GlfJTHVXGUs8DG+
VDSrs4aHrcN8TdTTvtPHGPi2/g2ccl80+NIN/4SLHjXJT//bFwN0qVuN/ZfBmB9ekslbfgEGINc6
USwm2qrscksEOKdq3ryNtMeY0rv1wYYFl6BIxFkTsZe2h0PQvSkaJLVpYFFOCsyABaEkvfblzf7L
S2f2NkoE0iXK7cz1b+EbG6V/9/sUzcwRTUJEI+mGPIRGWH7EMmhNjCcuAaAeJYlF2FPm9Tu65XlV
Jmf32F9GfV72EaIwLp+r2ZDgqQsq36rSAiJSfaPw7gvmlTHRBDs95Qpj/cUpFUJSzQvRHt5dMQpE
xZfV/5rry6nnVLd3KwRoet7QcKRMJw/B2adMIO86IkXnGUhxH1Ud2dji9xl83nVWJO3BpJMi1OPA
kCc/9ORI4jfSbM7R/H79z0B5evWuWi7c8cv6mupVAe57Jp0hclA9E3gWfi/Gzz5Y0FPhuk8DMrye
ARpWU8xwjdDH5SEWiChLrK3mQGoyQIxdc8aUy3Sx7EPKrSWw7yC44k6+qEi1CC7duxR5sdCfHgC+
N+GWr+PV6uwKGK3DGfKl3d8jTqcvW6amPQDEp+8SxG8vlPQhBBjDI1CmcElp6kfs/ER3R5jqZfPd
l9Oh0r1OsQuY9vWxpH7DE8oMQMMFlPxcKSZuwARManV9cBGBivkLUH/AbRepejbjkZBnRZUJIO9B
3DGg5YPSn86veRvG+I//aT4t8A9+aZrTeDV4e+m+Xp9cnCt8TRRrtLigp0TB8sM5BO3ONbQMfLY9
zQ4jm7QOmQgsOISKmnAeUzD80dbXfgIoNmFlFadAn0AKnf1FzVgnH+Jgff6vUuEhouR2EEE1xVjG
dsCm5BsPljxcrzeGG5MncRPsTxkQI0hzWau9DRUUypwunN4es6MwXRHnQhbVy84yE+AGDhpS1Py1
kmiwjHF9ee7YoHJZuVgkNZkEQT9iL4zBL1ygLPA0rQOy2lx3hRHeergzI8Sv8Kl5bG2uAWC4IVe+
SC44wu7+ipI6r9ERFxPRNTkREB3phaaZMbcFkwLf4xSClc4FVTTVqrOB0yc2TWoPlwIMiRpYeEm3
TQiMtErDfG7+S+AJ5rSR1L4go1SogWHwDGjoxY7uroCGRh44qYqHFnDneT7bXlKw6nvSlkRQDpHl
Tu5tNPtlWWLmUs/uEVijk0REpPESG6WHh/jz+UuLyOuvtajgTorOnXrWn0TUzlEcLsLOJX8quhAx
x7IpsecuIBTGBLwzbV5AThnspJCNtM7Q+GaUPBA1zspBXRzaETVl/RmbCVzNb/l36u58wTFAWho7
ZTxaTTLahtdeGFukDkiJFojwjyuCtF/aj8odoG3A+2l9VarVxvbIEqviMQp6ts1RjnWtXwG10Ww9
6LipBW8LuQO6+ab2MBonUyBhMTcmaYb9shjdhjat3m2w+jerIJLzShvorudZoykHys7HL9Mg08sh
nw1D79HI0vhXylscGkPn4IOO+jNMyBZgBna/uuUC1oVsInZMlA6KDE3iempOUqRqh9LdLmHiOJaK
Sp73CsDiPGVn4gtMRLc9XmoUu5gChOox9NQ2uw9NplbFZSgB2FY0JM7tgbdEjvlhScS3baYrsnbD
4eJ2aF95EetifI4Mh+Ab1y+axuMyb1n9HgCecJk49UI1+iibffLpRS6LQXs0uDXGNC13KBdqNuod
WhotH8sZLtgNeaUmAcfnEv+tP+sq5fvwO30HpMl8ykpHXCjHwckyWOK9U5n9rLSLmYDuAmUkquOO
2jrlUv5rKvTDfuzg4pZn8hQ7vpUB9L2B+XhCiM75vGdEG0jKo+XerAApOxrGnkUFhHUIYY9ZcOCG
98stXceNzfotyphhDH55Aq9+XEcYng4gaoOksDbXbVziiZn0ueRtUnrRTfNDRNPEpstFCNMuYs+E
6CR1VvK3+3vA6PKgWeCe74eRXxlczVdSvQYYfvpvxJno/A501vQfIrHyNtSLITmN7hTzDBa/Pm1l
LSTjCPbefo3eycZE6jpfqXD06LNZKYVCumxtJqylXKmPV4sm2T45ns3FiJ+O05sSO9699ZTSQWNl
p6Kq95kbgBI4VLBEN9CRrB7WWfLn331asPFtyabZAbzGaMWRx0169qEBg+ZfdtbrugPPIGSeqD2S
Diy9CtrF23BhZhqjU2p01mAUvGePLXwqTQZf36l2cex5FrMc7PZdT0Nu1ybsdAZuVy0niVCrfUO6
qIYXxz+CjbutLJPEv17tUKBWy3ThOOJM1w6Iuc+oDKZn9BH+iEYE8olcU2oopC9ypRb9IrOUUJgI
rtqXonBc3yRIN6wJr0J6FIDfPBq0OgVEWDdupMyG+PNfF4IdegAgxuxsaYTGYz4MQNp/zdGUH8zf
njoMOvmoMlcFdtvdxRndkfRc+88xGXsIWz2bwValdox6TXhAFQ1OqQ4tb9+ShE+XYPwhHz++sttR
NcAJQ81RUwPQFc7q8lgzx6jGqHo6s734fePTNXjH0qxG8eoAdSjeoIriuXmc3IANIzRwsFkB+weN
QWFAsbodkVvcs0SFvIie2F7O2OLtiBO8lVfWsfeClxphx5Ak5HYGlycOnOMrF5hiJbPiQqz68Ks0
F9RY6UjfkY2TMKQy8+a7X2vEMaiIi3TDjlSDnQ01xgpykU12bgyGvpc8LBJ3OB0ai35Es+ZfObIp
n0wm+SGy52etiQCI8I6yc9X5oYaO9n0eH7/Qw9QRQVGZRPK+0ZLNRrg202CXBpOg0kkK3Krb4cUg
/SNsGcU8C8GzOmryd1HiH/qlqbiEuqV9VgtzGGptC/W4JnP0q/Dz2hThfhJxtTT7BiNGoAHH55BP
dpIyilT+smM3qvswbGk/kvahc7msufo4mAtZwcPpz50YUDlRooADQNxTRonaBjdqD7rfisbR/xZ4
PieKnGXIh6JQJbBUBaSbMfYQYBT4ZVMn0c8SiqsicnJ520xt6/X57R0+xbF3fvSEXJKhGw6xfjMv
KATJpCVf4PS7Lw7GBN/HJ/I2X3DLaRqJTtNtNqEiL+N4/0dWWvde5jns9U2kqkN9xYGOhOwy7/m1
Ug1A7b2B1qGSS/sK0+mBkbn0P5fMosWipFN6KORhg3rYbqM8Yz2sINAdGGIqNfxFQoSL9fLTFJGV
8RcG80FL06+6PFhz/Y0Savo75c5ocoMyYke6/WoSGkCiF0AJaLcrafISCi6f7abYxr0YTr8iRP0R
KK/fmyw0smhSJPsM5dBKaNSjZmITMk6PdnJAqnrT3+A1CugmOPY5ukmRlG4QyA6ZAbxgiHwDsMkV
ft7TvVTYCyH6NysTYWzXoHYwpBdFeT/YrKT4UQIbPkyA6OZo0cbaYiqEC/8QfjTet/T4iPY477d2
o6SW0z15P+UHi2dwvheuw1MYs0+tE6OUGQAM46Kchkpij0ovX+lMhNdfPys9Aul4BN/v2yAxBYfL
esANDrteIk7sbWXTWaaJ6CC76xjqM16zyPJhQdVTItfuQuzvophn7zsNe21q7Hq92tWkL/HAB8tN
b9IBPbrgP8uZ2U8G9wV122vb25hozCH1w48G/1A3EU4lJkeW53WZNSTkcfapAV1OcYHjJnNJr+Og
nXXF+dFtecBRYn3FS96GvGx71ABeUWz3Jf8ry6vUVkiUYSXjBXtM6PraIZUVrU7EEMqufEvbc2ZD
rEF6o81h2K7HerMMWePKDp6PFMIEglmi9zXhrrBDUcQsZtOwZg/8yUfS8OArlHQ1Qro1LBN4iV0B
vPLH68rm1Y/GMnwtGwmRrtxcvoDEsLwsNLhezaNNtHzHmJoYsbhPFwXyfYOvp3HEQBDYEZ1C5PvA
hdFslcB7m3to3puqRMIpezqQ/yNIGb894j1/4qUgYcBM9glwV4H/6J0hyj9xy8FMcQ7neHLsyJ73
Wtu3ORspxZ3cy4HdSr0r6O4XshADDlLWeTYfRlM0iL/Qn5+ZvZb27MfdgBfqP/DCGzpAMxFthE4D
PLO97JcKPwgqR4xGuc26bcd8TMWFSh6c1HHQHXKqMwPxOqtTLKjrm95sqZnlN+IXAg8HYSKgR7mO
Cud6v7EgC8POoQtbtSok1GtrNtaZvSLfw7AdP3FjTEyuHlWpsokLc8RahPgsQWuYq1eukbyWvRlk
HJ+CxdkS7S5AFXn2ZCT2E8xV3mvuS1Z96Mm18Q3CY7sc53rC5doy6iO/UPFfaQ0rwxJ4oEMYjToQ
lTw133Ty7mBoGBZfgudvNMWxSShouDRcflUBHGx2tSlg3cn3QCtkRK4+jmVMJQtq9d6ClI4g94Rz
GvPTGPcG/FrDncKW426ADdGoQBBbSaLLGzbPOELyj608tpVeR+ujeu4VZgK6Zy0vEgoGtiGiQkpg
hCWDWYDMNLknmS71gvfUOZIy7KCXoigmg9lE2k0J/+cfhV42wL6rwnsX8exUu3g4LQLbpQxkEG9t
bql/OcOE9Fv9HIHlSB71TKZ4OJDeK6CtAmXuVDmaekKdaGWr4RrRuZchssWBAMKASb+F1MRqt8LW
0uB0D86b86gf2zY/7RZusvlNEEwUqyN3Flf5yk2KoSj1a/7EPi/wphUncuKrf50ibBCldB9LwL6Z
l3WdMOGNqCXyArjDuWzsAxsGcCYWgSYYRc0MChiYRoOmsVejA4RJVqrdAKA/wU1Vh6ZZE5NPTV8U
U9mvz9ArGo+cRnJkRkWFEyQ+5k0IyEzZ3Cbi6Qdhe4d3bmrbR6RsPKASp4DwYBJrs9VKgcoYUEQA
sdtnZ4wI3LAZlb7N3v0lZpfjf9YLULI05N/BSXhTvwk+ZkPrgO0KNCVQc7YvFAY3RC/YtLJJ3zbv
CXzWV7TfeVExjY002Zo+z81el6XtEQup5yik1RbQ3d6p1JQC2qC457FW7Ie/iMkOz6RsRHgL3eVx
JOAmb0P2SG4z2WZWpV0j5/2ex/q3S0amVIOLAxuoyX7yauz2yStznjMOftGGMnuRe2hQ/qlQWJr5
UHa0gzxDXofTirREgRvHKlYf1bPzdnBbcq2Ud3f62xoWBtJxjdWUdPg/jQJNFJh5+kIwPIIUg1r8
1X3t/zPYzO40ioxX7cNvWpzg3OSsQxTblheFTjfGymLDTaLRN8nGvQP0ch6u5h73M9Y8ZK9eSS6s
0hZKNciuJR4Xrx+Mww59matu6yUSKWjtqvrMI09FQonzmAQ7BliIcp5LnlF7ao4BTyKi+7FERx/r
ulQDw4G3KbJjhOcWp+BeV4X5jD1iUCGwdb7AXKDxK/wtjV3U/PhOr1P/Jkgn8rN8lJRa0W0zBwtC
0rs18mKa7tcSFMJPx9xjKpw2MskcsmOUoIR00EF5P+drcrSJcupO3EJhMA6cs/nFix8gdQFDncxI
riUKxy8UlHbDkwhto6qQbp8OLjU2KPxonW8CLG8RtUW/RzB/jjx8wRCFMXV40ne4o8CrL/Z2skZK
HeIAsYoEIL/Rjryl9ygaDjDGdQTbNcK6WFfTdSEztrJzQVjbWFf1bDrRUOi+2ZxGGnIA5wA4hUrV
2BL9gzyLJrdTdgWoftQn0gW5AfSuB5TK7kULwXBBgpfdVm6Czkr2+KtKVfxd+6q9KQ//QRl0JC3V
Mj3lLe/rOmshEaA6ERXtekh9AroADRmkZfV7rZQ2l4f3Yh+LPhuOZvnnvEx7kVUHUwHbFS4hg9vP
UpbKpLxgCyAIMqsx11tqdBDnLnZXB18GQUmedTkjn0ToaDoBT8/wYe/WdLYpDZO57mDr5odq/gby
Frh9VDynxvbW37lUVRFxsS8C38yhnf724M0D5AMxO7lrTIhk6Ps+TPwFSuavytr9i2VZl1HqZAGm
IIwxW9KLPZ152yBTW8bG6OBtxtNttuJ/eWXKVWkY7pqPqQmgL0fPkVSIs/XguBMSutc6CoA9hgFk
uNwYljkSdm/A4EqRWAiI5DrBlbsuGEp2f6js1FxaYbOwdO6OoJ4NF6XnW8vZ8o8lg0fLk7tWqKWU
6itD5SvY+g6B7+kSDWboz6CxdsZgztj/lcAJpjEPVzbIjKJ7NzSz1FzJWRmfOpuz5I/eoAJi1B0i
qkw1BQF1u9dx/HN0p1hf/qqetLrrig0eNatnheE54ZL0rWfcpXDLQVbtvayqFFdvVwCDqSvfIkrg
CmKDygQgB4vSWRX/OS5IrZma18+xQsMl5lD4fwsmWQ4b0WFMptRVzeCJfC852Qz/49cG2QOfDMOq
ck/rH81nWyDEDryx01pfvA8PFF3hKvhQG48ceXvuYFeFIcWEf86YzpwDxRl70MhYA00mGuu6mnUm
+IR4cihx9KHAcmZ6RK8MckGrHmRuB+ezITUQ+gZGSvI0Iriae2dh5s1/YGc63E4iUAnqj+kCpScA
3iKFjDKfXXtpXTd7VZ02YzHWD5tUbn/fuW0HJIKtE+ntiI1oJn45fXhVQeJ8dpSK4gbvzWmGqYmv
tlGqByQM7OcZZsZNpAJY/2uyx7ZHkLm0UrRs6WZdHezGynIFQ7Dje3IOvBRT7Ili0gHYjEWBOeSz
GPredFDBlHJ5D7o53o1vH76qE6a/eI5Oo1uBZfl/HK5auQM9db2as2kJGwnCdQQbZqpySk1rX15z
vbrHUahi00EtCzibnt3Bluw4RjChj2cBJlRS0EdrnYRNfXZFet0G5QAZtMOu25SnB3BtG1j6U7Kb
RQPhTDfZ+haV9IM8a2JO6tM1xfHGY099Gkl20Yu1DzKqLQgx4+7oU8r7jzW4VHONO0QhH/bH6q7t
FK6JC/SOHo13EpuMYLLzpwTNO1l+e8UrVyC7AxxbFwVEPFblbyd6L7n3FoR/ZDhAQ81EQaBSHRs6
M/FrRrggTWAyC2AkK96PJzggp4HvFlZggCAcG/Zye5ywcxMQlAe1qbnjrdKFZJaRwJD7PTfZzR8f
l+UMwkJQsskLvX2/HJwQ5DUGBi0k+ISYsHlJvtIR5SvlfvGF4Ifl/B+St7fc4Pz8azZcs8kFImZ+
ykLCtsqb0391B9rl6Y+y4sy9x8rgKzBgpGQ3aFhRojsEOFNfjUYCK42NHbW82Ke1WxyD0zIMUYCb
1jDHgk9pw+x2TiJ4aLjJEyY2HTYwuFvCQr098TR16wjz5RL48lk3/+7g2iQ7rGwObYLjlAY8Bqlq
Yq+ReArjb8d1byzHlWWHgJewabeWUdNU+cPMCRCkK2QTWvhU/ehlqHnFbdAr5IvwnHtzVs51j8yJ
EXCaZ7j2S2TUMdp0qKIBi0TgIr0/8xnYafAFd1xX+Qk0pnO87xXk7igBKRDMyIkXrTwYrp/ekpX6
4QoKWbO8+5saiuK7VEX7+PRMs9qYH7AJzw8OMdgWhTq3nBKSwAZtNo9sBfM5UjhoIeQ0dohYkJow
mDYu6WbSFcj2uKQ4xtZ+oQYECjjbUp+xah8TWvbFE2ajMqIAiXGYllGRGerG0T/OWIyre95Zn4eC
ji10j3pouJdGuoMm/3OyriL/+MkA9nEeEm9iUAZL8yqCCES2Y26bOUBMf2/gYwsG+vRnM1RJ1p/e
3ivGfShlJm7yd7gOxMCq5H1c6XXgOeTDTl01AjX/Oe55qGTZJuLaGcgj75JWBT53nlXQvd57o8Va
qVZ5gt0Za7U0d7g1LfqY8bDbArf0sjKs21UF8FYpQ7Aw8lPPreoxyJiS6hEj+vbNKXklyLVkXs01
5v96DsL/MXuGAyjsossqHexgXr1YpqbUfjXiricjmklsAx74YnMAGZMOaxXo1xEDHRqSv70CGyg7
4HTGqXyGtKqu67LroX5YNiASNtAkme5NTM8X3U8yzeSRKk2lCPphHfGnxmMrgfC2I9sNX8KLAlp+
g9b7VKf1qYEbVYyJWz8bZlaruzg+iks7WG4nXCq05m48fJQUrc0+Z4FhEVWREq6RVdQrRty40yyC
VKIsc4B8bMVpI6mBHyZioz2BMw8dL4YkE8Rjs/oJQfo7lfTm+xCeN1455pimQ++9xyBf9mKL05kM
nH1qhdXokqCXn3/Ye9lvP4IYDSETgR5m/z/+te2h4lSSp7DpwoA9k1IVmqV68EN9KQZKNojwfSnj
4jaoHoLNuDM1Gl3OlbvTrteq/7zZWSGnCTC/zEt0/syqpwjSQGFB14v8hnOSyo+GGLVyR0BQxJi3
7/+SUyqXIOD6v/wQO7rS/mcaYJlpwf5SNgN87y2VlnrkBILorOErwuClHtmk2V+vsL5UTFG/0oJP
QqKVwXVXZ+dYMsi3WRzot1xW71IHb4oXBvwrFKvOT+QUqINRhXAxRdVmN3uHZO1g/4jk8d73xUlN
mUnOkXRcFV++rn9cFqMszQ8JlELxobgmacB/dkr5D4hrfLZgNDqVQqwtrKJB+EUi1VXetb0qgAjh
yVoxBEkrRmDey5x6rP4LV7PhirG3yJSUQlP7Ysa8pQcpFujNlg8SEJfLUW1QtneSHbk5IWPvbAnE
j0GmG/luH4ZuKg3Z99l7/qyFxs83jTN0qLNSmQGXe1PaIyFpt92MoLFdFc5A8YpBkbQEXNSbuT4P
FRHkRg6S0trCixBT/74qmkGm9fXQC2J21MHbnOVqyTEQnZZ2++MP6/Ymcvw8NryYa/CWexwp/9zm
LFLg8U3qHU4jJBgsCgPtFzO0oycYNyMsGt6xQdHYOjSTdlllxRLv9SkFDqCMLCInnc/eKiz6tClP
wB+ZZDkoZWy/ySmc5XZ7nk8tTvFbgN4e3EyGVPcKk2zDjqs7a8mc+4gZUxpVTVBQZeSxGU3pgmnV
IWCMPTEZ6QofL4E4trUZSbozrolXrHf3XbY82W6LDhqjJB0ZU/CeUYBubQF5iOhEUR+d3l3BExn+
lcOyor+hV/i37sJESwgn/VZ5FZy9HdlnDzTs8eM19MWLoi2LMviDrglj6p9mmha84WnAGXdLJ1pa
SYAVYd8Bp0JvYZN6LQDPeMGJqMT+T01c2NzWg/PXSLlAURAwt7YcNpdSFtsmtOJOMLJFzxxiKDO2
5gXv08SKn0xYgcJh6HrwHFmB1z3WfNfyPJcaUogkMRg9+M6qBj34J7GDw2iSmWXUOycUEFTD6mw3
nVNo+PGksICyssMPqIhG03vOiiMKsFwHeP1vEJeWcc0AxkbRFOaYp02SJPV6qSIZjTPvpkgRmGZ3
/ZzKqcLLNWWyoYRnClzOInW2rQxKv9JCzKIKt1QlirjzqF/Z9+b4tWITy9dGneMvMiA0c/YTZ19j
XISsIaZS9q2A7AGurVYKXShQiSV6yXFNy5sy9AoH6xINroBvyZwW+iSFag+ZVcUky4H93pVaqwA8
iMpL7YefD9rzUI6CO+DhAx84OOxuh+GLiiDxCU0aCYjabUhZALrxEVQKQdvB5PcsRInF+srSsb8k
inb60A1KrhAZDAvT/iQquINN3YPeO2UoFdzrBXhj/Lrthze3c5+Q++rss10300HMp6WAyw7T8Vhl
Jlgk1YopZRpzpO3l/sYPNcGqIOHgoX4ciYIEeFbrQ3I53qrFFcDfS9Xsu8tjBoObuWqZOWEfpar+
VPMskgdQU5WzHr0hrfRoQwsLvzoHqWmbd4v95jzYF9q75f7wAnSXlJBbbNaO9MP8V+6afB15OgdH
bJZxdmMHb4I0W+umEaq/+6ddjm8+OTwv+Z1Adgfh3uvr8T5SQ/tN2BHOFVAwS1sXq1nXm1crcAA+
MsgM4HzCf5lOYKESWo4P5J4Pjtzg18g+uHTmAV788rkU6olHs6067utqKhFqMLV0EZutAw3nMU3b
29OX1CaGGbB7f3iKfjuh+3K0B8Z5qO6G9h4xBo1+Kk1PK0+LvCqHvIRExUdMJnoLZlYR7A8MJAKl
OJsiy7vPXHFor539F+KdyF+kppjeChXlglCq/xZ5UpL1GGl67JESUOeYrClf7LF6Bx0QRKQ5DLj4
ycUeKHRTB2Lj4KZDUXJqbjVgiETCRg9HBhAo7L0joVbpRqmXDtUMAg31EgCzgZmDLQNygF+gMKQ5
VJWrDx3vCHnBpGNwz6X1BkEs33joeBpJNYVBLqQGSOi9kQ4xAlljsGcrOE0GpG7BcxNTrvWM+BD4
y4611EDh3VacyFs6Ums5lCBHGZRAxFDl8Vxj3WKN7e0NFgyXwkYGeTmHvp4ErexrcDytEyZjfF/4
OgDcRukjUc0Hmy4v1hfAXDvAOKm6HJVvgzX/VxtW9ASUDMaE/oOleNT+cHosHq3+LQD4So7ps2JG
ZCfVQaifkjkhGXpX86Y0pEoQw3qqdovbiVWLqBcqP98a1GaCv2gNT3/ncl5E9Ssn6OTD7BnhCEoK
XMHcwJTs9PZILsYrjduUQx3FShAhHi4s/HYaoUe77slpOCoCYqKMACs2KvnHan4QTu8842LinQe+
2QSa3l91oz8SUz4sPQ4Sqnmy3ZRb42uqo7ubvMB4TltTf2MPJQlg+fHFE3bzmeWdQLpxGTZVYNBw
IbmT5jGmT9KVZ7L8MnBjjxxQQYWbHbiAslvvDfXgG+MLbC49HSehDhWSITMVaxqr1s215jiZ4raG
lyHEWzHU+bB7UpOSfTTi54zC2zWmThOGSI20CdasynW9rwLXPiMAq/wfPmgoxINeE/oi8JvPk+Qw
XpmXm7KKnnwSirsUHtHGPL7oV3Px5oiwIZtQT+scgUlXPQfpDfAXmp5807P4M870sbKmhUVlvWQg
InmqmijP/WKpmPFN0HXjzzqbQx+0OsT+5nMgDNVkjDjqDTLCBqwdNJMPhgyG0v5DYnCJHAd/Cj2M
xLoKReiCyHdQugpAwARv5f4Sb71IO5Ip5HkRwQQbZ0HFxDMT2naU2BqYAAyUdFzBiAwaMCjHcXvS
afVqPzseynuFe3HwIBvKjOEUAlCjh1wHVXFgZfIGXRdIkVyGx4aLdT0LEhfGI3eiZ5ZMMEPA7jm/
VeD0iQunMCA1mAkya8VsHSukyOnoWPWXVwEF+VYUXSm8HTh2ZUr0iSLZGog/EjYhF4sXrsHqbZii
FfLFccEJDXkAsWvkSZWFUoubPVTPx2poojY8pySK1Qpk6+dSAYc/zIyqZpd8oB+24BXwfwBM1sk9
DFpIA6WFe+sWNkXlu2cX4QHf97XQiBRSHuZZmU/SLIeMh5LXthOiECEvyRsuMiY7bt+372+H9Dk2
tWt7t3ZgE150shRtYSSDRBRdnRGs+h2KfG3EADQcM7VGXJyWRn+weSBAZt7RV3f4gKz3fVlc9tRL
2iW5G/bNQwo4zHDBpYWl+ZZwryUX35hnqvYTcXGgwClYgKaJaenl8o6xDOsxJYJ/b1Auu/VJTnNK
d0NSNLEEyVvARuARu/n6bSdyF9OQmPsTAwdQDkiz+LTM+3ce6EM61vhCeITmx4y89I6DiNnCyOZ4
2Jh7eugFEPSMkaHVqIaCltIOr5dB+5T+vOQSE+hSyNnUfPF9R/CdvC33oaDRQ6kCG2yC+ZbOBEin
oaf7ZAYbSLyOrUum/D5IwgJ1EzMXp5gTExpje+K29IQgUSw6rc98ziJRb8+tyKatyowpSm+ufKqD
xYkqnzXRDpEvbIeuxFd8CSJ0BwsePnRYyn7WnsxbcpenRl9UChXYoKNWxfXZtgWQyB+k8SGIHXD9
l4svD/FBgkyUg3PxwMKhmzy4Klc8VgagJbeuvn0CAbJ2c+hBbkq/W32DYpmFGUourVduVVkHTF30
BkIM7shsS8pmd84BrQq8Hp+Uxc6HOBFkCkzQ9WOL3NDWdADhOsDf9IGuOAYJCxN+8mNE4Xuj78fU
Rutl2HtpAettxl+0UOiXNrMc23ZXZpgGdQf/Nz+ZUH54O9C+85rD3QtrZcxiPS4jwvbfjfGnd8TK
cCKFTxkESHrmoS27Mdcp7Z6aSft1tKwAiKhImA1BvdhgjSocFb3GUac+ofCk/0SoN1p9YZ3xRcum
qG+MlJnPWUGFIwBWsvoRafhhERM+O2G4EBNh7TRgWPaqIcqLea9B3VQa8r5Z9vWe40KmT1ANoLLB
yxjLLZB9xVqrmzf1rYkHN08T5AUZbrDzinwA5bdFvvb63uhhDqbNcR+r1VpwM13jUsIprPe9jtuu
SsfswWsV5geip/27J6pON202c1YVSH3yIZVbvDzuI8xm0LAzRKILVKBajq7bAwW8yXdCwqPRdjAf
RsYX2BN9v4sXnZiR+REOy1X4rIQ0wqcvso5klfwW9sBHwmhybEt/CPXfkIX6xYgCb5XqdLEoLKwT
5g9g9eN2mUkYSkYoZnCyhCsDzL90OiHUMV9A8cf9U9PmGRXxfXnQjb3S/h1Qaqkwg5q0NZ4mdHaY
Q4aOSfF8bT9mo1ALOh/+kDtdT/1tSsYEQ+d+z9rMxMYa1h6lGVLdnjLrOL02wQYTbvHeBbgveFxd
gEi7YylHOgvym+mjDEIowOW31sKr01Gv9ntkL6rXz+oRHBpIC7ql+FzurpeTxVRqWdZkIGu4C3Ck
ZNREuFqltv/4uQy84Zo1NMUuKRJCsKGfXnfmgoQHVqJJK9Q/TTPBnDZgG88wLSTTb3wAbG/KyCST
e3DbQaYN6fq1w23EJwv1Y7E8qkPTsYfaqBGk0Q97l3wP+4/jlCsdW9f5AExuJ+IsNIrDrcadp+Zk
D9XJCTnzXdEMc75GXhWCSRHgbax+Kh9mgh3SJh4tE0jtKLecUYyjXmhUjepQSVQdE1VU1E02WkfR
Ue1VkODAxtbgO41vjATBF3GZM1IEP9b78S47VEyJhAyGTSSLOvD0zkBGZVk7fZJp3kkVZ9r/5b3J
iMlSZ6mr8BYqk7wu+7aGX6Cx3HJRc8/UfAg0UPJ+2zcovgrDJsHctc4yLljxNhD+g2frUV/c4qL+
EnGKVpB9y755JqvrAvwS286tLDnw5XSte9pMCGVLQSBO03FA2t8g7xfCbWcuoM1sV5GDgdHPnRLL
F0eB7ukAZ+Yiv1bKE+cah9JfzLA2Uh7X8luidcMie6YD37hoRr1Zh/YMtI+keGHOWAvvQd0CNHWw
gTCC7/2orKbQzxDhwXomT3CmetdMgo6GYBm4d1xQM68pmT/ZMKpXnpdgdyNCYojyk2+8JnT4BEGi
YO0O0uvzL/0zfY9iroEoRy3uCs00NasUpFbbrhqdkvmA0Hunb0h4V54cdPUGtApxU09h81ZCrZhl
4iaLTUTZ0Fg0bNr2Hh0FMdOWM9UxW7M8TzvSDovL6WSx9nW1fGaxk3BT+qeF5o9u3A0nohfmYCmQ
5L5OpGaqW76YyXPe3UJrOFb3SCtm6Mr+p86uHpLpmOSPCBMBnlx3X3pulETbZ8ub3oLyHudTEyWr
24XQLbn2z/okrgUCClovR9RKa+Xi9ds6ftkv/qE86S5q7/CasyJI1PNb1OwJiD4m0z6I0ULsx9NQ
jMNlAwfdls4E/eNNG3jQZNkYHdmJkMWZwMhKsUY6T2H4SHKjsQvHr88MuP0wxI+c7fgroMmao5rf
RILyh2hUgMF4SzOgQIicNW2brQJMr+EKQBD3PlyNQOcTErM6/VhuYBCAvxe/5Fnohc0e+2b2GUUX
ugpQ0gXmOmh4q6P02H3CyhJb8ycPvzv8/oy4F0cOc04cQXDft9zoIrQVXgHSRhhzKsbzc2wx/ECf
cK4YIOQLuWjVme/uWPewyDn3q6dPhFKyNFEJuxsrTy1PxNDX7o1HX52GYMG5qqWzNIuQg40XovX+
HWjS/d8gWM7YPlouabJ5lqHd6xYxNulVWHtigitzmdR0cBCKlY/lS1FIF8MzCoT54mCL6qDQcr+k
b+eESlAir2bGprls1CHtvzlz6nuHS/42JF8pQKWOECBi9zway4CV7I1u2iebmHMgQ+d5xaiiCl7j
IITHurCM+lKbPINo1vpgCNwvHlOfDvi9nU+aPLhJ3f7Vf96deXEtPOEwGgCx3JFaseFLBv5fcMVW
JMo8KfdtCNbh4XoukWsSs9l6Yjf3DZHnhBu83hpGj+FK6E/x+LU6HJTAVMemw1/NvMl2cCMi/EDd
UNRkknK2IuAvSNI5nKV1bYgkpTPWXdZeop81vILRzKhoo+rnhUUOi7NMPFOvk5eK/s7S3BfpyGxo
ipoblv3qMLtP2wBgRqLjq3GcvFtfYvQ05tF+PeB+e7zg9Ls48tygT1q7hFl16aGVOqTj6mVWfxMi
eH8zzJExF11Io7Thi/lHMcxDOvB5Y61+3qVGgo8AAh3seEaZPPNQOw/N8ixqkVgixyL8VmhzIXWj
PHsnwpESaE4xPWI53nXMkvfNIw1x5PJPzzaeVnBiuCILyj9gA7Zn2wSmWUOnwv8BE2A15Qb74Xzk
8pSRTELlYmmHx3Su54OYf5Vqc3hqfYzSaLFEwzBgWj8qYdDkN+W8yG+bc8QpUZW7sU5o5vsMIFJa
u4kSokFnluzOL/lw/Y/sGAbvLpLKjWXSVpBmD/pQhit4UotXAyngGewxQdu8hXuCHQx9A9q3MlHq
K/+4Iy6xe1uFsTKQX3lZoGTw/mpkx8MmOvVDhD4ZkNqz297nIBUt2N2rLZJqjx43kshLLe3tuVBD
EXOHC61kSx3arqQGbAJs4jQOhxRfShf3c/tJGgDKBCylGdwmW1ELq+wDpSjZuD5jazblAtDlN+eE
J3ygA2pAm3PsZYrbIvJTV9/bewLQqvqiCVS0/Lezz4hNrtMbEhdpZzZGJaRgCCHAyfBUHKOLVR3j
N3FJlqykQwQ3PEipPh7PtK485dwnDOhLVnqEajb03Ny02/iC8DkVgLAerSALDmRsAFjl3EN/l2Hn
uonmV133120rYXPp/ebt0YUv7o0eXI8WicJcGg9ItIugwxTz76EnVqb4VKzy2mN7hY0pO7KGnTyu
4yBe0+qVVkcVm0b3Fpx6yQtXb2ySuB/Grp+sy7nEILIZvhUEShnDq9qX5VaR6s7BWW8RcTc4EP3p
hpGQPiaHv+nuwtS9rkO5UP3rh0UXLr2bLkjeOFEExG/hVQfgFzLmHgNKUe270vtGXwBWQeIcjL9/
rGQfLWZxdte1iEAS3umiYU07KgY5dSN9m6Zxu6eWCBeTdY17AbCv9ljkJUbWxHOZY1F/hTjVtTC1
cT98EMowlM059O1i2tDCB0/Ld9WRtyENqm6fbOWoauTOUrDCxyu6FKeZm8VF/XyoG+kS+W15gaUO
OYaNz9UIHkle0+1S8P4kkmJyT2jSduVO8ydxxNJ7/luFvuNbUwYTvHKx8vxM1GGyvm4lZ2wvXOAt
QXvuJ53VHLN/+yCDg0zstvXWeQTtHZg7mK7d0PfnjLb7JHrAYYnlk6H3d7hOXeQPx4Tbpz4iyoHX
L/AYoRLVyk1hzLiCB9i31f+recExxCfygvijsgK1VkDbfEZW8JqGcxkSczTCtlVmAzzVWlHnXdmM
MLPEzBEotgC6L9cO3KfsyKY22sWxuXsE4EP4bx8R4A9T5yX63GHeswm5KX38edo7lS0EE4BrJIh+
sPeXZVm65058VCuCXPeDIqsseXSa6Ei9ZjPpV7uV86Wcru6gd2I7cIDPyWqwxq51GCAvqBiT183M
D3GUeAUfJRHqm13GB6EQ3dIk2sYNfqm6r6St+hIEZyL0tFVBnnc60DgFX02olg6WUFf7B8R+PvDB
+TTRWjInJ/XWVqK3y4Euz5yB1hweyrHtzWzWXAtZ3FvdMGAEbA/jjbjJbrg2UKdvGk3ggIrX8fJe
vJVTQHR6cWcBAza5iE47IyoTRztKhdI808ITwjuyavaDyam88k/n5B5b983xLOEuya0aiO/6V42d
P5cl+GWGE8OpNn0wQwfN39vq8SuEmDqLLyl4K/zfgIO5/2hTgftBrUoIZO23paGoi7X/IGWlAFaD
U4p9f71VDJLQZ1FJahFaz0RSkNSIOfDYWjxT33me+1OXhWg5S1q6NI5hrliullFVh//L/VmJFNAD
Rr54FAta2czrwfyzQ9cdOZgYYytm4I1m/gt5b1wEOhcGAEbwQjL8/TQlykRTgYlU3HXA8BCOczdC
WcsYED7RwKeb2ev5UCdJN64XZ37a7ytTrTQGnZ1ZfDfgUYyLiTHF8bfQJb6lqfmKgT7nqOrj9qTV
d7oaJofhEqxTBxgBYfSr1VG76tR/RiUHfYOLHkNIoMLmwknicdVq5SfjVZV/vhVLBl74GNnJnIqK
fmF/f0AlXNRAauPGDb2aEpOmn1SHU78eASkdts5ra3+YR+KzHLZPUYdQp7ltVUMyMIN4Imzpb5it
M1wLEp9m6fTseQKoH0lU9AAuGK7rH/ILQ0YtryH93DSOzJua96NewFVTvejZG0UhzfCyL64maZ0M
gopn2cBGEvSlcMQhXoUDDpynj90OLxjvXz2MTg5hw2eDpT4pGxlrurlOrerXLwjeYEwOc+Iih1dh
kfp16V0bsSu/OcvjPh+BrusOgpgKrvV9muWCCOxYwG9ysZKY692zj9DWhYm3QZ6GJ+Hyq4dovFXl
xYh1g42R46/f/LvhowvojyZQ4Hu4W7rxbKtauUphsYQyG400eJTmWRe8uoAziqHTkiT5ssR1cWIL
MqH92epz3bRpGc+wsaXtXnLx69xBbhOeyVmenQw8RmdoaHog6UfSLBerQovM2FH+H31CJ/3p/Hns
4Rf2Heca5KBXRjcjZflOFsWMFHEEjh1bOCmWHJJE+JbO0kH8JdO+3a/HLd8vAlIIjKde02eXwJyL
Y/IKHad5UwDuBuI19EGmS6rtZprxZbYe6IGOwSJBKMg88kazm8Fm9kP5zZTTl7xbZgljKlH8OYXe
08XLL/Z6ILqhJQTa2ZHkmG3T90jdfrd2ZAuO8guBX6VXkqPNTnJF4o2w767pLPQ2f6wf8M/vhIZ7
/ogtlaQxYC4qByij3FZ6nnieSINtYI1Q0zyX08XTfhpp/aFHPoe23vZ1EdI7CsdgZxhngM+UfJys
L95tZKE3yhefbAnFyMXxTpcZmLy2XCex6BJ6uKhdNq9Tep0FzIqJDLqnnw0+uAEMWZye/ZgEpCXl
pjFQetlJkju/MIqrw2A8aj98vw40+Tjggrw0dxSRqPzNZDQMFNFhLrX7Tam2fthg+cocDfwr6lFX
L7ViePNoI36FOcKqwsu8YDZBRMzTR+C6yz1GiG3keDqmOyenic8l7WArsP6L6EpH1TN0XoUORGEO
Zi0LZVKWTYVRak/Xb//cISBDhqWGc2uewD8hQuxDRN2uuR/xEQdGNI7fAy/UTDTp+THdvNkDXWwL
lNTXgBT3UaI+/fU49LjsQoRP/FMjHbWZUsSOGH5X2qOxN2Pqy8NMR+nBqTJ0FQGUOdS6iU21N0th
quL51cXp0VZRTKfc6NmiG2nJYg4riLWEmnfG+VThEyed0dgzbVjl83CnzX3xNufmSPbLwM4R04yU
CtY0S+juQSQMtmGKgsLH2G1Yg9sa3283PebQvoly9B/JXaz7IBJQ08IieJMC5jxW1wJKHi0P7NUb
9NCfB78lzs8TSzx5RKFoj0pkfKWsyH5JdKHP8w/ZX+wrakt5ZZL2Mah3EIEnVajiv0NERlRVtas4
ZsLYwDL7VG2Yz6u8sUjIbXzXY2Xl8sHmaeeYqnIozINFn2PgBSmGt4TEBZK3vLYe7aa3tHsWgk/P
8kazHdtiWoLmK4eEZcqpe51+/lFUUBg/AzmuEMT/drPJZuG+xgWdKQdkcvTV7fXI38oCL/jOIdDW
yW5Hf+ZwnL5uLxm6ArPtXBvxPnOs7lm0AidbTTbDZE8308WYXSc2pw5GqkPfaeWxgVHJaE1NC/Ea
319p9XJYV4V9zHVQXK2GN52mkakYSxXB+ywXyOGN8qixXS83xhAUmm4aiD9vYiZlOAy+2oHZZVgY
umq27I5ZxHcbUc6QIcQNmF+PeizzQp+RHxn4y+e33HURVaH5lT1dwKxBXWJf6iy3RznpAixfByK6
wbm7s1SP1fUhDL+K4KZ3/FMz9U03CLFEiayohE6YguATP0hmoMZ9ZRlrJrgH/fi/2E5v/a8ZYz6d
Ax9f7VmU33d68UywSDdhFM515oI8pH5Dvb6F+Ci3j1feyXF3idErq/r1+FYyo1NnuAeYI8gjs4Xm
VpNBhIHC3QLJc4uuZTsBC6OKa11nt/wuRe1c8fX1/ftTBSBhkLRuoV03eGtRsLcEekrbaVfzJhtT
hx65R7oV25B9rfXyjygiq9mPV9u0u+P+P6eH5padi13eE+IGlAuPlVYWJo4lifUyGRs6lQ7s0CHI
Wg648HDXm5rTjTcC8vOVYdVTThMJloPz+1YJyQ13jdL9Nf9W6X+1d2J4UKr1DazvEJBxUPCFyLPy
t4hqGfbMmU2cakjs1VIMOfXU4JZBsXeBo1Zh7wGl/ut9QN3+PT31bvSrhpXsY5tlt5hGIkYsRYSz
BzXiBwouEfs43WmKnsaBIXJozorR2UqKsPbxhgOLjbMHgvFBxqodgvPZisti25lIGn12sQZN+nrL
XW9w5muCWCfYu1U1/hDYq21+9K6CRDYbFxW3BBfH6fsMRK2M4jpZ9vD9F+LsJf+hkKhOYdO6UYvT
V9TS2RUf8oPrixiZdxBnEqXaWgHg12QNFcY6Ix0EeRI25fIWdRv8lyB4YVpG3VxsSna3IwUxbEGx
LwWvTzCV3BVygRg1gk0Rs2w40MqWgY91WrolGOSg3rTzR7Mfmxp8Q+WeOUwTSh4hx61CV18yL2p9
rqJMo58b6gTJv/WOPPVMf5kfmSiHExG5F7zvPuKwUE7n3cAHQVIxKLSN70wDxGhMnYH2va7f23IX
JvM40vrVHPekCK15TCBstZt1afG8H12057s9q46quuX8Vl+OZ8X7Bf4Z0qc5rkl31Vk9B1z3qFLc
Qi+rJQJKHHhSl1VszDs7OaimZZHan+nH85+NQftSpNoOaIhr7vYliqDoURllMqZPivY7kYeOFlOa
1fsps0MXsBIGm/yO4D7g0VZhJzyt9Pk9WFryb5jyiLnTOuCPnrpqwV/TlvHT+83XDC99Hl+lOMuE
yyqc5ciaqTCNGiBUBmV3mp9LZCH1KGHJzca+6dXUue1Nivx8xppxY7Hiyzx/qdFmUjmCEPElq3EP
m6JWkTvoP4q4V79tyBY4MsJ6QnLH2RokpIamNwkBP2wj0jLkRrSKt7sDYRGlYP3lkK9TxW/lhMhr
zQumoiHyxcgExyn1IRw9CRfXznvDDdtlvdeTU/e6tq7cR3fEkvJE9cjna6Lnyv5efP6x1TdUvnwx
eaMwIsDJcZ3tVA9Udrbg8GmTxNtzbsoABBze15EUfILYaJuF1RvsZcHhGQ43VV6VAB4wnAvPAbVG
mVQ5ulACZmLZHyITBk2HQsMXBUnITkE5LZLjS1w84eKohKcLYYUcIU4RqmV4DIlbENEhIodZOIsM
N7V9/vl66tM5Q0VLLJAYpK2ZCD7/jGZrog/bdca754FKBFP24IL4Ip1cWUNVDDpIBWYBoYaJg1Fh
ZdJ5zHn+8KtYbiQKZP75F1jvd7S8NLDEIEsE2IdS2psrT9/2dy/0fx/AXSIDpSscwX+1qhLWHPJG
5Ilm2w3yHg3DnWK+yrR3Sj6HReKAq6W81IXcMyb4GukWaNqvt7cRnvnemtMJV1shlENKBptp/jMD
9lFE0FNQNMuiUQKI6/V9Be2ZHrhhqr3Ct2aTKbUphrNthKlLg3Fuk9gZnnyhp7OgSFDO7Bv79gnj
a43AqTnS32iyZc0xw242o1B42XkBJE/ExMj8uKUJzRhBzme7IleMGqjXvoJrZXpibWocHyNBRNrm
CpTCUAMlaflQArL6K3bTnqQgORv7Tunn3SRSFU+Rr8NBpT1kQSXqVUbljVDJAq8CVMe3XF6ojrOg
KJ3mPQKYeCEs7EwtpgtNLQD0mUFOpvZ3oxiQ+ynbJMJ10xwaM9WYjOvr0KSlO4DksblafPiB9DaE
t1wSFXbMSf/1OGss6WyyElBXTgpFR26N02k0e0Z2G5z3hIS9NG1RdrJc69YX5kQCrzGObL/OSgg3
UD6bpvQvFbtMaGfIVSLgL00wX7zm2hCU6LIMkEb7PYhCTFxtUP3pHAXWNMfcPk0wHzBKsoCP4BUz
sft9+odyxZwMahyt+50Rvw6ZCRWYHr7lIcbGLlVhZblCLMz0/Eh/ZlFGHoTtU3cGiH1fp0znBIUu
m72Nj+VZmBludtimEJWfWDO3AH4Ky3vNhO5mPuxAPrvrQpURk2s6Td1v6KyGU5I03foDF8wjUz7M
WPuHpxZps/FfpYtvgz5eKPm21cwhxx1NVT5FKjf85cUHfQQOerV1mG7UGNp+dk7nKVL5L9cKo8dS
R48srLcZWaK45+d65833zZ9yYqKMh34f1V5tBSzXXRyz83R5VzU9S2GvVOyY5RO/ADBz00MMzxK/
G2WC22mKQme7LTcyHeIPNiHyMUW7/uLWHbPTrCFD+eKJ1jKzda8FV/VKr21qB+v1+Q+bGiKS3Ohw
fv+DvBS+qcN+WSIU97QUor0B0S2wLbKk7dH8THlTP+MXCCYPQJRSBZ2gDek4pYojFvMD9KANZTjs
WE9uNRuNX3F6KaiSW2IgI+VtqW6M2Jz6Y98JjCACLE6+EhXBPn1Ghda/RCqUQGF9vHdDUh+4Bsxq
xOdEGoEYWmOa5AkLRFaSytMXFOxm85FfBrog7Y4OueN2Lu78pJRUGZrz6RMbuIlUQ7VTm3W/DvTo
9nyuPzeglptgG4FIVeVJ+qu1lsUv8n+YbZYSWu/ZtSSs+cotZTzTuBnPwwllkEl/TqAD4to2acUv
fPO2pK4W3GlWv3T86TRPh6HfgOsuHLvZTWHPH6YNB4RWQeAEQAVbRp57Dvbc6fguqqYvNaygbXVc
2W+flIF6/e9/txOEuJA4NcfMlKpQpMzDbu9xsTcnaKVdqGg9hx/8v8teaVo+uKdS8DLSof1NC+KL
pWdvrlJS6NGqffOBnlxYb7KDgSqzQSECmjwWzewLtdpowQId09rA9tLR2EFwDAI/hAgSOrocFAh0
bDRMDi2ydeFA8fdAA3BAAeuqR94HPfrFoZuEWNIEmOh/1JqlK+P3pfC+SW9xAR/hZrCetdos0LEf
cKfxsLU/ha93wT/5vN/9w7huwVf7UyNsV/QPFD99h+wbq9yxeaH0PZW2Jf5Ndos8vaTddoZ+Exfr
Vc+PBxfyb8Xicg0KmGoM1p1D4oMvUHLX2HESlrjFWrl94SJet8GRPAylImNfDP16kjFHkhV5fCp5
3oyBZQpTueuSfeSByrEW7YpLd6hGohJu7CAFGqEjgy3r5PdFTBtVIEXZbY7urzt4xNg04y2A2q/C
1QkcrXQZUG/4xbGaZk/TNdCc4JgPUzMCiDmy6JFz2vmNm74T3nzNVCeo2HUpvP2mvsNoWX9nyOjF
gAIM5m2gQfrU9vRWkqmeNscRdT7PgHpiS1r8pTLhS2iDIYN0pv8ewB68SvB4moL4g2MegrSokOMT
vsE+BAEOSYHybnyidQ61YWrk3lvBqMqx7/6JFsVTK4YkRpq+dtkG4dVWQqpi64oA+Pc6KEg780Rl
5YgLCtemjpzG+YkOyjjm3CWGfGgF6UsYzbgRrVCPRl9tw6QO+dUb6AGAI4yxuo50kHyrs3kxQHjn
7jCt70gm/rU6z9u994afSTPlvMJlnkd/wlACQ9yPjXJ0G5pagbx2BvEfeqxIHSYVRpEDbiy3yfRQ
GqIMXSVW9Jd3bDxBq+PVJ4m/HHr2ujuvBG6Vz7NoHCnWrhRAWo6FackgizAJ8hJFwa/Jk7wqHp0h
4hZsRuvnLO6EkGHL5nf2fL1h9ST6244BUdRz33qDUv5Zj1LGggkjmXIZkdZANfW6GHoSRTHc3VRr
DSj/jek0JHaiT9bIB4uxDq2CaOyBQfZBwpd2jrW+6+s1oS6v8KpSj8mPw94uS9Deisj0lR8KyHT/
JWYTngAuo+L7vL0KhCVFlAlDAvHwP0jIYLLF3EnhtnKA9o/7OUFwj867cUgiFhJ4PofsQuWsizWk
mT+TDl8D0+FHri47PCyjb/oNpsSMXJLdaB2tcs87MdRVoo0MK+JRhjrM1z6H+4g8LVUrYLJ2gxgq
BgvCgUd6Wtp5HAcnTHxyIOhpm39p7XOdqXdaylIkEr6yDMw8DMB+SliG7MjFmpmaeiTXxmT+empL
UkRfdgZBfj9+pe1zgFlH1GTY5iLUYmyAuqTgkcHQ3aQd7pqPehvoxT9rFPo7WRodpJnNa1ONt5d+
zbCM12mwLGcgunWq2RVVw3NQ/iReuHjqpi/ck9f/8rUaSuQMHVhuLRBaC242EXbv8HDdyxQs22xT
Ypx8UCbMMcwdo1eOB97ExgmFlJGKKDL0a8yXw/Xtfaq9Z1sWrDoNN9e1PspXlPyODcwB8HaUxZcU
qMHOYvXwcnVAJ/trkEm+1A1wbOxnthBFteb/vkBEy2REJMSJz/+PHWXduRu2g39P6Fi6psDPFmKU
Rz65Gvr7yiy279T7PiaoemaHNQqVTNak4Bs8a/kRAlBgzjjPDyACdpxqk8v1LXtE4lOOoCSsVSwT
XxXb/zBipPPLjQDZneznTrEsvi9GZXAmotikrutkoQDRwLZO1GYIBMQkXcEREBKFEhPJyEeRtSTd
lhoGOSNqo4beuaKYTc1/oEOylBjYHXLQzfdOCfSxh1ojCKauOH74F6UZUTfrlMDzVUM26l5X+/2w
TXlcuGX2wJlIHV72ZnintY14+d+hB55dDBxhsFyyhFAcVxXEnKR0XGONI8994/Dvjo+jg3BD883A
kApiNNknql9D5DloQkVrwx0w4c22+HO7StasrG8461gOuYc6Avg3Kd+qo9oeUCi8uryCw/ClBCdB
oTvFctuGbCKZ30M404dKfbtqK4FSqxJIaFBqjclperKLH99kSql7HIuHMzaYJHNbKHhIOgdq6xeQ
4KLsqCTZWXXv4xtDuFpfo9yPl0lAH29HXm+kbnXCeP34vOMgGCazDJAOsXI3PuTeMZxKPKD6+Y8d
yNtCSqOdzgZs45gzDYO7pboTOj3QeO+5rcNa42iSdx0BjzBQwb6S1lD8xu6mDP9BjPGSEHrrGvBp
mJZ2VhhLkdIaldpWUX3NJ88a2r8WIR9Ac26XLa1QOpb2RKD1C9Gc1xarpaHmpB5tq8cj5By07S06
mN9XNHDYQZuAl0g4EV7DcgAxwgC0oHlZyHLynOVat5fScx+LYsjFqHG7MZ8LzNxxGGqPCJdYcxgi
rAIJY1dizJT1qTVAjKtqtcvWK2LQYCIx4kI/h3vFAmNI9EEOLcur4GSmZAtSgv9IUJ/AcQS2ySeo
6ojD8hy9Hfa53QYDp3UdoowqMKkmfPxj6J2J3BNdJLQqa4HsbOsYm1c0VD4L/IpC3X6MMwlyqLy/
+9CwpCePOc6MBZDzUstYaKXodA/9gFFVGadbLLG/BbnK9pAlO8WrOGAaPVgld3fkekzcd6F93K2H
torcyb9Oq+QN9G/+IoQLlZ69DvTqrJwdR+5l9RBQbVkOsqLn/E6BnG+o6psF5hE3xWdoMdIT0gM3
ZmJXp6w6a2VZiCuUfw7ux9mIr7jFs3wwnxBQgdweksW6RdYMq/zzMdqWAI0khwBy7xdFGxB7vpAf
ZTx6rRk/O7I2JA3//GLlAtbvMRgWOPMK5YUGVySp5/cY/GZ2lVIP3SBCxahCGrPEbfKCdhm2ZZqp
OFqLKcrmdi/m1aKwBEz96m9au46z4BNAuxZNAsVR/4z5/Jhg4mj67rCjR7rwZ8tckBowuvuUYOBw
nKZvA1se8OoqCUyY4o+aBu8RYC7/o7RHkX9T5kUQa5Hu6XQuJtl31lOAhce2hfeRRknKTBjIn5bW
yy4wQCUrtk5pqQM4tivLePl6bLPtkEuw7UYoH9KgiQa8p45pSXqotLC2Kg9mKvgxslJWKCLP3gle
pWMap1lY3MAHb8QbE3+hJ3QSEac46+1XWiT0MfBjxOt9XMBCfD7yVvELAHHDWuTJvglrqkeJ2rV3
sBTGwdTrMsvvAMX4k0rPjYK61tM0+ikpwGzl+muZSs6jE9vlgU8hlsy290WzURD6GREDnATR5hgr
PNcWAThNh940Bg72rBfV48xbRfj+eCPgFp9FYlgfEhApljcvsdt09cwpgtgtCjIzDOiVE3J6PaGp
gIWUJsukEeFhDXhDtsKRVNtOGaz1YyHYwz37AwfTgiqmxpEUO1Sw+92/KlrI8nFi1WnozVKRsJQ/
F21BI+Z/OVOc9/cK0ls/CylR69oINhfL+A7EotMM6NQfkpMJ2k7XDb/FghK7dDdJECjxmPCy2Ozn
l9mo+Rc9BiRd+tO34k37ryA2jiAuomK74+1O7OixogadkjSNGlCjVsNHZ4f+IEph+eFAY9vUdYkC
rmBum7gjqGP/0Qp0kDq4C0iAnQCrLGTqkRUDoQLKaCYaLpq3iA57wouDEthQCLsacan02giBCiT3
0carNIQKazQvJTapD2fWFufT6fSS6VQ1FtZ85lYBVHnL7cblyA09UANheoI8QK1x7QoIYREWE2RS
YZ+APuaCyZ/cOAeNOss7vJi6vNsWkWbJBfSIs7WqYfNB6d6cP+2z5kfWPKSOiaiahBt4sKrTbnDH
7AggolKFzz0yxU0kCUgHeQIeRfQSRs5A0iJ3w0re0wUJjEY3ep2rOWnuxfnopZwINUDowkNmelbw
i3iMXDdUo0gCGphnO4MCKOoJ3M69eJnhFVWy559yY2LD7c2Ly0okWlv5BBJnI7LBeKIwayQZmoq3
SqTtIVUNYGQSwdtatLgqbEedVYLYGkXOnGYTWbG1sYlD2zCyRRzhuJdZGOsYQJPnHbFfPkWYm/Xw
zBH5gBs5lJl9sjNK+2r8cOOWKpEq2wgxSMp70n2KyNonr+TpjHX+IZqLm3a46X6+S+9Fb6Dmy3cX
5QpK9aImRCjRoX+cWb39E5lWVm6Sx7njGrUFK6AbbjX2RDqZqhx9yRI47Pljxi1qmHoV79090xR+
rZ0WD+Mwb8NBMVLHNDIscNijYlMICTe/0tzT8x8lx/XdVvvAiHOE0+Xc/e6YWIAZ9eWGQR1u2M0j
hM+cFa7sN3n0C8ZuynGl+7tO/BbiXo8QHpQj3wCSYQCxojHp6UvMiKUQIuFHWlaMxdurIBCWJ0DY
W8BEfiW5h/J1UbLLUn79vqEPXdPkebzCqIMHVydxlkMGGG5yhDWriivN7NQQijkevDTviRi9gR5V
nTjKU43HY8IE5/ew0PXj+TIWKhHrLhEWEMVF/cj5e6eXwscRhac4y0cAdGGdd8TReTKN1JpygCIj
10c8MEUMFb3rvn/dKBHNOgGGthHtNwlnbmWcUWm5rkwlYRyynFWkxJueOB9vufXAGweD0YV7a0ky
HLfOFH+eLoKIJMrJxyQ6LxVy2HqHiJ2CdnROQt5NxTKuLJTD6ASCGCfOFSyEmvNBDooT1KXWbkF4
C1v6Qx3qzo7kbZ6tAY8siOraByhr6ZglAdN03TETlVlab4QKy6hM6QsYX07M5ZK1Fxk5RT8n0+9B
Sjx0Y/wQnDAdWu6mCb6KZ0aWs30wUwkLENXLLHlioDhjR94QMEhdnHnYaZJW9+tG6QW75GLCjAfg
cF3gqkRzZux85h01KTcQ76qb2srKtvLFzphTT2hiMyeN/ttg1TCplR/206cp8eEc3lnO0EDQIXSV
yM8/EEtYOEPkQDDTDAH/3eD6e0rrNfKxLKDk3ngvZ08KHUyXEXaUAuE9Fr3b4DvE3ArpKj50lJBF
cnkINNAjli9lF2CnY3NHGFoGTniHQyNOWODMTJzjh4NAlt+qDPb+JzvEcKkdHrEnqOfXJmN9jZiw
az3ZxSxdnbwk06h4bzmt45xFFy78K5tN6UvvPNVH5qzjPTr0f4eh1S8us/HGOu6jr9oQeSaEWdkz
8mH9ulRHyR8zSb3In/x9ZfoZNom+AuLyCuQSw4m5mEA5MGaKv31KmczUatHtVIu+7yRlVjYI54p4
CBsaH7EEwkv2ouD/kn5/sZ3XOxRAetDnO/1M+Ddfx7/6mvdGXEoEOlou2QZ19Mg1pUEEk/ThcCrb
EeET7h/jHi4axDTLHPU5tuhqDLGL+g0y8dAN4vFjSmu1a27FEzZr0g8kLzGPjRk2SC0UMvJHtQlF
H95YN05bseVXCw2mGi/+/22sMNWGeeo8Urqxl4WTUoIHnRm39gIL7QhjVMK1Fk68F9GfM9X0XPTz
vznW7ycSoC1eojdtlzq6YiZHUK0mv25E57r0DPpyeQDIXruJ3f+GqKmD1jfTCe6xcBKTAWsJ119B
Fz0D8J4+ZEghnpwDDfBINkAyI2gJNGpFAT3EA1ecvB3dtMCuW3FXCJogB9Isdv2D2u6U58D5YsK/
ezf9OQtsFl9qoY6dwPIpnxcgOjVSqbRY9bXVO1FYt4yv+I91gIwCJPco6QM/a0hwCBoTGWBaOalR
H6sDCBGgRgnWh9sVSanZ071pNI5+iYg+3NkqPAYq3w19XDaGJIDuaNm9TBdelrMhzZ6grzfY+SAM
Z72B3KOqIqqH3F4nVgFdjaxILberz2rnoZoWJfGUjvgAvkDrZb1TjsLuS3TrF1bLxRF8GEXS7UBi
WBQRPuvjZ6j2toopJZQBPWb7BT1wVsVlW+4PKP7vpgegXoFXM2m6Ysimy+gQu8HndXsWBKcQbLaZ
EhrFxj8g60WfBAdznGhmwf4osNnZc81yLceSWnV+/ihGqF/a4A5w5AAXYVO1jthonrFDcM12PYMy
JVm06N8+Kvbivb5LZxy72p2X2qb3dnAV9GyTPXQ5XkKvXgV7An6J5LQJI4lY52hnozN+Cn/PT+6W
tKr/k7xJOl6MO+478Lape11tFOnFbk+p9Sbe+4ehRhzESNjZW0YkNof+7Vo+a47waS+fEyn8XtRo
46km4DDYCEIX+l6dN1Wd2cj8Y/EopBsXGCmZ8XicjEwgPKzGbpKlfPdST8/Ks2Atj9yVnYPeCw3j
dSeq8I/KHWCAcE5sXDVn+51QJAuKAu83pcLLtqZXbbcrJyZ/IVtEonpmX8Em1L0taccNDO81nUvk
pGcZGIbt9sdH7rlXfnWQMmjO6s5yhyUc6oVUScRa05lCGHpijP7oDseIZFUX/E/EdgPopSorItDh
XMOo6gnBjJn5Tje4lRyZHDdcKvU3IAAK3eIrwZgcdL6kXWna86aKTyAkUffp6B3f9VgbBRUqIeVl
q6b1Ds1TmxpDMYRm02OlZA1ghDzvFLpE5TvfmFc2P9eaPayj/C3bj6ntEJzemqKQp2hv2haeYQ/J
Igqq2g4dsC/Wx6LYKltjQ1vBwoajy8n6CO1qxQvFOlshmBAvvhsF61WTC5MM1B4I5lSDzFoN1zlR
kpD1DoKK7XEU4e1Jo8S/8kqtjgNG/uE6VAboSEr3lGEcaVVto2/HVCfOkGZpz8w0hzKDnUuHTBV1
Sj7GMZXHZvLBa/OT71GYofpAJMDEhg0KHvYw7/c4DsDqZoIl7dtWrHHwosheimUmCw82/KxxhgVr
xdCCHnohSFBlFOmez0fNM5fOM+WcObpvy7VoC+w7/a4PAL/rFzXJ51Xosn4wOdUDFxwisZlru1HO
J5LQak+oUsaPlJgkPaccpU7XPy0ieNx/7OjDdTRmVCdN1GgDzC1AWH6/rJHkjeypg9/+lpdz8X4d
UQHRfszVcRCaGjIKRI51pGsjqsuZZh+TR/tlMRHUx4tJrHYM0Pp1cxU96+I+17k1g3qy6502z8Kg
isqYnM6UAObnb4Vjb8cPYq53N35BpzZc0IzHWin6kdOML3pdnLxMdPwscd0tMDdtCzRIjvkVunNH
Vqt8bbI0NP0/19lZvkDwMhfte0UgzdApNWzxsJYDq3AdivU/Kqx3xITFuGNKpwfbvCAwszgCUwJW
7A9QlmSsnT9z5scjwLyfWdg8edw/5Gjv4YMmwXCwIg7BsBpba0I45MQeQP2UvuarPcHNlMinHWkz
Ky8rj83dPKAWQDbHIonePCQH8LnkOtibPU9yn60Z7IMBuM92evv/26cbaJ6OAk6o3ERr1y1jUA3v
TJ0z2C+7C2M2HsCeLGOvbqWtYq/Qh6knZ8pyuKTqLrIYOpKIPVOpBw5LRx4KsZDJnUb8eboZVcSE
jY30mL0aLcsMjio3JZZbh/l3Me50j9UUh0j3R+jil9Ilm82SAgVMuk6zTzGDwvfDld3NfrzQuSyx
9jCXizTva8lSEp/DUV4VDbH7X25Mhks/JJIzaiMI6Ygihp7AtPs3WUrrEVSiQLfmIfYgYWCQlN6z
6KUW0Dy3KpGz4EPqgAgWDEDjQMEZkHNRWTmy5ISx+5jOSjM/DUQAaw6drtcxfh5/RpcC5YwabV0A
uZsXmxkXJJfPiJE/HqkZigSLXHbm7b7HefxZXSlKsthKyzg0V1DDjJiRUio+LvBZRgYqviMj0qsq
qA1vOaOpZZ/w+6ULD6E7/vIU9y2Oy0+XW5yuDeAbsSSQTyT661rs5C+TgD0eZE335+IhM5ZxnRTS
rlwnyV2la6sz3MP+pY84QJGPfrGZ/P+yPVZzC/q0fg84hvdyRjDTHP4a8jNGtY9TsWbf1LMmXUuV
oDbBuau3YLINwZb5qK1cymZCKq0ZBaIiYmww0yZMOGceKFTeLFeZiUemvqABI1VjgCRAnaQLlc2c
uwc1eouio5T4odQhVCf97aaRu6iU/G9oUJCH2YiSoJpp4z3nGjthb7ihdDnavx9J3xC+NQT3g1PS
ezjOu86AfS3S2CpytTsREYaeRC0VKE+VZT3DK8Btm7yXod4Re+yCYZ7OuySLdkZmAp2FoyQ92Nn4
4SMKONgnTuRvyQGR3h6S+JDSTzUcgjbHsZ2ZfqAKdsXRMwnzSOrb1EBZON7Tw/G3dPsAIUOEm52S
VUW7yBKtqYhPOszhTsYffTxrcL1G8LIlGnL0YASX/xvxRFNUB1iRlMrfiEnuisZlMhyjwjLeZT1t
lLags4aXEVndUefQKDgIB0JVX7eXM7JDH8hLt6gJY6tCJFRlYzPlp+eaOX6CAWF4nktCAUhvyvfF
QQmPi5ijoDeQHC6QZfRWVR/V5iXiPygB2djEdUjERBEQdIFkKB1Bi3fq8Dxn9/yyU4WP02jcTE1v
ST1QYOR2rK8Co3Bx6nzSCIwo/la7HeUCAAML12+lilUt35XqPZCaifcaQ0K4YigHkfDpICtG1l8p
KjHO+IUM7EFCCGRmg76EnOf9oZQrKaKBdVRiAkuKlzVoInEeIpyQ78PpU8cTdAB7tPwwl4JwcOJn
1gqvWlGUeorMwI203THUN2i/asfAjbPB0YQvqQL2MX00buXxfTSvrbBdlktAA1ASyvXhvIHU5x1k
MzLILfloteaAZhntERWr4WVBMOw6xgiZ/pTVxvIVrPJlSUdnt8RC7LXij4jq08gJNFFmwO356gVP
vE+RGCLErKVsXo7G0Vj1rthCsiI0r+FILsGW094BCgPVCg/Tvd+zMBeHhndm4bAF708hHsa+oj9N
8RH6SIn5N6LwPQiq5O4uQJCVPDA+Oh+MFs4MRXOz24iRNOzlrR1uRHYx0qivbimpVls+ryDi/jVW
vMkRZSOo2cJpzZ3xbkVPYKl1IdV3JxD60UPkD3rpCphnIkPQIhmfbfw/SGXEi0/IKn/O8WdTUXsl
JeO+GIh9GAoxvG0Fm/GmcKxKA4Ojoa8tCoLmzad8VqrvSwWTh2XrVHfn/xKAiXYFqkoCssEkfMQ1
w4SgGwtWU2SQ60jLEG5Ax5IudrpmND5hYANlhCw+n01XoQzGxpw0iX34ZR4eiz1SCLYh9W8i9jZd
sKyvtmCdJ5C8yvUlAflhscyXNp/DRtssNzEcPzEPn5Nu5FdouTe/hKMkxZhc7PPgb1HaZVK8nqbT
X3RuIS1PrVhYECgu0rkmxUmiQVZ6blDh4gU8IPjCWIEVqkFBtlKPcu/1pmdJMLct2bOjQK+0Bb5s
9QyoQbdJfZo7/3wVVMxwzJcwyDMuUNT+EAlLycvstAW6R14X0P9XuvN7OjDaVIQCJSCDjPS7FtgP
MkY/xkB/bJnAskYWfG7YswO9PmsTfbQ+avweDTqlnkF/r3oeNl2FWw31vnQ5V2tpPZOT79/Ebxcv
EAr66BaVzklhFVuY2s91yIXRVNvwBEHLvGiucl/2FAEKs6y9vPpM/v3iX6cn6qQgFvVgdnX6HLde
n80T4SmZXJF//B5OAlQvdg5xas/wMlK7BcqCps1/moUwYddF4AYiQmr4kN9ve2gpah6ckqW2BHFK
XjWXXZdzx1T+6hJOk9O44suqQdP2DPEvBQ7SBcT2HrBLNMHoyvzLAq4n1NzhGBurb0F+2RifgKMD
naRL8l31c+rWe6sHwLahZkqVZ8TXPRX/Ir2PXsqrlA/cE7dugXqu86zim+Ggp0eRDgUVAfRmCNfo
oM0pg/kwfvdI+SSwg9f0e3Xcup8soFGI8nZTgC7IqMJqNuC1PduTSLrNZmPdi41hU6Bb+2xBKjhw
DuC0LGipHWJ4rOjERXm3j8WMVoAZCCw96jGM+aujWRD4UfcDkHH8pHc4K9/4JRtUal6sH1CbOz6S
+l0SzFxQBro7nU1AYJGb7aYTciq/0MMhxv4lcwhOq1l5QK83OfbU5D/EBBcfc6L9flzKuEg+3uZv
e3b+xaiA1XuLDBT6wA/muDsHyyadzdLTaX/Dalu5HMuh//zmxlyazTsf9LplrbMlYvSqy82nwz9X
lMI1+tsowLczWr+euiXv1vy9AHrABvvezDdDEMHP+p9kNZpycMSxUOnxIgpmfocrfMboTLRGxiDI
pjf7Pye35jY77jZCMEuI/ARkf1IM1WTdXSFll+00QOvTxIG14al3o273UuB5TXHfFeohyddilHNs
vVnVTunAqKTj2lij3aa2aZqeiPNDYPz4rB5kMHNFcS3WRetudHZgt8sQZNJzqs6MH43yxvKZ2QvH
+cT5nLt3ZzFwms02KWOih4rvYKciI8h6qJpsL4XVY0nR+tEArXAIrUgd5WxEUDIPRDEywSbwin3c
/YCPpz4ZoR8vFQ9A4YCRE9JWoXiK+unaXf1DysxXosuGWM/IPnEuT9QuoEuhQPDUbsYQD3RpE3an
AITO6p/g4WN4L/PXyW5gpmBHyK0fvmmCyQJavqGhrYyeHfWavNTGcg9G5O8DmdFP/lia2rxOMyRK
YFUdKuft6PcaBwlHT3i6RKPdH0sEcGn/5uhwWttMte343M37fcaNJJ6gaXHuf33n6tbfje567JUK
c7kkYvoTJEjxoN2kGn75aFXumH7SiWanQeZvfo66j3k97xNnyDPiKAQWttvvSQ+4CY7VT5QDiZf8
6GgNSIWsfiSgF7LoL6uO7vrG+YYJTvtyqy7FtMERFYBPGwxa7iKDMnA+9QD93fa+nxKybgckxUx8
XDU0P2iFcAX+9LOVUCTMs24QibH3A/2yCF8XSPY3uyM2nGCDupzZ2v1LnetS8mFWKXprVlq1qazG
VbRWdJ54snUOI9+5Ric7P+aoWDagGvs5pHtVkcF9pCkSweTG6WXLDInpsoKtKEnt1+571ZTfpClp
OF8FjxbP00WBCN9XnwwtuwwUbU9hR4pGnyVFmYyz/IbtnZ6Jq0tuRkPQlofcOZ5Ya3WYeU9G1K3l
JRp2eQ3aAy2PE4eFPhVzquKxdXidoZbmmZ94gBovbLk4zVm8iXZkchU0MBBBNoZBYiX7HyMpUa1O
Qi1q1U3Sj8eBj2VSrQsJ6u/wtBnPaANlEbrSSm08dwue7DbulsZCYgM/qRP47O6aSYdorKDYI2bl
yq53I4ipx4EZ79GUTblAI4b3iRsWXBUO3WQz5YpQhgAMrQLg5xnNBkvodZ7d8Gigm2AccIfqBbs+
HsENzGRzhcnp+alwITT1uRhrpdFf+67tJPjo7W4Gl7D5qB0+sJSv+9PdUKmb5P/jokoidq83mAdG
vMkQS+ROiqPF8DqwJBqiOfTtQmwOTAw5QeMiEkkS5dkRB/aYbblJZNoMEnFx0BnINX6OgCiS5uJz
6sh+x2G+1tjkZfJHfYGnOIEU67C6dQrhtbTZoI09fCtpmRbWOeCWB08NKBPkAUKPf+uxAuI0BaMg
+TKfdegI8Z2UeX7tI27W1qUqlMAVGOr9w0XklwTZUAgIoAMAHcZjwMjLF+8Y0uimCnFjGe9FgS1A
Jc8ZpOtnr6bjdgsK9siz9I5s87WUdkKczxqrcfUFtk51QPV351W/4ral62oGI4DLZcQW22wLTnfO
Y7VWxa9dW/O29a6YXzD0pU0ICm1jX4ZGw0ItDLiTcJUjboCFkv6iygf/pDeXgvqVC6BFN6qge9ZI
qiIOBhi9/JO2bSthh5Vna7lMsmQ5nTv0eKpZ4gYMehhhhCWk+kgDMA3DD/uFccNWeWrul5+xKP9Z
tu+eXMuQQpbdB4G/6IUr4TnNlwMxlduBhbPTjf9kJv7c3de+grQxGjN6SgVTjLoNtehlAF3zVmj6
af6IFW6K5ZhiQMU3Ob3frVV8iJirnrarrYd6XROIYPlWIhNcdLCMK+shRQ1Syio6TczSzkPNqgpc
XFSWceEYnkH+535fx/8GSauh6lOOBwDbutuwnMWGNwDOvkNtyS2G+sgMgZ7nZfcfVp3IsHTJD6Iy
6BYLpfaQkYzDqgp0hWBGt9suvqfWEp2l7qPiVcIeKgiW9e12NSoC9dnvvFoKsMmg+qzwZ/nPz3p6
/kgc5/VvyrHMbnfiPwpZY2Acscr0cqNBuwN+k2rSUPsnkZB0Eg9onSGeWrtVx5hulrf3cGt1piHg
oMhOOAY8I5UY39vNbkWGrWOVh0S2t76pEjhw3S8HRFd+zwzaIQyyN3Enh0+KhLwTdK8b7bZqyFjG
ey9Svq30Y5+hc8nvK7OW9ZevDi3zCoVuOmf2PAriquU/OSNVjhcQO9b0AnbnFmH+Q8tp9zEeXlJq
rzhKFC5j2X4Jta42bxXxr8LqoBrE6kzpkOScd+3V98mjNzTG7eid7FQUpWT28r4lEjgJ3/RgXLFi
F4nyTW+gtIW3E5JA39xffq2q4jeHtPAEvV/qHIcWI2qF9F5v9V2llC24LwNguRGsp+nFEDa1GIsI
1pz/ZzjMZ8JoV0KGEXk+CFuvJ3HA+uyaGtcHaoedPPVMx7LmvNUWkNQjwZdi1u+u3OvY+fJbOrF6
6P9AJHIlRV7XsIP6bRi/t5B6duYyToL2Mlu+RwrmVAEL+5OZK5l9yM79ph//EEGFJ59YNByuPnDy
gK1TaMcTmgFeW8Yc3Zr/GNQXZtQGGiONBLc3gP0t1vIVV8bq9ShMaBw/sTus05fPBgaI06gNyrLY
AIP3iEu2Vpui9900wgJjmF/aJQ5/3YY5QwhIjhyP6Py3Y96euQQJ0dVpF89s0IrVGnKaIT/ZBr4k
cqznVDoBVDZd4m4DrcEh54MuvASiPdKPDbdzCfpwzroP50U0AYVqWgHTbpgi6YAOAK5O0RX+9t0k
3f5bn3DiIhOcmb0HVy/MELpDZv8deI6QQBXqPWtCe3mRnrX7w981w9Gl7Z5Co8xCSIC7hJ8HFoHQ
4E43vkA+zB5r/JGjj0si9xk6xLvD+O6N16F7swJS0WCaTaZG3fMpip0aCdDTOMqOSdILmqBxzk8I
L29ovL7CbXx+VDu5v6PEn+okeYQ5DSjwMcvdD9UI9sEKLzx88q919GAw74EQ9wG+5yUKMp7uv/u5
mfLSldHgcXBQ7O3LkHIfQP4SSIKxPSF0r3qToOJdlOMrUIoLDw6GJJ3UhDe9h1VM4O0k81wJ21ws
/hLxwPUdCnD4RSls/ciDKQ3FxPiu4sP5Drrs8Hke3kCvV8HgV4b6ZpSuoWDsL3TClF6Y0zDQXJoF
jJeuyLYb0+/SMRMpqgk4m3O9GlMxMXLOMtBlnDjmUGp3QS58JJIRazHQvy0jCRk0EuBjUxIy7Vg7
qWp4bcY0KXdIhzbrEQwalipC1g7AS4vKV4abDSKMpm1NnO4cDXg4MmVCg+VZBGyEg3+nVR9aHFrD
OBPxahpnoJ1g/45uzCiKvlGDFzsWV3WWcJ8Z4Xi/xqvm01uJUYcVKbwZY1QTBf8rnJZDAqxjweBd
s5cQ9GQunN/RLSAeHP6p9PVJjmaFhH3cq2IuFl1LLVmSB210tZHzhIRPY92V1HVn/4NqVy1tMrBG
D3Mto3lNfO3mR1TW1qyMEUqf1dJ3Mr2HHwjufFX4P0PyUZCv2Qt3R5gQ5wntHEsmI9oF9vwM/gdv
CVThEywXofNZJya2bxfMCk5xt5IZNAkbDsYhgxTYMrY+sIZ12/loP/Wat6+qbuq7FwCh/jzDbm/N
W9AdgsX9qAH7Bgg0XFXbFbUXhncU5oWIoPAxWyrVBmh0rNeq63JzFshlIe/zd7D0890NITkHV8qT
U7OuK704rzaKMtgFN+9ZFS2esIPKY5XO4fnS0rd/Flj3LT6Snrwpz7/ced/P/qLvY2OTSD1IvJwH
URbMLyYBDD0VEsNlrWsCXi14O7kkWWnZ/J5Dd2zPoh/GqrXpdqhTmv8OLFexVDGM+xOewaLGjCim
5YdevmGi9OZfZL6T3zhPE+4/KEcbiPeeZms48p34enjYIbME9Xqmp5Ej3lHtibltKjghdCg1b53N
WnDsmbURCIw/SARs75GA/5kvKMrmGmOC01z3+x8mP3SbkfHspN1I7GDMRbmhoJxYB57ESRiTg4F/
n8IiEemTig07X+JWaPvukua8I2WhiNWtYQTOfbuif/mnGKLWmWcUnmsaI6KaWQU2TjF5USuuGcSi
E95qzrXCbsi4tlDVORfOUdF7zU0N8WGnf4W7x7ktwRTB8xhQmpvamo5+wMlmCPiFumYCxjxnKRxN
z8pKKGe8tnGwVctkYZI65Qiw8sJX5jjlRv8oWxjSVmX3APZlfLyWx5JLCRIoomS9dHdtU8irE4do
75pwW6UrYOAjL89DLSvyDGko2I8X+NN20lgqEgkWr4LVo2VZASNFR17C5POn4JSTriEjaeixbuho
wG3a6lIOfKWbwrkpt8snClWf0VH3tIk7j9xMhBom3p6OmxLq6C0M6T2/lswG1O0itW8D/lonLcIW
1mGhlZYoJ9mVWQrFPT+Gl0XH8yrfJqhUtV+IZmHEVdiOgiDO9WVSEyMv2hSiUWOgGZZKnqqHYtU3
NfCtLmV6DdGtqf713feat/W7puCetk5prbV8tIoKkNKs+vwQOOf0qjj0esfjUymBy38oGrx6cWoV
Z+10cJDQ3KwM4DBiZmrK1z31b09xhqJroKrY2EXmmvEnJvacbkNnDeWlo8L5zQWeAVKs/nl0qtWb
GRQ7cHIyGiFj81FADorrTPaNgsjSLsJwGKWZ4DR82iPsB5zgD5hNU3Qsch1MGTZf9mWKWz0UkNab
y/kDpBLreh65T15I8WBBYfFi08OtBOqXvRb9ChQJtvh+Phx2LKMeKTuRwifgwiJSPR2Hm+enybDK
NP1cmDSUQD1kRXiMYunKtBHgHNgyHUc1USydzvygHzv2gpzvnzLVuji8bnKM13x9OOO5441B8oGt
PWjvpKozNDorIWB2rPFR5js042lx32P51PTJUJ2Jn7cLTbtgQ+2WD6NQwwaU0ysg74vFsaxOx28C
Vn6SnCN0bSZx92YW1P6zOZFQbvs3WugDQltVq/y2kzWyf+cF/c4KBHZR2AHeRpG/m1t/wj+9U6Zn
yMFa2V7HuFsJREKM6/VKJOqPEXBF601HRUk9yyCjBt6XBwQ476OKQ6W5ZkUIV0Vdds4mOvMY0bc1
tOeUkz8OOVcVdNFVP21eZTq5qrq6u+cZYPVLT/HsmbF3OewDwQhliXIWz2y5SY4eBAEHnbnYGGcL
GbqVcwXVLPnD5Fj4IBMo/PO2zMZH6XEZh08R8dJNTjAbTIt1e2//2EZH32BrNNC89MA5YYyDh8qU
8TF9p5HogxdfB2mD/2OJ5PfEPxeo86gAQ0etHHWKHbvLpB4MPU7soHZZJ+ZmlI2ByeJScO5SMjT+
x04UecPUDjLtAuejLWjF6/loQL27SGuWMoDl2Bl8eETTwft6MJpbvdVJulFGivYd1IlN0q6yqt/7
HzNxETU+siCK7Spp+75OfmtjWJ/GOEoxZ00zZATjOWaLNvTeGTnwQFYW9i/v/esjbbAhdXVMYuvV
EsHHuMfzoIMrNlTBN7KQpVwTkl+O79A0Nj8FvrTI14Tdzo6KM2rT6oao2cuscloYiUQk/nIydJmD
6jjF61vofKi6PhcEzvqLQudIh3O4A8s8alk1UJeVTXM5Xq2ZULraLLJYl4WWtxc2JEQJZ3YnkMGF
d2wCzzavX7OXunn/9vYZ8+CmTPKwfHxBX6blzxS8N9UEdaGcA5f8pb+FV4BxgYQdijynhRkTx4V+
PczY8ZC0ZQW4g9cO9xTzJRZ8JIoQEoM91iOSelfqOLzqn5U/Lb+1E2yPM6RBPDJA0KS7UgHXHzVo
6aeE36ewcHoJBe966yy4Nxn73XnUHiy0src+EtC+ZDhavj/wsjqg4yObAx04JsfisyAu+ffCNwio
t65NgArUW0oy+3SX+ez7EGC9mM7XMxQeK8NqXYvgBn+kqx+FW76uD9CyVN4Up85g8V/ifhJQ6nSF
X0GiYM0zoQtjs6vfQ9rw+6IqkUT2DBoSGF1tsf8pfeLl3T9lAb2j50IgCQWe5/sug54Xi7xvpfoe
qSkMW8bvcNxqMxkLiNP6cGgTxo1WfH8Ceybhy4CmbbUpSvoLQcKyT7DbdA0bWGiEXLAvZaAgutb6
bCJc3sdjBOkOnPnYxaWdJQ0r/iTRL7rtP+NzmzQhQJszFr4bHPvBfCwWY4dG525OgT+Vj/Pfn6/o
3+Rcd/S56XVNV/SvRiZo2iDPRAvXpbrbREVybYBVIVRc3PYDU5Eqoo5/4fMZRCc9mvoPblh8rlX0
5nKq1aVpq0rx6Vl7v2sYGhssQmub4JwovGpTuDBEjth+kG5ED+d0ZPii8zrDmmPI7R5SKKZydTdU
XEhqC5MmAFIszZ2MHMgVYzznSDO+d03Mow675rSNGs0x/dGS/atGEfnsmwTIQsFsJ83WjlAkxlLz
/+MHAnen4V6OvryUrnfrQx5HuBOn+VpCDfBYcC4wZRgoLlRJHPm5ZqGgygpDulFwmu6nzKheOXNL
70iYXeeYpSlinvqAAQqpRI5zhLhIY4CQixS9aZsXUZkYh9zAwhvqhO6nEKFNJTQZQs+SPU3w6n3I
byrrtmgQKLypJYFydWTE2gyREYk86Q4IkncKl8YT3VUfDSJmdTJ6ifNd1PBIo8KeCVNmHXqk4IUp
oVHClqIHR89TgKDFBPiJNGYAH18SS1dOzjFIARlXGiAmODKjNMKITrvizl73bkV0vNunkasKhrmQ
wTh+TLEdPzEnIz4YG84lBY2EFNCQZEpcnar36LoF92IPQM0gcONI/z3IrAKc00bU34YbPYv82Ts9
ceMAqy6lcTzl9S2AA4uobYyYDIgt5iqWKdXw8aADz4EEa+9vIlrpEiwudgi2v56VSCWPbLJNtGu1
Kr6LqgNl5rXfGbhAg8rmgLIxT3b4EEh0s0Vxaz9gpr6THk84ctacczPGi9suu/6LGO1dooVyL1kE
JBVMfeuG9oM2hGIj7OEhWehptLH5/Kz212xZnOyUXJAqHtfSTC7qLZKt7+dL/VUM4n+p3sCZEX+I
eVeg3D3D9vXY8V2TDaFm8GFHVMiUvvJVcq39YCJ4NZjnmp11/K4FsXqLWtJsh/pWT+DwbAEdPfIr
M7cXfR5Py/RXVwZSaEAIHLZ1gVTeHxGyg8gMPDJqXhQPW6t7lpU6jFng92zV7kANmRrZZFm5EV7Q
wHiIJF8y0XQ31yCfs2ksyH5BE+d3ihblkttMC3tTTXm/PV3xfzhOjRVdeETzodjJfFJccQnfsxsZ
MnRAzbkaaWHI1SLDKBh8m3BN4p5NM4w0TGMoqTDfQmx5m+lgF8btpR459ZTkUJJIuJiuy0Pyxb4g
xbMh7AWxIB02lqmu/qJcKoE3uXMvTvPaUhmyBIZyA4yJajtiNUJaE7x9CAlf2yjzAf7prnsqBGuf
VAF3mlgHUFCtgX2pXtMGiFX2RLhDYrSJsaxoqL/NfkY+UV2ELxp/zm5U9OSVGmDnWGOZTKNW9UFH
Qjt5wf6A7E+7Vpvqv6izN8kQ3Z5G5lggmDMy0HiENIcsu8weyDLdv01xttYWXtcXp6zH77/uD+jR
AyreZcj6opZM/sdzSK7MCNM7dlPiiZORD3qXhJ3yC1KVWtx0ZXpP1edBQ0XWKh9FDhCtEDuPkl2/
aTh4qJve0i2th6C9GwV4/I2+wHD/LxbjLdjokzHp4Ji4oKvL25bsOvhiadfy90vaZ5AiiHrszKIm
cMScs/zWRlp8lwOj7r+ppFZqD2bdNS48Pp42Psr+kIwu4yJ4o+OoKjZImcY4WeBJ+KrTE8dQ0G6G
PPmbyDPa2Q59X19DtZcwV7J8iXgS5VAsUUHmepHR8sLIZRa1qazZFEQJFGTj/xkxourMBnJloXxs
kRGdUAvzJQEK1tqgEzfxqmabzXx1l6Jw+cSRII9NNMTXEsDKaPMM9hP+13+bXpt2a2MsLIYr2mmF
mn7vC6vU7JXLRJr27lJKh7XJkmg8B3ZoTHD2x4y5zLOaVf9ENv/qwF5raqm0o98AmijQpldhxTtj
PRsxOqdHSuxhguhKaGiTr6pP7L3lmrO6BC5KyzAWNuyuIXUdT7tcZLIKvbK9UdjizEKYxiLejRiN
S8t3UnYxZjkxst9puO1HzlTEvNQLWplV4g2ZzhvBLYORTorbwfAjSfDX1F1D3+IPfp7yv791962Q
SXDVbOGK9F3jYHZWzEUEjIpeeKg6iAXi3WYTSsAqoUq0Xp9V6a8bKlJhIHeyPxeyHtQ87Bwnr0DG
4373Hk0punN0DCZ+jpxw+7gcxjjtjdS7ixvg4HkF7OJG1TZt7ui5oJH0/8iWCnrLUgmtRUBkwQf/
vDx4q+byR7UP4azGLhjr3NgKRaSAQAI9QtYbqr8nzgpksNnkbYxa5RodJX2cgHZ4C6LnYno1C2Y3
+t/gKN3Dlwfu5ekOj6aTVGnbX5KHxdmsZj18pcvk82zkgRKD9gSDejvoBLFtyzASRns8nqIhZXZ8
sOTvyoaiOo7QR4QU2/KnDXZc87EgMOPg0/5NryzpWcn8BWVdD6UZ6Z8TCzhYA0WDtTXfhKBGebUL
EhOQx6FKuC+Tcs+CnlldYn0QK5VQgb24Ljkkdl5lxYMSlJnW/Zye0Y2eMWhmBlJu2pkgYlObiQlh
vKIVVPsyucIsA5J3ByCrBtpU5SrFArsMbR15G9uDagt1hJhcquzq2IguI7Se62E8VZSSybJ/h6ch
gGo0VQkqmyOTbV5jye7221jIUFkPrBW5hkf9v33HL+ZJU27eusKD/DnB/UFuRy/otJ5qN+xQSQsg
i/Pj7Lfg1oDuEPp7ObVFlrjnUM7Gvcd5iopEvFYef2oStrTC1iN8p/vmjyzgQ4NgFPRUp4Jqz9sh
xyx83ddAPpu0GozH6j7y1RRhB3dyDYZZ0Iyc6IydYA3OIWLUsmzHOBLJ8HNRJPh63YYFRYz3hIVy
FVLWwZNcpULt5M8bcE6oV0AjHPC/ZfZ81ttFtnnFy1Fj2GNq78dIzFn9niU4lq9UYeewmkXwazz6
C1fxPq71Fhy7QvQUXSXDHo/Xo2bgh0PsMbYIQhZ5V8SkSpGU+cJgX9n4z25IlnU6nNeTli0ULwHf
wIzWj47p6Uheb+qhsWDq2jV9XiLyzQtAqZSvzmcvgh9YfWMzqzQ3ZTi/VvYzSj9Xw+i94YLMNaHB
itx66aiYzCfL7NbhFLK6GXbfHPXEbFJmyrNHf5reYCXEX6XZAYh64dKXmaAhCQkbGZSuYXVHWD2i
5EehlzLjFiU5YJ/HE6etYS8AztJW2GBczTd672TZTM+6DpUf8btG2i1SXfX3rI2pHJMcMKPwOwtE
dAfJAFpprysi2x5jfdxHiWydPcKgax5eHLaaboen9pRpjmNzdH0Mcm8YMu8LubPOd1q/Rd2GlD2v
kLsz1GnJtbNFx3d3vkO6ZoLV8T6W2dW+AUaNrd/KrfNK3pBLcyd9XLDHC3Y2EnK0tCH6Feb/NgJ0
THPBUs2SCAbkpunA3kPTNzIqPoe3bTgIc/QLSScdaI/GuYMSsret2Q1dpnBlT8N33VOnG37Iz+0b
7oNEZojfXSpvYK7d4My/uOOVen4tEjakdT/65uBL8V4a7oAuSMXfgq6uvGyBAhyMxpBryxYk6Sbs
umoPQUX1vJ4ddbaG+y/gIqnjcyvJDLuRRO3DFdHBERYrv7dyQJNmi7TtQRrbJMuw6p9XHBsaXyTW
5HtLk9cdLkOxFe6mYjcoiApnvwJwdJ7/6NSakDsiNp4iAcdZrm1bbg/NB52Jhc4QOGo6FfHMCTmq
sjipBMc0sjhidXVVbYjoQcXx3QUX1m5ZAZWdsNEvoGfuYc7iWeqZqECzHDO9JlXq1yZNOVimVjzV
TykNAfCW24kdUmTsKgoIwcGojoWMV/P5BORgI/7hrLFyZAvcLX6iLC6Q+lsL5aEKCDGIDmufcPdJ
Id134oGtQNt1oVoDFFK+E9rbxleR0wsRQMkMSM8aoG4Yb3wj8JuamRgHpTWjJZbXloKHJgfGP718
5t6bnBc0dAxz+aV7P7m6FjBogaUIkRxVM+xq/pYn833aHk+UOsGTcJBf9B0h5AFtmsE/830oVuoQ
hFf059jwRDMIBct4OUhLe2XKederxrMQOeXo3L+yzE9umM9Bzp4NEDaiN7DEnH/PGZaLWA4m8G+d
Q5PVEkZR3ReqVuwoT71VbvsRHVDfeRtwykhsBWn11ZEV0Ui5i0b3lYGFuZKH+2NaapHxrizHmNDC
U85jNy7lllZmVEdykszoj3opEW7R3qb4Ii2v9gsd6GNaNRCGPr71TzY3egwUW3GqpN79yKC6cd9U
ZAURafViLlMAXx4v368XnBRr/w81vwT19VlfLnrmk/JQA13CT5vrp/+ymZzNgBxol3zLnYQo4wad
jd+UG3N07EdrZLeqAmBjeEA+fbfTTS42QnnZ4c/hKpEiLcqKDr6OizswT0owu97tP7riHW1MYL2t
KirakHyqRfmii0eYW2jiCZ99IwhH3wJRhnLJNefeUMgUHFEKjPSunm3fB/rtg41azpTjwI6oBovE
fJ5dEL2U/H6/5XAwVLJZ4/LEi5NBJE7V7HtYYRXSkYy4bhbZtPf+Xeybomw+7iw1SDXV937bp/iE
U7/zzHIQWddSLbPv/Ql5n30JUK0yUH5PRfV44om9YdeTXSDDEF01z4v4v8IZsEl+a8h/2SLjHE/R
x4D6wDjhPGQN8iupXq6GrLcH06VXD2iNVDunq4Zam1JcjJqUyM+yaVG7DZwsaN6kvlYkg1YpuH3R
jGHB6c6+WhSG80rcWxlI4kw5hrFVs/MV6rohlP+mWKMPJLll+Z1/Ys0Onl9eiVhqCyhXmveEg8VT
xaT68JuPMmM3XlaEyyEco3MTLunG91kcinfZe466IBN14+QUYXUuKBrMi+HEyayQyFwxXmSP7m/H
uGxPy34xihbDlWX4thdXGd5t2iLLXDeMXgfBUsqS7423ojrUbcSdyYCbV+mhi+Pns1Fhrj+8npoV
ZUuC1ml6oJHIyByU9F4oVo/SGZK78G2nStVMTmfqC/anLkt7b6SUU/0vdDkAwQoIz9U6FZi1Fpel
qDK8++jXhxKhJOU6ICEp9aqqKvY4dOC76z/tsQzpoyoFIhn5S26zvB4rzw2EqwJwNkhf2VproFlq
sRoZr0HKaLNMDDISVTuUJZR16CzMqOekRwmhBx3o7SCr4ti9shzQ9Lp4xLgaZ7YPn6uZncVguz+Z
PEjwzvKKlexQd9kOZqqTAr5eSryPhbhFJAW5qZute16yVvvcWPcjgPXa+Nr7jKARJa62ALSOppU2
EUmbqm0DMcYocGL3xA+/wZK3KmAyc1KKc+UdQ+wtcxU8IJol81fWSK6QFQ4pCdlGMBo+LhMXZV59
/ku8iPmoT9aC7Eiv4DBqnR/rodkV4l/3T4UUpnQdu0VnCo2TNu7z6e/JHgOaJfKkOGs9gFhYjlEw
R7WeH8Ws/tcnd3fQ1YNxpQq/RfmyZMFfvgELfp4DW28WkGRsa9JD8b+T1gZtUuSsj2QZ+vsSqO+d
936jdqMeWPt1xIRjXfCAKCMeBXq/lEY9XX+pUMVZxVojMpBjDMlB41V2CF0CorWeqWzAcoPcqH86
5mFVFog/O/2yqHcRSMcQIoDTYkV8+gZYsKV+d2SmUOJl7N1CRk8S93eHfLO6yQ3esrYMCU4ErHO8
TrRn9Tox/dZk4GIxS6AAqf2kRXvjdEX8RKq+fOOuJTyRXn0uqbzLeNgxa4KVkunppLegn48Ki3e7
/7nxW+UMmnTGB06PPELSkuczkUAALyiyheUWw/hCFjqH62cMD0wO7pyjhtj+EP6C1PbHxzsFfgBy
eXlsvCHLXrzKEOCBEzQ9iyMMT7jqCYTb9MwYcwTfgA7Zu8iTSBQMSyovXfdycJv9VmfKm5GxMdNi
bI7qYRoy9Sl3c8P5t7aEtSZuxDHCOB1MYhuThkIaex1f2mZd/1mJtVgmMrfC1tzgUqjVQDoCXelg
fpn79DWeVWeUWswHT2jUd8NhvBCFsNG32lMUOmvq4eVkc0uwFWHWfiCg9kd4B3xgl6a2LPBtio+K
3JW8C4ZzoKRfPk3XdwK9F5DpwZkN8Zzgg/sdg/WtA8qNcQ9K3R+7U7qi9kBrMeL56hRw+2S+Fkx7
Rl6IDsovBFDKUffgCqtS/BHgrgoqIekz7dnWLXX+rA/flWko7OW2+p88Pn1CD27c73ahawj5AfMW
4/flYfeaEQL4pY5TwL4donnTmW0hVwEEa3Kvi5ZsUEAQc9xX2ELBZN0CJwbfE6CnlUsHllt7iVPZ
c+QEMIk296vpJJ18YNRxX0d4RFq5kIlfzIZ3E00XyjE8+7FxXEklRVpG1PqXCkE6QnPa97DVfJja
LqoQvu6LpK2YABANJFVdp6bg0h4Z360TC07Fn/bWH8y6NrL7N+8d9vaGy0LRxNC0qZ7ATd6HjKMi
PIZFDRqTQXQjzJriFgArEqo+kGIv2g8yazMMFKP9Gc3m1JJK9haUC/suka5Fik2QDCQdLIx3+13o
mRJK99Szc7uMPv/WHIODpCtlsOBF8Gk0cEK8cQkdIJ8Rup8BOGYRy8hlA+kTeKevT95zSOWDjsT6
nz0cXoNj00C+OND1jseh4mksFiGxZ81wzZENtrBvki3c4CvC7zzxu+A41wRgx5BPmQwRCF74QCsP
xmCxiN9tlojd6MCMK8g/tvZJsB/LiXTFlsN9oMKJN2rgccquepGNfK07BQK/GUUUj4KKM80J4XJz
wqCpfrpJssm8HZIyQwBriC0jNAwA3iU6Uxsu2F5opwsW9Xm2wRr+PO5cYBqweIKpCW6Z44+bWYG8
cOPQ060OWXPHFYUa8ZTdYijgIKXf40okc134mjQtaBQlBFM3IofwjrFhErJ3SnpErWuIFFsOBOtI
6TBNbNDDver9StyXbpcVPLkB4M5r8mJcyyzitdbfIVdbYSWHtzCqOEzbpJ++isWFN36DLb1HCxhF
WgNK6dVFkLwx9tKhxQDgz0gqFXwwOmou3ryqxzdFpcUfiWaGWkpJI1lOlM3hGJFiEbgUy9uKLWQp
IjYfBkh/SegLJcTlhRk+3U8TKDhTpi7aKNDz370Seteqv0MmTmkOauLpNJCMV6AvGJYrHNLvHZdM
yqKjBWV5yWDBDzwcoPYbsvyksa97UjiUJoGKxQ6GP1PriIpoKlYlWeZ1N0HkgqrZ2rADzhwpl8mp
cq87Vya7yh6bXQLwHSGXtZZnTTkXEuoAlelj5kTMckYkKkHthdNMNAMriF4C+K+xTDejBqCxQWOc
01UhJuNzslpMgQntzIujDxsJRHIcaIodCExPQ4LQO80hc2iaNzcNQZYJm3iksBHy3+idZS+qKPMr
c5CAIdovAXreeIMSM7n7zcvE9zguNKVr5kWCIzO2v04LU62LXGkXp+8duHpEpVl/nOdAhO0Ik5n4
RHL6UxVL6tKg+f3j8aISX/hXbp0+SV6PwfZQQDcuG/XIZuio7pv+oQTzaSVURGOgzA6IXNZTCYAB
m3sjQXAPWMvAR/bNjR6uqSKzdSSgqXxnyubbQ7xEn2o48SqyPVuM4VA7iEiqP0VJ0ZFe8HqZZ4D+
oxMJ1bJ0eZCsAH/BgAwpKNmWqWBZlO5A9c4vchah3VltLGQGlzaBOM5xOXdPaulhrs7cHgjKELBt
rihXGxxtqO6t2gRf76dYW8gkEykfZt48Au3GIrTUxYkC6Bf/f9NgX0G/C6c2prIryVDnmDHckoP/
45VEGp1dDPf5XenQ2CRWEZ32aTsU+oiLzCRQHdEMyBP/d0/1SQsnskE4DYZyKc149z7UlCvxaUfs
Vf/h3rxAkOHyDvNi+V+xSTBUJy10HkbMIbGatwnn+10njlvOM3U+rl1JRhqiqGeS2Q4tlu1XqJq9
q5bDFyoOq5S3be8yUJa/zuw5fMom8StKxbNyRUEK/Yx80eoFmgHRY/RTUEFqUb1/t+kVFd6dogyd
h/Atu/U8Gb0ILs35hUr017IyAgrQaQ/zdzr7EcZ1GmYlE/8Kcy/px3jvYmDByIBmzJFsOvEDihOn
gZMC+8q+cONApA5HKogu6hc+6T7J3ur2d0Aw6kWpS9gr1qFTvSdIbKdPvEYUJzvXc570XiLb+MC3
xzIIqRAqUMFhxGkZmp6IvbB1IKJrvz2ZCnV3S7P7OPtYfT47S4NOuZVq2QnOQEkn7MKXf9mGoTzU
tcNnCANPwrQvNz6nVtm789/J1aWKTCVl8BTMNzQWgZhBmZ/ZpNK3cyZU0RY3hMCgqqgA/YrL0p9Q
kZ7/VZgi2/CAcUqVTUkNlTntHN6YNuUsdnPTidMI/dCg6mHyH3dIKlyM8MJlUgXkHYmLfOrHTRUp
8J5oySuD4wve0AkJsSFX1SGknw3swB9zBt90ZSTNDb7TkOgjzpfwVfIev16v2iJtP6Xi0qb1H0zL
dFFm6urNwD+nOsMd5YsmJPBNEY1ctNfNy0E+O6gDD7dMOZfQqz7gaqmdY4pehzq0yZ+DfFS1bs7C
0+FlTaTbPlbe6WEQArdIRl8uhSb0KkCVLpoop/pULXvNMq9SKlHUPnkY5fP0A8banOnnDB9uu3Wd
s1xQWnf5ydr/a+nHDZkQIN/8jU07pgjFJS6z+iQZl09pekH8E61t1loXuzO9H7Zcx2UofyqUVofg
to8TopAHNsqby/9eHXCZYmATk3jyuFyh2ucL+vTrrQIofxuidtbawGCkT1V0cv9GbocTFWv3uRvX
PuokQNwhYwALCMf/bLi0jStac/DwxSXXNazijAU5cqLvC2IXUIih1+y2vo8oiOi/6FNgBCLkXFKZ
OY9PTPxnQIuwn63RZaEn/8NtBMrzOMiUgAjcYiYT9NSjA8+qemVmdwDp6znjMayPvvoLGn8riWlx
56RO6T55kjLfNNlDgq7r5aaPOzHhdhQTFq1nVOTP8W7mTxosLAAhUoiAK1JxI94Qm19DAKPe05aS
PxwvD254UZvvrqCNg4MluiqNF7zDjyHrUhax4Lzdp7AJZv0S5JNGpi/HwOU4UlQrb2UnMqLssMGs
ddNIsWGBs8oGFImd6BgKw5X1JokTu81z70UrvuK338aX4xt0PqfqF8DUtau3qz9r5vTGglXEJruw
KCLM48IXdhUo5iTNpA5nYurw9iuF7KoMAXzWs0E+8zustge4E3ZDqRoeZRAorAK6o8z/D1Y0j/0P
t0OCj0HmkWI7QXhgahbCZihIG2RMXfim9njhGPn31Q/CgdZuhEkKolyBt6ggOtXSY8XAM/GhOdK8
xKqNxIQjqdwK4mQAcDrtrewVI2/Ap5dHpqkwUlyzVpbHqy2/JU113FbOhrjzAJjwRXxqIkbJsfVu
cFXWchXcaHs0zo4MQjAO/4PBnVVid/U3h7sM6NiRX3AbaSRYqqMIS2+3RPVvWwZGzBCV5tOeanSg
Hd65L7P/hgihrC+SgjmqxzIljbS+ZAZ4W6L/4btcHL6P3II55ICSKDZLk88k3YYqIJvwkN4vwI5T
rNT+TBR7C8kETXXS1KjDvyKF0w7Ov1eDUAT4KQxkyb9shgmEiiu/cYqsClVB6HJBs9hf1uLWZg58
Sqwad05qQwiGgpdRTmS4iLMM00sk6M40VdT7qODbGBt2nX/pve5dS/2E6AwyiVQlQ5Y6pvwSgeCM
e/i+3OUMVlNKtEV0MNw7tkLAZYUla3goAjtKoViYrClfKIVr0kmHh0u5YvCTQCKsS/5x2ZiWIxEx
ffWnvvFmrNTdmLk+3fae2zS1PDSSsr0CmMYVKezCvEncTCzIaCBVMbfcfATAuthlnXnpxHggP6Sn
8/w6E3G/9Mv6fy96C14gVEcun7KbsWX+csaIHabkTS22v19cLBkxoCQFg2dGwCH/6nnrEw82rEb8
rDjrHjEu9fzppDPiFOYnizjBgEzl6Wy6+7AH3SrFSh7betipl1deks4TZc2guKA/w0ThlWkApdYb
OKz74sim7Jii1Jpn1XYc3ArxpeVFxX4l8sNfG/NDWYcYTPZ4KKb2e2MysjQWV/gMxJXkwWN+vDlH
0Cfda8LMXBiMJAQ0NnrMymVVrL0Yr94AvtQ+YtUvN0PWjkvAVlZV8EB4wu5cphfyiioRSQJbLqdF
mYN8EYF93f508C7blluWoTYXVIR7YhL45fnvZA9yOdppcuN2bpOPtHL+jhvMD6trL1Fp6LNsh+3p
bVW4973kEdRIm7djt0MlwtXBsDLB4dp6/8Oh9/qHIpQ2yr22ceUR5OgXIR+zM4rE9doTTmS7MJiJ
MN69LaUZeWz7V/jG7w9guw9klL50gLOqxJEf2EtoEQ6u/X0/VRWmZzGxii1yXDXMYaoKrPG+QfGG
I9H0XAfHX+J+3mbKZFJqcQBgZJNIt73Yj5sCfLsEhwjDqr99Ck+LDvVcNmhQPXRcgN9vGYqI66Uv
cferY5pEsFl4tXpgI4DeW5Cns5kXMjY0XTbPFBdnVOKrqWpoOM9krAWK8OELm72wL+2D/YrZBH+Z
LLNzD53p5RydbkGW2WW48LnYwLUyae+IzrA9o69uzsSIwZFMzji/rx9QYzvoVZTGitd33nXgnzQn
Yeh/KmhRHxjdz5qfvXuZTVBtuyfVb4w1D77F4F2vXPxp0dj/xXyTasnL3GsQiVxkrkvyfJ8nIm3u
PPJpbdE+9V7DFCPZWfvK96ut+9JvU6stpeplbPTVRYqdUf+P89EvDtWBdFnJsDC0E+knYDOTtkaH
GJByfRITWOvWAOIM7CZ2SuuE+jT12b+lo8jF0V25HckiTcUlRcjPHCmrWf8ItAQu7s3WkxgMrG4m
yy4uOsP3QHTl0VMjPv0dsGanzeWVuMzFX4QUouID4AZn+rX7K6fkuJcvrxVXkzzNiDkrR6STOpWx
LlMDMMl8zm4Xdz4+mNRnJ7a+k3t5P3AsosOWg2z8MI+vpGZYHkexoHseWybW3u0zUElvDoVzxr1M
wpTwMAiZfWVKwe4+tFLcK5IzQb1lmcHYN3arxmS3OgYsfVuHs+/z92lIeIQYmGGaVC4pj6HAUory
bCyK8ceXkwMij3kAWoADhnhqI86jmX12xVUuRSrjeGhdBgqiw/2JNqDPOz6nr6UqxGnNS7jFB+ut
1nXO5iXC48GJU4cFQyUatyN3vyHQMwjAzuz//N6jzLK2AqkmOyIxBXqZzTH/OPrkkP5R+1OjG8dO
fuH2rk0v2jc+jl/4tALt92Ja9rMl1FBePexO0QKmEDaS2KH3mN69Hg6E3dPdcPjxZgW3swiWs+7J
wPuFT3kYbJGCKVNmsYA2jgQFdj5JS9uhHDCk2pD7LoZjRcYr9EZd//Ns7P2ncpcdsOlEf681xxFs
Jay/cMuj0hRvj54EOpMgfFphW3NCcpyQ9b2H3C+MPvMnN7nk7laXNoskcmroyQyyS5f3c2ezjXwj
4aT6VQ7MGuSbfGsAl9m/WHKDxnVUXp95Tzkv/8sAoqK3QPLtNW5hZsWdjIhnKuwTuwp7eo7acE8P
igmv8WB+YQmOiHMVncbOjUCg18ubouYzAJ5ORmWFeIrs4dWeJcorty7EmUDMZdOKfWbdxVFpenj6
b70bmWvnepVDopsk7PqU1D6YwF+ej1ktJprSd8TPGN8gWJcjsUc12OEXf5pfztjWyBI40DWkKhfi
qo/LKxqbef713nhx+Lr4JHlqCHFGfnkptVHSNXkY2M6zX6NWHzJQy7rl/2yL60IZLmuHwBj1uPi1
XJAHyJsc8FwTJaUbX/T/ztwFsCimPAeBMJe+AMRkNYz9CxZmaydPevpGOAuWklgl0cF/Eao8ID2w
RuSqv6l6g/Mg6xBe4hyneR/ez63tLTmWdLTQ+QSJ2f1w1a+l8O7A35dUNdtGCnFkkVbj198rj8xI
hcTnLYnB6uEFww5a7x5bX0TbYZMWqw8gCJL2WjoQlklxo8VRz18v0CnQ0jDLgYjppKVrV27GcVjr
/RVV5QPtIrayyoA5xaf81Vna6j6MXaQcYus9rNCwkWrrzC4G5FbgCxmdaFoxVXtqPhESjoyikO4G
dN8PlVQzxz7Tq4UxHmvlcPAPGsztLUt4y3XvD8HLVUv5KKFakvEwKJObwmaSl/rcGeAXAUSy7mQN
qZ5SWH+Xh7cBRx7Xhx+AcM1u8IZhi7jHtwafEeKIMgO+n2dN+eiZh9VI6KvPQihnWTW6wFfsA9oP
JMQrdYNh+XxPFrHf60a6RWDvjwJbn8uWhpaFa8O2bvm1HzmjvwqcsWYq76yAvY4gwpD5dNu62HBZ
dJ4A8OfqKSoxjT5kwx6G76JMtkH/0/wWY8iPS4HKXPKkJ+p88Vcry6yESGvCu5m8pKSuSPAoGJn+
m/p1aK5+FpWxR8rbBFONBwf+5LWPDOdN7P5TDQj4gFQC65cZuCoy+PAsQNErnOsSu4TXevzbQ8jI
/qtlKVT3w5XnEFIRe/5VWTFPHX0FQvTtDKu+KpJfCwRzTBVTHKiybTb3jT1O97Ny0eChMtYmqaSj
dzmB9xv3GLvTX64RjsILxMXJyIodEKhukMb9Kp15og97ms335iLt692Y7H9JYMw6Rhf2Q+U+y14E
r+mM47KIFzp4qhwrT+/OyhExE2Up29aqLCMjtyuAixfabBP5gmi7jPIeY7bygr4uCtRjZ+9cxmqM
a7oJQtFixhhz/0ZGsOpg5JEVLNlmXSRrbc9k/6CugRxRVJfgZDrMQNKAopJr17iZNWgJM7eFgkXi
hagoCYaaQ3nVIjhJD9dUzATj8DG5qmRb+0rrItAdqdBE5Q0tVqwJUqZt4bOP5GexGsUbQDZ4SPyu
W1bKZZ67xewEsnorfY8TjoZ4QcSaAiPDXqwDYMsSkTwy+N5RFz7M6UAY27PLA2lPltZimk0r0LfD
sRqj7UHmNXE+wXRLt4QDCzWIGzD4khKkGuCuVVzabgrSkGp5qo+/jJOAlo2Y1lQmydpooX/8IPzb
hlqJIdVZ7dWfZosOOrOqz2FNp/VvNgUmRMjpBXufnERBWE/uPCu76TE+rfZejdUPakMCaeWjVCkE
g4sDuAPdRgiH2vz3r7ZxTaQrrznpQv47te+XBTJH0F0Ug7I7R6s1q1vy1CHNTLxoLiy3GF4+Cy4P
lOsrG2TSkr1fWuo1WO2EF1gaV1Q64+k1aDRtLe88pBVNg/Xtvzu9wFlcaS8j1/B6CvWBHFDPo+8c
Z3MtI2VV4zGYOUR0XDSLLzmxImWXmPAk+uIonTvfhjMorYBPxUq8N9aP1hXiS/59TzLccUJtfsHX
ImvkjBmSIyUg0x/qE3w738k4mrdo79Ve0FyB/Fdc+BNKRoyhRbwD7s+aLQUQAvIyN61onfz2B+XI
gVT21eTfGso2qBUb6J6M6E2NxHB/OCe4X9o55RMMauvw4zDZNPvEJeZ2cWL7AzijMuClAFTg3IPl
OrzjUKLBeLGi9iHEIb4Zg1lmqeT2oxmZXOqoyMTGrxWPMhZBrihjA/dU52Yedri2WfEzCxpIrzNO
SSkrmNj09Sm9PaqA00H69l8NXYCptQ+iGNI44KNLZTWMiDonAKLC7qyolQCEqb1Ecp45pRLs3RFC
TnTKLjcTJRIJuUwo1J2dPcDfTV23hDrIANt6pCXo5bWnTFjsyZ1U8baEsPkWsXQWhtEL35cFmdcR
N9iajjI5Teg67911j+BnCM9xdDtq4FFhVu+ZE/rH4gDdDqODy0u8aNitBZx/ZTuaQzkwQUEQIwfM
7AKnI0+TFhxLNB9oGdWsiIpvWJvJVdpJ0y1/9m1rFFsBq0E2Wc+PwMyIRyA77Nx9iE6ioXeiVC5/
dzmgFEbbedNfGRLGA4S+491GBppYU88Xnv4IdSiCCrZWlwsWgQAbNKW6BZaAeyyIfLHcAP2gA5Xl
O3EFsHIo8hFXSJQEj2+puNRv8CdEhYimipZvUBFDfKxqm7VHYdxjdhZJrQoXpeRLDd5Sm0RlnSz4
cIZHnJGCxQh2WBQEG0Uf1D8BIPb55A6OfE/SaJOAtt7fYk6HMXnWNqc1rN4RfHNDz3fRmqJr8rE9
yqCbzs0fgs8FNTDniSnJug/hhLtNEob0YY7OwV5k3nIbyTE+jl4nuMdQaujMYM7tW727yx41jATH
OGFNLIvsgLtGxL7Ajv345b2cw3sJukQN55Uphvts0U6huV1CT6GWGzBLQxb86bFdhPy1lOSDUg+I
L2VJt9MU/OpRJBs4+v9FLP1LbNunGBPXz0n2Poa+kMyImGPHD9o8ofdouTtFHM+MLgv/EqCDPWD0
SjaF6Nk1WlnWoMVPJm6VBGXigqsowWhwMTrGLV9aaDbfB/Zfw82IcL15Sriruh4gXAm0J6W7Sc82
45mQ03hFMytYxrafCbVkuYTV6zPSMeHWIZwPXA2CeZzoaxxZQgepdOuGFV8KSAKCMZ1aLELrTG9m
Rupbj5gBYbBDcuAA8/1vJFLAdzM4XpgpqrY6XfzAYo7OGrXLN5ZoXWQGlJzc4Q3+M5Bv1tVr86Sw
y+y5PNpSDcFO+HEKTu2Jbuq7b0vkmg5w/JYgDDS9lH8IFfwkEsGwpzy2FKdj795i66XYbrs2NavN
MhmkzQFjdK9XGHObUS3zuhe+IXuDrjtMwsF1VIfnnfeuGaIXmLmdYgppsTk0EQfW6SdMLMtrJ9wr
Fs3pAgDohjnNHBmCn2f9job6qs7DPkVGAl1jrjgfiFgyQ9aTTQdqXpdcf4s57drWXCVwKYVlcRFb
5AWqeytY6duZjgCbEJ0RCtX9qSBfk1aJ79E0sD/E7Z7ZDJfh47PXXJnZK1ftY1wAq507BhXhJ4UM
3AlTuSMJBk1d7WMw23VZPZo20ZbTyEHk+vb0b17dvsBv5nwGDNvzLO/+xyEJUWgsaWcD3buML3Az
4WUD5L2wdsylzoUfB/jhvLG9SseT0of1ix4UjhSL1BfkYDFlWSxNWI878RgfmBpnwg0B/t3nRGZu
2B/y92ztyCVoj0NJScaKajvKbheR8/lkYdy4bpRv4cKKhIDqJiKJHT2fObg5D0zxrY6HZo0fig5U
7zYIzxt+FwB2FaP3zHRGYK5J093w2GHJHBgx+lXk/Kdbeu7xOpqsTjRZRzv2Y211rSSq1TCssEfL
oKYHq9vRGsQZfrVDFyGXRcqsfAhs2wEcT/4wljWNE33Wmwy//CVMq33pGedNJOIQ2/IbabnsZCVr
25wYE9LIYxI188KVSzuOTKEYRPyh+xiu5S/cOKxJ5z8aMlY4Dj2jJVS+zvIg0Y/hX17y6gZSfUOx
y2g82mCtRJ7SRPvUEPH8xxbKM9BV7WGXJQAthxYdzIjUpdd6Raz4O2lGvQjTXaKlDZW0oaDNI3Sc
NqZwp3A1+oHLqqkpmV6GH6FhMZZGDrUO8Rlk/Vo2A3zL+6pirLy1R/WEW8yZAGXG4Gk1bRsaR1zQ
gupYmMGN8ZqOWfdfDo/FFYV6mZ2hJ+IWf6uggF1Qlop4EYZUbHhiYpzhRQIMu0FuO2e9PzpMTA0B
kBFZO9ce/4BhbrmO0eMfj7qStCCFVF6AmBe/010BoG3jdGXAVq84109Zx7QloQOINNVMp3S5UYLh
3Gdghggy6fGfWJSG65s+ERCSq2ZwnyuH+vK8cAn79FK2/grkEeDuZTaQejzkD5/eYmq+pOe+QitZ
Z88E7Y/Dum/kCQ2X+j5WDJEblWjXgd0sV4vb0DyeZmUWdJMa2ZVXWHA9fJ2EwxL9txMFQlvPNWYF
KC3rs78ND7q3Aq4ZFOSJpXAfpn7h7F5boQf6XRsaVyO6YIQsCuRZLkfvsbSRmw1p1THigz1EjLCE
abH3JNQkqwtlo1vlYYDeTzFXnhepa3Su1L292bcrW21pq8JVFBjmWPD8S1pa0H6pBus2ju2cKM+u
KIOMach4gpK2U9lCiVsy4suU43T4LQDyAvp6BYNVGsT5JFsOHrV1ZA/3/P4JBt5KSxKQuhbAugbm
lQCFD65X3vjWvmYbe6wWme//Amb13rj4Tfu5qQdjazO3b/4gM/uslfs6HTU5ClUvaBt/fbwYh8AB
pQdKqcQCxi/ksQlFhWFD6e6n0JCi+n2w311oyM4lxSZP1jUWKDR9oARv1Whp/bDqTGPiiyYOdvOz
U4V40Ng7shgHd27yHIzcGimO5LeesuVveRUGizKquBXFqpvmgneilqK8zwl43CCGiczEcDla47uX
FqroOZWoynyzlgYb5pWXPaoOdqAvC0EsNqn+eUTkw7rWNi5tq+vshQ8xo3YHtcHFMxn90wAmMsD9
+l2wanDQnptMyC0rVlvDF5EzZr0r7ZIPR56iOXH5+FlrdPc5cG0wIHjvYISIASL9PE4XDcr0YD9Y
THcyrRX7cxxajur7orn8Jx7Z+vEW8YOqpCZzxn04er/JBw1hs5GXfxrPZvHy0BigcrRhuWmmZ97p
AC8SyVMlFGEQW1k83k1YBhOPPHeS2aETeK9HIHtYFh2xG/tHWCz8V6pU+gM9TBVLEkL09VR8Gqwg
Xe8y1DLnJxaya81BtDaOQ0xqL/1eK5dN7CgsPWNd4IM6C37aKBgXlblQg+YVCpIv0OT0hd9oOiay
zopTDxQeGswatru7I8+0dmupOfk7fYnUUn9eaq09qEh5w1Mk9spKEmRNyz7lLgD67EVQrlje/Ck5
K2YX+5woCjZJhb4bNAN4Fb1WnGE9lOn7lXNvoU5RNHNoTCE1JzfyAsqChhiydKNYL+kIy8AON1GH
nVv63v0HodU36CqAye4uGzEJUN97tZPnkxDqybKesMbt0vq201aOUkkqTnC0MU42JjcZWWJpywWk
eyaDaeeIS89bNFaxOyj9woE04ayGgRb2yfTW/4ZdPBwMS3tRiss59R/FjCJpK+msEOqgQ8pwa/tq
OfNW9706QasYhmN3StkqVm7as64TZ1Z//JU5kgpMYgHy9pbZ5444QP4l8TC3jVz6/SrDMf6TQlmO
NtIdIlH1TnWFKGZfANdvoLWvmsYeo9tfR32coqvfbBsDuNOvvZBlwHOG2uZYH9k4QB2aPrlMpo62
/mw3MRMTVMaoVQ5tTmpUlEDp3Z2emEBtGvbcPqqpT0ke9sHl6YrU4BNZYDDavjQtnFtWb9QrlvxZ
mFiL+v2djF+mr69ee5fPDYojfBDhQ4KorqE03/8xptCh5rEJBolPnmYjudP//EW5adeNrM0EMqVF
auk0+Cjv7Jn0f4TQ2PALvugr+rES0xVQc8BuaSWSU132m3VOoMNVlRjo3XNgAhcjy5PVu2ytm7PE
JA0nnhAPANHSzKxSwaEPlr4HBSqx+104mgAjkJWNoq+79lVHsj/I42pFc24+yONdfxocJK6xsPcS
UrbF6vFYwqxHdEV3rkgXzcHMg8cb4jNbiwUOy01ll/OU29PctEvbMXdpLbOIQeOwQrt1mtV+MLa6
F48NWnEMbTEWqaBN41ubCQVeXXpGqIelWqfCkEVPrroHAbi8/vb5KtLyzDB6kZWmDYjzJqH23s9H
4lj8eZOFjiCjYKsgewIMkTdSB3iEUNqMwGGHJtXO1kaZ2PSEju92qzNCsgEWJy8VI0rlk/EeLRZ2
vI5i5CSIdw7lvT2o24sBL3VaBNZ643ve23WwLLmd9SevQGI6kgnWu5x7K8Dfi9be9kD6CrSCRp/G
tkc2T24RunT3GOH1LYrdM4lJQ9GRWHTdv68mxuzgQCc2YhIJsAX8hKcUqWgPWLXY23cxCBzeVm1E
I4bZbghtTYXsLIPYz1NHKUAv6qYtjKJmrc7/4eoU/oUFT/Nzmqqd+eoxhoR6xT7McX4HaL9/vHb8
wZkTMTGtQUMsP76bQ0wuPlksATmYus/a4acgf3N8VXbPhvozXcoEqUxZdDcbFNhztQuHy0Kkpigu
nZaCH7Jdxh2TpG0leCXE3WVztPaMrSf5Fcy+3gpzxF9F6PA+VDSNXLxiqk+sJu5SKPfky/OG8yU2
06h2vT4rlAdW0TlTaETQbJp18H68H8MbL0ePXxmg5L6POHH/GNxnkSaYaF6PKfy+YqIbTX8UH+60
hB6yVRn1lm5Lr8wBLOIDJwy/lsvpY5Nw6MKAwy64yvXyynlbFuHvIIab32HpMDdYz2mEyJaT0bu5
2IO2HNK9KnWhAEE4f7gXdH3rvPNrUXDauF79KSPHmveo7qZshOhVTShPPEeDHQ9NiHPkTMpLRe3/
ktzGqhkTafo9RY7+pVj4cuolyZG/cAtQTuBPq5m/XNnKnRxZC20sVuKjEWPqkckqtKrEECxTMTlt
E59c3S7GlyM7ireE6aN1oZ5JcbZwqvr37z1W82IjNUuN25+NBOGMqr9l6hW6x3nXTCUTkzOqF2sQ
BKVeTJgt7XfNO0KGSQg0vHKaYNn32jDtdp7sX7dq8m0ekv7EThl/qybgzimGUZkt7nmwvb8LDpOV
Fid+gHVsP1+H5jrp21FMDhxAYTMs7+Hx59HuC9nWljy3CAF85q+NxthGb9Li15og3oINHVshGmI3
BGqVWDslGrli9U68UJbI6pGg0iHIEmBTaIg1ItnMtpg4/VCqUJ6dimVSDgSHqMKgER0DcvyB/pf2
6QAUawcOX+n1AQSsNuVPpXzoWnu1maEb06JBND/PFWs82Q89/OuYlkX7Dmqxp5kvyxYGxjqzlZI5
+aq5FrHEH5hwSEvUPArTksnlrdXiofKakI3PAUQ5T9u8V5+RTLLuXHkboYIR9gaFYyji4bADxBcI
WPv4z6Agq/W5KYC1iCy6VLdXtDsN3dOpxdPqMCJtHMSoRWvsN2SjTTFBKF442HIFrVMweICignVS
hnIGz7nj31oEZZK4Ri5Ty/B5lAzKCYx2vg1Hgd/TLODebVnydmDVaKZU6YkHT/Pxnln9+Aqm+J1u
/XudgH7dreFkyj3ee0ocg1qomhAP9kUna9p/qm99J3fRCum23OBxiv9t6YhMgQGPLBd29YMAMMsR
lWccLjRlh08hM+0HZGkJm/Omaf2oYyKyxYYmGR5prUAfjPQzTuWjs5vmI33V8QB50I9vtVAtCIz5
AYQ8ZL908l5qb43Mqpr+lCvk/hfgnu9gzT4HXD6BIXqLUSAjCXMIHuhVTsoUo4robBQvHOM4/rKE
3jL974TjHh5f2dvOzglZfrsjBwu+aq02/WinE/yy/MIHhyI7NRA4t4xs8XQ7U6Yz9P3oqGGJ9rJl
3KsngvlxsSBKJI3vs8zBubtxMqi51DIMsrCDwqVNIpn6x/eJai3V08IrJVbk1GpH5trgQKdT5MKE
kUcP2Rvan9zhP0hHVbAk1gNiVRmaQbDYCsLMbjpwgc9lBQJ0W11q90TzSgEahZZhnd9ZPr0NAghz
cTShm1oo5f1Glq1N0TRSKcHsc0n39t1XhK9kTbjJE9XgfjcOfV8erjZtSyfYweYVcnchPS0bVt7N
dUROwRuHKbNcrifPYeDVrMkZQJ8H5numl2JR50O73e465KVcT/DzNvwz3uNPMvV+ZuMAZ7LM4+U/
ari9U+xnHS31KP8xuqWfxiw4oHzLfVQvlZD1G53svjsYMzle1zWPGAo/oOYB5xtWnDM6m8C5QiTm
A2sIgtLEtqTus9Sd09e4pclFK5xgklIvkaWjV+ttCzii77CzBz3cYFkIvaw317ESF2XUdEzDIkHF
HP8Tg3bBkiUGwMvBT1DR3q0iQbObP6bDb+wedmiVoBr7TtWoboJgDVhAdf+j7kcDUFtAUGMGECRf
BMnIIUVHRw16BS1QtxKZvSPsToASxElrUQcM7XmcXi2y2oYGmXIryKWPpfAz/8fspnfKYEReR4CE
N+HdZ6mSAGxQ47I7PuDwDYg6cg4b0Pw6CmDP0u6xfGPe2a96jeFwdxajFoTRD13Qwdp1XrTMUk5/
LDgH6eHZJFfsQAoLXvxBRjWofccvW3lk76bW6iyrC26++8xjWFEsB7mIa+kz1WHMcY6jQG65kqCT
7+eJ18ljU1LZKYntrPEv8lm/akXv9OCWUzM3dmPdbuVodB2P5waGGm4crcgBFSP0XztRyXX3n0ih
K6tgMwcJituMLkeKBewuk9xGImFh8stDIR2NuRoxGDpqF5DcTD1nCXGs9iXOXOtMibqNcxQvfCrq
1NNF+ezZWmC8v66y1PscPwhdljOkpj4d9DEWUKKhOVQREEwl+qAzIaQ3lcSab2GdjYfUQgh00/uC
FuEmoU7G24aWSfUu5/1o+LIZXy64pOzuxnPptS5+HCSDksmgWCNkO+u9iA/j9VZm9KK4r1J0J0tk
Br2WODxkgEq+Qx1MqMQI731qdXlutg1DHL2bLfh80muq19CKmlO1SGjvmSbWOhXFHc0rpquYaf0M
m9TNkrE1Ixv1Ze8wzubdoPMBTN66CtKJ7bsdZnEnbDr4UKVdorcof+WNYED3lw1TP4dxsHhhKtWp
xnUewjeUAo4zUOci2rBsdnn/d3RZSzZdzOaZjJdxKPmM1DwCmKG6gyvHTDo3D/+EbylFOmxM0EW5
P3KQ6bPZFH+gML1iNfL564tZ1iI3wa/tIalDJPNZJYGvNNb4WYB4LMfgJYq7a6sXzuUcc9XodxN1
gYN43Wx8H+VKz2q71srJYMoMpA2DUvsGGoscBQkXvolsYUGqOMaL7D7PpUjaig8sQqvTphPMixIA
Pdld6/BTENj0Ae/oIXY3JftVMhO7p/6pinx+GiFhuPlP4XWtwVUZriAnu6+0f0neMVGLxAqAgjC1
LcBTwV2r5+ragwfRq2vqfp/8qfOJpZGz65ADMv0R+CrqyyORNRL9P+5oJPjNKrwe7aoo/VdBB+Jr
VxuQbvNUyIVgXxtw+qtvqGYKd92B/uAiUs7k4+d+OesKH0Qzvr7p6VGAA2PqPdTHO0zzVbjO0JTK
Frp0SgauPLyKkf6IwcqLQCRq0UM80c0OXFyMt7sfA40hOWKwByl3NLUQyt3B335XHp3xpnF+RSo/
jzONsV9zgpBOR/pZChCvHHwZpnLbImotbRZVEXmRV7AhmgAh7teYNKoWNBeL2/FodypDCiVnarME
wO8Sgd2KykMq6Q7FWq0znXmQ03DQOmVDQEDedG9Ee/CMJtuHe7RBoVpjfjeKHd0aE/PhmPNf+ksO
Ub1Ri9GZ9og4Qv3xNrJZjthAGIEoxtTdvDO6G9xZv/85zO69DMN8+9T8DLq3XVAd7XeM6LlFO1+t
999zs9WyyoD+H75SFMnZZRJt9hfDGbDz//k+NOCvvuYok34pmeiowK0WJH0A/OnZzehsiCJXqoga
A3Xof2thaZ4XDFxcPQyVbdTsmXwVx9kE05S/+tQxWjy6sTLnBVxZjl2dFDTcJih2wZfUeGcxtHLI
13xw51orcBoHip9rYoV5cI9eQDvypBGZdGm4Hsi/u7/JjwL2z8CAtJ7GfJO/Wuq3G8dWi6GZYRd3
7eX4185GzBKWq96zvCEnsOh2/YCqS9s9Eas1apONoHiWbxAgch1UAhZbUVzrA27Og0LN7IlYxBiQ
9vXtzXALYpqIL/5g6o2gnt9lcsdW2BfONBY7IUsDLfVSDr+WuP3qz5XmY3RzxV6EXfoHfY8Hefb+
EmQp6wuQ37ujZsJsQ5c+0rlQUrswN/C8nVmf4UFGvTQjGR2uqi2NVhktJGnh3EOHjyhW3KwDSUhT
vw637bnKttLahQwCyDSneeul19lMgBbAZYZNGzWz+nDp+EmobUMUydkm8UkQ+lrvr67ZY8IzxcX0
vpLoai1or6KiUiOimV5SInJT/H79icc2Cdf7IQ2wWiLFBzJjh1eQ6aYEnRY1T4BlfXTPII8pY2E7
PuWuyHmVAQNEa/e4eQiDOYZncd9GoIPK41ckwL2VdqVGqIDmTafv7jHwt8UgjkMWW5VD4i8hR3P9
FqyFebVnw0XtDE2joEEwynBeI8WGhtEa8uaTSz9M+K6Lg7RC6BCR7rAsgYLC1znOU4qVCVTQgdqA
koTom/Na2bKsEEjVWL5rtNw3kgf1gv5dxkMyUzWlbyzDL46nAmW9mZOTDEDj9FSvh41iCk+azRmX
lgzXz+rS3EZP/+BfF5SPoGm5JwvK61MXwaDrOx/2GeY3/WmqrY9HISTba4SuZvnXRa1V9qs4JNZR
zwttVpBNVNvknF1o2EYMCsHopNwwaoVDCQ2V63StbVkM4Zi82BL+ycP/li0ap79z+o1z9xaUEcQ8
iHG2+RSMWxGDNzT8prCIVINc/Of2plX5T2oKF+6OpW258vcBJ8gYUVu+wxeRRANlRmkIQxUWTj1H
MQWnlzbU/yFrzKydrOZGNW05V/VlUzKJ1mXYGNCF+U8EWwlLdQcKE72igD0zFvYHZd5aUQOIs4Qq
wLoDuYK+DzjFla0qrupqnoB0y8GAU0MgkFRA8LCq8ndjqFDXeR1WqS4ynp+WdElRsgYJkDrirSKZ
pxGFGv7euOkHPjCOlhQp7NnmWd/aBR5zKSf7JlJKGhoHzSzITXPfVhGpNIs1EJmmCv0fqhLBonvp
rm317942ESnPZNaJlQVL0+FtW91hHRWg11aRoQJKt20Qhlzh4QlE3CB+S6rY1oT4GsX+FXSUGEwV
SX+fCMCc56w5o2OVUQuSMCuIaVXfKy//smrxFVk7xpeW/1D9UqlDiVi+eOxStY76jUqMhHD5xNsR
G5vaMbnN72X9pJyGJoF0maSSeT3TIdXkz1U9X4onS8DykdD0vYXko3IoR9ZjliWsa9ckfS/AXqhp
iY6SVP8xth58oITOqDA4hpYyASEz/xU+pyzKMUwjcklIbaoYXUveLHrM8jZlBVl/QDqzOVu0zyXV
tIsQjrmIdfI0XG9EFOS6Q2E1o1cUVGT5+Ki8W4XcJgupJFvlbGBZMCZYh6uVWY8nOyRi7xuxyuuR
VidQFdnKt3pb3Zd0PSY2w/ChS4ZpBAb/vac79O26blTDvGdTAuSxMlb/zv/8PvTO+xPz3xQvlDQG
/RqMmflHsDfdZqBDKd+wcw9KeysXywlbN72NYMj9sp/rTkpbop0Lq8uNBbESomXOwCDTOfZ5Vzv9
gdir+jYcca5dyF6t7tL4t47AruUxV2ZPxpfstf5vfcmmpj5uVZY26+Xn5EplVqevL/fA0ClkJfBs
l+4RUdnA41D+jiibjF+ZQul+uF4G6byC8b6na/ONe6Kym/+niCLCsmA7cyd+EK7dqVm2CVL4zDpg
59BMbgZ986AxtR1xrB0O2hwWi2PGpZz0227KYv98MmuusojSge7m5SPOoeXfRl5YeOFRlSSB1AON
oNrtIqfMTTzqAoI4h6MXVnsXG+WCuiYfQtIoFYxq6PEwqCroUozs2/n5vtHuZSkpvCWD7xz4gOjg
xTpmKRCoTgAqflyQjVHFrP98kyQaEAg08dMsj+VsvMLL9+h2NXmF1BKtt1sXqniAZ6zlGgh9AQwL
lTehC5KM8p2UoZsgAysgcrCKj+R9rJ/zPiT2SGRQKmWvk6OccU9tCZiqHBIjJmW17Rydsi8NJFan
7ZFrQYWzVFG6qwc6wYG8U/YcLbBcERLaeViDqmpkylDACjlySX0ba2RB9cz9VJi4hBnpZuFVokaE
QVLVehPLp0pTCKRfVPmtMzgxnLO9mEFvbNysh2weFd4bfhDfj1+5CxHhHZiGP+mtYwSUcWqL8QMU
TWbXC0nIqX4vcOSqJvcXom673Y9p35WGS+CExYghIx4yP3+CkHx/aZiwIFsYrvy7J9zfo+3D8mZs
y25q7Db1y2VP/jiECaVHq10Ff6g7cv86Rrw3sX5RRJnE0vZScP254adiNYjw0mVoQ7HLI85d8HqZ
2ra89x4Cr5Z10qe6pGUWkIdvq8i7XgY4sFX8YlzC464V5u1Q9MJNldTyeqiWlPSqQDMcvzO6UJAb
0K768jO41H5nq4GpqkUyU3sDoa4fHhepE75PFjEBs2B1tqSH9YGKOsFhjM3zbwCbq6wEJJEOjXEJ
xVuoYHVIeKzLjsZ3TR01BtVVggaOtzn8M2z5K8ejvAayaDMLr3mBjBkcOej+Rzeum7RqnUW/V6a/
gOiXNNc1QJoqGAGdu/efg8ry78B2IRXcIacmchDbGgrDfq8QDHj0e84YGNCvtFpw1jMV5X2PFw8p
NOUtnvwvRajNmiAQhm87uObdgokjDlbfm0jwuIUl9rvHnw1xZ0/jgNoShDkRG8PcNlaNfY2XKPch
VmEat94/n5nzYE7xLCiL5wltnNI7WgFcFeHHgfz9gXH6Hc7zYbllJ4GtzNzmQsjHJazBjlcyN3Z1
H7av8NtS6QEPlfyKrZbzcdYAiFndZNC4F+vmi0WFGFDParR0f/1trbVwQITvqp95X1kf5ruBH1ud
ZqKVt36zqfuB/qfyS3v4+ZWlmQ88+xLnNu+PVhBymZqgTj7kYb1lYLbdnAxLrzg2+Tfah2eVbqPn
djnlCsYvUsoqvQnp3sgseLdxpuPTsv4hgOqTvvjp5bboBXbZO7i7e22LfsNU8W8J9ssdGR5FBooQ
gSt5Dn78kH4krx7sbnlRZaCpGVsetRQ66M3qiJ71Jl2bxGDNAc+NCzZPZjOZ/JKATe0fAr5uXv5R
QO+J7MbnwDMusqNKIFgd0VYOX+MiwADaaZAmkh6WbcVRKN8JKl1JgK6ZGZ5VweytesatWDeMCio6
I9zYBG4EdNNwoJ7H1cr0n+32nJfH3a8PQFTuQPK0TBLCTtSbN5+Fc5WtMArErLEbphr/xqBflze6
8fYqJ66ksFWT+L+nHVG/XlEQ8q2S3X7vPLpQBYuISjEBv1RLG2+7hJ3C9KGWQ9svM0aOIkrTEntN
WQcs/ZnM31SsZyqhE6t/iEpzCiESo8JlzUYCJMnsh37SRydmdctZBu4JMvHvgDCvSDZ0cd2qFXoE
LA8Jj8qKWqjG9YQDbyG8U7as9Wp4ArncOwMR6iSh2W3TlFLNpHbSK2yygYWQdRulv+mPUNUgOoGI
UgXnUkoczLirPKCp9oLm+wJZA/WJdliMcX63ITsHQtS4tE81qLgXCokDXs05lFFM7cEok1aQyxfi
/byUjLRakBjkMeNJUPUcNbvQsywNFcneYxULhxqkUo0U7Y7nRMqoH97vm6un4SmjrrmzzgNsKoty
0YLXy+NLXpasfg6VKPIJ4kKiUdRNVkqZIZXaIhtTxeED7L0eQTVMnMUmEHhN7zFN+7m9m6h++ZfY
gSBSgB/k+cw9gl1q2/fPslPpIz+gpT0Nb0nJlM/62NCTv9K5n3+AoxCW/CerPxwF4G/+nf0B3Jfo
y9MpN0hUsAwc0g9Dlvh5UlSPBRobVhMHCBgurVWkQre7WtVz/yDeIKMbP6LYmz/G7c9M4R3d2t0z
h9K9EeeA5SXnnNGWJyBaNfqK33xlt3VpJFZ4yYQGUbdgjEXM776qeFSZE5GDVeBRtNfj4AlMWwvU
wnokAzv8B7+vmZfS0tz/NqvHIq6S32h8dXN9LpHhRh9jD2Zt+Z0VTypbyLtQTHmsBN3/2rJW8hQc
kaZXDt9shmEfcvgL++QZJUlXA7BvgdeeDGr0cBuGlFaa9WmkekDAzX5VCKt2W4qlWwOuEFeqvclt
AGBfrWy7D22cy8q9y/gr+Zquyr9GrFP37CVmO3FYuDVKQiuHOpTB3OEOFp+sPgmXDdsqsdcpMHSe
9UCsJPPLjhkq91RoRZLxy3Or9B8l1q/AwWg2gZQwn5iizafrkaiaHa/mtbwXVI7rlciPL8cwBzqd
Egm6gXpwhOlEpgq+fAne/uX82W/XJwKV2YuhLYanyyaEeKzFsrd1UWtz25xOqG58+GTz1u6GNZVs
qa5iham0R7TmZDhtScupU1OFHoZm9igY2KxGLCve62KCFinWjXVrKUJhEmbqSk9cdmWvYpdn2OEi
LHhZgfOoBPzCWj5ptHq8usCAeyr+fZEHafJHsSZ2mBmmXx+NJgR8ptoi/XfurMlrydCI6eB2dlkM
xrVToB0nDr5Zog8IQo8sKUyGkOVmDcErfMt+v0xa4pfgwoHFmgjnxcH+SugqJf+jyocvB2eoWLJ6
rDplkA8Yh3iJJnnND0fKPs7QFBgpmWHVdgKDHzfdyyTXYKuA0SUWuvppfEdfiQkTX6IWSfmdSuJw
uHDC77rXDKtZ9JhFZqVDCb4RUUBE0D9rTeeWllLjLUz1DffZhDcFWbGx4FgdQIUrQ6otCFFdWa1h
17mWTzI/hW0Rrra50KTGzMrXTBxHOCL6kg2JXpb9iv67N+u50rBB8HvZLdPkNw2XxXnt9LbfANlt
DSoHzaHi0vKuO+42o7Kn+P1DxwTQGumT0MkZemnt9Vl5gQ5XNcXe0oe1hk89XzAsiNehkLbD26LZ
Jy2Fvc2CVjKTd1iDN7aRGHWnE99oYDngiYN3Gk3HXl7xQRS5+xFHxVsaGAZnBSnm5oIIvEIF+AbD
yQ8PWqXY1qB5ZBRqEeTwEberHm+zzMXQweUyzzjD1HN1QK0WfWnXKdI5WYobzRApoyQzydR6u+1N
/uump8nCh66HESkwTRtVBxhHsqZyKyxXufjmtZMPugLr+J9B2wJyAxfpfGwWzXX/AOq6wyt7c8PW
lankc96mPf5+ZXvA9khWFxIsiLyh2S/tS+ATwFRXpbwbvMg2fkvn6u4kp0WIrWo+U097yPlKFByA
epF6hiuXm9ZuzxT8qLiRN+ZH/KtxQF7ZZwkUcmepB47r1YfBNatlPTV7oCwbUhcrK+pgIAE3IQnb
bwitrJOxDeOJPpDsWLxFcQHkXduxMFSq5X5qHpVBW5+gGRufJSINrb+KxUPJswyWr+ZRjSP9DDtb
rKkmVDBcgFh7IXj2w9XZb43nobsaJBCgyhl0mV3KVVRUErdjj3c3O6Ga9/ZxaU4h5Y9c1C0pWK3z
Gey7LYfWVD2RSuqTbABYAbJhb2dgXTMevf2NqZcwwtgOMEZ57AhMYGsW3kUKf7xYPSc1MN1sLxWS
MmZJ0zV+1dJYOnfGoPtUQUUgNIrZ0SKyCccbn0/uhkQDssxp52qAxmQL8jYUU5+mFg68qZ33cLy7
QkqefieFXFl0UDAt5KwYcM3K4DuSFG3EZIA1g2YJ1bhDA/pEG4o4Y1s1asrRmi+QEnUWBLYt3qSz
2rFxun9cghmrruk+fbdZKDq3dwfU+VZQfvPkqpIy+/D/k2zoNFOpPm1CEuTBo91wQ+/erkKvBxiK
w/63o7vDQdYVyqfKUyy1HsilbShfaNhMzEcek5313Lsu4fB/q8XilQkijK1wTfAZf3BW5tEGt8hL
WNoceN0iwq89FEuHBI044sPw5NFnRG0MAHUwohicWOmW9+AWDVxogHcSmi8sAkmNqhcZ2FJXWC81
KfoZimIo2r81lyJQq9f6+zZFrC1nZJ8ko3E229jSrJySKR7uiE4QvZs5wDXkF2OQA7RCP34Li6xT
rmfrO9gVSDG/FK0dCBm2RDTrd/OOBs2eu4vjt3FWT8QSXivtf/W9yBf1RF2sjcMMblj3fKOnFNGy
jrFrhKUuRmBtP66wQtdg0FxKdraiYFbvsifytoA8yIGzEdHqMWcY2DoxKo2skBoG0uyUQaXavD7r
Zw3DqCK9cxIG9l7WbcMfhe3vlnVT/RykeRhgtZJYSWusWOTlyJ0dD2nHA9Cta+FiGhxhpBGzHEne
oGxPb96OWmfrP/iMaKzIZi8SXHglTMty0rQ/3E2mhHeoBW2rLWLQ2BiONTSVsz5b2HDyQfP8yGXj
b9kkVzCcMaKMu9gjghT4/3XYoLxBGQgAYBMcIIhVvGpqjxFN/oKHPoGHt+VKTGBhdxCfN0Wlnvmu
H/O6o/jWjKeT8QL0Y9T65EXiktleeUeck9AD3xldR6SQ1PodzFSgGcPutRYjOusoBB85jO7S3JPd
EchhyE0K+cMgsUKc5sC9q5N1l84xW5lRzjqG791jSTXb0QQrnm7Zhj+WoFzKnXjAvkD4JxNny0Pe
CNgsrHLA/E2IXuWnpIOmVekc1GaA6Z5OoLZ5PYs6uXM3niGSgfF7nMBU7dGIruERpQd6Hyd32/Fg
bk5hMoNr2ID3HGWwE0w7ZRqi4lzY/6xtLxalN1HgHy98e7dX40+Zk1CH5Tw0exShbiSFZ3RTMbAw
XDAnjrCkHjNeh9BjX4JL3PhH9yTTBGKXB90Zuk7/xymy2ZHcJaqfiKYlpBAwRvmhIzN/w19Mb1tN
RVaJ2dR9SRrZqdzvGXXTN7cS5+/mfOo+Xs1PGSWRZVHRU3HcstKQafNnkzEVA4h5R+iBkOyafT6P
k7XQpntGNyi84mj9HM+qCWYxFz3Vfk3v75i0ljcGpvJ8lmK5jb5wFnm3FOXeCPlN/jyHCw5YIyrt
BcX2i4YXM0uy5kVbJtKaPqr9aegJJdMQF1cXeTyl4rwq1hmxQKFUf1GAoI2nFS2uIXyVutXW/wnE
YJlucmn18YzgjWBZmpxXZqTaL3EolFY9DRvM4DyRaJr9hIFOgQCRrD6cKrsn4JSVwETssv/U2Dc8
aQyHtv2FgqqEnVYE0XzY9nLPFFwq0Z+Bvh0fJi8YB7YW5fiX6wqytBq4gnw4wck+ylvLWf/2278j
9Pku4v5zwQ6sJDUM9l7VMS1p9tIbdAY7eHj4Koy32H753y1jsrYiGUuutx7KV+D4gnXnE4BBAtxx
aDtcMuVbkctJhMY7RbM/YmliNjLegwO683zhl8OvVcM7d2QOABrj5GIMO5WfRbw9mHD3GQT4zZB5
cWasw7IvDhrZZbo0jyg0tu+m06L3qDDY/1qNKhhbGhPEAcQ6LA2obvEK1XVrFKOk8oUio81YMWuh
xcVJ/G4VpHL52ok2dVE3VzIc0JyOYX4NbSS26IdQ5V2GY1F1uOU4nkV8FSgqLiaCvw37QhsTXXF+
pIoUXDyggg6HfYxVMJvA+OUfusfvOiHmLNQW4IKoJpgYt31X4S/5BPoEDV5G5KcZozZE4A+w/Off
SRQ35karik07W/K1AxQrwSQUYesEbKf0LgL707LmycH/XpXRaWk9bc+v/Ef487nOvQS7EUq4iCfu
sEFpXe20Te35+icCnjdejAa8UBfpwoThB3jp74lFEkvywnZXgMMqZ2T2+w0r1S/y0gLauQLXJtic
NzFzCYrm2X03X29BnCVmx7qoAysW1tAPDFqlbT8xOf7tDa2D572NN7iHLn0CjqwNdk7PpCNBDFqt
mNnLfc1p0GS9zXoLY7YZvV7ntPPzt2xufElPzpFtDL0HZcYDxAwMChDQuf6uwPcgI2vtGSL6AlQn
iE3CVyLxuDTXgaBMUxgA5yR4fndg5kBz1UqLCLgXWNn1qdHq+4VFmCPzIESZeqddM1R+t1FObYcI
jSKYVj0EoeU1YL1ZH6o/+EfmdDgxR3tGNJVP2ghiSWEp5bkmMFVyJcoitYb+0PyvziV7GyReOlYh
a8jJXyqxlRwfbbXK3CbDQ1zUfdmdbZDWVvtZ6573mv5v7zSUCQGd3bGqaIgYlVbL2rOyt1K3CeuY
zf1dWk7wvqZ7/itZsBkAg5CwKxRBmGO4ixif6ECpU0Sy4G1L66aMH49cviMvZUbuFutmm+w426vC
Y6esBqmBSCxs94RgbPmjQ4Qz9CqGOS/fdGLf9ysMzMK/OtB+vnS0cZb9nu4KR2HfCwH8OC3UzsI6
rGBXkzv0lIVkWzUuHBc2QT2ERvKkCawwBd8utgf9J2pg6S0vLhoP3j9xAIjgNc2+bz1Xfpnb6jkO
N9tE3XypTJvTD4L8pd5aKUH20zuuigOer5x9qidXcH9MTcsXmUVnu5VVumvWx2hG85pgzGyUfwBU
nSLjJUkk9/Z58dEZ+gX6oCquevBuw8QbAyyRkRtA9UJPSmXSWVr9cJDjRs6ioENK4NzbWMbe/GI+
0ctOmSEuf4o0lOatRzukDyZRiup45UatgoTH61dzJklmV2M7zGTLbjyL/sxbBXVgiw8oTT1lAKyV
a+K66nqkoJ+AAZ/wGK2tc8Cwdv+fZ2d6uGD7dZWQTXJ16CiX5q6MsJGKDNz/aWp5L6aEvbBWiS9U
YsgU7vXcGFDALFq6vCI356PBKmWYIpfw5g13QsobKwqGvnfyiQrMl6ESNOwu8SWSLBtcLL3+38ut
Bqg8koC2/w+dEOt8FPxRHRALCb7wX9lzxvO8KtFwLE5vCZ6US309SEVg/emy7fKSS+T+lz1P2YcT
dm2tnR/jristPZlZjAwFG8zI7iCpxmi+JwK9iGh1C/9N8OsaEHqqxso/2LcPnK/wuBu8ljVu6lt1
G3V5+1eL5kW/ucuQAwsLEnMUqK1x6bQXMertRCNf86x0OfYY/8hkIA3v95RCBcjlPlVl+4vSkDzO
JLjzs+F3gdCKStU7N56roZkwEJKssM24brIgWdRUAOs8TAS/qDmbDK3dP4dT8ehDK4GXZE6aRT2a
uOXGH3IhhjTewNem0B1YUIEIPLQ8rWKKpNcl3IVj0yBr99BlsfXY8mefWnesJc+7y0kkhrHU3J44
hgJMSEmZFQ4y7s2/iPMS8cDl5KEyK/IQY3EUwOe+XQEeFDbwfsQwg8HRUfmWEkD/C+OSrgjPs7WX
/oDq//DSZ+rSDDQrU44HJdrBrIShymL+ZifidYn14+V5EX9K1bbmW0WiN8LiTXLx9wLpDJp5Lfc1
BE8o93muvpmyMzVIIpNaPh4/vUZzESpVFpxrlIE097DQNCjoOjo35QgOWqluUiSptSyLr/7N7CvF
C3Xj065kK8zm0VnMtoi61iHHHKSuORdnp2q2YqTN9W9eM34Fs8Unbf6WsZNtOfW+KnmAARxPSNiw
eyu/+BkDMxYsU1AP9bHh8ISxs9vWITuUXTu4CLmLJHkKa0aDt5mW/XNwPvcHBHk4Yh2Ht7fNAOq7
FxRsGQledRI1MYn/98rqqe6YbxyIjUvVLyoILSF/Bd0bnOTrV4s61bKjl51X11OVOX75KtatgW8l
a3wlgXtVOWfGq8wZVgnYHhg5hi9vDiGJry/T78Sm+raJpMIwwYUrRgbogXhaPLdm2+FOiAJIHS2d
JOzJvV9ilznIneOvplMct5aHZFZ7wP0wyZ3sJa22AcN9+GlN3oPcA8wi1cEOot+Q11fMrtr5cvCu
FWyABOgjcSdBn//TBUvmxJZoBQ8kKEbDBQa2VB84hQZeByTPw2W199pVaVgvqRIPFst4h71jBMTz
CyJjkerDrdMXybhoAwQCRVSTQzekuBcnc0brs4gLmbPNU0I/nHC4UNjYzt7wbJB27sDgpDd8V9sv
6877zYfvEAGcbzlpUEWAn9sUP3kIFsuuJX76ctwqnVgrqoAjmiPFkEltSXwcQQqLt4Zv+NAc6utO
K4YdVmMw1WTAeM2MKlKyGvV6tg07j2CYOSeYTecBECsAzWECxbu7FPRHVGGb3VpXrP3KN5nDHTKd
p7PATg6AUilvtfpkf1V7dyFhbwBWoURmDhaRM1v70kVb3BFYya7cQE3kGUVmWg48v2myZJVQc9wd
c4kKfgkpKpgisMR5SOrm/J4QuEIcRX96CuB50vWywyqS0jflCt8lsMGka4mDgqMQ+k6CLW3Gp3z2
6glGBhi6Jt0aN+LGnub21To3LZP1TByHCC8y3xKACruz6tMczn4OJH7AlQaoCoB1BZmaWSaVfBv/
0cPdf4hemRcdoEEy/xr59RTwt/lbU9PiVdB6bodOCTs6oeiObAzyV3kM1Wms7F0szI7rY2xJ4EaT
SKCLak2SDNqWJLAexnfMkaQJm9qbuX9zTYwkOwl63OVjY8ss9TDq744vvYVF3Vrp16HoXBegq4OA
Vdv1sxSr5Dy/dg/PlF8sem4ETiM0bJdOHDNa01p1ucRMAdFhlQrYAcOmHSs4Ort7WXe3SaRWkuFo
Pt577ddKt5Avs3Ro/jAtHg73QrF/a0lPtf4WoLmNaLZhOHYuauGtXgogIf3xi9zfsYSkBF1oM+I8
dtTQIretV7dqgt+qf2af2VfPQ3q6H4ft3eR2rFB9GSlF4Be6fHRmu2YiqlVYJflA0O0eYplOC4HX
dVJE+s9Fe5ATgO6TnrD0Y6QAb2qVTAKfOBdrZUPLgt0v4w9F5w36C+GFShzyiGikPhMUAIPP9l5F
4j/dd9TdV56U48qnv9ZUYf4QtV59azYtSqHS3bveo1NCYCBC8j5zzFgmxA6t41W8lsASAEAiJFcc
WYkeNIpr+EK3FNCXuhyl7WW5muWEipkGt9sFQXY7Eq2fY5cFH1iDU4map/LUkze6KV03YdGQurkl
YwdPJ4FJNDYnID52DafFlXFKndWXwzwdM0i4BZtuIJNhZ1tMCyrVmORPXwOGOW3JfKrgcrLkUiaG
fx0AKPylmFNeFAn/SI9WSYES4mCjfa2Lr3WpRJ4wOgfCnvNaD44xR4KmQvLRJXIvPNcPc5a54da8
p4wqPVpwXYK4p1FWSV8YU10WmtPyUMpxLfd98R8qZn+NNPCJ+0xQiaG+mTlKnnZ2uwajmASW/+5x
JRK0N7luD05nRHZdb7XjrXkYYljFtRluuw5YWahFIO5CBFGFNb01LDmSYxRGOlfResYVCdxtBhN/
q7B6WTujqKaLVYtuwaAkiNprAUiECBzEAh+HZiYJi3sR/B/Q8ayRKSfiehmJwQKFYGqdnoxkhV4O
e+EqU7/ZKonv4YyIuJC22UUmvWNsMoYgkqmQufXcL5FUlmsCRX5rgWMRARhATFotQMJNCmY9ln6M
ghb636E/u8ssD4qrxPb5hmvthkhpaoYnajiZvRKXnOhzahzE3XBxjhN/c4NWC491Uskf6D/ABlHT
/zAC24RqkLljFx0xmtNzP/SXWMDfXsikI4yHxBgvTuX0xX54Eb924kkClNKmvGqC/tvEUZEh9ZIo
ZdLk0KTt2Bu9aDHudsnvDb8lyel2yGqI9+vqPTo/zW8omi1lXsZdTSky5bAYFfG1XgPXBXKwCIk+
KOxjZafAhn16GwWgpGvTBIgqCxU+6IpxN3aahWTS92tTrPxoPo6Agq5P+lCBtPPxA/ptp5GDV/n1
OWRfapMbHnRQ1/d+9Kttp21rjh1RHPi+ILCHhFBDwFCEwC+DkfiLvh2E3ailXRTNopwaI51m93pi
VmWST6wIOIRnhNCPkkoh366KEDyMfuOApZojxVvgt8npAjCR064PUqgKs8vewbP7vnvq3J1kmHdN
ak1VtPY0AS9kwmAjAd2XZkvLwcApmrvcK11MHWnvpIKZZyqwTmyPFVpdu40NdoTuKMjxysfUpBV6
q0aocrY9adAETHv9onNVGfptmv/c+jrvCVMlzQsRP2JmUNP86U7yWhc38lnRcLcqGhPquK28CXvM
tHHjLm+Bfe1XjFtAdKzKYJoDCtdEEHGeSMcy4GKY86zwOozyn5OzT1inAP4LZ3VDg1kiktWxvSWl
hHBlHtszB2u2IsPmPqvNYlWnTuTzxz5WZECD+Yx8vU4RLdedoDQ1hhsQuL1Ni0aP/0qPXE/EKhi+
lXGx97kl2aOolDdGobN9V9CohspGoc9t0iJOEyNHEnn9C6RWsSPbBddty1nJu0N5OE0Fs0HVfUaX
K0BRLU7KwrbFKrnKoAeEaDD1NWlxUghwIUU9iq51O9pbb/+7R9YFoWGoICFtHY8i4JsAH2eoCPZc
1Z2+IWorB6I0kLU8I/F/QzyXy0fAmwEN+N0mvVBvK+RTMPmGc/VMoSzHrkVgEjwjP8TH2OZOFhwl
HUMyWUf92gm3V9VodKNVZaVnrZh/ajB01mHojSMKp5NBoONASrV3J9aFzQPGSniq9WyXW05Ahblx
0mzhEvJKfquUO6hZoMXpr8IISA9NBZPZ259QMynJssYGuUeye+9KYZvsdZgH7OZpQmajsA4VZ0hK
RiZu1GA/4H4Ggj2oLMx17cqCjXc0hP6+8ci8e8+AZJDnh+NA+c6CIjwDdre7tHrHWWCK/fnltvKy
7+pikN47CEHpitVKDYkKnefuKH8ZGeMj9TEXhO1l3N5KPo91UJW/cIcn2qPvC7dRlnLhKJdW6yUE
Taqauc/YGCBmgNBcdfDAjX8FG9ZKhvRgSSu2fIibIXga/zHjcZFpk5WkhPggDyLjdGaUTzi8V/Si
TrU7C6ifIR035YPkvx910B7oCaeLt/HG3qrPyPqTfLXwyxWS/ZK0APufi8jScB8C3THSGSYStm83
7xN3wv4Sxpu7p5G10KXssbS/ahkUX/agkT+JdUwu4xDb0D4WXwuPNV0iwYaCaH4nHeMgUvjJ3jmf
7cEQeBlyIcn0T7dopeZ716/0JUUZMuJSlb7W5jK9T9IcGEdDgnkTWS27lM1UeBo2PSb/Ejz60flW
vZembeHKPk3RibWAljkS2o1kuS24CLyFwBNnhA3zukRwNK0UpoTzN80AaSIQDY7qvj6dYTXIytWG
p5ai+0VC4mQ8rXz1Y0hN7Eu8+37e2o5nxPXUN55DM9rrQ3miezD24zWBr2NfamWu9xIOJnmnvkbD
1vNrse7gPyiC3ON0ZDrQe3PTWNwE0jkqX0Yx7IrH+D6cvJ8ezMureoo6bpNbCuxS/Y70RzaGCMi9
fNf1b9cY1S48Da+Jtx2/sToCEMbrLihnHbaia72w8AYeUNpLcPoWvh+OJ4JvCJQhszWrCoUDqHAC
xnh6XAqohQS2WZoXSAwyR8bsBAbE98LGJXOKVt5fTSrKWg0Bzb3UJl8QowHg/dD98R/N5IWoxosa
qDBibwtQ7nSrSvG+VvNvwevxjcKZ3bNYgHyQR7nCfrC9ch0rRfXfnRAQCQgaq+9uAGU21aQuy+8X
kcXLYO2PV/lqyyg/2Qeo3K2J/Ik9z0wwC3HWOc53f0npX/ehIrrWNNoeHTvxLiv3xVRWqnhGzr/K
RTnWyUNu+B1QMElA8uZ8sVHRr5HBGR/shppqC7Z7NDezgDJ921NKfTRiAT8eyqOaWEQHuulUi77R
Kb79Qlj9Sx3l2OngT1uqUjNlsTbPdSGeN9B+a2+3m8Govw4mUK98ySIuE/OSmN6NzalE4X3XiXQz
V7RSP4m0vLuhZU6P/xllDUbe/NfkiClMLDROxm8SRygLpI9/JJ+yhvqnAazL/bzfwYo/MeLy3BkR
wVk9EeB6gAGkkfAbPZ5zgGrH0u9CjmuWTdYRYAncewWLM7KUD6CD3GvB562DrXnXlaBzxNrz8T9D
9uD9sR4tU2dPy0hHl0Eidfvp0gXwNoaDUtSTodTNfdm75arSb/oYnuJOY8xSAQx57ToKceOc+KkN
0iA5dB/s5y2+XL2XCiJuP7ZPysUbIqcRpksZD4ZtUA1VJytF//F21ix6thhseKtQfQwSDlIg8xRJ
pJ4q+PUh9fjjlV64cwgEXGZKOv+g39jqQWp2izW0YR0atPQkzHh93p32RkjDJwWWz2dkoEe2a6vt
iRKE+flNyI4nBk1RT7Y9T7YGkl9iD/yyRRrWmXa5XE9mWcVRs0aw5biOpMtB7rrqX9hx5wOq1W7s
odG6m4zdNVN/eo0KZSxr+MK5dS3dsKPyil8y20ZNZ+hGp8Nwucc9p6q57X+EgY8hAtQpFLSSHx7F
A6QFWxxnf47uZ8QA1A9wLAbjCYFNG+Xr+s5vTFVagM6gkZgQvZ3s/GVnArT9htjaSPECWPWLDwnT
94528QisVS/fQHhMqxpod5sveoDdwuC/6LUPnsdCYvVVVN+I8iLlXTO8kV/lZ1Qua2uDwF9CWbPk
/7C/15/WkMyxRINgFIppjUcv+X1TO5p9uXRDWWdbN4Z30hyEhFlREuTNyKsRo+CvdohhzFzOKjOl
7BdIwdas5gfIC63XvkK3XWURoPr+QUixdo/+SH4g0kmHhaz1wqeyYGMlzeYjRnNBAU3391guOqlB
x9kz3gqrDnfpc27Yyk82IVrzBhyTtLKyuLG0GqFCUzaXRaoag8Zm5a3Py8jOg5yxvKcwOeMA2mMa
AUaHaYGmsbm6G+Fi0XEKajyLcVp1VqqqdIJ0SsBcqsg9sJNbImQPOIlWs06gfYed06vqv/qwZ/MV
Gc1gluuG3fPM8UksBeyb5rD7Tgz5t+fTrTCcIgN9M9DeAc8AksffBA8ofsB91dJ0Ystqimj3nZgZ
h3H6C0pQVElvSlpoGD6GwHtMF+bmekXwJTXZT/vRwzgKO93oeyL0oGSNsMo8PhshU8l7j+QHNcBP
1RI6rM3zhq7ctwJj9+6HxIj4eoHQjmsJmYTlDK3YCPEP8tWXstL7IMTrVoXleeDtpeHHBE077LUI
n7Jhnar2hU1bBf8guAlVZluFcNfxsy/s8SgS5Yyi6z8Rsnmn+uCYzW54IAPCOE4K6QErMZerKBZt
3Jn/NbGSjP2Pf4iUOu1u44vCHF9eBuxRTmCM481dseGalL+pW1u3XdORpxPq7rXCP4/CtuOkVSrG
Ga9b41ODLEzUel0CqIGY4f05eEn3/hNvmZs6YO/VAOGf/yiVkPnbpcRUQAFCSeExvuySnm7xtjzw
HWcjboQjqFfkNcxw9psqWewhwTQ8JVvdMcT45HDsxWMkgIKHgfAN4iEBtlh+oOeDDoDHo6dKJdZy
7lyC5b9ypCY9s9Kpo7feRb5ZU5Owq2oE3Fyp0eOOEQc6eaJO24HYFXs/sy4H+vR3qFx/f9GWoeLD
pj9NkMhtFnXPwd0Wq5Z19saC0PDgG8ukGXhECNVFHRTO3UIFibA0TqwdSN7C5EFdNr5RJsD4Om65
C0LSlLuB0PxV6mx2gSFz+7zCWB+uUfHGjdTcOs36YJdHDToYlcg4AUzqx2OEpdYpIXknfKnhDeDq
syX87A1Mtsq3VUrQg65AI+rc/GMHy0Fpwjqw3gKXUOHhOHKBYTeN26bAhYuakiByImrbXosIZUiU
O6E5eKyv4tpuS6D9YsoX7eB44Ix2P3FLOsWVjwEnNK8RyCfBthnk4dVQFUW/e9SYt9ZijcZxRnEg
5dnHx2zCkrL888izDRkbofJBCoIiA2dGsWtW8Q7L5mgwWxAm6TldCD03rBoHbE1Ml8BvvQCLM5/K
wxWYeG1jBjEkX3bGOBxQBjXzq+xUBIC/jN2ZmEaSz3JcLZdeo8e/boJP4cKtCSha4VWaQOR8HAIm
lfOQ0rH2CWE6X1tM2vwUWDzsy0nLVo/CM7HNO1TpeB1Nnw2QsY3fxj9yQv05VySfq4NznvINWKI6
tUH0zF6Ow8NagGglMWn9dM2kmVTCqiFKJ8lj0aJrUcbfdZx1fUnyYaroCHIYl34tTJl7sBHWaKJ8
5gw+4co9+oVUplBBncF905UkTBv4yKp5GoN1EzsUBsJyYeX8kcEQiWsNqXlYMZnPs0jgz09xIRJK
660xT58nuHvjH7DgdCb8ZiJToXL82vP74nNXheHX+jAsR6f6gk3NkmFQkVsOd48qal30Ow9bumtC
/G7VWC9WmJnlNFM68WsjKZPvNEX6ongDoqEMtnOb01TK6s2jS/+clkPQ3J4d398s4PO6lTk047VL
4LBtsb1XaXwNHkC3LulOac04G/2KxBYGTqylMYFmtHwuiwPpC+fVNmHTuHpvr8CvUG/Ogy0gpCGD
5XYKY+tdfHU8rwWAy6DsjCLn6XIO2zDbp+6/IUHX9XzFKqbwMVhDU9HCI2ROrWkAWb+3MWCnm2EX
rTyp7AL7sdqfjxJ6SCPbObkxpeiS5O+heng+t3oXWoURtd6I6/jzIwmzrk+4ad2dZxHTv/3AcGY4
DmyUy3JpBDAW9Gd1LR87Ovoojz2qnYIlfzQTajo8+rtIMmx/HDnAYnWFRUwg+F6pWgwvz9LXVZ9n
NweUPu7PHGyE0KvIjLqYpYUddBhZaHNd6MBJX7WMmWRHdkF2si0xRUSloUllju0VebHKClglnwUB
E0tuHAlMu3B7Et5WhfFl8cHR+BMZiSlu8JRlwtwhszNW8iiSVDS7qIFxZ3tPYinAJnKyNZIF+twg
GVEMqPpfMpkQNkrCmpZX+EvEIFoUuFQIX3qlqy7hEepZnpSyi8Yg1JDiMSvdDCPBvKGV4c+WPg/y
KGTU+7Nw9pAh66ZuMspyaqoJEdZ2BpuGocIfK9NI1+KBeZUM426glxduB35HDOBe5vaDb6mnJA+K
vLW3hhcIjID4SJsOW1pUbEK/KIt9epqVJLcpxDQT42hwqxAm/wSIB9g/0/RGTTNJO1xVvSI3ujm8
si1/SfO6hrqg7qLGp9NkJANcfIBULCCW6aM9e7ExCMDxWf+mswRDFHlo61Nl5YPzSmu5ItRY7ZgD
T8RaklfhffLjOB4y1uUvhYhHhbVGS4eZPJbRrM7H2gab8VpcVCCYthqcTCIafxqSHPc6E/g3st1K
5PIGJrr+r+uHMWV2Uu/j3TSb3mKoyPPYteGxNB2/jquB6XA/LWMIkSzzGocvdaTnGiWtL6WFQx7r
JaB1KsLzOyIvv4BP8ODF7aoxatJmQpsOWps/Bl3cczQaDV9iZRS5i1IGWX0JgX5lthQIbCMj60zq
Rr2A/zlFdW+sfpv9xVIwnlL3PzLDhbk6NWLjqAleMV8PxIsENjSddjXbW9HqJEtapSP+JgS/Id9L
Fv14wN/hbh2y5OUwf9fZ/D+n3uQntDnX/o43g8HPWcZpMfQluXp625nq2Opoh0m+vIUHm9lbZTBk
9TeIZwGT1SXFL46LV/MkdpCzc39sbeFFwX4i98nFJ93ruveub73wjDCSyJccH5GDT3p0joo6lR6r
vpb6E9ZgMxvNt1Fij6bDwQyXcFtd31rUD/DWJB6vb0zHa6XWFzrEXhCNTj50NpEwmnb7JBP/fRNt
mdJ7VFHArBYo56AmH3JbtgP+mf8NlYwPgXSVcv004PT+RjWWFNkC0TzwO417sxlwaETaUL50LLH+
a7AVqs4DxPWpThkiJ1HOuFyU6232vKMC5gLtkslhyaWwx6+JwGHKqsj6pm0wtc0Rl83sb0+OIBZk
HygFr2/3+w2PBpCzrd9bbcSON58agFTenfPFspeqvxzDqNNEml2s81C6CUHMbD6O1TXqwdrh9QI5
gh4no6/KzxT0J9SUwfIUigrWiJ3nDOKcy9quoeByU9LRyrnOlOyyMKk1MKLp01TsPvzLSwZ6T8nc
hkziIxGUZIRjaCFxIixkHEwExPTNTf7gcui6mPHPSLAioFYJObSahF1hPYxlrb9Gw7j7YzlfHcA7
cDarRYh7bw+zMyva++sa2EATXnS2S++KAv7HFRTdaztQu7S1wjj0+8moTqGP2imRGwrUUCCWj7cD
jlw5I790GBKcD8eUgwQiVBwTz8W5ZeK+acx+oOP5khzpy54XkRuxXk0lEkcoY5K4VyA1iaS/sjUd
zKRaCfkXJph8a2xX5TURMNUH6SlEJWwMwZVl0OqIoxxziPEiEg/vZbmFT98Tjo9kFt40Eb13Vdy9
AuslanZYivdgRIptve3nlFfFPRjkVeRpmvVrQyrXSyu/gFl+yqpaeaAbjmdd5ZLYElZnalj+rOXL
fLKlX0H1FFhAzeamYeyJlNOb/mwR19WpQtAkrhhuxH3ySbFcMRbzq/xkZrIMjiAoDQOPfX3jCzJI
NLqJHyTRZtleEMCW6CsIBzKiSEjVTBCrCslvNODClR3Acdznzli8YklYv0L7g/Jht7A4D2KjdXCV
7d4fLPqqd5Vz9DVBksmxiBG/oz3j75y1TGiEiRr1FmY4GHkE/eFIgzjGC2eFe8XYV/kzidYoIuYg
X+QXQX0LZ4ZEL3KTCrzinqn0lAOd27RM71moo8nmNYfS7FDd1BqHHdLBhGeyBgI5tmeM7iRZrmGP
cE5q7nWX9/dRLpur9DPhLe/mx+1lhrxoZEjLPww34q7Q08hG1ZiZHllnQdRB9fmu2MersnUhrEtK
ZTtoccq/fIeBkiu9lQgDyBMWJYXjvm9wb+IZ6FCwiuXxhY3PXdt16h4xGViqad5moU7PaorQqnNE
5i+2EC85Vuv+Am262Vy/sxlMElcykR+PMiO0xGGCXg0kKgZttEZJK+GUuxTXWxA4382UdlxSW3yV
14JKcUYAgsAkP48aYC30gxATzLE4rbdWxLuxGrDMQi0JnVDqn8tepzWO0trOyBSSW5xhaTsOki2R
H4ymcRblhVQWx9oYN5yAPfTcfGEVnT76LDKBGUzgZcOrDGTAGM6onM2O//iO9WS/1zE58kVMfZsO
argGQ2cLFbeGzGw3HmaeArPQn5mmMkmiWV0SU35Ml3QjygA2R5Kse3k7ZOscyExfoJtof7c4YYin
C2JZbHTWCsQ2LlynjJ8iINOZSfEMiKsZ/aHLlkI8pybd76J9djJYFuY8f7RuRGmhg+yVmI2xovLO
9MZeShLxvvnCLbHfOjZgDy0TXXcAtiMkv7hrwGzcu3lHeC982fyUrB7QmQKS8GqpQRxJAodq/jBy
6D+tjiIpWQDGTrU35SkjWuKxbU7N2wFRpH4c/ct5a2FCdFz6ZNKnbSA2cQXaP6pI/7zDJCoEB/Q1
d1h1fEZXa1r5u1U2LVTYJmRdyED1EkXXXALa55msSWmuyLSNSXCmWHUfPdj25nDE2Lw3qVy8/7ni
jP4f7ZmJKE+wvRHLeeqH07BUauXYSJ7WUMDNQilHmghPWzKzuZB1BYelMrjWoNtay5FvTZjkOGjh
HomOAhp34dvPLYklEuql3YnUp9Aan69XLsAzWoFolopMmh9yjJGrVP6qm4iZRRcwGkjme33orxsm
Tix6pvtrmtot6v8945omSXVkqLqZhdEtmeMj0V5XKDgi9V75jUEcb2s7TBWupuQj9ApXdGgbKlaw
wSg0Pa0VFqz1r4OeVqhAPOG7RkNVKYId+4MR9r4sceEOZuLwYHUXqA9NxBfP92/nNWzxHEVZWOeG
f2Yazc/xJQG1mdgP4AUetoOTOZmctk3rhydzX/xpt9TzA7i8lXyfMaVzvRLKFH17eJRXCAYDUY1W
yrxQW5+clpUsg2llF1lmdFuiCB9W62AqQiqbtWYOpMTgoC3OGtdiftJvEuR5EW7kKEekI6PH7NqM
FdBFVRnhmCoKnDfoQZjHBOeaG11bQyBqToVexeQp1G2XkMsrhT7ZuUSun8ZvRrj9PYsoXVaQ9g13
6kjbApc6HggRbt0Bij4z4x04+v4hQV9SNuqx5+d/bDQ9P+Bg0PswPCESAUeSIvlQwxnBxsNJEbnA
uGN1xcX/g0J07R7ubGD1EdyVTwRcpbUnxwf8XjUuVdxThiwT9PaDUmZhFJcRJbi/YlJ/iV0JEOJh
ni8WL8+6fF8XZ4pTpste+1874cBs5V/D6DvGhwMOMXBXDF4pIZQ+YTaWfNDmUFk+d8CmnTena3QW
w4rSBUxSktjlcLA2skgAe3A5v1aBPq7nBYubhLGKgJu7a+O1PLkrxaX/G4tlIFcWzlwncdfl2JCr
ibB3wnCTWW9vxBIZppxmOQIfhNzVr3f+jnZZSFWECVRrRIyH6+Rz85p9HZn+d846gKa4c3sP03rT
ZKe7t5tB4CLn3zqPtd/AoGKM5+0vRzl37vSybcjEXV8BTkuAKHps9LS+KBWqihsv2b0a0VOTO6GB
ZOxRClXRgHqfUNoDKUnHhoNJzj+KSDiF3oxA81QqJJ4IX5RoihXBkB/NN3cejk/4rpytYN3VUrCZ
G6uj+0+XhwHTUSokC3vUiSH/VjC4GmG0oTEuSED9O/HlJu40mWv0MEkgan36X5v+eKHj5sTjszn1
du1709HhApAuXIcw2qWHzYJu+hokA+yYxg8LbW5awT2k19g4jRR16L468VvT5z6w6sZRed+RhqlC
Y5Vs9Mi55EdLmn1vZF+KpwdVGOWlmfVn2cggkp9fg0bkLhkBMO4/AvTAvBotoIfcOJQ7MilYA5l2
WNbXx64JFeZUxOkZpNAQ3IZ3ykmwtA0s6PKMBLUIxWxVhNY5KSWVEiFSM9G2s3QJaQE9I+ZWPYfE
uiudDFOTlA7TGQCl6Ji6AtGsduDx64tMKkVpg4njvrbjVetZKBVrFCVKYtbfZil4+GaVJ9NzwzWB
7lITXnbOLQmAqRg3ZtbftlpaHB6PLzauwD3OhcyA0aIm5ucYY33nlADjZAFXwKc2yKFZJR+6ZTiK
+Vw0hxLtvcETJQArEn9hVFD1mnhy8AbdJcomkRCec5FUc0TpEYhOkUZjGtkuKMg375b9yg4twpgj
Yr413CFLVc2nLUhuaQzHpcJxoCl7HBBwzJtmQ5te244Hwg0UhgGUxW5I/iQLi34cZzO6f7zi6DUz
yQh8UWK1j41tLXjHWmPLKnvlfDz75XGZs3WjS0WAiFHETua7kaO6g8VQb79bECb8IsPZ8z02P0vl
ERHBLG32kD/oEA/rglw80upftFxktTPZfdrLdkx0217DPgWzNEFi/SMA4clu7fdkpwjRJ14Y/0eN
/8OWsv7l3OjQkc202t07wMfJtYdc3K4baR2c4RBpcAAk0Tn+0tm9oOrQXxJs+jzKYFhzM0grSwUq
bEMNce5j9O1CQK9vtWktaYW+RzG+Itel2uJGHrkM9hkgmDAx0EpGc4dgbVCfVpx6xiAE/QQUl0Yq
qbhQ4EaqH325xbkSBXiwcNWgMKdDaE/B5AqoBMe2duvhjaeVCB3A4w5UMd6JXzTOUSp+75yJiJpc
tzJFYaodJWPavuujWwLpH8wul7LiylxCKLyhpsAdCBXlctdGTnWnKy8VAOV2lrIzuBvPNDmuEE+D
M7rsW49VacEHV+62q0butieHTTu0y+lt/9CEPbZ1EhWe4RCc0pyj9SNaAYaqWCmyf8wa8dNwfjzH
5YD0kTeadaBUb2Rqm29hXXB3vhHSbIh0Xp2qI89EG1M5bhp6b3mc6a8LNgDYRkwjjZMhZBEMCmc3
W6V7zFbrORZEP4QAoVKA4cdO0DCVH3y6ck4ZENkyRhs69syq27tyEETQucafV4/n+cEpDIzany6j
Mci4etXx5Nu8QDyC7jUGaTt2JvAHZQ+ndB142zJ0iQAgRMANis9Z3ixJ3LRxwr8iZU64tgII2k1P
muncFBimhMNofrjYu84I7K22zQ69+QluAhtmA4I83Y0/D8rbl5x+Oz7yLC+AFPesIO0Fo15WWEVR
gQKCfNdfr82Fa2AWULz7wwFileGaySIcT7HgAo7WkmbhqdXo6MqLfmc2NWy5hj5hPuTT/ucAD3Ii
o60yj0VOIRnIITgzGh6humpxcosbj64JAMPCbEAxKEtpUhzQQOga1blP3PS8h5QF5kREqQX0jVyS
qbq38fwXjH7jB2ieWx9AjLIXg7e7oRz0/LMzhyC4B/BtuUMIOMGSEE8R3jSDJ0Fhz5sOkfrlO4bl
CUsVhENRHrZvnCXsfMHVnrDGVDROn3XOy9PgLej9fD6IObuJs5qSLeTVwY0yumb9NTHA2FKCtH82
jjNKyW9dqRBxtrKPIRHBgoondneKOlyks5Z7vapF/HCyX8vr4+1sOx4YQ3ktrd0RU1CNF4nNHZ9M
IEZGthonCISNk5R9VUkJvkd4IzvVLRVeTUPJk64eFLjZKt0fZETghsHqgPspFESZWw+hFaFcvyqO
u5q/x9VKBXs2CqrA46rUA8QADGDit2L2YIX1n4moeq3AxMzOSicHquXSAzNnwv7687pYp2qrbhDJ
to55Axi/luPwj/3jjZ2VqctUCd8mh0l+X8r7z3MbsjCA5jO7dkjWDYepDGLh3jn4l5EWI1UjAA4w
p5anuQIPT9EW9+uGbQ5m7U66i+TSU9rmatbOvnuHrT67yjzwwwHuSfO1OivMKNmWBS4JPj+IVZ42
NtzIEvsIJ2pYBslzxTpfVaRbDFmVDhyFWw0ZnhBLHMnDJkcZ2Ed0uwRru39P2IK6xmtFzkmOZm5x
lfJ4buCUl7jyVDlePzamvXkcUVJRo3SZjFy64H4Decem7Q3PJWWx93iTc/GA0gsWcuxYkagIUi74
Ntboe7O53p5yxjbd9ChCRBnDGTpUWYfXykVPxaWJYx6UVhy05FGq3X0k1H8xsdoiKT5U8ahZ8uNR
637eTQiS+M9i/htFUBJmnCY2m2yRdumU3Loqxxx/M5QEFNPLySrljK+q2U7jhGainEd489WNuean
RssxmJVB0kJW1FE8eWP5R7i1wE1mx+TmJRMGQaXn/2AFddBTHAdDTDvX7ZvWVTBmz1b9F5gJb5Ij
+VSPuv+N40xo4abgdoK0Fv0007uWFZ4tLHx9/oi7EszPu8QUdScmZ7A0S5mW3J8fwwSPgFESWt05
y/blPjAaHzMmbN+c6t7onS/IqDx7EuTAr+MfqhD/lB4lvSlDAA8vIz3evVIrwAx7VkOD3G/2JHJU
VA2GMgDqdw94nJgwLuy7T7MC5N0CHzgg4hWBkq6CJCXnTWiCelPRzBUa6GH0zw2WWnFqhuEvMpkU
3hAsPFu+n6BfZO7nJKNkkqDwyROTLSDVDOAijcKJ3qbS5kernvVjS3a2H3ngjayka8csubEZwtlR
W22+fsz5ScJdWgdMhUJITZXoVKU98kltF3tFGbCNO+Vj2d0cVg6YWrncNnjxh9yIoEYCeF8BO+77
eU3FIuBArM76wW8zaxv7MPdKaUS8Je19bTFTuTgvZsY0TiNFBQB1w43SSNN5oPX89WwFVIR6SYly
uoAhLmn20qmEZWdQrPyz9iz7aPRSGSg+h41PHnJvCKgTOZvCv+XOcqvltpogMImhJWtLu99OwZJ7
M3KNs+15AZsWbL7rgDrzU6wwBEpx90JzbmcsT6jceYj9ygJJa8+GJ+OWj5/ZI2/zIDHPgVNQmFoJ
OfWnmwjL0Fi0aWkPKMIz0xE9WE2nUZINLWGLKQCU1xIeWV6JQTGIExmu8SSyA1tfA2Bs7IQcqtCm
K/CxAUs15jrDLP+gwL0HpMOXC4+uF0/d8mesviUHjzP4iFiqnmB16Fwxb1S3JgJmpbmiDPCSQpwX
1z0xaibXvmVXcfq4vYFrXvLYigZM3ttbUvCn84sGTe5Qmamusxf4K/6h5EOlfhPtz+YCeIBosl0I
Bhuxw1jqnwlYNRCpYEJ74Pg61f7Mir0dZJbAm5tSJkicXPA370ompnv8mqEg/vpvXTeOWhJL0Yqj
7OS6twQUY3QYrg93z+5CQxROc++ReKGlqsksqAOrLdJOqJZJwXVpb94J80B0ogEoHbgP7SPC5Z2U
EEFC7e5yCOPJ/E+ATMlLKkkW9OzD+D0cSwkFh9SF8Y8b6CgETUklMQFGvgIymT/+736d+6VBJ/uo
gF9ZBkU6m2mgOAARJcgIpZEEKOFrLinaZ5MEzWoyZDqgYbTdi2j2lu1lpVEKlF8Z1kf5d+3ir3af
uSLwXxzagXYdSlfdr5/a/7zt0mywIW1msYZituQjhv9xK9i25TXbQ/QbRApW19t6TPViHTdhgYK1
rXIoPxZL7nEMWZx7HkZWzQi7iWcBB0qSLMpMZzUCNY32v6duH4EBdqO/9OXLXHAOimIZs0qhBFZm
TydY875t541r7BBjGwoKMAR1lfS0ePvdP8jIN+xCjZlgLHFodgFl7rV08owOnPN6DH1EVOnx2DRP
Fs3vMNcmYFjghFZ0KtLkHQ96XLhgWdoJYGg2FXiZZCZSyN2rBLLewFdcoK4UMxOyzZhoVGS3Qd31
G0DzztOdtEWrohIHwHFqBVHd0aifgj7OZDO5bcXdnkMSaZf4C96gBXNx8OMNJawpRfzHk9QK3OJP
KtGzDiz06GWOKfBw1tyDIkU/1Z4PUeS6DLW7waXpMA8HOVAjDaOrIx3YojYCLJ0qvy7NdezEJRI2
gE8b8p4tcFiH02eQlsm2HQkGRekZOYnb1qICOwmwOYaiWBhdh1JlB8e0SlUvfexojv/MhScWqSe3
ZTdkO7NhrxY82aSe0HHizd1mBLOUtc0rArrAgpheNnP29kZYjHbPaN4q54Kr18Z2tI8WYLz88htG
RJH0UBzv5X7WFQPaNcgvv0Xn6WmgefkT9iv9pzIwaQK+burJLAbyMqneetlEjWmr5k68+MXDzSN5
Qhvy9KEyVwPDwkyhzxLq2Qwd9OWmeL9nF7WqgVPCl23a4AGJLsdSQskCA6haHhq9l7zo1xLBvIyv
2Uv2UU6sZdc5Sgj5aYePlsnfhenuq+7zTDHfTGpllEbjFkTod66niRcyP7QHZAmIT39d4wLVS6sT
plPKdW0K/OC7iYS8/LD12cA1H7v+624FqMmN6q+K0qmMdXxc4oLRH5PMoHiE4Drftz7zofWuhIOA
Bh8f8nW80zm+4QjMi8nmZ6ZcEZmD0ULHqRP0cA54wQwbOfSo0mkh3zwk4JFjOqdP0tFXexgavcI8
IzToshCZcgAEr+fMTYzrU+65eiSzH77acmIIP8JeqAC3ddsST881C4YGLC43xVXoPzfhqPMnth/R
IKWIANIJkYM3RDaooHrTqxdP71BSzsf53jY+CPouG2Q9qxO7lYXmC7Tub1AC22pYHifJjwLrTRR9
LTviexLpB6/uRKWHovV8sdTKaP4OvNpI3C+mZ68BZMJbE2hobWR2hyr8f1gR+pafsX/dt7If2v6P
5H7sPb3PX2hlfMlFIJTUhB5bzDPjTXlef+3MIAz78mZHZA9a/6Md++cAXx3WXaXq2hgkB9wZcjM3
O4K2fo82r7mfGVDpGbiYhUIzI8dQtrZ67XLHEPdHCIx/7D885A1heF0ms3YV7/ypF5W2Si6Fkji1
gU3cyaLDlaJwDqGyGITcv4STp+1d/Xz50jnW8Z78pQBpMTnbQSmbUbzgeHThMJLlMOYXMIVIk+pW
t8WQkGkQq6NP/YWbUCuL85OfbkuozYUl46pG0PIOqwvPbQDdOiwtbb0/GsH1iCDZEg+sMbeqRq9D
DBFtXTdaART4LPfEPlID/i+cVWbpW1W1pqdvjzzz+GXyn8oHJ3tyZLKLXom/8lvfXwt5saEJQrtP
DreKfR7fbdkI6U6hu/502HdLEYP0lHiF4GKJUJo0R3Gga8KeOlpY4mXj/PxXmj2pBzuBwG9O7j1n
pPYpTat6qsO47lBSH5i++rj1B7ZzcZNgkhQfQXehGxVKtWiZsgkdfNGYjJJDGQqCEWHV3ZcWn6e5
EHQ+YyNzrt0uWAXdOqu6u6ucAGSeuet+kTd4+/LIdULFjOLRhL4RDhSMeFWB5WzwsdL24zCCCMq3
bsrrxsUNcV7XiLHHCZ95/LzePZMgEYGSJcadTRy63RmlIYj97kft3G/8GAhEao6YFYgBP77jOrPt
Ln57yQP/cr5uWArwGIfHao4vBH98EqPfj3TU8stEXpDeWVIh+zN0bs/n7GQVeUr7oGycpyf60aQ2
CWbXhXgK4RYv7ndheU9x4yll0ZlntZkt/sNIeRc9mHggRQojP9KzfqXp8Q+WXyHOP4AOZ2zrLcuB
WVaVXQi2yXWEZTcpHJkSXCo1D1QQrRNJPpaUbBfmR+NfBvGl9g3FHZT+NNj3ZgPa74TqLnVxCbwu
2E8PMqh+M7XqOvFfCWVEF8HVBlxEOgt6/ssMoT/UAqLoBPJwErw2pxahY87CcblYVY9bOi+u+oai
w/cM0s5hlC6yK4i6i+FNYimwIPZXx15XhOqOMySxIYXBT2mWLtLyFQyilI3VFctWBPzjCX5HLo4c
08FVhnDSg2veufFTLIdj1VW5JtzfZGRMhhqBVqcpemxdPCpoJFCH4SKoisOxOcBxGJFFLSrlitIl
caMQk9NPWOnLGHyZmza3s4WxPD/1wMc8H2Qk5997mc2pGXIQFVXTc2IeMNwIrWt+FsvyB917Ru0p
0/x/dl8ftkCLR+NIRUbgANhLzMBonOdo0KDyow0IHMdwxg+Pva/m7tzDOXb5EK9BjMuCBorRTUDU
RtVfh7nFmE/AbirGzmCx1l4vMhyGmVXrowi3VuJEpyNRujl0fU8DcZD8++V5H4OqbfflmJ3d53Jn
95m6WUheECLA7Jqj25cpF4ep3YKojs0uXFUfpoV1ZIEFsdr7BG6+0WW6xVJtU2ll21XHw26rsLji
mxJ/u5KO4P0Uh7FDHgT1BX5uxyvqzn+Xlf+cSZ2DADxAEyUgg0pVmNi3WMOBBHuHbeKaHE8ND7Hz
NYdOtTwonoaguoqx0He4gBDeHJ/G8h/pIlvkjTkOy5sueZ0oxMD/6QHFPfpSJywwuieJiOjXUTae
JPFvA6ld6c8hfSWUwxbUq+mPBFufDUu5Afzyv6qrgS0ix/6Tj40xLORjs/jkQaf3mXtScRomdGxk
JdzhZzbUj9C42bhs19REHs5p2Roe0SDToG3vqAXfmjKHGZ2lbbyEMD2YbHGugeTyydt5elMoUx5v
Av5jmNMS1mkw07HaEOyweZrJN+Ts01P6OzE+pjibYuQeXrgEpBOd/acKoFRtv4ZchtJjr2SdHFr3
i3IgXqZ9YMLBuFQyVxGL6ZbaUvF4poq2lgJCa6yeIHbTCsaySAI+bnHMWVgsMjJqZcZM713OvOPy
+3FQpFcYa9pxBOBa8gl6rxV4DzRS4mN8mkOncImfQ4EKwu6Xoj4HGlDHsxMJsKP2VUbyU1Teksxk
iv/0GLmIWONjVHgaRZ/HJ8+xbT8sjkm7D9Sk18txf3dY0pw95vigE3Xdf1I+aiwWv/6Z95leIcfb
cNJPdR+LNMLe/aSW1NshVpulczneH3Iz0QwvFBf3TzmUyheS1BT47kChY1zqtZEQIt0gMKfFZoh/
SNzOsYbpsTj6JlR1R+5D4cPY9UM3OWnECIlHTAZ+rt95ogl3qhl116LzaU67+hNl5iVOozNVf6Tt
8ZjTI5xVtsxjKRS+pBJYf/71rwfHk+jk7PjyDol4fd/SRBorPdrPzKSjaVW5c6LfqBquR/1iQ8YF
CfzaHrK7L6ozooXXiyZTmmPRKLEr7n0ckaKFbZ3VTNfugm2UfR8Dnudnu3dDNlZY03kKMmZuNoO7
CPDpCYjkhMRy+lbVZNHH1ScH46bcv+pVrqPq4hMyhlMP434XuHjsnLC6rkk3jLk2MBCoQt+nnzj3
TZMM//3p9f2aPsk1GQITjZQPP0YU9E+e9uoQhE7B9hwouEarxaPtZfPWqxBJXl75/R6EDJNCjCU6
W1UAIFiABSyB43TQ854tyMv1mqijXjPlMUNQTyoh0YLZbeNrYilqh3OCcA85tyHANl+Tv96bf7a4
gwzEBpeminONa+HehmHLE+nFNQf2A/fafr8GXpYdjY+E33uhdSwxOaO5DJUYSmo+zw7u1aixc2TD
EB1Q1ZHAW2oDGVf2NlN4aYZh2IcVuR0XY3Zj3ayb0ig4ZW+hgDO9du3SL/gPWX046YZSptRCH17D
VmO1XsxEpcnCN4IrpOuDMbz7UppWOatG+c03a/n84R09wwM97PmqyAvZ2DEedKKt07I0QcjeZ0Dx
pRcl4a58uErvpR/dZLVWPFAEM+vsFz8j/82vqH4+KNzMZj890HVc2Hkfn/aPo6U/uTbO3XJCdqOR
Qi0CXSf7/3Riacv/ZR/BA9Tr4snp6rcqLxNKdMhlYGmM9R33NFbZhogSkPn2dPPjttfkE28tt6zN
lEjDNE/i3nX8gJCgF3w2vaUP/plCdlkkq6oQluVXg0S9AHJ56//5aKk4JE3NfTGBqURGVi2a92ZQ
lhonZjXT2olDPjaNc/uwgM0k1NxFUMskcIjS6X/1X254dFgx/xZEylF0pNfsUsGjqPhLZO8/Q/eN
+mPmx+fTZCN2LwL3R889CQocayzSYclJmvNnP8vChiGJ/9H6YWCTdUnHjMGgV3+uVgOLyEOi/Hl5
Xad+TWDIUY2iHzsC2btsQYcmvgNAY2WBkEA8IlY5T1xuRwduaGuHaLe2HYW1FdKxZcikZMC9S4z/
zqZeGlTrdJkJZAGDdUGYJc0JF/IgD3Puw8h++2VqWmdprAAoDxKnydtWVlyXu8Sw1X1CnJ+q11S0
/SjIDTj7IgdbqTvI8tks5SOzNNPlU3KQ+5Zuuihonah3yuJ9GKBHBJODK5iAMODREtPJeUMoRNFI
1sKxCVYFXLemGVzeOp1eb/SpIq0I8o6KPkB39uplffd6l+WzlGC8kBECOSyvf3V+CQczb0qC0KNV
ju7DRKu9tbrGWlP0wHTESNgWP7VD6QnYbZMFyihwU9mqcunr1iIUcQQNok7RnDnOhfzrAB4RThpD
GcLEk+oZQNfFUI9R8ze9FxYCpRp10nHE7WzQd0tG5GwoeBPaiaToF9djRbrlWCTs53SVaACwV69T
l5Kzte9wtl3vARVX59cnaUqqnZC/V/a3uaEakPM3t44/FugRo6YQQWiD12JUZjLdQy6kfFrUcnsb
DHZL06XNPiMefKu/muF08gCpddlc14cHk0T8mI9QVUi0Xy7dqyul1Ra9j+zw6YQ8LWPpjco4E4Jl
I+/C6SDjfYudF1vVChTrsHV651+kQwa+GGqdMCuAJ796LXPAA56VbacbC6LLSN2zWS5ttnqPqtBd
sDAEHq4Uqrfsz6YTYSDyJi75o+l6OHsCfExL9C8fpMz0bbc/JtfxToRucqUmkLFHZOi3mOzsZM8F
8ONKTvQcDOJLMmJRypCDDTtnEtGQNDzFX4rIeieQWF1NfElFACGAe9JUFNehXKBTQyusyRUc2ALs
g4FyIPGKzJc0OfqBzTZoy8LhgipbcXr+sXkKLwK6IUYD3tlio3qfMzuvFL9OSmB219AXQe9XKQxk
RnvABMzi4EFmFySexWpjwuwaWiBnvHCwplDdkrXWL8NUDjxSNgQXHMiN+5HQKOUUhOKuzpLlutQa
nuLFCiNJKcjo+lC3tNx7jt/nmDJaYKP9LOkaoeTp1EruEqRbNgR207SAJ/b5RlchM+THoOTNdsiA
Sb+eVus5HyM3YEYBtW8nbYl6SgivPxAXI9cOJxF9lYZONi+O/xAQ6nDBp3VVwaCbAKAPxVjSfnpO
R+bDcmESrHiH44PeAo68QAV2BStnAK2lMjUCyMboNB0EJuMIlQfBAfx50OqQ39faviT58/TLWKPl
D5rGgUcN7Sy7Go15Pa4xIFJvXlUmHwi72t4UHBA6ZqThnlms6vQ1E/anQ7bFlA8Anap4jREOzrhr
Q8z4V7j/qQu3NgSXT3bSmxgezAjd/MvNORs7HboInzvWEuHwwM6I1BNzalBVVueM+FhL8HDp9jmm
cMKOu5Suw00Aj3Ts5sm0ldmNNFMP11tmmuTfr0VvPVWAKMC8JGrRWTTnxfy8FQZneVwHPVR1yToM
mN1hzcMGlKu2+HuHb7zjD7jHOFfyt6fni1JShS/jGi6hBVtigXQQcaGckPoa0lglKAHwtZ4q4FeN
ISTP6Y08CS6byJBhte3fyvSu1oOjzOtHLO0/HGagqIfIYO8/EOO+DUDWFdDMPu8hx3AGH41QRPz1
ybCGMHPZ3XwRLlW4gqrPqJUcXeZipjfs6lklRJELqdMJX/Sh4HRBuQ0cv/8kqAHn+HxDzPkFHeo7
pPMkHrg020cxw8ssroEKKBbzRxMK0eEBrHLJQvfmreB3YZ1qNoFZan6Bi0f9Kc7U94Bx9XnUMpnS
kbCGUgaKL6Pmz6WtY34eOa3sTWyfaBlPJLLKVEz5ymRJvKGFa3I4JDZ/U1s25a/9Ruq4pqIdB0Jn
mk+4FHREL3E7hrihyaVvn/CnHnI1d4xEX9TWKp5YdTvPnMFOoz+t3uLTQBl+12glsfRdI92GA4Uy
YMLbPHk8vkypz1QUpxufO1XdQKn1/UrchxI5p7C3kBWyYjp78gL1GX7cEuG9gzoV+kSo6Lj4mQhY
eiZUGbICUGHjqCTB4ieeEFWQBGQXcZjHQ1H6Zs+mhP9Klt8n89zC7Jk6EaOFqPGclpTE4hrQccD5
6v3kevO7LYr3pWOgoaCpFDokZtD55ZGQK+ODNEjVGdkJOhZ/nxLUmdD85GMbXkCqUzEhRobH0IMs
mG18gRKJ9N/xPBNPR26G525bgkEbbJrUZwJ/CBG2mwimTRRSDRbV3bnV3OOPSsFhg/6Tr5waN9Xw
GtSQ7BsOzv+4O4AWJqT3HmMLCbz2rA3XtGrd6m10w3mrypctNu9Rob/Jo9n7nNTHOaSbQxpEOr7r
vIK0Cu0/tnBX0nTDZS99HhwFc41YYU+XlBSzQ7hfhuglROn8rtbMFpLuPlb1GaU7IG3bx8NWLXaI
GQLJzVsV7lXFKnHCSUYXkvWU9/8YHN+iX0egJLDBrMV3mKDVGEY9s/9oBbN2bQc62DS9EPvZPo2d
c+FHd2g2q+YBRNF2hQZgWTRR9hxd2Ii4YwLqKatYSoBQULCUYzy4ANQOrWAt7XXjBLY8hJKSx3R9
o0kWie6Yv1uMucqTYqmU9M6l+1dp4ZdWcIKdP4+UHTh1RVX/So/8HFQnYhzuJoNtPqGOpJwWRF2Y
e4toZ3PmOGYqdw0pwipt1Qr661Ji7vBmUC974FTvu+hQghhpYVz6nFCq8JuM6Ce4nzhM9uVpMPdy
VgNs/K0Si/QiFkBHAwDd4qEAyAlTITmfom/PIyAwKhy6RdgVz7t1xe2cB7T60RBcqfNIx41S+jeu
+Pv7vHWEKqmuxV047KShs0G/Ek9aDim8VdzfrIsthr+w/B9UE+19r08H00Uha8XFKkdO9IH9v+GZ
XeBhz8mVe/0T6icFuCchEblXbNJker34o4dx0e5OvAoHdB8bIJtLApfNW9J2M7bxb3FAe+iACJg8
SC//y3ftHX/lZpQ/fL7te0mHjt9ASZz264e1DaDd0+HlmvheKQxz+J5uz4kvi0hUrgI6LbdZppbv
opt6Ya3EQcZMb8jYmmvlZPBZKc1PgmjtipR8r9G+kDbiFpYoZ/QoyWTQlVxOSTsfQDL/vT8hKzKn
Kl+4jh+HpmC2W7LLvtJOB4OznRPJD/fn1g7preQ4BLSMqq3gTSGZj5e4vl1JqC+Z6PeuTn0Q37Md
IGN+te/qmUb7FVQOEECqV/O5JzWn7XPBuvRro/UYKd3JdzIzLMp770vR2m62YqKJJ4majNBTUeTK
ESo9Dyip4+AYs6aoQcn0fmWzEQq3bGmSlP1mVcPk0zu3CkkgsxMRBXwx4PY5o2rt4WKzQOnhKtaG
OmDrSBiGkZSCViJBtUwU6/fWdXVWJL4fdMxqt7bfSkQjcPt63RDQL9NusZ5NnWfiTo8Usf9w/OQz
HIAvOLovn3FG8ZS1R1XAQaOA8kb0nxPEFZQnBOQ3k1iFCCcCPeSOunSz5KnrPEbLdsiCuLHsWtEm
2oxrZ39t18oP3oIGoADBNTY/8u5j6xefMMChdONJaJ/m7U/rtjeUuhf4DTRHpsFOvYI0rl9Ws9H1
x178WswLQSYsf+ea4YP2X9qU+2C5VcWt+vqVf5mVWm1CN3NqgXzyjQrIIZnNNKvW9PFmYGUAg37U
P5lCgf+/Xd5Fa7QN1gmB1t174HV3gnCNR8y3PwaMszdvrImUxdfEyBztVE8zlLLUHoeOceyiiWWv
QoPHU68x/VQmcSHNSZsRKNBmmplpIIgz620UyI+AQx7t8o3sYjiCq6vokZauhAZzpyvCXC9FHHLu
DhR4RPAv2SkW1HnKV9EKxmUyezjZaKdBD6+vZgMC9ZWrb2YBvwuKFVAK/oSZn/DI/4RpvT1Huu9T
hRberl1Q2zOpvqIpFIhjDWdLTwVDGqQaU2/TIllfTyM3GGDCyaIPEcGGnFOae4jIYUbIzGD1OqtX
X5/nKzl9edKQnsjq0Rgqqy1nCIwTZEvOHG/clzYTp95ATN958P89Nfk3ctn1LUkOl0dw4awmM69n
M8nl0Rdhz7XvXbq/Nje90y/gjV5QCeGUHjgd3GDPxsKAfTZPodWr+2EYDnsjERNzDU0GuZHb99jC
vw9tE3yFjvKUxGRm7rCGnEpArUIeVHYl80Jg2O+UdjEBDG5hUAyuqB+2lEYppEwA9WHqaSRmb1lV
woZOH7UkBXtNFj6iNiT+L4G7iYerzaq7h0fxpYyk0a+Sddi+6rpe/MWJ9g5a3Z5aIKZ1HKOt7RDq
w93t/RgdMARdlLMDmtKzHbAhnMuZX2e68eQ1l7/5wno38DHxTWj/odQoeLaDuI9u7hKpkwMu4kex
7Oc4ORrbOX+u6Wy4Xx81bZ5jNX7VLXhTvKUTHA2CS176XFJsQkGgjsMdwzwyv9zKlPH/gowPqTKT
a27314lnVSzOO1WWqP5f9tQ5OLy0ZRQjKKr18LykNTGZSbiu0xPO2kevbQ4fdD3TEAjf80xu17Ao
mPOtMa5sTvdWwyafWDGj+mG3B1pfNCxNP/CajxhfSCyV8UaFSKrGH2oRJJIVUk2+GU5Du7Sax9N+
wgowb3jz9f6z3jn+G5qBpLKQPoQOuQYhLoHQLlIVCUVaOFBthQfkuElppLXGkLR7zch2CaSF4BSc
QVRqtw3y5qefTmSG0dwv0GdXHQkypNlOiuh/lBBe+8Q2OURsnqPxMBL3WvY6vfZ+/z7VuDEaIn69
AVziU7Pbt92S80yGbH1rDy0nklW1xEO8vMqGgWdCa6/WiVD3i3VuITwNHX/M/TjfeOPJqu8B1+WS
d50X+/P9FF1sHLnbO7azRDvNdGUit1yJgBo0WHgceJvTqWQgJOiGfnntSFW48fcKAmDDQU00tQyS
uVTtG3bDEdoFbeS0nVAUUGXfT2SUEfYb6u/AiwWjyFdjeNFNfdtBnFi1MOXvN8VWmIDkCzYhpZ+u
xkhmwU61zzshkQECzXQsJiw9NANWY571eD+GgZryI8F7KO429tdFkFhkLo8CrU3qK1yb1bCWyO//
IvTtbycPkYa9D6mVLnuwHBLYjMexKSD/CsxUUFwJQI+UWMX0kedHeRLPbhqEQSbIChLRAYm5pFdj
be/YeETsR5E60or8l0gl70Yhh1fJOxqtMhUmvJzTB955UXb6pjB+mv17bBbbhw+/RfnTvMSSOiYG
s7BISScuC3T6ZV7Ftrz4b1wFCYA+64I6YXKPLK2buVkw/KWPUq90JZzKB675RdbK57Wq+JozTJ+4
jZA0a9kzInIQV/DejX/nOfsTC9qUuqltjJZrzMI0rftr7H5DxjX1l29xmVk+4QT1J+DCOwudx4fn
91YK36IxKj5CpP+nKOFC3edKge4/dhAdBAqmq6lOqRc9Us95lQ821Mtk0R+CFvZv6bkDksG+lnoi
do7KB4BwzAUCJDAApGsg9KtTIIU8zV28LQ+hFS4FVC1YrF4/qhAVmjgg6INZtJs1CBxCkmFjZ109
BBl40KmPAi74m436d7/ATSa4w1VSsUrOZZlnHeEwc2B3zCiLbR1akJp+4UA35QqrLYNBgO94rA1v
TQHXjnZnmT/Tszf4pMqnMY+P4AnYk+M3VaZeOHILXVWV0UNQl5YhXsVZpvL6abwLNuYq9VxHAC4L
eCAIBfQgvYri2i5jRsjwhiRDPyhnhRJRB8Efm3VUVAPoAc/6oJpESXFX8XXcRyBy8Jc7rx9RJ2aD
V288ERpx0m47lS0lZfXaecBqYKHHVP+Ts98z6Yi5Bzta0T/CJwN9jdUMtICr4XbCcHIqke4r2Xrq
Ock6tgMvzUsPoBs69A4nrT9LAWzrBb9J+vaILEKbgGRDNrNBb5SWhP0neUiDMe0E3byw/BheSv3d
QUyyV4yySveQqGMGb4nbs1AFUW83zX4ljezR6ViWMmpUUO6RMuJTyHYJ1yt/CzHQUg9mtOspw2+T
3DWfoREWli+0zrYMm+qglducrSkoMpAOjKtDCal7R4TQLJr41u3duvGrKW6uilAOYZ3BiF2bQryY
koNm4QbkU0fB4Rjl86lwMFDz+xZ0v4IetXYs8kkW+z7qfTWuWL4ncwc0htHEcRMWSYGuU35QIqam
GLrX2gIdvTK1A3ssnEOOD+qtK0yBh3PH5AghUSdlokk/0cyaJOGPJE/TQsd5WFzxNc/ofQZwGrwp
eOTvV3v5MfMeUFXWdTumAuOJhaH3lhO627/iCxn3IOYHBVzyk3ZlxwTPhs6CAn1OzbF4h6JXJfDP
3UZkXsQl970SWikEurz5KjYc4syOhW26dmzJX7dcVGr6reQPsV1d2eJ+vIadGyu03+Gi/Q5A2tUX
IbNJ0cqqopU+53/Vno5kMA4PFwpNj05zYk4DRxNsNMQ9OnCSFzdpcmdWX1NplQK9VHsqA3L/4bU6
GtM5VeV4kcry/0V9N58a4uYmXr3LlJHclIqFib+okzx+8VuhFFA//QffWMxRQLrH2FPQSpG6KZdK
svJX/MTDOo2LZk/3XY52ytrLTwQ2U9Vu8qariIQYl8aCfYMd6saNxSe6blGwFKRsEffafE45vDwj
SnFeEMaq4s4U1PMK8el/bUytV6X/OvPzc+rSNHfImauOgzkW+mT+Elzb4gL1QXtc4pDP+vDNOnTD
bLxBdrHB1xiGfa9qPIBP2e41RqDT0t246Yz09PdlCoBRS3zgoOEiAi4uIGtKg1/Q5s68CVm6Sa5y
jwUfJBR+dBN/PVm6wUswCWvW7gt8QjDlhcZnUIQ0ks5eZ6S2NjZRAwG0/oYbvp9VlsYVeQvLVtBZ
qMjjbYu+96XvVR9Ncqr0a8+GCr+d1azTfmNQvZEK2ZjVTMw56W4owiL5rCEHQKFGnbTtBh/OnMvU
QLcxMW+4ptQwJlNcm3425HhQA1fPQge68ADTHcDChq4eKAFXtCV8JZoeNSSiMPe/wey0yqUQHUmg
NWVOdq00XG8FQijtr9CJvAjN9mt5exugjymW/CpAT7lOVQa2r+4bCPqnxUxHPcQvreX3Bmq+aKql
AoHS8kMaM4qlPi4CZq5ktTw3Aa9aaszG+ddi+bc0WoJ5A/J9Pt6FWcHsYVclP9fnuNE7ZHfL/IM9
hTEd+IMIR69EjvKBCOPNwXP+RKzM7+cqZvucDiCAgyVEfpBXqmN3xIr0zf4x1fgWmt8wBpR2zCxf
Dhiq8soELgXkSDMOP+qgYAQkVw5I8TBrlKRN1NBRdKqk70hWzdVpDy7zaw/WFkr7dzfe9D1mRMI0
j6H6YQ4Rch47OqceONK6xuymrIJxOec9ZkSQuoUO4ndllR7ZXb5MqGAcF1nS6VCOTsg72btVI0kC
RymSCfA6/w4ZagdD0IFkQk9hz/F/4dGrDTsSyMBjiwAVcDVo22rLPYo9yR12QulJ/izOqmY9sKqX
59LPJno7EJwA2NYHUQs37vTcwFPU1FTMuEs55i+RCmVheRpYoGdFp8acg/MsfqJFBvsBQoiyF3U8
cbCCohLEQd29C2dsKMGhQFfkaL3HoiHtTvtXu1JGZaruq1XY1zIk+bYqOpIbPFC37nvGbvElYTAQ
pZ58xDZbwPMg7M3MT9mzxPCnkSQ2p2Y+oeZE2cNI8dDHLIw0w289kcWZsrznLuwsVRRCtZFTenWc
2Y84mye8QTFG/KIULzt5V8kH9FfJ1Ho9KPWynLiUwVcQkGqI/UdbW17uqO2CX720MLQhAa2lXsO4
YH6wW8yqHIrMEAn9wXyqrENjwQt+dKQR3T90Jouibnr+hVV3EYygjY5ibaxB8wGIrzZN8yFZ7rdF
ko8Rx8DXGwvDD9hcW12R0s6MxMyN1gAFE42VD9wT/NguV6dUidHSu3XbJjVHJBZ2CQYeUv8tXqZP
/YMKvz9op7TUSnIKGCuwy3AfdvlU8XpuGFqPrPy5yRMQGzvtPZYMbcyPhA7VkHCRP6MZuOJR+Hqd
CDZrDpxoUvrp1vmWjgfG9oiFKRc3Ycw7NKHm4+2Ae4AkyDpp/389pUyPambHX67N/pKV6X0yLCye
lIaLgvxCqAK/Go1Ge0A7Hrn74PHiFTqT/gU/+LUsgkoYC+QOhgz9WyhQ+2pMOmog6uDjnR1f+zWd
LYks0wwJ8rx8jZfADPSEEJNrKa86vFIZ6ZjZ65aMtcsKlKwKTs+/UMwgdWsKxFd5ZeMQjh+Z0aGp
frTUs2pYza+o6Ze4wi9hCtdgNh3joeAr+aCJdofDNGOen1hvyuf5ZJvV4AAxmJxzSJoWew95P62S
xHiC7sDtTTFIHRGuDugKr3qr18Bq+jeGwakWT9DFysqh8qREyG1wyy4JWqkNI3EYw8ObnqP1rMA9
gYMPhnSykvHSQ8Cz0hE6RvUd6K5PVYoc2h0Q6a4KOHfrNUJA6Om2qcUzmAb5ZiaWScV41zhaxRy5
XT6tNT9rI6b7+9LBKLgzE4NSI0rd5lCBYyuw4PX80eAscxSM4OXWlcNu6Qwi/Z2J8+oO2HF/1+mx
5VA/7Pnt0F13tGdyQasmR+YbtOtpuFJ/NkSxobvq6nECaENIfCkJlMRWZlZh8fDJDcJUIHYhEuVm
FvJK86aYUMgB9PmM7RHqoWdiwm6rTG9GhNyYmcCk6/Q/bEFx/pFkQbL7J8P/5g/jAI1nVfqdOrq4
7B7wJ6WXgdH1WldJjTXT5r9lgCVsjrotGP4LJlZY4UUfaWHa+Ww7O1PN87Q+zL8Edz3epspBMbRn
NLuH8b2hxQeo4JISjnQzosPtdAMYj5v+EcLNVvXyJiumDq/S0LHAGF3sbAWSflfch83LTGlxDPOw
7YZ0l5qvqHw3OXKosALp2xlBrfFxGiawvv3H7UROct4SJHswMM++oyaZN/0Jv1G1R5/JlOWuhljs
hIDxI6ZyK81GfMHCt47Gg/+Rqx8nlAU1IaM2/lTLKlUEkHKlaz2fMfZSsff2+fV9z8HVLbIDZZNk
a3yG8HveClCEFVhtNgvBaTErSHvrGt9/2RAYenIGKYVXLBV72bXh4dgdCXqAs5ekDLbw9WnRAob7
eQkYtg3RJfGGfNRjSX/KHd2FvvjsnMHgrMCVjyv8/KgTBl3/Yc8+KHqpSky9aYsCmU/FlzjtUFr2
/6SWuBsYvbyWFJLa6DR7NWebx/UDqS1o15dd2u7riRLJkrv4wU9qpqozFVChYeGU39MfZkZZeXfW
gHhP8l0w7O5aCSa0hKZmGK1B+CpAnumuTfYvVS5D/SYjCJ4O0NwFDYm3sfIxoBDCtkT6M96PvXNN
+zOvb5gjKmUTQsptF8e4hWNYVDvNKWb8QoGCgpk4zCMmlmTjqn/yOTb5sj1IjXlcLodPfqgc6Dsu
ECDOOwDGfIZK6uHUq9EE6FNqEGb2p+PQNuL4NjsFCC1KHqlGXu9WxQ6SRHAdX36H9A3VjkNJtM9d
8pxbmCuGXNUu7oJV23FCHbEGxAWbA+XZjCAcdPYidHPuq278kbgqQeMSRx8VusyptAQ8Ytptwguq
/4qt2yW9QJRxqDD6ra0pvDJ2SmrNTP2PJOL1XEyZ4pXipA/xNavBesgqHbipSi31iA07Ax6Po5PQ
26TRCoFAfphw9kuAsEGgODbTCSQH62JP14HoAXB1cwYkrAcD1DNKfU5dpSZGyytHNMMUu4NvZivJ
hecVeLzrd+zD9xAFjhC+GBew01nPAI724dvjeojArJ3Qesxa+hBC5EZ49JNXhgDX4wjfO7Vl6VvO
orp8JRRW4ZqepSlirwqct12AbWb/xjz0qFocT76Z1XDl4pQEIOJcBYpAADyyp4g7WgyD2EEkNBvz
9lIfo2ZSUp/ymYchpcM9rprHfos+0oAjAfHun9WpzKrDW7jqRlcwEx+9yMWctx71n0h49gWvW146
CBZ+ybdmse9WUJItKVljh6v6i/FFGkrxq70pYlouICFQqcOpT7GpHKzmRpaddsysjZaFQUsaAjIv
3+9o8EJn8SU/SBEuVnoKUAu3fEc8KivTvry4vCQTY3BhzXCshTqbC2wn3D7Mhwif440iRoC52SVA
zJs0YjzFc095wBTh6AY44jv1asy9ClHAw0LuAVVT8IaIIyK3GzNbW87TdEcgEeMSHKyEnSPavikn
9qb9A/KVL3XE/d9K+juBrGDGtp/V1zqL35C2SL3uaJalqlm5BrGIUF5UJ4FKVcxwovqhWjT0h7jH
4T2M6R/TRUAb5CI7cNN6o5QD112l7xm4M4DD0R1oSJCubKLLrxFezE0LiBSD7+a/gVW61yjk7Xdm
F/6GvUQcUvRdQn6Dboz5vwYqflX/12gz8XLroW39/7OcthYndX0YIvZWbRlwOnuLe4IbvqFbWUTV
PNW0hhmhq8DbiUabtLaulukPSz63siA1T78YE5snJaSBT8kiYeVZqHl53EQHY53hynq4Wc3VC9g+
vBVnw2MkN9+HI7H09ryoqHXIL6AlYLKIGl59lrvbJTvjM/G88DnMKggHr2yZRYRdMOqHHViKXnHe
lcII47CdIr+4MyPrPmB3zUMWK6nr2vEh7LwAh8q78E2TGh1Gpy4g+RnAVK5rgMENjN39JS8A2PDs
PybL/lnmqh/jTRfHXX+QVg3gcGwO36aIcdU8Nm+wf1Kp9Qx98qbAGYLXE4UhO1UDIHmEbvepup4z
wGCLJJdzp8SyyxgoIm647DTSQ+fafxsv3saSu41D7bGOqkR0aFDe2QPCv2M+THqGGSTYH3quRc6c
f0bvbgxeBJk+9bK8y6unGG0OYIAXq9yzeGw9YscWzToQn/qnM1cwqdqFs2MY0KZsmF9DU+Dxjcmb
ejhnIOvrbYR3EBqEcxJTTqjeo/sf4CQppGzmPMgXfTFXvtMjuxRr/EKKfY/jk6JxoMLMjNhDlVsw
CHDj3FDmUnHEC//DRW0ol7YEa5Xnhpk4Umd/aVzC7/tI7ntcq1XPQYlLKdUcBfsgpPcGDMgd770h
BhDeyAArdlILzeN037iZQiSb+gDG8A+odtUH9hDgcDTb5ZxOIhorYL+wiL87Tk42XB5i0/BGfIOq
D1naQpoOoTjHNcjp3SkBOq14k6kEnELcqT3UlU8/1WhnoBtA9gJMHmzUoUXxwXIyRqbCbqxNciKi
is1pDht0YxKntKtEhd503IlZ9EYugYF57lBTlyqJQUeMICb6X5u613p+71YPnoKVe0kxBlcbeDyA
e8+fiu5JAbSvDer6UPPlXljkVsQRzwGgwMyO/5G5g2xsWafR6Fx0LxfQWe5fJO2pmftO4s3gkssD
OUibffbbiFjvBgXPRG44y92Q5qGxYopD4D0R7UZyMendcJ+74gVKJsDHmqPbV73e0HTtqv0A9zGM
An7aDjB3PzRhMYXm+a/o10xx1KZXrvChnEahvAiVCdnMMAEv7z6JmptY6XbNEFcIlwYYSKG3kypL
Qvc1BxwUX6dvvJuYaYfd3HiVeeJSD/5UPORADRABKuoB75pIqLlKP9nAImguXhjUXY5M7S1bzhF/
rLOk+mPaTzkPsIs5NKM1rN13SHkyF2J/bFKo9oIXmbffZaXFh2r76snAjB2iyebjfuvLGnj+fnMB
6XEN8u9kHLadt/XWOpierpNXD9Xu0nOTqEin8MyxR07YQiGaSFIWMqt13b4HaF3A94joMEz0pzjG
xF1ROQeVCERwARroKdPrhFE2ULAJiAZHZzvC7dBKmAaba54v8JLM3Pb5cveMwMap/mXTMNt3jPeB
D25eYpDvGZfemGgxtL6Tz+R30e2gMItZgJzmlXmiJkyw0xeKXR0AF8NiKp1ixng3ffHTXJ0/ditX
1HXFkhQnLLNeqsB0n3iku8N3ypvHHlWYQWZZbxSiyhQSb/aaKFCKbTG9eaqTFPfDNyAU5gWBRsry
L1AsDgzLhLM7inoIIRz1nwzv/KZCcy/08nPtvxYVSuNTnX8vDLH/Y+Q3yMuUVcaLEX25rAu6MUcg
++6bsxrRQaI11TKL2BuJf6B7nwKW7aw8BTDN8VeLidG33f3OZDZk3R5LxFVeNkD6oAmsO6E79ecd
di15jmY8lnF8itslBD20EKFNfbGWgMTzdHGF/W/rlbweNMEr6YVcQ2Wu2fw/8zLIa+MdJ5D6MKnn
hEEpX9/8UyqIdF7bzQpZnJ+yzOsJDIpNmjRmhX6pGoFWOSk8Kyw0U82Bv5o7LXqNlQmc1+KJKddZ
58IoEpmwEM59gHW8rNnSYkaLUfcYQa9HeD5WrU5HwrTLBdfm4Z+LfJkRa4PIH6ZEZdvIqGCuyMia
aLa2xHq1ZxlRoGUA+veLh+PkXX5cNZjqGaGC9dmWOl5Qb0aRE8NWDuUzPhIhG/AwBtOgKJ2JePtp
NkoJX6VzDA7hidfYxDNF9D6brJwNQ4AmkXbIhWiHXazrRdwGf99PsAeElJlzgGKvcvXRQgpu/pXf
DnPrshDGBlO6z7gjsc5Tm151zkydN584nFr+P3Gh4ULpHAdwadE1Va/fBuPRxpZgMkz+o0W+Y6h0
fuQ3VXY7cSBfogziymUic7vT3w/uikQyUw8NOzAt/1eTNB2NmDzQM1YiorH9SDFy3j8FGv8nv6LT
rxiTpbdMw6H1XxMJeA2zn1cf/PEyESjOJhG5hUdm8dHkIJt6dBJ5Q++DdgP7T3t+JzDht/j0rxBi
eYyvvHFFUCPhmYDEAJXAiklhMooTbDDl4fayxxHwrByRWzBsSJNcOfhLn/TZfzMCPX/yy6YnXrgi
51A4RkG0T/1lH4+LJ7QKZ9QT6RBBU4G1WpHZJjNqdt0IrdJZTrL2a/bC+jxpUCiU5pmjwpND7jrI
ux4R8bYUMIrBPlAPZ1+X1a/pDvIHxIDWIEGFR5tckCPQumzUEC3Kj8RJ/zlVMsKPLLMs5wffDhNM
fgDWJjwqS/lncW/J2tMPP3hWbnCxuHFmugVb0eWbvCw5kEMlaYrslXzuZPttsx5SI+GZlIPEODcS
5gJHa8Pj5KaTVjaH2zMtiTdtus3OsO2i92RiPqPnQYmgdsNCOcam//K9wGaTcOLDMTa5Yk+GMP3s
EbzTJ2yNCWCC32Ditg/I6zfh6fg71gsqkdFaUk6FN/TeY4tvzjK+gLs0s8IgtSm/BHhiMySQYtc7
JxaH2GVVVZVvTmezxvvD4s363QhpR0R12HeA3TuQol+CJwXS4hG6Est4SIM92poqY0BFn37y6vrS
lxZj+8xQWOVBQJJ8DUUKWFPQ/q7j9N/ngPh145/yIvBzUMw+RlMCNWaSl+pA9sKOHdPGAlruOjCw
epy58uj0wr3uvyi9Mko4Xud7Xq+0wWqTnnsaE+WA9atbHUB0niMCIOD3/ZzCMHoD9XlqhNjjjYG7
XsZzeF1plAD8oR3Q6lWvPL60BgDangOHLAL9HKGFa7pHMmCxEkuzqwcaP3wcQRxTMCc8vkBJEleJ
5R0KTpg8ULBdV4c+Twgq1lViVBkxZcxa3c83xxzhyWBsAwkiY/3HebjV/UuCZHB2G0Of4LAelz+x
Xq4y+al23uamF5ftQqkqzopD+Twa4E8icjbo7+kTE4IOJYPZebW8MJDXm5ZJFZXH08K4iCh86yL3
8dH1nvSmfpfJgEo4eE+jFIufYLU7lsGPel0Vl722A6soa5OpnH2s0S4NdiyUKHaZ1t6Uaolh86kZ
sVLaCTFMYOwQc723crje3F6ND5KCmNzynP1NxTtmtWCXXmddFsvKzNF6NqAo3xtRW8k96pTPRkqN
xi8UaUxwnoLsxysV9p6Xni1c/JHpQfX5wELKhPjpSATqdF43i+CvDN4nTw1bG7hpyT8B3LUAuGtp
dOMfhaGvGKvOmENxfWcVilWeRxTK/qsKM6KtvcghzxGi7LQ+fXbSMUHWrfoj/tzXO+T+RsBanEXl
btbtvc8ek+C+vTWmH4WLWbyFM6GCwNCaBhatKvd25vuaSnqU7yzwk/XjqV36cjocJ+ecyVFlHa97
Sgh45Kcu2/lj5W9ZMXmhNSyntaHhL3eT1aOntBp7qy2d4Pn8hFfhvEFtwCKi8BZ8NDmSNjXCUglQ
h3N1z+SVAmyrqJWtnqPgyQQ+6cpXWgSUYx5yLIgGHHiPbTPKDOwEcpXAlGIIUFikHCMVYXYqo87Q
POS/ChIqRh797GN4SlKJDYhHrIu0YDkc0+O5ys6VD/T5Xx3xJBcxmoltzPbHjXmXXewo0mDq4tqJ
23+POzblbpxFCw9buUzedS2Ay9087rO398cSjUT94vC9zD815CREDNa71eteBq5WFsYz9UwtD7tq
5pJeaBloBkL8DEnexh/G/6llkoyL+ynLCrIPp/eGrQmkhoBxoHLBz/BUGjxGFDYgjTfNwW5CEhmT
A2FW6t4/uMOO82Po1auqc/1G5a2sjog+j4136xTPK+lOQjVGNmpv+BsEKFjF7VtGuvYtFoDOjQLV
q7+CVR8e226+1R7qGV270BhNpeeZjiKrK6uHp8EMYwiNxjxS5kiRKZTfefWuym5rB4+Evu7f0/SV
2ZPYXDhPfK9pUIuDcuz44UVHnEZOfNVVJ8a3PqTJiRVxTh+RgA98N9IhLYeuQprmjcVTRxj+DzVJ
KBMDyI3rFiuyKhY4jSOWQhJpIXx+rKNzek5b/iiPXFqGfn7fifNaFPamE6QyEgyzhU77jB5m/Z33
tpqr8NQhNT/6hfqxzSmOFtPa54bwUwEVtIBDT6bW1WtZ4kyqw1zhbyGnbT3EFhdU80UyC7lF1WFJ
ZkaJNmaYUHixTfSnIae9KdjomfSQS+7lDPBXBOKFuzdZMZ2uGMWsawvQekQDMzr1gFcGY381SKIf
vB/nvLiBtrh7VRm+7d8JpHrXP3omJBqdTKsB9Db/tBcXSRDtUqx7Mp8XAqtlNfJP87gKyD4eJJ5c
06lEnqQDKMhtpuRMSgvfKRrVXvVuo7AtcJyZ/gJ6/y6eDcwRH2O9Auj+h28NHNH8qQpq/jjI5hdP
Ew1B86sNuP0lJkDs+KK8HbUl+7xJUnFINPp4B7Od6eNATcEU8ySa03j/82hX20lmnbsls+uAtu8S
QtPbCPeGWB4mc45F4NWqb79ZEemxH6GGbOZCbLHc7PZYbFLyKvCKmD2SXQDL9xHTn027bjmadQ7z
VNyZhBI+gBF1+TNYTFTJ+8P6OV35uAzT6xgC2cFt1Pp4MC6iA/rIf7ElpAOrRicL2VSfFhD4z7R0
JQyB6cUISVgCGsD9vJv4iHB609ky3mWpPTE/EIrYlrzeMXICYLEtaxSggT2HBhvKFmoLA7zopxOL
cJXfHwyrGsIylNZSNJ71g7jODzk13G2yzNuyswWmk17Dxikz1wis+lGomCNEIrajTmcIUyhPh7+I
n1veBtQuIQXHtmGsag++6jFQvPUkk0skHA0TbA6Kn4txzQ+2tynIPlTKQb/+NnExMPOzormJZOJy
bL519x6Zan5Ks+lIPQbQjQ5KoPNrsBh2GQdyYOgd8CV4fqkIailnm519HVtKPZfwzUxZ2EfqCe0k
HCdiqJfTzMytQgl/Y7gIVA9XXZNHDCws5/daXc8hnMf/657Asaa12vI7DrkaYC8sM5bEDA3RjlYU
V/6+anxsfXlKy/SmCWBV53l6zMbGit4Rp5QelrxQXP2qqfFSmcyq5LaHiO0++vEc343ADezkw+1C
btonQJt0VPCz6vdbT5YjUNzav9B5NhNKtfM+Qi4Qgm0jbWj7YDKwP1yIOcCaQyI2Eanr50g/EW3A
C/lEcXaWNOZdOXwniLOrW/d+w5TpHeuyIUx7o8/8ZtAe4ZJgXc6M0oTZMO454OtHfaFIaVRXQkwa
7TCCpsEzVgJ35ZholLgDDXn75EXc47Y+9EVMtEYdnt6Poxec/2U0hogeqQlN1c2KVmPHAGYUlwLA
NZDGjHD4N09u4A9sEI37BaSz8YpnfuIy71a1hHYSK9FrFBNFNY9yFgnzOGzaLjkFJV/ySyHwZtK1
GCfNx0AGkoOeH3nhUGo/zAJj7cjiagwGQ9DuB3UFAUU8art4JFBdLbvKxJoJMoNdCN1KM7biKJjS
nr66RMZLwcF0bugDB8MIlxWUQNUa1gghFDvSEv9zNSBddHe+8QyhtQVNWlM5YaCw0PtuWSdc+D5c
IPQL5bshdVNAVhiUIVQX0He/QVAQlieFd8ZdpCsoKyUOdXpgCsPI7YAMPPJtTjvA8VxtzHIOeVjA
szcTIrdv8yJ/MpTKNN4TsNCiYLCdfH+ocoUepLXhgVGJgyTvMMzfrtD8BvXd3fibPMrWrDzzUCLB
mvL3OFwexY0x7xv+8rfr455w4IrMAR+e+DNOk1dr8StguW+vkrpithkWKpOF5+AI5bZljKt4QcoI
XW/vSP2mKCymVFXY2OsXpZM1cZ3QK+U/pLZjPKzBSkdOsV5kXZqaWuNYhwk/81Yrx1l+RbT+7H30
qlCIqrtf+EMlT+iV7w7/q8ENiXBL+4LbEokGaCu/asrUeN6f+UJLEyD3BStOXq8AfdGU1uJjsqrv
YqTCXyvDvnufFAFxcKnma2kuQG5IxnBzYaBiPa0W8jg8Jhm2pkk62VQWczHDAeUCZQbQso5jMyyh
nxKDLlDDqb7ih0GHi9Xn2qK6cvBzxTo25DrXEYh8vLNmG4Xaleg+Ye5vnXdiv+2ZC2ssKV0daAMX
WOLqs3VVtbpg8yjfOmaIaMtpr+cbjzT+BBTHeAYxODJ+Oo/ThUFHnHYaHe+QedDZZid/ulsViY7D
FMl4K1aEXjM+EF2XpK38Bp35U9LAYpJFQZ304zKywm4XKpqUZS87Sso9VMzBZuMDCKgdgmmL097S
TEfTApXeBftI8gWhG7z5JPTpBLUPuYdZMUVrU60mqWgiI3z6lea+AhdeJlE35hAiDFAxodGudKyr
kmjggT3PQTFjVtvr6N1VB7vfdHbLXOfJ+ATdjPpgH97U4J99hp0ePeKhtGgu/VV17ezBd0Kuuf4y
qXsAEGiby+NdNx9+piyfZ8BXPXzBfoVP6X+2Q/ag3A6aNNuFwiBfdZvXavhX5qtX5uB9YsNjRHdg
E5abc2usB8ANBR0QooCbQmx7n5U1RtIhORLMUCJbMI0aQu3/vT3nR3R7zIZzwKN+EZVUvfby1wKu
0MwbRBqubkOwaYkXSf2qJ4fWwD3V/6/ff3I2GpDk+2Yr6LYsnD/JLFxwgudkZJ3JoIy8BkFdX2Wc
7hC58607QmNcr3cvhMMOmRg4MXlVoki588t7rgpVpDw/pRAXum49x8h/I21gkrnArdHQUew/OGiy
Rl0SeGxey7JM743CbvJQKWO9VsBq0avAPxOKYDBJndu62B9/QEErIDKCVMitgdrAto73+JRhIg2z
YqzO0ymlt9v4A2ywe1qZmUSsPFACQ7OXxqHUC7/wUK+tUE3reBdFHUExtcljCBoLAPgXs2+C5XDG
c/ppbntbTEEZcMEXzznyYEKy7AMpEjLnkJetvSyFJRl3D4vbJkOlho9H95sO5gxaPOn1lYv6btXH
f8Bbyy941ND1oGr2j1XILn8Kdeo1DhQ4x6I9blv2x/HSK5T1L5qhUIjyvNMRjUs1TFRLKlx+PlBU
P523TlC4vsDcLxz2sh+Tr9i35zlg1VM6XK9hCghDVt525AZly3UfekpRQM2D1tGLSd7WLAfFvtGD
ynPq4kZCJSWKcRDfju/jIaYdhtclXwzb7gmjQvh4EhUI4UPfg9aTHJKRLjUQ4ksl+KVzOU5ghm0V
Yfk2V5QD4W0p2P1Nj/3A6juYP9E2+K72WmHndlN6uCfqExYU6Or/HwH26uspwXAttWISg3J7lPUr
aNg0s5EnfAUHIav79W4puEXl+0ikvsotrWhnQ/JGs7qd21dz86Q2ViRVBpC6OY+OONbOdthkH8XO
4utcF9+XrsUVPDX5PL8GftosqqyVeVxAP+cWfrRusc1tvlu7v7JR6APCblblVwQmD/Iy/vN4Yxk6
SJI7Y716RmwNNkM6t8Ojnb7v+4dmtR4eaPW728BpJwzGxPaAdC9Gh2qsC+rMaJcCwAUwfGwbgyIS
GPnP3TFgjTd6d7mm3Vldn2Wn2G2v0LMVJ/3P7AFulwZIEmsXAjwtKFpbp2/q3xTfyGy6xf0ePOCV
MfVcJdVwy32tjsFd+Yd6RLzRaCByhpOQ7IH8y+ClKndMrlg2UKJrkbD1+1KmJ3qyiGFvAgd/AfPc
MLo5R5z6vBK9cmBCu0hYrl6c+IWnq2Jkh/tB9SI1Gfoaa/+NCZ0O9nRGsBxr3sOuFQMcH3I8G3BK
2Bw7ieY4kpPpa4HNSb49zM1Ia9ki5Q2kHfOhTuKxPW9a6YRLKLFaE3pwWFwBg92ZGuReuVL+fR3n
2gOF30gLzJB6anO786C4nCeq/gR2WSnD4L3ovmh9sps8WoCO4G7cUg4E/45TrJrq333j0UliWOm1
MGSddJZ5VWzPNKvr7+8EFyuhizsqUX91XfWHhfgVMxigkEWNbn1rMK91R4Oxi2Hw9awbHgwLXPBF
DvPEYziHaZYLIiVWUUP4M9i9dMJebBnjE9vTCoMMMQ+kn3DSVWjDaZzdZ1/ocMXtFDC3yAxFkJXX
cjdo5nLeTEkQb2JzZF3eYoncKFb8dnPngLJ94VWowBJqgEczxCXW+FR4ok+q/+/tnOgkI/8IWbR6
iEHSF/0ivN1x0VhJWdiWY20ys9szj6YnovlFp/k6YcYUQ3gtbYCGmjph13uCfrT4oONEBKBHYsIF
Xx6yKOlC85BjYaE/MKg6jxbHv3d2EqFuIoyA1DJOAn8huPVAOdFrWtS8MwOgrt9tIrzftTbalLbM
V8MqD38n9tk3qOIN0TPdH9U2FdQbpTw5fSAwfOxBtgv8SR5uHazwXIDYSD0RxVO25KRgz5ItPZmh
c2V+ePrVzvGVCK36gE3EYix0rM45lKxoJcV35/s7lpt7qMunWA5kZlcWSgwHjIc3nC2xTfUlbu3g
S5vKrbXiL2PffHntMMJ0YQFnIiTaHfYTQUYPapuKWEYUsbpkJrt+gcUdc/vefcTk9JqRRLR+HvfP
3bpB0vGiJNJUuD0/nDzSa6lHU4VhSL3o/MTjMnkv//GiN6Y9TCtqnV6/8r1bv+S+BnHYfUkHKkjC
5fu6HYr02GxtXBDebJ+f6NC6VIXYf1+fYM0XArYGu/C4wIIpWAqG2I5PblkpOK7poi3TaXxsW0Lb
Uxrw4upqWOOXQlF82lI8Jr/lf1josfQH5WTpRoJ69JjPw2L9wCu3zmeXsFuIOAq4LkpaCARksu8f
LijWLY9/KdoX2BoUzyj0REc+ebBikd1wRcAVx0GBydlLc7sRVx9mHWd4sC0MpCKO9YflkkfraYGC
5HbWjYuFIKtsVa3y0+JE1garEE10CvBxDgbP8zIlVGB/jZUFS9JHwNBdEYiECvGfYxOdzD5OutKB
xVf4vOtR3MnZM4lVzMtneKD11s8g10ZVt1hwxErsZkDu4eWrunUfyFQEUIIPaW9ZCLfk/yfaoRhy
lsQTiRkAFbQO5OyJL3WcJXnenpm9BRA9rUWBXSu4XwaDfgkTTy7RApCCDWhWb94jzG6K4PTJ4Xd4
S44RE7jVAX2heYIzjdA4o6HDofPLShy6DNqJvfgV4Y/oyTjnkJeqXfdPhlnrVunCakILGJtq5t4L
jBdEKj3dpN1rjF9qOo7uuDTW+k9+7TBjCEN7Bq8zoJhZEJpaw/OOGNYjLWqRSWT1Lxn7Uu7vGzOL
+I/TUJ3L2UAy1V9CMzDuKf0Le+4Up5UZ4KkA/ApGjSss4dAxj9FmiFdQMtEDE39wbbtFjaNTuiea
+8aMoCyEKoqTLAREXAqfP9hefmwrFO4W4Wc/JDAreDwICUIEwrR+DXzRRgIvzYnO9OLJvo2eN77x
tThHUeBCIWT4eNSTyIneonAOFFQl0KrlZoFRvxQsB2Hu0rOwU7hMZbsI3KhnBO10eA0mHiJKx1ff
MziviIU/d66G+JX3JRmOT2PuPNqQMazk0krRKHqkFwysR1JGuqpF+KNG4e0D3liaLMi6XOmoONdN
bUjKS6XVBjcryJo0V/XjPemV7kuiM0ChyGRgaLZ/AaCMuYJIYzH085+YEMTsei0EViPVX01qlkZA
rrc06OSI7NhF3o2xNB8zJ6WaQMzBu5iJYBH82pG5WxPeSQ+jkdK5oA+yvpGDeLhHZ+ma6Y6sBFk8
RmuBRztdIM97oFr1WC9YNYnIM0J/tWjLM+OuDCkfJSONaUBKVx3ThoUXBLCWcS7Q5FEeBNGuPfvI
3C7d61dXMEwWfVhuv/R87FM6qp7bliXGIGKlztLwXkuxUuvDugAMqaO0ukU3M5Zdnbz7EsaQ3oVl
h+JnQ3ue18k2VoG4Ni/ZcU/2IErxpe9PaEUizkjHDJBTQBSElDIW1uJRmN901VXwVUWkWqBQIJDE
2b5vEVYdvQUixlVlAkHMHN0RPmvx5t9IiHVqtMMWKGCN9OwEC0G+UuottZqVH9SIATcFsdBhUPNt
sfe+j3LJfXPrql4BtnhvqY7SV35Q3C8foIcGvSH4XxPbgEOQTtWRTZq3v1j9HXFSunnh2RV4NR7m
mjm6noaaLxLW+XsvOEkBPL2egrGrfXEI6Ols+DYEOOY5G+XfH5gMGNxf6KTYGT/waQpXRy1BSN7S
MTW23CSf6SvQg8ufLsHxPxc5DUa/NnEfnu+dzdyp3tBGp05cSS5HGaCU/jiK2fTrLeOlNuPnCnz6
jCx4Ul5aebwYVgqoP1kPM58ltUg4wlFZJT7qHU4FAHOXCjkEU4ZqNpTxNSQets8bvkHfBbkMGZA9
NKxlzSzU3BS78UNTYcVRDswtywrpBtGNH+lvuUkBbH2BJG9WEXA5es/kbU4nrnHCFVqYf7ij/8mA
9NebugKZhcOi2m6P9Z51C6kl3YZbXTpNzczaZqoYlFLYP6x8YeBjjeIukWNUmeuDFLTi9FZXUZgr
As6Siuj5nYDKM2mERTvhdOVhGU+WRwoEjRqelsoumjOPPUNmajYakBpxbGglPHKKf9yZX88f8fnX
jbR5dP+oUk0skBS2/TmzI6E9WETtc59pPvdYE/h2KUW9Fcd6z7BHpScC/DBkI4g2NVYJxgJfvhb6
jzigGP15VDdBr7wPWj6SD/ZyG6h244yGi8dnGOIyR+ReV5CblWvmFbeibwz+TWceC2zvG2enMHHW
ezogcygYTEJIhP+nF4hbl1lI5LnGwpFxVQxIrxALFpUre/umdpWruEmMNnZQUitA3Ek8edfbR/nb
jvVLCAs0sY9eJ9pmK59tbK6gK61fXki7aJEcLPPugUv4nYHg45hFYBUvmTEE60qOHmy8amDzNBBo
iysK7UA831BJSahGAwRO830SKys7ALFkxoZAgc4I4G6wG92ldDmaXWg6b9HWnJ5Nmqf6/GQdVaVo
KkqEvnJS3LgaaoZuEkg6Cq41DtfZpNRnRogQF7Ibs5mkYSqVi+tsLCZahjsebsT3GsJ198tOhOI9
b5misphJzNzvVfhp7THGfnXFXcoMbbtgD1la28gU+j0QqM/o9vhg6hqe3lW+eDVbGXCzCq1Oar9v
ckbt2ZIbl5KTkgGFTnP8b20b/wFz+hkZ3wmd8BeFVi9+L/2y4EEfIpNVGwdLTdueZGsLZOnNdene
5HKAmPPXcZ/eYHIEWNkGXAJ9MrOsLUvnUY3iF6zAsgPh9qS/H4ipXRZdajKAgt/oykm+EYH4hJxG
SUwzSLjET2OagPkPkolJIn44WX3PY0ziTT5ZoAek5l/CYCv1M9ZcIgZj46J9FG4xAELmdx/NY9uU
1oP2FJZtgXF78MmBILFGf8dXPHtGsxlL/vaEoBp2MGMbRoeSbUZY1BGUuq2rqxJVwMZ2USDkhBIr
CZ4vquh15kmlyJMQS5hgDcfaPCxtDl2XLpTLl/dPoy78K4gLV9qMd2JEc8m7XNrOP+gel2yDb/hs
rj3ouNyIbME4ATEJee+AfrnoxTCPmIwdHbFn8U3NJ7QwRFP4aLJyGa4T/16hiNZlpsvchr6RS1QN
IRoXyV790rlzY5YXtG6VU3ZOojcT4mXPv00zw+PhSBdCyUe7bKnrLRVprFrJgvqrPqyzGUaIMncE
JVp3GRyTHBmLc4olH+DisZ7pBi1YCEDgF4eM7+D52aZzL5lIkNSNIOx9ctT3mm1a7G4RUF0yO6Mh
VCe1Vd4BeigtavTAPMl4yX39p2v28vIgaW6AsYkNHdAUccMxQj7HTTb/dSW+baEzkRwhFeo+BXYG
NWddeiDkUm8Aw6sKk+xBoJWb8fZ7JPcq3hXDPdwZ3eyIXEkuSkFbfVYtj5qG3xb2Wc6nQBiMr5iy
GW+AQzKO7XwSRGPLvaZd9CzPNOYicRZ5z8haEAUZTntKjIKk5r8Jb/ooAVMI0zk9omMxt1ICcVi5
4kSYnr6KJMME37VUpePuBpCyrZGQbOwMlUY1UGogk8KLoC7GuOfY5gSH/OTdzAjbQpucORqeZeul
BGhPkVO0Ugd2PDTd1BgKkgZizMpJrnAHs2A+Z4wu0f4E3FmlXROnF7/XiAuecGN1qJgu/vXhnaVJ
zhcSaVSs4WjP/S/wfA8nUmozxT98hRbUV/VixixlJwD0eFKQtg0kt0eT0G/n9NIoR4lAixF5coQE
BWuTflDvpZxn53CAezQwv0mmCTQoeHWVYu0E3ZMCPg0OQ/by5/rFUXIzPL8gWezHrXcv5rEm/uNV
rH/MUbg80RPkJbFX+/742ztcfG+FqELYoYQ+lmmxHutAT+Z234G5+ov1FFF5dL9VijjiS+lYYOzW
4i/noDqs2TIDXmR2oTzCL06zsxb/rUHPbVTSRGG3dyLMRJVSy1uuFpd0non5A0JagFE/GIoPfDUB
afxv/bX2JDvi1Cb7+yEYvABgzuya8x/FwAthRuAeMp/6inWr3szzq61keUoXYffGWcVpYDsa3ewo
Jb50Cdcn/mbBdenlw6OuweBht3Dy24xgob2jxc8e4TopcGPU4LARw91wo95tCbCT0CpmpnkLnN4e
8IurIOQiw6vmgmC35fehX8GP9gMCp0u/O+hAj4Af4CLskXnzkUdlsGPK1Vn0qAox9hSKC32Fhq97
v4QBag0GjST59tgDSYRBOaYcFPI2Rv6bzRClKCZzLVbKzPRNTy0Qxj0i7TbxCKpCyCZP1EgxxTb0
rHYZXXP7XtYK5ZcSAPAGpVZJ+/RSkVfTjAozR2Ekop4zS3vbCpqdWY+LdRqDpvCAjIfQE0YllKno
onR2GD7tT0XdhCzq2gCkdhxFKC+ACjqo4nsYAuUhtfs6iKB6UWdt2PkHU016etrbpZ7fZyZ3CebO
K1DD+k3GEutLh95S6mX/Nc/P2SkBMNOQq/tQyGAD73cEruSJlfbe2L94T9EUh+ydpQ1yEl4m+23U
sl4wXnukmN+IHMsWKG4l1J8EiJ5evLd4zy1Y6rT4uTxQhA9lqEl3RbpYUsdQUp3PmI4NCIfIF743
tHGVSCv0JtRR3W6/krXolz4vp90wUrmZzpCifOdRIJq3NluhYzYm9mpIH2mrbWvAek24g+NLtW5c
0KZvkFRy55WQaYczdACg5AiBmHtkYD7isBGXNl9elp7bXVv9+rc666S7oh3KCmtHtK0rQmTky8dk
u/GF8a0mdWdTVy5ii86yrpzabjPqR1a5LBfU1lByu2ow7cxyTi6mBoHhtmeVRcpxds0p8Rv/UMlH
UngAGGtxX/GnIuyAv4CD+pSkWD/zm9Q+qLS9wh2CuEyHdRVpFy7Verph6Jbzptm7tr41PMeg9/d/
/xUYjulZm+oOzcEG1ByTAZ0ovcFloik9MSTpKJFpvjz5mrdj6ehXaVG5AHfENynFAXYNmVP0G1N/
Gctuca9HzngmoQifDl1DLGLjsmkL/FS4hhQrpd7o+lbNG3PsUDVaw7HiiAD6ovAqhXDZrbxDsP74
aPbIEz+RnLeTLsK+AsuOteyCWTUedQRg2n0LSAjEsgOLlO4jGZFRCyRHvubBpT2js4+/ExwL3V4N
dFmb50TGs7n8jAzXROFDzqMQUTkL4jFgNfwIqrEfb9AOYZSDugYUuYY5+UJX7kiZFHzpKMYlvlNg
UkSPOQbwKXvT0itOKBHvhxoYvnVGbynt29jCOmU5RtUCqeCCp0ds0ruzYfgDGOPhObXxpIGIPGn5
xKfS5+6i2ANez2RRDIjwnY/ef2LiGRSqt5URD8V9G8meOCZiMe+Rcp54or1fYdlLKPeJjSD6v6+6
chtVPGjF8/oc2ZeemKo8i5dP+1aZRU3+DPdzU5H+e1zTTi/RHpia3Gt7L/d1T8gcWhbJiwcLXqiK
f/Tmb7zD3nO+TCAahDDe5Totp3KsO6zjG8FkBaxivII5UJktA0P6nG0JhGQIoZJjRF0UIe55O/gI
x7bSOvo6KzmxGBEbqLv3T7pPN85c6pmbdFanuh1mlLJadt6lB6QCUOLLRDPUYEh6QeXYkK2DGlTf
PQEj0xm06wraMDP9zeTVG1iRnxvGCrzWkR8DGLpbMcd0pMiMQ3bqYEuKxpBu7PwSbR0l3RKe+sw1
O9WTos0D8Ovl7z6Xgou6OKETj7UtKx9Nz+0YKODsVd59E5Jmh7duPQfEnGgIZ+UjSkWloeBzBWgK
pm5U1vKRl0BUJsxSgEm84K7ZU5RPjatV4RKAyXEDKztV76jE2OULm/kW660tSYVw08G5ehpYbror
ieWuXT5fqWJNjb6OpjsQdEvQNvXSJVfoAtHfdWjTl7ovOmPsJKlbWKVBHl97MJHB9QhHIiUy7jR8
bpmyGGoa6G/oCNLylscNH5Ugz911unpLwFf2YeZ7p9c5H8wgHENp0TU/7FurhfPQYSnXj6f3Mo3f
oKc/aQIntBnYEMcGapuwug+Gv0aNsen1lL+bQE+2OilEFMM3gkbTBs727ExstB9/XgXISNbPT0Ov
v2ankXdAdWzScI0r11IuEwPOr5WmceJaCS4mkLLvr8+eCcDwSls+DyH2Wb3I1NZnCnEZOim0LG1M
yxB6l9IN4uo1Y67jSVF7NU7TTISOhW7usvVQpmTIJqT50Dw65uZ98Jx8zTap5+uuh67t1bVfQXBQ
DxcnCf9eNxtqKKz5pypGMlKW3l0XicI1bc8hu9iC2yaPkkBhcjDC/sM8aVfHGXX/OJTs9LmTl72p
Oy/Na45i9EomtICLnSX1lgIcCAzX50/NRER3nCKeGd4zfBR6E38gDsDZwTnE6IP2QTfaS6OgHVVd
EUqsHH1c1MFjCwW8g3WlvdaBlhgFb5y5NHOxeM6DTYZZYFOP0lMBSYNkZjXaz+vxkR0XyeV6VFyc
wo0nP5WL0+fJzKWVJziFBbihbdYrUCemtXnxH8YurlkzVFX48865DvMQ0QEtVgXKhRhHKKlracun
gNO8knZ1R/F8JSR2vygcxYhiwlPxiY9dVIXgBCX0efnetKvM6bOSfgWD6v4nTZHQRpRJ4X1c0zld
4kLt+8egBBk8QuKSx0bXB+sSCBxOMz1P/RGLlMQSiBWaZDuycsmxcu0W8Ty+IGiDRcPpn7OMNVGv
AYZ7oXupzVCpUxQO1sZc3bQkyCdxaTpwOe+fwvx9PWcpZVpgP73qcoQ5AQjTysFJ1t5OPl1XNZek
Id9hIMeJ9BVja2EQHMHQEFKZ8jw+vDAZJe67q+JuM8njmfykFvW74X6sIbqhqAF2rgb1JwQmLK08
F+eHTegC/B1zPRp1S4Rztm8Mc31qmp8Z0NXYNqfHFd9w5l0AwZ62DN1d8mWF84jtkbxhFYzho78K
CZpJU1q8Mi1U/xVLOpAhWuLHhSUZPGHkVFlHD7659PuaC3ToYBJTbKOH/tOf5nO8yWB63L3OZC7o
aBb9IW0jX+e+5K75Z4X9dNtjkLTNF82pS+C7bV+vEdtAYBV5+AzjeVtSh6uFI83P6KQzobfZkQvS
YN2Q+qZikX/bnsBiFfssfPbH55WzTlmPdub/1QxzTZ4pBRBWs5ko61DPAqpZ6P/Qwza9+XbdnOeJ
AZoi6jQAp19AowLSycNrKcPxGnjHoYujo8f6LNvUntiD/b2/h69saCSgR9U+kU5Yy2sK6CiZiNwd
E2tFrJIiboj0jQZRuTPA0dW1MLNy3bkaq7iTCN1RNK0rz5U5ElITTeZ7CZqsFbWpwQfjw2AL0ygz
WmiZKoh/wLzbFfttWWs75XOMiu2rDDuhyV5PmF34ygvgf+F5b2rrRiVpqT0KNOhGJbInv2pyReIv
Cnxzecapl9o0f9oEmIyc2ADBapRkXYjnfLTJ6nKKm57s7bsm+9pgrVMwURGLdlcQpo1B3To1GOly
arWHXKbxJ1w8sLl+acNC7jrPGzV5oWxMw0C1InX0YqVkU4c/zlU0uyI8juk8+mGtHa6X66Wxx859
DyCu+vpn3SkEzMiH4SKTe1CkD25xIcMZdHlaYWHCo650bH5SxYXWsGQyc2QSwi5zZPdNGksPbbc+
KT4Bkx8fCZs8l1hKJoHxP++NeK4jHMab3iFkn63ZjLoHMORxy8PgI9psB7OPzgagS+wgvMrRTodJ
o9P37rKJC5eP1P/yWJTbxtl1EXqcvSlAYxu5k6Ix6gqYTQAcWT+L2Rj1kuh7JqIe+DiTKntopuD2
iE5nkljqm5al4nsUeKY0c2DByCUvlbkN0vKh0fMJyMiMXaOHx5qGvGYOM9U7rTqO060VzbKUs1yV
3+jMurXW5Uak9hTDBalfiQDuU+bfWH3rlJfRlTpxbfDXjlw1aS4qVAQWtITofWnOhzYjU0j5wNK9
nIbV865rdaVmgKVak50NeU7FObxUiD92ldbAKReIDya9tuTOjK0JFk3HAj7ZYzB2T5McEYkulPR9
YJ8KOfVI73H65vrsG7MedHPuO13DHyxh1yCBAGD0Zwby0/sYyLuQ61A/5m6/+fyUHkecqOsePd/l
bBRGHQBdLbmbw+Q1Diil7r3rv5Uil1uK/QaXoy9IZicyRLxSut9QB3dL/QRpx1/BOi+qNHZYfmQr
yBDqDkQ2G4N0/cmZmdnslDhE51yaV+aUWyW5g/zr71MuU9ZtS3Sblmsufwp2Yk0+yJU4mhKfLx2J
o3OJIcppWq02TjgTNSnKVJ3UoiuRfrCCLlHy9kG1+5q73tPUaaTPyf0wYnY24TVbzFlxwCPNt8Lj
KZgpyKfwMxp4UVBcKtX4LKQgo3nyaOUXMyusTjYxKvzJ0UssoINW4gdgl+2/9dZ0mlJOsPXx+vM+
E+FWTYBH3lu3rQJo3Ge3p5JtuB+eY7Qxbad7JU/Hx6PiD4UwNYImbELS/6UNbhz8CKYSXUR73U6f
hEU4IshiDkS6oq1MuclSdsyj2kZhwYd+Vq5ZGqkyuLGcrAAznzuISqa469Xc4JBCkuPtCbWNdi3f
Wd7Wx+EpwzNPfUpIfBb754zVFT9vOIrVj76lTjt8wTik+dFhAfsejn65w8b1rdBi6LWiKSS35rpA
5J0U1FS5I+Y8rdNGsXmQp5+wtbvNFsN6WatpP824Q1BhjCUVkBYhw8Un9QkCYpJFY0Br1i7EsBVd
gW73oJ5A3zFOZiMwL6VdQT2TGZg92MWkWQB6wVSYhYIt8jxlTP9g1vgNe5CN+B6Th3paaOfLizlh
B6QEhKgV5t7LV01imrwMCL4xX45abATAwl6Q09sW63z1j7szl/dkcM+JVFn5z/SYu5+7rn70yemM
SMzNqZoAUV1ZX+b8za0gmf2+QNiFwR8Scvk+jSI1GoaA9HAw8yGBZDcPOLZ3o7Q/9WaN1ROBcuZz
c/ai0yxHCEp+FWkl7G9ZY2W0m7mUTGxCiCBF1+ztZ9bUk9I6hkKLvpa9calrWa98YgzTfvxK2qXq
Ta58zPpN7I7lXJOTioJ0Zq/X1oOCX/lgDKingZi8ush8aTIHal1BnPbbIb+fF/aCiVlIYZNuiUGa
tL1Js7mYyfQP9UCAlkaDf0/p2DCHxncid99+x1tZpZqekXlRh/ChSzeN01s1dAokqZkakqbWSKWV
0bk5lgsJFbaJuBP7MBUcTqM125WbndJa7CNf+4yoIknlzcB9AiAzYqu1hC0Fu9ZCsinbeS5HQN2/
5NgmMf8VFDo08ywsNjusS+j2+PZfbtTKE/rJQ925ziO/+kYlL2Jr1eZhEBCmb+jTXFX7C+LiT771
YaoKzN3qcnvKL+3AS9VHny6qvdlQI2px86/FUOLvf6QBu6oamAXJbO8pV67+LpYB4cPrTg0Ww6qt
pqNXqhqerf1sWjINZcvO7xoI181pKRoSVCR5dv1KyPkbtNkSxRF9S5MtbTYGHLZ5SjA1MOZfcXCb
1YGDp4R7oKjT+Y7ILGTKHSpUtlNFYd2jCXX6IuS5aUCAgCY55xztLC/yxllsx/AVAXtio1UeiSLA
YU0CxZKQzDFgDUYtv60CMNb2IJAbEuijKTX+PdQCVZWrXTGGwGo//wTKvPPksZAKCh3Wio1WEkXq
5LD/hVKoTQ4oiN3+ItXUgmRC1WcyM6xQBz4eane+A3L960nvJlgFA9mw4BEb4VnxLw9JUhDYpHjA
b1b2cZUfDOMk8sFpLZRITWtxd+VIRUDMHBTUUPrYt3nFn1upazuuIwjqXHw2MXKTnEXPvMLmpuPB
VR+8cK1uKOo5rXotzBIFSRzZWh2GK2en/HY5cl5IHScpj29wDNKMcFosj6G/aHFlvVwibTDCY3M1
s39mOpVkx8OofosnJp+T4MHSFKsvPP9kdoB9TcOKnglVOhBTZR5UI6neIHTMq1omisdh+zQAAzVR
0GadfB9TaCOhIupXngnmWMKbTllCPGdgfhKlJFFUhqpmykbhaYySaNJalthdiceGyeihu9p70cgo
j3nKJujlLXN5EHbwLZVVfClAUPbVew9TnYmzPkIanN8m2s/FV4tTAerN1UWophKUjbFaTLxog/jX
9TaJaIMHp/U+RtoRN16v/TbntQPuRDWqVZ7BUKwyzfawzmJeTV09oyE19UsF3BBXSlIGZFuN4dbB
hnzmiUFb9s36aCWpqjwhLGdxP1fuTjtGhP65Gj7/TrJgGjFdvxli1KlyStHrxdkT3rGL7NfSb7vU
pZv5h+jBzYGFK+UtkQ/tzUT0KqYkHyaKHxTcZ5H1lNUeGfrJsY0lzAlkORB0VXyme4pOlhFWu/NU
CxUh+FLLV3jb7WUQG9l0EbCeGPNJXSBCgLm5+kCGOvD3B5SvF0lBjkX8w2ufgHeaEis+06JDefMj
PPoHVoi2iVcXKBQ2mbx5k/WQ6oylhIlFNSvYzHmx0EUf7yjGy+T7lFC5a+6tBE2DrOrEyptNHYfc
A6mDUW4tZMQSUzHgvAKGVUXxiSfrSXQWkuQzCSTnDwYAbKh2CJ7H9X+M90A3WG8bxtURSfjYa5Bc
wx0kK3IC3DydGQNjB4NdnP/D6lHN8WlIpJ4nU0awKp6laYnUpo+trFQiDAye3lD8KzyC95zaaciz
GDEariG8NKVrewuV8hhJUiG/eUNB7M2IVhqFXpN78oQSKvld7rAlf2ZNcpk7I1pXpOSupEN3P4V+
LIPdbXiTQeg6y3JCuaV83q4UaD11uFUrY8Ph3OdYsoHOCYJeYqdqB3X0jlgBLRVO2CYEdOxqby5U
8dt2Er0s5pak8G0TQ9pq7XGfvYHhatYxkJBHjSEOtBhLFEm9Q4Ot1BtYtse8xTd3LavjLPTyvFjN
YWatHbROOuGMy7k5ORiwCJHJiVaTnhnskmGpS6JqaHW6yrjB6wCn09o6ZM75NPNJ6ssJRxjcvxYw
hJjDkzuzoKxNxQ64Z/noWhjL3MgXibkug1m+4LFZ7SSsO+w0FA9S7nrm3EDOpfAQtjA04/jjurAO
ehgIJXwyYfaCmShCO8RNxSuMAM2wRv4voUd/mUOlpifheaxqegY9jK6dMhC9VvpipH0djtmutg+k
wpWMWABQCSggwXrSTO2K9T7LpGO5bdSwhiDXm7zHHzPhhUirYWbFZhPpOoC+4xWXN8ZySoQoVZJi
ApUXhIJSOSz2+5cnSCOVDy8Jfq83mbCV/4cncvwhiJ2BJqyHyVEhPDly8v0OF/E9OQExjleYiOzH
6i4KXx7I4z/J7b3qXK3vCFGyI3hYoNjmqlhaCkajSOjgONoGSya9FUi72gYpfVRTldNDvlJAoyIn
MM8wczKAtsZavFknMlDnr9ofHGYCZ/gcfkJZshot4/Co4B/RzSPkU3R29TkKkDB/jMmWoDnh8xdT
lmSlwtZSEzngoCefbMKBoXnmmcxsF/XPZMq8+LuRtHLnXwL3suiD+/89NPq7wGrkEH8UYPhrLDDQ
t7HdSAo+Td8hMr7/lc7Q8cSMTU0aKlEsdlKXH1LFmBT7XlChEUtMLw+P9a5o0z3n8GWwqy/5qSn1
BTtuJDIktTm9pMQzCL4nIXa69B+TfmntoWj6ZCXHKJXXcU/xRVk8kv2Rz5NmQ5rWk9xtOW6QVVgZ
KwZkp4LoK11pxceCuGR5K61UoYfb8AA8dj2XnHaBOwmTSghJSn/xrc6yzn9eGxmwbCKlBMlHr+8i
3Ms6mWDh8xyehDw/rM0sBjjKP/p1UGXShkV/DKkkBjYo0BqP9GAL/aZBe3SX71vybfalezuwDPLo
JAOwOZLyXRZs1GEpvJ19n6KdJ+laNy47XXRWAL9RIHUDqpq7VQAbr9rjTfH7oGumUDwS/eDijhWh
jNm60p/f5IaYyfyh14DvymkcZ8yfIXDfQ1B/uTIIDaBNzZjPbMAjvHu9zTQI56Dm0AHom9Q+6xXV
Ju5CNQ0l5KbkcDJE30o5XCMj5u5oy48r+S8MrcYMEnSa7hju8Zxxx9PIrNJ1hatgSA7oAzCrV1qP
yQGfzXQtQYfq9fCNnGKETICpJ4YWhv7AhBpXTT6zyXyYGweKHfDWQ6vyJERkAN8PGyagLujW2l1r
HOxW41gwmxkTTTDQ5gY0z8TYXcgv0wZ/4BhFFVZzx4fdODz1ltLrjzhrxZApJPIkOdnJd2i2eQmW
KzghybDN6ui1AcvAVF/sIfnRuS2RleXbkaHD7D2uu2bSkqPZsubt5lbpRrI2D7zHSXPQczIm9cDV
wtnXD/NwmPcjCa9ibB2CfHVzhILhGm1nJZawezwjxem3xIomrtoqQgueu1wEFt5cceE8W0Xm9s57
HiJ1b7rn47XFFM22b/yeUe/XLCM2u3A84zeB0T+ihjxPqms8yJ/gJy2EZghYlXK1CD5Eog243+YR
x66hNfxpo5KsAbZhaN1F9RnlYVtL7HR34w426CvNEnKwEoNfM/R4cT9bhPZzN4QDyr8FBuhuRKQM
rf9Kd6Z9QGmA1JbZ5WJ0nn2t1Dx/l7cU0T+LnoIQuK4vC384ffb2yuDCnk6nxzO83ztDVMZqYou7
me0NgGgefrXvxs8szwv53Z87FGH0cNYMXMpbDzLm3UB6Q3krWmNQP3zdx6RpE+VAdtuswYCr0TRM
JnNoxauyhvhhC6M7b+xE+PoO77+40NvndffyD73EA/kIOp5bnABVohRuZJbbl++WIPHYvD+7T7WH
WClpsvSV43++VYGK/9pEwhPUqtg6JVMFwpyf2/awRpVI7//LX1p39Yf5RgufFvqcCj1pR4ODXeut
49lqdgM6qcRwgW7lJ/L8rj/P2NaoNUIeINYHb5MAvwQxKoT0X2tV3MxPso814ZiWp2ehWaX9XTaI
SPisgmpw1OyapERAfKTvs6TWJpS+LyN9SeipQxReGZk4Rr5/7ccYZL3QtZA/3It191C7e2av33D/
1An7SzPSWdt/bexdX+vQPkyHUgYzCsCERXTxevOGX4R97NwsPt+YK8U785mMZmzvXbsfu4z8cJeo
BAFgMFsp2uVZu/8DK1R9+IgVReD/BUZha6GMEY3+tPISTFWts7qdKouViVa2skOMLZAHgI8nWiM5
S5p16ge51033Yg6dvGJReJfRLawCD3zrwAPeEFD1sX5lZYp29/MLohFTdJlHnnwzsyoIzDvWIRLU
3speYAASi4HgXdZcAGTMXm5NwDvHSe75hk1f/yD/koDCTXJVvzd/AsdV7JBXDTej+exB7VXjcrW2
m/E59xmVQi6mq0k812OWAHZ+/9NQnQbMASu6qGFkiBaEoojyduC3MKKMJF7j+BVr1TuGrj9qk3Kp
2QZfD6gRa00ulIeb3UV65ENLyypVgkLq9GSA0jLw5lCYkpLbdeUzA3Mjiop7FV03Xpudv8ZSGjJT
tzPNY2ssjRfGYqyDNb/si0qiIHXVqiKqWRSB7ieSOSAnHMVEOI7I/mTuld7ZwcoVaFld0mYXgPUH
NtOiesZOE3SMRTyPyl85UNLp/m2g3l9b9dzgdLST0+Ar0zognmClC+T1Zg+wIrgIxuwuZxYvqn3g
E3u+UaNNluoav7SKTYpr2oDz4/Vd1ArqALSjZ5S1mO/eIZw62almO3k5FoWXq5YT6HibvAXPjXFX
HLmr3QFBHcfY0vLDd0Rbb4a4CAwL6Z/n+kzDPi48g6XiKLS608CddbdHxvnQxMKi4hsI58ZO/Uus
01NIOw5gb3FjtvoSaXvwpkUxsBEktzhGd3Fi/HfRlHUFfeHwIOV/tsbVlSrxn8VLwaDqh+3K6D27
FGMmKnxQTbNCYm0KhoUfxwifzAdEXblQx/D69xQJ8A/Um5Fmwfp8zgYulrjVHsPVU2D0jzAMvuIK
aoGluv2zwjvUuJbr9yjNqheLMceZCsho8+QKREO5eDZf1poOHI5p95YcF/2U//R/ghHCwKO4L6e9
EFgxLSm1K6BGLdJFLqsUgIhN7jaeDiQZGe48Vmc51rXcxE03i6ACzF/tnIJaNDMQX26+KLtx6jL3
/fPZb73IH+2Vrd5Rn/IWbrKQVz9n3FDM4YJQFP8cBOAv1IrUcAl0tt1bo3Hne3YEn7BQF2IoJGHG
QZtRapKBaVr9+8C6bR2ro5F0dOUichWZHAswbn7gsjH9c6/I/gXnGzfTshhnz0n233UVA10+8qU7
khYyCbQPJwjpPVQzFR75gE2rX5WDtZgKqlioKPmB687wrmsxsn0nduxpIEW4pHtPbvfl+3rEEKFk
IUkqI+s+bfpx3PV9EmmfZkBKBf1ByVcTFvO6u6GhQtRT6JPWfaP0aKiSGaNnno0OrvDWZFnStOyd
dQl8TNabScNny3VFWq8fU/YZWhidfwtTTTArK9L20YtlQNFIp5cYoWmSXGdnao5UfRI3oqxtBnx3
OfZ5mBsSpQhavkKO/HISZ84tfjQfAr7Rc0SbtU0OHGguTgIICSbAF4GrJ6peYQ42vYaDSsxcFiYu
e4IlSYofjl8JsoST2ya90/uaXLcgr4oddcwaGobfcr+d9WxyXAepwVTQ00L3VldqKIJpbI8Z5+Zq
IUO88gvetIBCVv+tBDttXoxTe3JPKEjXjmXxpKiWQeh5mEoBZhBhjgcTlIajymh6sO+/77O/Vo6z
lOlsk1AXTwpag38xi/S8Cr2AQn1NN1I8qkBU5CFGHwIwdohC02t49ahBMrUC++wk+LzvQPpyytll
71m6n9mNwMwIs5knPS+/BAmRBVWaoTOIF9QCh4bSfuYZ8Tzw63yEGpsuvaY3SEpDEu/MwWuDlDmg
ozIrAilnwRLduo2L9M8UdG1qRxgt0a1+qDD2IO4r1j+dC0K4MN/Gq/5Nx25HR6bm+2j5h+yitTFN
YZkiJeRft1o9+y5k9ynUpCC0ETTJxMoMQ0+qftIf9cmuqEmHAsHfqr6fr2ArXyFacHK6HTOA06Bq
1VVlNoyW8FrKaMnopQe40xT5mr6WLIgaYRnbz7pCtImV8uIlj6FN/jrhERIgfPBndQQRyVa5jnFJ
rsi3RRSkB42E+Mnd4kqcxzWjTGGpCtRR1nXT1iSzIELLv9+867pyhBmqOGP0p4TXhHcibxqmJEAD
urRPP1RPFuUgtdWVRHP5mTFT8Mv2vGia6danDXpWTLX9wwrmZ7CxPPGxagul79iPNfF+GnnAD8JR
u1qzfxy6z2k0m2rT/gcszdGdRkLqV8Ue5ehniwQ0mojzCeKrUdbodDa019zTkW4abTA5Zb0dmc3h
AlqOJcvLVvIrnM8ogz2hMGCXZAzrtFmElP4YI5FjO3AYnysFOrUNNw7tC124AZygxHQnpKpQLdoF
XUY75tZaPvGE2PBJvdpjjOLfSraZoR9hLFH1MzdHa4WCz4tq2tAKiPtAAac8CIx+qLgR3Iz2AUIl
e91JWzUIivPaB03RqR+OC63qbZK5BgcJNNIj8iMNzonrrNMA0iffhOZOtzF+CNDsf4Aftq0Pumfd
y8Fa1wF93y5QDP/MhyYjxsMf4Vo3QnIu7VN1p0nhUlnrtZ4FWva5oIE2i6QanLiJNracnsDYXwb1
rDnlEg9oIlSB9iOa/v/oAMuTuD3Q9Fw3mekvR9Qailezcae7SXV43mJuMnWm5Zy5R8+EokTVEHpD
OJrlFHgelGEbYYNL+VPcPSD2SpTA4xGNqG2Ytsfwcs99GHi14a6TFJ+X+/r5tHmW1GE+ygAdvmXs
28cdQVE71bf+VxehTGkNFzOiM+8vCdKQ3rGtn5B7Dc8Jog4CT2peeguWgcx3J/Mwpu4fX7VZMvvg
Ect63DSN1y2IkirrD4vszCxOTeYkgGwog0MTlEIyPL04GqglERJCwyaa3qFDkhVdXem4rWl9OYSp
BnGUixP/c5cD+eRsEII9cCrDKdK+Oq43exO+67lxcsQym8/64FyUOFjbjiTSZ/V2YTPf2Zin21AB
vZtsuzD9m2Uf/jBreQACUu4RrCSRksWGqJgeKKsZFMW1c59exPRDZujWty7bJwSw1u5tcx9nPzJe
Yn9ZQtpdALfFEpmhziWmoiVw5vN5U7+rVkJ+lL0Y7QxJ4CJVB22FQHjIuS0qbDhIO5czRFOTYh9E
lGOf88+nv1jhQgQq62SJCcy0b4WKmzDE/8zI1nwjS5XqsypZqRKTWRU2fc7UF9z/bdsslWwbzUQ1
CCF7HI9vqjTM8cNOGFFbAjkYiau5LGTEsOdgC682vHLmOhbIdOUoUUuf/qD/avA5oKEW34jHAExv
oI3ZBnuK8nCRF8zQwMllJCdf/FI9vGyhE09oiUZ172zEcU2hrCi5rjsOg7+S0jtXFQGN0ZKznlIN
gltlK2R8zfuvGxyVEEhDdr0zLg0e9hELzDPrLVUHpP0xC8Qd8otaMyo8dkRZyLHMj3CGpU/9fc4v
zKs3Wl5abmidF639DekViU4qMy3w0ljZcFHbO8+nx7oMHGHNU0swmAIN1dVpmSZnIEmablVCVOv4
k1c+5reFpn2HOr+BuIOOhc84EA7DQnHAniU2W7GnXK41KfpUs4e1Ynaf7KEROsK9zJTWT58fg3xg
YWloPhphRtPgn4YGx/Xswb5MboOpMKYGUiYasn+/pFBTjcn4I3JPEv78Kqz7T+mPe4IYrrcBY9A3
hO1537dXyET73i9uig10d1ULkdxnKEoMSZyAwjBHZpTtU01I/ZaHYwlRnveJjclJYy6c6ZcXLntM
5LnsbLbNrII2PYK5Uj7fBBDsNjXTZTCV1kNWXQqhFTiuSKkgvz9kc2bRjPVlceEECV/x7gA0eu8f
+fAp+4peY1wGj2vAJYHrFT1irg2r3Haf9E6jImOSU8R/mfjiZrm4CwqnZQDIxSpTtaHLOpgZAigl
r+ggwfmJRpTi7jC/I6+UeUm4zXgWhlzrIq7UchPLdq6Vj+HBCpFjtRtaVEx+gRmXQfsn2JsjZ7c8
/TdZBB6c2HOj1+IPO9LMtiEFrRAB2tjdBhyRcxW8Qe2xfqTnkboFQa+nma1+PZ2LpV6S0UbNSogc
WASFshWsAFRcPUwNCQzKveM/9lXw21TjaMcyncrQARYiFa/ciJUtoI4V5Qil6u3RkWz6xGot4nc5
S1b6ez1WASI4p5K5Mhc42txPEIa1CemUBGnlTuiMcC5RpxCf40La2ViqVgtSK8fDuWcRdSbu5dMK
wYQCcejo4bYxQ2hEKAmEP4qrGIrXUrCeeFQP+zxpOl0IRXwOqj0kVokyiF5QuZgdVbc1af1IlKmA
++gsNbTEZhb0w3Vsgt2GMlKviNwud32RTTSnEBzetwb4f/Wp2WaGcbFEOMWZ0K820IWHfUtRpi1k
hTiAZTUQQ726bMqlvUJcYxP3pSQZ6s0ofsyJuDu5+kPT6Il3RmxhtorwUVVwsGQO9GNTaCbyjFZo
dgYcz6jXFGwqJIj9RLiyW8KKft2ybdOx1O6yZroFufN3ZIN6ljJaGTOIsXFklEncuItAwz0+8X3O
xqF1gr3+qJFUgdcn48Pw0J8Re7VFPi+src/yLQzWHi0R50jt48B+Zm2jNCgzTqGT0rONg08hckEU
UqVOkyWtLMG9YLpJSxzVIMvOLft8gfpBrAaya8USY788KSlgzvDwxoygnedPA2ZjTHP1S4yx5SvM
44J0olvO9BJabVB8OYdUtOcXkr32FI/v5vy1qbHp7/6KaebAXSkT/BghkkbMa0uE3FHErexvKmAO
tca1ooSueqgGGD0T5uLe/2ygbc52heSixOAbQtHVEk+3xsWxGIjYZLHUpwUouOVzWPQb7AmhrsFV
g42pivzc73Ns5G97SU1iOOwLa6dXkBXnpNAD+hrgu/8DREz93aYjIyqzTbWvVizWFcxl1af6LvkL
ozOe4vcRWgGSob7nwQZtQXzjMx2FQueOIbnhO768d9tP83f5vwtzLTarRvHqcxY0qHUSyaZg6I2z
nxHfoUJn1SWrKrF7A0OMSp0LjCH4V3wlBYUUMYc3Q7JJpeVWxfmnmHhDMJuX7JYUP7Uur8OpEGVo
feWVEH5FBd1vVVCvn4RZ+YJgkPFFvZ0XJ3lH/LE1mHY4k/XPxP1V9QOHV1QIDNI2r3gaOrtnJiFl
weZ/fcfV/B5QtCbbN6GEL4SARbd5vnnaCtwealJjN3+iR12nvr3EnPVP7lAmgYSy3DPX+afbYK+j
uivMFl7IJn6dfpOhmQRG4qDMM3hawhrYLc5jN4UK6dHn/fr6MHk3dFP5v4pgOlVo5qOeoswpFmUw
mh6VmSYtSPl5/ia0IXiisFr+pwXlo5wa1f2BdqpMXEGCUvrTO7Ve3g1RtqOCN9MwCcQfPgHO/aOL
MkZbddFwQSvwIiTHE5pdcFWrE5E1ljJFNKXO7wDnMALpbK0fQqjwKMSarCdmUhSdOF4PHTX59c9L
zEmhJDMxDSUKDv48DKimbusBC71+RZf5TAu20ZjuseGiWdN3mW0xRvaI2BF1h/bds2ZYZzKx8CJ1
E2D1csM5XZWG0+VOXxC7JHDB+nGPYwVqCCS9yKU/EyxR13cL9gjVpfgswYwEvVVrozMxlwVSGbSP
EpjoDvGzvq2MQhNnxWseO06t2IqXOFErxZ+GHmj/mkAS5Ue3khnMVXhQVZQwSc1gkpYI8lDjFxFc
PlcXBZVQzQG1TRNRciOz37bYj57xXo72F9b83C/ySYEyElWjd50RtD2yjPXIdvTMg0vwz2sxH0up
vJn34HgWuwmP9PjrWfFWNh3HeVHPfFjVttBLSHQXM+6Fmp9UD0ESwMD4W0cXGDjIdxyzodgHdLHC
I4WNMkb3dBX0h1VBG9Q6mZK5GD0tbpppcsKtBqoyHraAaEBSNrwo0K88vTCj0qMgcty7MfNDgK4W
6eVDAyHdXJtgTQ3aaEcchkdc0iKvp3I9zDP6dQSYdjpjoeyb+/mD1UjONBhwRZBfsR+sVXdxMT+3
aVFm5xOhsmfYxxkO5ly97hkuS1JmzKyv/lP96jVolpRX4c4nczcfPXuCVSC0HvrrzTk9hoWLgr6R
LgGwRmXB0InaoNUX+j1jDlc7gjHz+lAfy3J70ketUYYLBp0Q8PXLN7L8iifgvMat/RZPhERDVtj7
cXPpE2ThneHJg9b56zCpqCuAbFXOagiw/b6uYW2yUrDYkrNqBFgtPEWIeFGLfgBmjou1V4Y7I45P
Zkr8Vwo0Lc9Ysl+GbXmFa+tEiB8hSlDcFen4PWCGvU/pfd7ELky4TqbwyWskRx0HubXwxoOQPfW0
dpKtudbsyonG/ShZUb4tHEgWq+SHCIzBuQjLSjtFCyNrjN/1/h3xF5l25Wnnd6iRAcRlGiKb945s
8usGghpoTqG9RNELrAaVMHpOlyn0eGZQETiREFnNE8m2P9QJ/SEzIPK90mbGIccJX7hquNa3KnkN
y3PdbncKWNS4BKcCYmK8ra9SBy0a5TCBSMDsSxgxMElXsYgEI+LdO6rO8bpa536WRGGhim7ASVne
YvWoCeAukd4ktQcf7Q9roDuMj7s/p4gUM20Pc6IcI0JIYl+MDWJKwC700iYQTsT41kgPM3IpwUO3
T9QJL6md4sPpMeLkwtNT1ZWY5+HZBHE3x/dmk8JXW6Msw7HvIPUHP87kF+nTEo1CXEezWzech75p
Xaw47WeWT/a4M3b7sqiPQkfxh9x642ryvOGv1dtSJuLOrAmpjTGl2ysAX2jt3dF0zcvEISlIm0rZ
SYJhch9nU9OIVMaSMf8udFEtrk8vwWaEwYS+zNwYIEndMOK42/wraO0Eu5yOIvbkbzQpOjTdwoaS
2dvOAa4wBPcDTQf7fsSEKk74X/IUx7T7WQjo+6QcdVeg0CJ4UHxeOiWJLePY8xV2T3H+xrvuLosh
wc9vGI0dPM27jSNCL+3jCUgSMfzl7Umb4cYryWRNwwnq3VqX052msGnZXBflR58FiGwiTJD7nPQy
jCDlXJnhneuWiAZiDJKDxd34cdsSbM/sZJIOVlo4cptKq+D5+iRNMuNBu8Gg5WibiSOERxXHc51h
39U+4GIBvdQyWrGEIwfWdEBnueTkj0CEazlyFenlrcalL0xEIOwFzpWVKC4iFzgYtiL4Z+S1dKQJ
pTnKnsdt7/91ZcXW2YvHeapy7KQbb/+iOXuknekmR5QbMW9Gbg+2vcWuWzNu8J06V2+KO1sQGrEt
xa0T0zLYmIUkKTlQA/8qJ40RVtOEukerz3/fcO8QRWvjSYRxfQ4+nIehWt+vwoYaqEs8pY4GUiYP
hy80hQJR0NR1ZNjjEHRTJXBgJf15h5eJ4GgW8vvwz+Q6h9ilNfbIc2AUdw7MF4GZYZhafq4Fq2qI
tlt3OB6zkobJu8Mii5EF9NplrImmwRTI8zyzaFNQtRn33oY8uRm/osMqCK750mo3KEFkYC7c2MV/
tSI/0IhbOTaWYv7n+O3YLU4oSG9ZEgL4LMF45egzdsLQmk9jA0M6xRud5xvEhYJ02N/Wxk+R56IX
NLDaN8kwF2qRX9QarRyvjzmTp5gR/Rj5k9zKm+1SFqOCVOQrFRdX2WZTPt+BO3VmOAb04gqus58Y
3gTJ/eRQ377/rmKdRBsFAvOs1CVvHYnlQkMtxV2tRORMI8z/fdBUB/rUvq+jnGb/dt4M32Z05Rqa
B8ZzjhXEKSx6XDZ4Ob5e8Vj1O51x+G/pj8UHuC1NdcDW7ConhGNg8T8dGihw1dtKQMCHNd9qlmpO
SKyfbNQLsYzidsRgyXXGrnZHJBcVoNyt/IvZprqAX3qbLDkP1LDeB1BZkCCG6BxAbTKkHcaMMzTH
5TxWXaOnL7TqFJVAauUSZlVLqHrqqe187yF1sqTceNqR3FbW+wG4H2EKrdcjdI1gdLqy9oUX8gZr
g6yss3aAQFRFCpTkYBBcpUFP8+hFGqGirrp18xPukRCjn3BQYtgqIDQzXqnaeDKlOvJ6VOmQA4Oz
F6jkFQT9d3AqnoIN/erCgQq42QK6nKWs++lC/NlU63ThVm0kt9glEovBJM5+jZH4ztUZdPOqymQy
S5f4bjI2p8L/lDKyvtpDlwH76cXGqdWpJYTm11gcN9W/kemrLsod3tFP+zkHRXu0+pwAaggFRScb
U8tslrZ5QyzlCbnxum9w6vyqSNlAseAYCLtHL+pkffFanN9Omn7Ej1nutsk2Bk6ALNCGydwDZ8Fs
pVfKlFA9ZtO8xqGBA3GmquLBJtEjkwvC+S4JGByWVa978RoYYOZpDc+XjOXQ8XJ7Ow4g09trbk/g
sHu92DuNEeMz2AzkuUGE4Ljisc1FiM9STESGO6cLs0YNoatTaCi6CmDLesfRpsxgOxkzQCXk+hOU
t9Oh7fYRuh+mgwGM7kMPYCncTkrv5wBqeaMAlkfioSkPEhGLEZyAIdKhqvjSE2GK9QUx+v0VnLad
znI7rWdpTVlh/tldIxTWKZGLIHXlyNi573t0ULdVfsBx2JXkfvrKp+u0QMrS/gaeSAYi2Ic+qiBu
O26wypO5mWMWsxRy7AWHTQeb6YVZU5oeipndQSWilMwXyiFE7Z5/jONamXbn6wnwD6HrdqHMmSNy
sOwCqNlmH4+IkulY3LT0cIOJdfH8VUYuz9IGySaW83amgUM6Bz91+XIPjMv80+zC7zOSRlHpVTgZ
tF9RqrXX6+gPyxr+vi7idEo1jUe7JOwmC5XUBHv71v7ONF7h92bKhNF2+BkNsKcXb3eTDhiU+j8R
oeRKG8Loj3ttrJzy7Pvyjt2jyXmryw1dxH2IyAelTEaYu97qfb/0vD0bwXbneFIkrW8hto7N3rAm
BcYLzugfk02q9e/m8zZhDMGY6CWggj9ZfUt9zJX/fWUPdlTtIoYVtIJgm9TfnfAuOybYyC4rh4MP
UZI9O1m7BsxEIXp1ljFQfqpBgZ6UjQx4xflVJHGOz+9peFpVgY/xIiEgT5s7lJUv9ZZc3QFCVF7i
QxrAC8fhTX6F/JFaFAkGrw9L1kTGwZDi3alRhhjKfEcI4HFeq9ZN9Co46EhdJgTrtIKPz3+pll+t
a1G1DgDaphspgII8yQ7mZWrZ2fWKf5Fi/Fxo/9XwBH1HFpo4asPHlZoC7XrbYdle9zrEDRs9Vb13
1A/Fq+hJTptKw+7QkdaE4GFDyfCoV5ZX4wkSLqe6q354uzl2SqXlX8SBPA/gDFGCDnDs6BHngqfh
FgJfbO5w2OF2r8d1Rcq9lovshpqND9MDjxYaAYfcyLmW7p/P41irMdbEofsQctqsLUVvVr9FI/uh
NHM3vwYofkqQowZBwU4kj7pCBtgYrFFnmBbsMW/alKsixpR7qjBHz7o/YvvpjBMYK3GUzYUG1J6W
AiVXVMruKTNuyU5nSGkfYrAZZTGYePEH0KgpOrTOKUn/Yb+Z0H0+EqMzo7Eu0Lzf8bREiKLwMhpw
EcJmMd1lh/Bkx/aNH7BBd1Sij6S/PDhPrVijWcJ7sJzrM8S1ieZFbavC2fHduh50G2yV66+L5JId
pConiF3vvna2L29pU6hGbKXzVzzQN2jqfoueFfOs+6+WBEk3N+YZ+kNpJ9S80aR0dGsWLcM7ZTsi
xob/KDo4SC9XPWZkYn8PAFDTCNZ5hd4mC/RvtkQpKt9SKNqOvMnBycY7Q8cJDXzpnHp5nRu8LiU1
elt/wG/TmgqILsuDV1mzhdE2UizjJlGC7lCBEowthnx+wAXBjusb/GD2CDGvCYnDNx1ZOOIdAWZN
2BTZ/qVMyrYj5LbsgnsPlMpHmSDmezr31Y7uWnz1JhjTxHyzhdrg8gu+CAIMg781/lKWiR5eft+m
6pNqOl3TBSciLiqUY2GitIpQavjOyNmP6UIWnEkW8bR58J4ffrgJ3sr6qw+IIMHmUx4+7hLoCNtS
j6uQFWjXZQeUhr4kiqrEP2+9tY5jCVT1IIBIxSwTBnCrv+aZAePmVqgijGMuw2EVgfeA0oLIHybG
p/5pX+7HghMdnZ7F3jIbQ7iyJIrU+FF3fHOrlN6ohF1GgcqC3nspn5BBcGwbekaEPK2VYd1ZETLk
6ElO5NUL/WSNsv/D3V5rXlqKA1kUuqpMogZHrUDbwZiVp+f0fQxEDXSzXZo3DI6Fysv+orQNBVZD
rRdpV7sKwRFRRUFqw4c8HZSmlugv9EMhZpsqAmjHE5Ai1EDPnsGR8sXPH8x5CrJKLiKzE0uG3D+W
USq9rbUDEQdofyBYRH7nuG/bdGqJe85kMMcmmerAD6CAhKUpHZs1JZoZELVlPm+GMgygtnNA6nyK
mGaEWsSCau4iK2kMuz84wLNRryvMIsvvN6ucESkoFGBrH1sWGYUg8SkQkfAA7UKlyrrxMgfYpgPG
XfrWlUP0yjMKXPNG2/HfBpy0sd21inYZP7OomlY5GGroykITz7EAn0l8Tz8tbCcaqiHsOLIzx4XF
ZYESlWGk69A2ugwb0xwc1Xy16BJZoaRD/6PbismWe2fIwdNoSWTCERykr0/c4+1Nc5+HUIP+dflS
zVXo0R7SWXQ3oi8sHoGU4EtOMHPlWav4lfxvU52i/gMT4etr+PvhHWQapAsw9R1NE8bo1xN2wnUg
Q/TzZq9hR2w65ArW04XWV1zPBamnjrZG9/f3fFpCs+wOmR2LKj2CSEQgHDQQTnilxnQervy539p6
Z3ZXSAjd4Bg0Sj1FztW6mbqmGsvvrczjMTHmkDuOyVSakumYeD0K/QDXNJ3NeB2g+SbNogbXpo6o
itLPW6yysmi/xqaFULyP6IkEUvaj4iDuSlXTCfHjxGXRU+LOEvqTCxTjLO3hslGITyh5N4Ak+aKB
x4lEzvnGBmPV4wVup7gu1bk94O4xl8/fo+n+u1Z/dyb0P413vxgeK9ST8lpNtebuz//V11S6WidB
IB5CmST8zL4pTrBrCmyB+r/7X+HXRdscsKraHxI/seVeAoysqYplnSbrNAnIX0TlvycujZry9raI
TnjtSvZpTAjLPgH6QMtas62EtXduTYhbjYLHT/YQNob5twDbWs4JtR1LeTen4b1fiCMLjNvBmC2B
PvJ/LIr8IuuYKXE7x3GNW4dbagyO2jrc3gwKKNjwU8k+af0M7G3dAevc6T9qY0G4AcVIGMT8OWE3
9uAlRrBDPB62vCjENKRCJe38NcLwYcCkndzxgb81I+3QP0AGkRJr1YAPj8VFJ5kE5GuLvM1RMe6c
QfIwLh9JqEx3odiGtL+zwdzYRih0nh/OjtWp3xTo1rLLW9CrMr/VBDrGylrsYKOteAKcjRQw+Z9E
GDUPgghOCY+oqKMsX4PQ6JDDsn1pGrpSC7i8zQh5nCOfWT4m/VX95jctyffguCjrpqOy+lfA5x8c
Hb/zq7mwHofKqUdqwYvAiegilJ1sdpZhz+FZKj0NYsMmA07VxaCykrMgOw5T2JCf1UpP1MGlq72V
oMJN0ri/BgGoSK7bwU1AF4HxdxWQoU4rFWZdLdh1yagSt6WW/RcoM28VmnvlmAbQmw4nUcoqCwun
TqitrMPk9LEFwj1bUQtguv5TUm145FuM85FxY+soYtgUNljaUgWzmj5ynf6g69dA6BwQfgouuzDo
on1z9Oj63vEZs21hgEIiMltdKSxpSPC9XfN/Z00jUk0pawk0DYMHaPAXj8PBPnO7KC03yzMPmNPi
3zkCbBfdIMzNXLIGL8kjq953+0P1Aiv64PtN/0LEhYForqG+hYvhp2OnCM+tkPjvcDwW+K6Dm+FI
kNOXZKUKtK3LvCAzvjCjMSR8Cg5nxJnUyV+Qr3JMBMgMhG4k+5aciPTH13Luv+E/hFJAJvdRKLso
RQ6pNfKVwi43waiWwkAQWwVEV1cgjCEWLv9u+ju33MBEUNGOwhFMLWgITgBQ5ekSuUBqr9jNs9ED
GxZ9oIunlTxBjuAXbsjXN7qstpeMpBzL4g8UJQacvS6jV55BGHVRSTcKI6fog2+GvgzvR73SOYtG
XQH3elY9t18FUA8R/I8ZcLmiG4wkUFXuJXvqG2mXG/bbGVIcktDBZw6Wh1eU4aR4LoKw7JIqqBkD
NDXqu0fwAqVPLGY7pGedXUdrO3OaRJ9qvV9Qysus0lEdMkeSJ7clNlNvGEaB5QjLUftOoeEQ3tiN
s2lRHE0FT08CGxavZ8UAotUBEHzhTUBHKFRiQv1RX33SrlL+RVJSpXaFGgtnFyO50ocqkabWTdHE
/wZQf1SkqM4a3K+R4S5qciplC5Y58e0supTt5yuKpahbkTV5KjsthDIqoA56Ahxis/067OK+j2jX
AVLaoXFh6BUgACpcbtbOjTD+X7g1tSpD3xF6KcbhVTkLtIsWcmb/RKw3AlJda5RxsiZcB491ZXuS
S1pyQvXEkSrUlhDi9Www5ZKL/ZvP/5vfVaVjr4oX3UalASpyXkDR7fdYRZgA2u7z941D3EiRBVrA
7J896qPzCSBwpUQpA3LQF6kv6ihfipBnm1i9gq7YIF/fTv+1A57lnmE6fo5B5mQx2Nj35tUDvbyb
05MYVV2nKpBDE1KtlBtS139/ze+Cu6cSdLetbP42NUTkMAepVfmOLs2ohPXDttv3pAOx89E7FrSh
lpXvVbmWQKEKzHfB9Iimy5jkFHF2bNFCSOx2IQXwkEtu+7ZoEGjtF+Sh3HgSzJCUHi0GHW2NiOzw
x0kG3I0KNktmxR5ygLiZsn3zun+xPWuXiEccn7rzhcAlS1w2g67lyFoFSfg+aswiKDUbDdxUq6+8
xWJV9fSIkm3bkuRHFQTqAxMuMmKaRX2mLEvGKBL0TyXVCRmCFlxBEYkxTAbzwyB5url48VTtoKWT
rCYbXbtnky6nTqQ6ShLaQFVXZxnMFvzdHxIpsdMzNkZ1kamQFJEkUHvII+tz62bGgFVfoih3mdEZ
B5A3Jeev/vVw4I4Kp7VGm4vHvR094k22b723Y+/nJbavFg9EwNrEFJGqvFRqE0OB730Hcifx9u0D
ojd78mSrixmNsQ/d7bslTL47wuuU3fZ1l4op4QXTD2nJxNE9FcKzGIWnMyjNQiL91lYYD8CFrfLH
NCu+/lMNqqPIy0Y/iR14aMKiFrtRw/IJyL1QVQSDCJsBgwf48zBi72mYgFiNQnOCjw5VymsHSTdj
xCRMfnMVV54t+Iq79olzF6jLMH1A5Ac3lO85W4aQk5n1JhEj4lDWgggnpIQljK2NKju0uIYR3Nmi
v2KG9/tqFTcRpKGvQ8ICtuBURZzEtCHumESNwWEAi19lVT8f6BtwhgKZfuz3eWwaJA3CqWmrQ/hY
zXJoZi1EECpEvmnLN/ZP468h7HXE1HL1MFDOo4cTubU4JrUg+jNGaPLYPU+PifYUUBFPVRXJ4SWj
IwykIfR28AzPqVrzXNHGzfN4r97ZGikg1H4HU/e1PKYL5JWn0chTG8UU0HsducFKK47DQRhNU8sy
KWYcVqSvmvk4J4dYfcMm3jdV57LtNHpyJrsj4e5sda542eO7wGijnERL26GXrf3NVLYUTskJ9rBn
TTHYhb5j796EOrKhbN8WPb4qVxb909OO2vxS+TRhlXv+NO1bgg+QZdbGo4TMJivXqf20CmA1OITH
0qN3hzEpiIIagINP2qJOy/awyUEM1UdSiWOTSfeP3Mq2UzSdbRIN7pFz9T34DB9/gmZF8wN6YtKa
D743G0EBVmpwYN2aqZyYtnAYw2uBA/P3HTnyqmbC1iA7a87nkJ8eYwvnfzGYP6jYS6i/vZ4YnaLF
2bwDLoeIdfBTNRVZmC0nscw9eWCyEVjsDQEUlukPBmM3t4TxaXigSVEDZiqIU9WD3Sblf0bYp0yf
q3FhttmfVVVB516e4VHO1ZsswBRxvmiB2adKDL4FJJwtZycNy+FpAl6svZweBzG2UqU2a4Y5W0aK
PJ1YZLauj0qM8yy5Fat86DqqXYfxBkJKUMoB6yXPto5Q3xSsC+rKZV227+8JmklVBwmf2t42wWMR
BpuGAfza18v9tjPdrBnlJAPAhiMES3OBYopdkKeCfAImfgnrmgYm7gLXzuKQcRRUmfTd9ysLkQgX
WYPhBp6UbPkRKONzgqnBl+dbNps4LiWOVIkwmsbFHotncv0vuVz8Bq2B0PdNyY2uBeB2dxTO2DDv
q8XYsnQTAyDYA6EvB1lYD41myDbmZiPJ5rLRRGiBRnV2BB45yyLst2JEyAwqZSeOnsX6+znhqVMk
PaOsEupXHG0Nqd9qn/DfwCbsbswdtLanL/k4BLOvKYTOuytcuNXKdXv5GDhIQNzO5UEmde8Zy3nb
dapo+sda/OR+F2qAktEKA//aRXAU7p2m8o9pB0k4wXqGqukCNY4tUJcoaq4oRb/FvtdsyGrYE47D
hsJA3XPi8wuupfeVWO7gO6gJrZ7HnyBSFFyYMEXSQJtir/y48YYwPykOrpsygeu3tYtc4LffxovP
Z8Fc4s2KQbYSFGo7dfuTvsLuPv3Hf+Yc7BfJ4/M0DZg8Y12GZ1n+owwKPWXAx0kW6czQiY6fBFtd
mWESE+0tTVdcZHPIipTgm5mgm9xN+huaZSiitcSL+l5sNpzP7o4dRMn/7gKS+9yzsb7L40FCxTNp
N0ds+dHJfQi8D7k14mJEZFTUedBSQt5XWNZhyGEZgfTYN3R+UmPSI/b7E9RJ0qKbAXeBV3CbH1Gu
v53HoqFlXJ5WuMxOTht1Skvv5GpfiPr8T4ybfNgKgstn7iSgBqIWBc8tmtK4nwiOUahGKjaZ96/3
ezkWrZ9cqCna4fMDEDJVPZBVjhMMjoTuPkJym3BPXDPZ6yeIXeKrJ7gCxOk5zyDJKiD0uofHGkp2
IkD8IjHw3kAkfMj+hqroAQo1qkN/FfpWq6UIkG2yRScx+tlaeJ3N/kW2Pij4xNdBLx9RNHmef6oq
NIjy7TMec/g2ssp2QJdvb/SdXkXrUH22gg3YhQoOcDLp3BAXMSJ0CuzhTA0hEWdtImqbAFCIf1jC
vRyi+Z13+lSAfAChI1RXuLcGZrSVGO2Z4vtIIlgy3gpRFPxYermdM3fuyvPjvXUv5sh1NyIawBtC
DUCt3xzXX99iPjX+s7z+PEZPDWaFi0RhGrMJz+gPLwl6QN8DtgfDAqHvqXdWosafRLKXuzpDeQiD
FMckT0qGS7JKjbGey9Asgi+HgvgjuKSlu+6SQoFx1CHcw7uxpR1bZdg4gnhZ+bNttq/yvZ8J+Xj6
iTFX22z/nzBfp3GqPcARjK+8HT/5RbWm2QDSHNnxaAlNk6o3shDRB4LWgHt4vCCbHgfztZRvzfRJ
pK7Xyh7jOLjtv3Aj6KJdydbt1OsZLSzb5/ugOIl4kdOp0WurbRv/DXhHLnxStz0kgoz4MRXpRK/t
d5KLIS5fT1kDOaJRXvvx4f0A8+Ivy8Xh3K34gsJo6Ex28FVoBcZWTIabtphaB6gd6kiVTG+pyrVo
rQJbVxnkXRs0IGNGQhQFyT5GLSJ0AwTKFeilspOYLm2AlYkKNzhUTmEbTzkZNCTTlphvso73y1Mh
QOKVwsp+xVf2zkbKGtqjx3GxcekhT5aB2f+LRAca0DE4GzBTQnzItlVT9VvmDrdt9KJE8EKpGbFh
RcOdqkrx2hHkQNyGOpV6yZ3O1TRlymRgeuspks8CXqC5NG8huXNqdoVbAjN1K3slfWXHkAc94aUA
qTMhuEfiiAzA+pyDKbUERwSTB4Usxrr6SxLu3Nn3p+g7Zif05A/NAbmNLYZ8+/A3bRf2+pCbm0C+
ZYDwMsQ3b3YanwLvg8PuJyRf2g9NnbQ4A8FcxQU9vJ46Gmu/lJr+fvWq8Rnodot5eBT8QAzWKVEA
zwTs1dp00sbi17IqjZhPGhbNYX/1ck8o96Rb7LkIdk4RdfviotxBS4uusjL5WvC46B8Yu3qmGVPz
cxfEYAqeNFdXDFkWNKf2+g1HDlwi3f+Eht0kL8kVjusCUUQkUtp6M1XnAbOF8lOnvKeAOfFhapZu
jxcrrVWd5xHYNSp+RvoGnS7oC09HTYD+mJcsp/YJOR7em4hEn4ZTUwud2lPTGFIH7vZJ6/KQtIHj
JMDQ/fUL+xLdVIGIy8q4QrqMej2CFeoiWDFvpupp8zqUziPj/QPLgfgOmvxttunQUYm02t24zLG5
fbbEZkWk5wN0br7IRtJKi5NVchYdapcJBG1rH6ah8OLvotWzjYX72Tj1RRb+K9WmF4h5cJC4Q4ET
7rJpDaGUfXOhr36u7oM+XWq8WBobmY+W2tny1Bca6Gc+W9OHGawT8aoaN+sHlnUooq/ZZ9sYyl6B
Lb3cuOYlcbcDKrbjdLgeq032qHAeKopwq7Quk/2sJkkoXfc/0vZ3yDom8jRW4I7mybAW/JUTHJ3J
+FstOLSSxTjvKxWHNHUsWuv2BMiTLc/n9EjSVxONNGDHrQOVU0HSdTffaMMe6vh2Y83io1T/iUP4
a8vU+w+0Fat/bjwtCk6FA4lWCFYbokxQI1BTITl8dtwXHTKLdiK31mgj9ime8l4y56TD+lyF9+js
VXJlBpjknu1Ej26yMo0GtOE1Cpnp3umQG3O/xrYmgvT3FwseBkeMajN/kHCVE6y4Yo25xnquQYiX
JK+UtDrgaP1qTosIYWtyFslmlYZ/g5p8zQl6+MqBe1lfCohpI76wJNIF+G16FJFVdigpVwgsPzkq
dcPQmoAY3Psl5JpRIhnlS2VtvdSw4O5VUR2EUtqvkNQuvWmr/AHU5r3lnS3UzVRa4Bzitxw4Yq8E
69yw1U8dFECBcXV4rTGRKglkFnXNff5Bzq8i3wiBReSYcvmzJkLCGKD5UQXEcml3BFqueAW2WwoL
jXSw8dipm6OrNOEdH7asrJCwBn74GzBsNVCgio3uTr0CaadtyeOMZYTiA8ypFw0lCoa02fLcXz1Y
kdp5jJMMuRJwuI+sirqAGnh+IdbE3JnBFynR4Kpt6rsyxxwdFmboUfunkSMKGYWPJxHMH6sWtu3j
61U2q6NTJ+PVp/UYQSwSa4y8UrZzzrppvayapFFy8+r8rqpLa5hNqt5hQAnWPbQ0/+bsKIqCXke4
uYqHhbW3rBa4NLbzaILMHN2pmllR/gPeORt3jA2qgVamZwvOQLRuudQu3AA8eJV0WzFf2m1f9RkX
gy8UvcdEZkfNFYT7vkCaPNcn5564M7vc98idYTyiQ0JO+dHnu/XMmZOnlLqOACcyD7x0bfiZv2vx
B4HTjMkuLvjVRlhxrzbEn4cQstxjzZzr8pjzd6LVHaYvq/5MMJ3e1y8F2aKxDuBemvVoztAVxP0p
4fe83wFgSvjdAVbKG9XPqIZye1dnVy2Xo3CD6bGuWEvj+MXPgoDzXDIygF6CR24uBmYj3H6IJxRP
NRVggczJSYRsOctWG0U8fO2C/oeqvin8AHG/3yZb6aI2xIOPkQs++uKsjQ5xUECgulY21gHGbSUv
fC047XdnsDcKeAwbndnJrHv3Ncyx+4Ur/X7MVYkfK/yQopS/SXmUwAgxSdlgvOFzteZ/Ta1QtANY
iqD9sz46rwNbtHX/n9MokWUdJ6om8+vUwOBtolgyCt+iSp/SzBmILmQ7nNT81m4iNsdtyTosMI3H
fsXbSnd12qHaxoCf0Y+1fpzXLjWp0G0sjacJHB/XU3y858J0DdGcF4NlW2fAgW4OduGprXHpRJHo
usMhFRoM3ahiXRbq5mRj0wLh6rsrH+RiXTwN4OxEQk4IzZmTK61S6jlXLsLpbenlgP0mMXLnuU3y
ocB6LcdzHxZOgYLL6rjuel48M0NJXgex+qMCCxdkpNrHd0fMW2bo1sss92e54yD07WD1lfO6O0NS
Sp8Z5YHGsI4YBc5AHPkBwaE6/o8Vzv5YmYk2OQDEfr8/OMn662rwnJy7eiHVWpRG0SnOINOuFCTb
1OX+a8SdFnOAbxGamdFF6B482VXTvNEbc2tvAl+sCMHs7GX1MvtKINjIvvuWWmwPyqBTIdvkZgdu
bkq2Ipo0GuykSFravnO1edirXDN1BWInj9PidLMx1V8iMODxHzkZxnplgrP/ebMImzLmIpBqp+g1
IdKlXdgtQZNFhW6E52guzWNkCknXJHgHkEjjxXHCKStGbXgONkGnc2wpEBd1xhtilIWJDurneU5Y
N7twrdrpqlPH4oM60GBqsDRxsUgdBI/C7jyK10uSUT7KguzzsACz9iIoBnai+RUmr/id7weWqHBP
XZhjEICiJ8+yQRWDqaEGyTnJgZQBbmyKlxezO//1ziegqpNoVwtemDk2VEtV3qYNljP1r2OfU1jb
QcK91Cd02OzWK3cxYLJ6Q4qzadF/7gfLj8Gu5OhiAS8TRqfBzICmQQhD66REus0ZnTfeG2NdtfKX
f4JarBy0DdP7TsJJDG1dkOFPNe2oMjc8LCpofGf2VYTkvDKARefj0y54wbjrOl/9EahS59T/1nO3
Z6FZN/i04s3sZi501YEEpgNraa0ch2uhbisAt9LU9UhAcYd9o/OEQ7KdC15qInHxParlfaFdWeMf
7gq9i3YsDQbezclaCiWhBcjynrcxrX+X+dfGP/u73ZENU6D5y/eOKh3udNg1tN4jnFGDLgmmOHh1
9glsnv1RHy0Jbikk14csMIKzOijSBQgjscceVTzXTA+YPpgQ3/1UE+brLCmLaccD2pTsl3Cgm71m
4iFcmlMYM8gx/oXmoF5/6+CPFsVKTKcSXlQjBCuXsLs9oIvRHWutYtnzlp0Zc1fQQxuoIqpPLkIr
65zkNFv/IHNHNrx3eRDlQpV/BA4YFDZeqbCJFncdGijGk4g8Sq+nn3FDT5AVnYAqxBx9R5f2CpjI
2GjJmFNsa1euRYShuM+3b8KjznJtOLneZ/GZE66xXb/cWLxVwE/0RjD4RHdJupwsV+GgyVvzBTbE
kuXIxtaXmUsLt8Hkw8eayDqDOqZmpFWB1PFpkMIILnWeVj+oePq9tP1IaqpEO8NrQLawjo7aNrps
gdHhSX/hLFdgjQpyZvF8nUy1GOp/rMg/+BZFD9EAXXm0e5VUQU6IsTM8uCz/VF/gsPgm+9aQS9AE
utnEduWWC17K9iHYHbfdlzOZvGnVhvx2i2cq6oXPTCe8qJEWlGMSe68FS4YEdnO59mR+ElWS+n5Q
sEHSO3XD/KFEZEjLzICxKSefcpXdE9kijc7MObhXYFpfhRk0D8BXK2pMrWH4XM5YoZuGLgowyw9u
6F1jfY+YANCJX6YvqYe5H35IED7eAP6tTTDB1bX50joUT371cAc7EHghUU8+cIBmOJeHmN/UJ6pO
NtJhubj7QzbAkF80aQocUFTsaQR6Sk7zFDSBBP4CB9ycbPzhl0e6XkC/u3dvFdYZ4GRQaFUMZsnE
HWYlz9EUzk5qkV6afi/HzzMaVSSv0ToksE7bYmfwsv6LHkOMcI/q5jytSy4E8FAKs1AorrdSm7+c
sxqUKjuRdYcLlMH2wqZ3Cwy3WoX87E/ensfuJH+Bae3tQcqBokx8KwScshCTW6+0f9CZPJp+DZ8Y
PYol1ej1MNl9lKvBVj85kUZ/P+jb3vJQX1glkFASioB7i5+cHmwSZ2EhBPCBKNuNnaJJ/Lgk+y/s
bezj2D0oVi6jRa3KS4PTGCDcvLZtU0uxcLIfl7cXJbl5FBMNP+Sz73t176ZdmrAU4P2QJ3RvkNBu
5/aO9S/LTlzD0A4piDTK9CUAs3QE0HF0On6FHtzVOQw7ruYTFg+MpD8Cpx6wgZOWxOMo9Xd5Y+84
OvYrBbOKxH/uEMaXtFEh5roYfGT2Fkw2H/mdCYAKI98qa+7T/887XdWCbdf8tKkWXk8xqgLy9q1C
WOPD7QmTSfa9ZYTRWXYjJDj6j1M+Q0Rl/0JlDz1CKidAneK+muhyw6kXCO1QT1L6oLqHmDNUBLvb
sAobRB7XVctZ2QQgq0b5SVB/sU/13jIVLtY/xN/vPcl9WxojLgkpKY4tBQ/K3v//6A28SX4GJ4a6
F4koAj+XEkOpLA0iILRddESW8eEr4sf5z/f/kwSbGlqBnWliefBl174Qsrwnd9fk/OI2I2jXoXkW
n0Q8ee5p89ZOPL6+M+DFxXBuTgNfd6B5jMP4PTcvksewxN8NDhpyKFGL6BVfrN9ZycPKPLVToaMy
i/cJkg3vE9Pd41HB7JYUPEBE1qJBhMFS5tJvfJPSJRiV4X4QR0jHjQX6sPufg/EyTnDxtsln13s+
fsNQmsxDSeupQOCtNu5DMy7+H2VIyiNY3ezLr7hfxJ9gOJFOj/IadnS4bwE9KXUimRbcjdhXBqLn
UlFMlB6j7X5RZQFXXRb7yJBthEtfB4uCx/+1fY91+ryrQSLBAOQIPNQwr6DfEo2eHx2rDafkQuTg
8/EKh1RHG+E5qYUacb/h62Z+2OtawePWb4opsW4oF75MXEUB7MLDpLv4DTxr1sVvS7JjwFc3H6Og
gntozIr9uFq32pWYWXaveSGndGLGXADMVRYKSbE87HHWSARAt3RrELztemQzSCiUV1K0AAO/3tl/
YNcBTHHxphlAPgCSxjEp+IfkeQtV+tAvtw0Rrhd2d076O9QQm2P4/OXE3N4/7Jv3wGDHXVDW4C8/
b7A7fCifTc8erOD+5VP39dET6oONlB4zIRgGu5h3XfeF7AaNWIt2PHdSWsnx61NEZrfOirL8VmWq
uRhWvSvvP5AwBBcW5tk+zh7pIoE7G/hH49PY6bzcDJfu3G39ZnkvXoTZZtRIIDEMXqBz4RLYBhbH
BSUySU7/lS8oShuaBKHPYl/Ua80CWHw80SnnbvrrBOPTkQoNnjXKWZaAYYc2QPnlO0JVXqNJJ/gJ
sbbJMITp3FHnapRN5Q01MAQ6TgEdpZT8ZE8MvEdAt1JphZl8JwpcwYnI9V5EHgH/Ik2Vjg0zO37s
5hpdsidTPpicZ3bHxdPIDChwt13aEQ5c9BCrcr29UtN0ZrUug1eCThEPS5Ra8EvHF5e07WFeZXeg
0Sk9Z/hasJQc+JZv794/hAoVn7Q5E7USJ20QxtGCgDu0N+2t0Qd4L98XWKoRBzt9js7/pM6Gf5Tm
c+Suws2f6SsyqSBdMH0nwMAlWDODsMouTowLhFTrItw16lKipxgFytOk+jbX1eR4yl7csbo2or4t
wAR/qYxhJYgCSyw2On5L6TCyTOejWJptwHuGPmadLb/GbJjyaHvZQoy2hEWAs8+a2tSeLyJ3InM6
ZGUazT6K+822hZvDWdBlahfYjpWtpKyE/QQiNzdnXbOw3zA/n8xYNl0FMERAF+oQT6l0I+ttICx1
NYzu6EhZkf/WCClx+ppU85KI0RMbGVYm3Kv83DrxRU4ChwQfKNTWlfhzfHeQ9a3Wy+YImlpM+58H
s1e74nZxjCUZEzUry08sW3Ujbz/cBETh8z7nGj2DjdsjrzHQWfmBSBTLfYXRSuDSRGQs6/XUlQwX
udgFcrMKLyF44dkgtPRr9vwVQCZDQzWwnEyXZhGZ+KfblKck+Xyh9GBFAxjol4cirW9es/YRCQUd
W9RdLv9sTLKa7Q1xwp7GrD8Sz5c/NBH0/haOl+TfWPBOIfk/UE0ix6r+WkRPFSfrLE4iA+4ngkop
c5WnnqpK2n3hzORq76iiUZsN4yptzkctSPdbaF+TouBx9lwYZPtCgAH4AamcYlImm0L7y4WscDzv
zkkVlLnahGuyXNO3wEa/KiYjErBmDNhWOXfVenOt9aA452ugKFwO5lCB6W7BG9zT3sx6MYEfI9NY
q2+y9zha8i/OELlrxn/GX6Xon+q3LSBjRf5rOxXzFrFF/2QdwX/EGiA/KY84Ahkd2Eg7D/0JRWgf
VQxnBv8/bAeMn6Fakldbx6E1pBkJKmCHR4s9JLvwTOji6i5I+QngASokBXB55GuDnGNfcbVH7FOz
Sx2g4O2XUIgyn4S+cGpflbzEcSsS0mVEc55wRd86uaFOL7VuPh0ghXM3n5/bc2ijj8iwWsfRGxbN
h+m6c3uT6H0huP9eeMfQ0NuGVTaZe+ceBoErWhkkSyFS3QAEYDqMFO4E/C2iIo5qK4lqTNJNfVto
eixQh8bfb7iK/r4wUnzKCXaLGIV+R4x7UUKla4G07BZS9AWRo4j2ItKhYWGM6svetzKy91J2Zali
kwE3euqs2cWy+h+ivVGP5onxOxjYTtNTfEam7co/ZxDCg4MNaGKYp2k5VfVm/BbMti07NXbmXOXV
A1mbgWHKA4j5LnnKRbXwy9pBkNPAq3mG+Kpqhd1BdAjvuxr8B8PE1rmAicvhtnMBjahhovLALVF+
CxaeH4q0VXoBq1HhMydIB0z8mE8gurdxzKe+taQledQehQ0QjxZTVetMZuyNmV3IZdC1WPARcIA0
62pCTVa0mikoKtKZyVG5TlrXJLYpjGVzsls6w6ZmUDunWHjl/DYnv34U4J/GC3F5IS4TIsvPK4A6
T8PCWA1kvx2jGxHvvM6pY3BE4BgYbobj8lhfUptJ217NaKMdbzmDv+0jckd1vbqvmhWM6d1d4fDH
v77NJf3HzBWygSFtZlMx96HMwMsr415fKI+xfaXL+bmr2z75+ELSa++cABiBly5PySsGz4N2J02l
mXwmLWiUvWZn4ZO2nzY4aEQx0OK6bZ2QFV2klX+oDHFn4Pn3N6UZsqL+lY0B8AtE/Z+Km3pVtIkd
TGfXjNs6R9/Fht3UZtlZhYy14NUVrc04EjJMSQRPxPRVCTw/Wyx0CBequGDv9KwVK2d62QMTB3Vz
HGpv5MqLKnRFBCbmhZctjYGRFfNVfN6sRYNbHYGxnO3YLEpx1zN9yFEROiGxpVKEa9G8aILbD3HA
y9Zc1RU6DJIbgQm+MdPZ+v6E88m6FsNZgh/a8SctWWqqQYjLtUMvykCasqFUKx8Bbnpyea6HLPc1
Y0ugYmAIypL1av1ELpQ3cah7e/C6jsX4vyGuDoqJKPArCbrqkFRhhlhbmZ2ARBFGCJ06mFhC2LVT
Xc9rNlaMBx4dSyFuyJZ3LX49uD7gPRRXgohoOEssXWyoszuoruKY30NnLe85klY8CXses6ZYOsgO
+5wf6tKEzPvzlBoyl88MXrwoJ27ymXDO0mPoSr4Py07cP6UfoVjyvMAF02nUPgwPCF7VyRqmjEAP
q0OErPk3nC0DZ6ui04qG5dlYdb7jRfJd2xIgdmL8dHqwGkFbugPQpBxvoIDYbZnXA+sEK5NwGd67
7NqtUcHLspNrhjnKDkeCLGrqgt4T6yr1dwMafOwGK7o9T/UPXPJ/0jjlBrdyNzN1H0QbSCaShQIy
FdSAr5Z3JrQJ6wqxpfkNu/46dCm+VUMJztflty58CtKXyWtqSMJErfLaXzC4l+etcNb0mhn1zcew
ysRz/a7ODeboGbD6lboxHv1uFncJHS0i8WRNp8YCZkJvS+JXJERxrRnjEAIr919/J8pML10GxTYt
GdMHuT2Q5vUkHSgHwFOVW+MoT4B/O+vSYSiKCgHU1Z4RnzVvA0MVN93C+tE4TRTQFIRKW33IMgq+
6YfFrfe2grde5zb8beUCsLbia7s4OsGY4QF/rkXezxR5/rg87suh9VfRCIr8itSCn9CHqRKmadgj
hYALYIKkmJ50LW2Ggd3Cb+UoKmA9pm3JdpKWGyJsbo3b0mtpxoUJ0Ym95P9Cxq0SpW1ofYbpR2N7
ub4ZR7JkfCyyCIKdtgg6BUD3EblCZKPFu6Js+OR2K4qNigNtPaHQQmChU7Sy576qKWzuMXq03A1c
HI/g8nWvrw2mrc1fhpWij2Nf7ZOv4hSpAOp/Ne5NjTRLG4ZsK6SETUviCtdIibcthFsvovL53tZK
/f0BeGodsCEAwj3jwD8+hoAEyCE81Kd0YMU2DBAx15KT6+Us3+J1O7fqTmbuAD//fEoQpf0ndqFf
h7REbq6XSJlgUeY6vjmcMcteiHyxvV9U/K6dGJDvMXeReGiUZoeZNvaoKHKgojel+627hz3KjdJ6
ehczdsXysQakB/eyLu4OVh3LhbWPesJdmHD9q62DvA21N7vqT1gX5BtAaRYYSE2S1jzlGh8gDseD
WgqXGQUu697wkqjiMqMj79fMabdzR3xha1SQKPz9ngfkRWvg2CfhgK71HaaQonbvSBhZyW+RbKjp
mumIquK/aW8/xvtBmUnndSy8wY6FaNcoricUAvD3PKB1nvxrCITsKRE/QH2kaRfVXv6oHk4FrboO
ofr3vDliUFkKTQueaBwQHZQZwsxF/0FF+yxia8GtwSpnN2kxMrjJm6pbJJNQKGpKvRiG0fBke56X
0w8iCl9dLBde87xRequGGZ/WUAWCa8zf2bsFBzY5FHIWwy46dlkpD47EqFHuG+eufX5VHnNL7jtw
OT5WnUkxG+WG+j78HC5Byb4KkDXz5OZgQR1cWcpcibw340/HSTUwGeV0+cpdlcPRYUtG4ZYWGU9N
gUnq99xSZSEPXpdVdCr7CYt9CThXV4W18mc/YjPJfn/kU827biit8x+QXXWLgU/oFZKjrgwV+gJ8
p9rBdqEqj28vYLJK565KJS1ACg0t7W0+umeHKTSrTFwClHUy/GcPmS1gS7MZfqYtqLt3vXkYl/Jx
hOEaq1U4OtT+1wYpKAGdgck+jSdCzmqXKt3VjWOXue8MSeO2Qv6HsMYVZUEyns0F4p21PthLYKq5
kfrTqOn9y1rc6BFImGte1QpF5ovs1Z7thnL6tvmX8j+wjxFl1OVvz/JANTNXLvTwzsNuyRFFvPVD
pKxB4DtD3cNoR46PjQmwJAdFcpUHjGvn8+Kn6TGTkFdn4tROM3Zl/xIsVPRxIlUDpwB3NjhtUqWT
oR+8jDlGqk13AjmcVrbY0YdOeceAE7fush1mSxg86kM34OMCIVBNcjATMeJ1rVQl14TG0YRZh8F3
ibCFtOeDJ4Ox7+tYJqL86aE1B6QWJYjBU6ZVMhePOEWkCnme9ZfYPgC7dVx/rq8VGqXqRJM4Y796
8M+XuRXGsx955kGGgmTKqjxlHO5qGRhGKgprhnT4jHLE52W+kyC9pZnfcsZYY7TBlOHYlTqc07xj
lPEpaEKeN8tPcSt2gXxWBdXmRR3RemHQmZnwUSl1dDCgCThqdM+Uixi4plx8THkMXsC2RsMTq6kb
wC/Hz102K9vc1WvWHZ+M7FBj785u3wrYOoTZs7oFtucyVTz5mQUXOzr9jKnoVdwzOuCduO/zp2mS
69lAiv1Ve63fH/o6ooRciZieRI+Kb82GCOxgMJhZijFsV8Y5RwZqTu71EJmP7PV74UkiHhInZtcm
XrytJQRcUhUT/t2VMX8g5WAUnWfB0nvsXI93Dw69Gec4SFlXKDCNmt1dDFzxkO+t5umw7O6xZbUZ
uC6ip1tH6xrEZdnR8ya6cdIP5Buoc8U7rxFKZR0kND8+cnZhSnuKhbpwbpsXXtNBsI+J8LkNPd1Q
A49ttgVRFfWsLYC+rKcqNBxR4CyK8tVgAc0Hd7O3YJSyt47dirrNGdX0I84CLAWgPWg+dkw658Uz
CA6qK3WdxBbmGw/miZfHpHO7nTh+oW3C3sldYPussnwqyZhK649SLqsDziIhmtkL6nweO3uoh3lF
s1Qy+Q8yp4kH7iWs1TV/PVH16ny6tgBL39Jw2s8HAIG/BtMwwMbPS/UPJqKrcI3TVBMpXlTvq++M
74FbcZ5432bxtTyom2mx34AiFpbkhWs/4F/nJCirztyBuaadB37iW8fPs605NSPqjR4lw9I+xmq2
GR8INky5IMSnu/HuR9xnt6OyGybDWWv1EXl7oQk4C5Km57XPdQsAIq0okpD39ZT5RlyBJNjzrE6y
mYap4VVjIBIxpVHv5GLQF8vl1lfXA9dALLawkIjdKO45RaMyXnVz82YemTpieIgEl1LyOmKFivs9
1dT6H2clnNHDN9cyUXzZbf3oIoColxOPdt7SQEvjeS0uqU2y/JdorBiFpgrEegOPkWrLHn1mmWpt
dvHSslMBfwzzvtFI35EAKC3v9Z/Y0SNKVmCRBANWd1pgeF5wtC7deUzwu2rcGkVVvRgd5MSygL7+
FN1DFD/a/ts3pAs+0CwjazdWN50oiF4P3yJT7GOw+VXPMSlpuX51lOQuISJzeLxjeR+2SdoEUNXp
dOQY26RG6QU1v+P6kb8KFIlg5N1YoNs51WtTgFlZW8HGxLP91AGuRlUKFgdFYQpyvQEuTSEeBE/E
aCXHTPwMDPLoTEfNT+HQxEF6t1zZYhgBrmImZ7uXvpcapKsW+JiENiKBpDZcUOYDyIP6RPZpuR7l
eT7Ub761n7rb8fDXXm1f+RXXuCVrq51c7cQetYZash6iyeyYAHFNjXJKrzFsewzlLHqvUvv7Qsjr
haUgDhARPgj174K5f/E8KkUM61lve8p03AEFG9iTZMWRiSof7dbckQyZwyt6URGrBBwu6q78WkkX
RKxg7f58yfJmzEzuNoxtSET0tGJBXCQJS1A6jHCGPFPQmrvQzAUC2oul4VGBY9fDhYS8eHVoRBmh
2SdJcYlb66NuZ4hzOjF8WINGa/QxRVfLk+oWLxmuF6fETCLunPoLmC/WiIyGKqE8HB29k01/0MDM
IXHDEbs5v/tmRSEw4dkggakrkNXkjOF9tz42lpHzuPHfwSGNt6OMukjVLLNhf/CzW53gwZCLhAqd
5NiZ4qMvQopVjyE/dMEtKisToaYSKFodSqr0lqLOuPghY27H8Gtc46oE7ISxqJU9sdTJEn3WVRyW
sXTA7eneAiovxlHq1TjSeBHkk1V+8b+CNn+y31c57zWO+8m4mDTrMCZod6sF7BEfB38vKF0eu31w
qr5QqjTuPeyALuLKBBh5ktfJpN6qCBFs3WU6aNzCLcR4igJdi94SAHwkfxlvOToRQsBnMogtLBB9
Lk1t7Lg391uedHqTFEb2+G9X+EbesfP8qqC9ZztUe1Y1zenb+Wm+jS7g+p8L4oo2mGipmJY8Bs+4
qS/nEwL2ZU3kV1D6qNsZZ3TkMttZrPH3EF9uNQxhbrBFmXCEjRwNPfX40LkWN6CE/uHQeJpZG8hl
9c1ZcGwvepQZ5MfU/h47T7L271JTYqt5uLSV+y6IGWVGES5TobLAMrZInC+z3NBbkcQGb0DjAFeF
cbt4aK02KOfZ39AZf0yIrsAquXh1NkpAo/vpa7qYnAEZxWlMKkZvSKuetSDCGMXfOcO517pXiYFN
A8LC8RXsEW9XH8uBLw3ZVnkxZFP26lq6Sq4l6LCDaikUsZd5fS9Ww2MFI72pyzyFvwvOIJQsYMmy
Og573oR+AlfEl7FGggt0nKJXybmJ9AaUwerJVE/KMe9M8BHfd5X02FcL0hOu/SGEn7xuOzTrs00D
iTt2wouLQr0daVX7PRZs16txTDYGdVOuucJ2jtzKLDTDXPg3Ch7wo3pgbQ5qHNSTsG6Rd4/Svs/Y
6C8fpuUjUryi5s8796E1/YVBMNJttB/nYhHthHiKNLbf0KB4fO52d8KwfnDH1RJUYPvyq9z2RI4I
himDfpnOPPIbINqPE3UAFZhvp4TNWGuHTT1mBKFCA358VyZqLJyD4H5EUMu161eiE4lL0gLPomln
1oxvE3qxzvBDy2A4fhbd2bNa0K7V/NjA7H3K0y4mm20FoWy0v2MdUJpm+y3LpoY4mrywThlGJRrI
Ow2fpb6MkCxgqyASbUsLjvualemLX6oYI7X1Wfc6Lrtmi0GnMIUzEwkzq2D2RXTJU/Fhz/Az3UAq
lBDG9l5MxvJ820a5MhGP7SLytOSbacCbfLWOU9M0cCVd0ITENn7Ch5zvcyoY451VAEl9vMdhSDdz
uxSLXCoT1lBXfySZIAhr4JftI06JyG0x1bb+IHQRP9YIW+h+a3MlEKnhdWH/lt+mf/YbvrPvHY7D
sM6GM6+XM/rxHLu0t37wCXz/4l+Vxa2EfWhGpqtSlMCU5xMA3uyVUURrJalRRQUpF1gSFBKUri5T
xgwENkga6KkJBWzfiGx2JrHQ1vic6iLF5fiI9BBn5DNqf9S/tm22I0uw5kliT3ij59JWrc9k/ORy
6V81bdt5Dtg8t8j3z2pQDWYhiQcn5w+i/sHdYpC8NPMYME0nx8wiUo+YfvoJ2WOYH2jSamZ6Eojc
45mjiFY3IwC2RTJMN8gZ0hNqnSJiof9TEp/umTu9rjHJmDpz80kJcePCki5b51c8pCoFTo3h9dFM
x+RcQ1nQH591U5zL5VWKGg7kuKfO7r4IrJG2j2p+afQM4/uIDBkbq6dK0U53u1G/Y8yJ65HZTy6F
v1WHNEBtwHgy2H/GHt1ad6fFqOcr9SqPrjzFh8yddDWieTjSotC34l0/vg5XbJWUvg9XLapsnJ5b
acSpDlWG7IXBGexwWbyvKChP/H+O9Oik9dqPwXj3IbGlkcgpX+qv70KsiJLHQuuAS/Qf6Qo3LAok
s0vEQ6MIX9YKgPqayobxvRbhVmsttgVhTtbFejHfWS9/HZ0DT/rhBwF54u2v88nch0K6cH9+7v+d
yR7iTmemDXrZkdO7GwRnNIPjHSNDHx4Z4U+gDk77v0GtCQtDUXFSMc+FvrC0kjxdILvbjIB70tgw
WvZypE2MNU6TYWB30A81CfPny/X4GLVImeC8mZ839iWpRn+QtjSDxTrF9xBW/Zn5TNTUp90aCEXr
J7/wplC1+Sa7HRNVWjxUjxJZjgUI8njSg1/rN3czBJYjEORVOQysoTEVjf85hDvIj3lVWY/MTB4S
2BTvtp7uYqVhrv3uiGxlziY6lzJc2QEr1/bU/1u/PfmmX2XNuudDqOVryf3qAnE8M5IkatP4KTbb
l4/y45eXHqgCHvWDA2yn7XYR4zUpe5eg1yqJTSt3zrzMztYQT+VeA3ANCj8q/pYoexCg2l2s8Kzn
nUVBtPg0f1jJ1YZjMF0hxNVdzloKRrTQNtJPljjXlpVaqlZMC6LXH/zvGSc63PEbE0VYuU52/sYD
k3JR7Ynbd3N7qRUArOR78rgJXFOiaoPsWGiN2VlgLTDiyosw9iehVCDGfaqqaJNUSZ39k4kf8HjJ
43PZrLoJ+YqZMaz9sS+801eHEosr9/kuzC02/dIpeHmWDm0q/CtKag2iw5vwXgJHT2/V0PiBomYx
vNxGgU9HNgQQscmsU8VjiJIfZt1VRCUlHA2DulwECxRU3xbmCtWnVtSmWvVeopSMIBnyM0QiwLL2
ndgLRs6CDBZLJtflLT5476HI5tFTi3hPkZXN+E/FR+Bz9v3NDi/ecRc8BhdZmgaaPe/y/Dp5TDA6
wjK4Fz8xYxDAE7Py3B8Bt1K5GiF3C/YkJKdtt3ffEP1k/QQYtMMFy+oMvRG8xIOP4WGMU9S5Wm84
Sjr18/Iy4pNt2I0Jd40mjCosWDm88/nm8bUdbTExXxqs1dwyobkEQ6J9BLwgwNd8P0Go8xgjMAcz
oZhuYY5a2HBJUosEownBj3stju3x1N5+xAsDKtgbfocVpTNDYWOViiyc/hMFBGKbdoq85XrmA8pd
uts9+Cm/AR5rktdA+vfNOa7rDnZI6/ke9++nbQ0A2M8fz2v5uQtpgQdIshS+cIV4Nu5/KUtQIADP
cEUfgObu5CmC7ICD3HR0OGs5NyF5z1B6RAXzZX+o4gAEHL4asUo8Ngwg5I+ErzGQf9HxbkFD4R0A
fHOj64mKuo+GiI88aFCCTOHGuKeRLhyb24ycXQa428S7hX7jLTpUw80Fj+BCfzVAWVV67tmFJKPj
TsuCIUYHRPR9gw6zemA9fsM4CmLMW4YmtnkrIBCrlBtP9XZFR7/ntxlP3opX0e7vqMoXgtSb9TJ5
179kJGFU4APxgFyeQAHbBDu5L5OugRl3UduwrRp0JuQfPYjxsd9haksxfaDrCbGCctBmupSfqFhn
yzrxu70WSrhIpQGQB08VUykv0sQnOyaUzMxcnkTRSIwOtzvMK5wTED8bXV3eM1W8AXeG0QHsX+ar
YjhwN+Cyn8tgOaIry/mvSWrhQP1ISr8HqFcF5RWTI8Bf1KLrBAYzTt/Q/gkz9apzl1+7LFdFOpX7
prDKIugBp5uCRAjfikMS6T7/ztq9xNYmcaqrL8EFkiUrggFI34jXzlAEnC0iHq1cQsAbtCwUIhWe
Dk7bpuiQND0wztrRq9r3Es1QBvehKvVByDcLOtWiPPcymSu45Ua6fdsojaufQPI+tQEeyNg2Hs3Y
KXuNaO+D3P8tXImiEG97VAcj6xfkvqrpRDhweDrUoWUdkGZ3FGbBwB+Jk9m1//C72ohJimhE263T
Txq86fqa1l1Wf7N4ODjLQhq3Ia1nXEK2sSkyaa6bIMPn/Q4QmfY5lMXCgZ2sw1ZUtOsddx4BGoPx
BMWeMPZhNNcFmNjb3oMjlfbT1dxk/RPve9GDyAjxPd3SFkKMzh2aOc8YCvLuAqs8/eQWAnHPBSWy
6gp1SSaeuu5Ak8/SGDTXYDAfNi2kvS3yskG9zIjyOVYQbRw3BjbRHUTN1+RMXM+sLHosxj92hrIv
X3cqO0N5DBWdZhn/PBNFpFM1bZS6A7GRBXGzNK/A09L1dFv7C3tFZGHZoczUPqQfro+5BwcMuexx
036kbwrmGUlCDSLu8ywtMUaeufw/5DFdMceVNxBQ96myPDvI1or730S4vvkYjvp55OmTxlRDn6GK
/RMawOk1zul8zBm3phSitL5FGmnS2eqm1ARhgB425zZS74gQAvhxoMGXp9WLa2aMa1dsM/Nen65J
A1RQaRFCl5jO96DEGLpz5TgaXeeUfwYuQKYJOO3APiLgrLk6YOAmo7VimMb8BwdmtEG4Ustv0rSt
dcyumV0rzUgtNZwWr+YEzUgJ2ItpDUyunmMlwNYLgmIOBHXfREmW0KosamJR/hbc3w6C0iV52QfH
Aw1uzFa0lF2nagYjdGoYk5phc5MCXdGpwecqDMkI9HoD4sFMUiO8F/ZpIYNOuldEQK0nzGuNysvC
wdWc7LwKvFgU4T9SyakFmzyANxqO0C3EPvOFM/lLItLNsVPA43PqL3B3JmcjxXYb9ASau2vK7P2z
eTIt8VpvBnW2TrJJ5oxupQ6EDag2lkQBCMEYT9JD9Y7FtIaTabB93Ju1iIYLlETtBjDsToNkPM8B
4kg12wszdbur18WK9D5EsXgpzovAB6cR+yJfD9EGjoKKFVxjAIj6YhHBEEcdD5tpbQrjVL5WHpwW
KykoZl8uj5cC7c63bbe4mx9AjSbbcI12ZMZw19tba5iWa10VlTLA+M+cGLJI2zSKHPhu0UPKTV+6
5UdmIuaIedmL3Z+Jou2IEmH5GNL9/S7I/b7kPks2vU8ctr8XF78JCQQuuVAfqGdUlfHgalkVC9dG
Qq2W7u8ovzjQy3qqF8bIXChNbfAYQXUG7xBa74K4TSDLjuhtLkRj7VuYtXLEb8kJADopzasiogPu
TQYcMtIfCYb1f7H1EJP5YVyskzDQp1cU3Ii1aJLnHkTmqdnJs/n6awUnc3EXNEsm1TeYA9mEyXuW
7fOq9AbR7kQPSbb7m7hwg3a2gV3Ye5VJ11J5tAv/mtSDQG9Z0MMFqQNhWlqdc/hpKOtvLLtIULUH
Zbr1VVXmCkD9Kc6uTalSU+fycnrIpmlZTDtOULhrmKoEoOqgYaumL3X87FqNr9QsTCr71WX6i+sV
EBS5uWy9/Ia/RIw4+m3p7BtuuX5EInIRS7rcvglJTL2k6/oEoTRI2z9SNAqoYQLQk+gUaIL/RTjy
ehaiqQj7JPpXitOP+R/hpp1c5QQ1RLJZMXUJYSL7jkWUsPMug99INUoxNuCxbndERrFeHepq4ctk
cNQ2/UWHWGuYstc1wyMh2DGcxdbcyPyE0+P0P+7g1xUCgnX2TCD4EJyjvcxBFFNa+MHKc5CNiBRy
E7RPNyBLBUC3QSxJKymK8lKn5/aFFKBY2KLMuTWn3SNEWPNhAXeDC4Flq0hAaaeXZ6mA+uTDVmxV
B0rz6z70B4QcjJybz3mQyw1nFujFn6ZLvSqCBw4mK5+2xWbGRcRId5DKfWXgZf9X2NE4B5NXrbJY
1+iD6i07J+YTEuekqb42xPgdJ133S+2/NE+xTMoeboQUAAzrQKF5Pkz698tx1wRFhR0z8scVk2mH
INY0A4jpQrw/CWLsidFtYtZaM4vj5cnukWhsYsnkJcQO9U/dA8DGrY1eIDcR3AeWo1yc+vyObgNX
5WHlXyLRUImKl2Pugpmbb7hsFknW/v1CqvtNcgFIftt0ZVxzsDuSyYVvh2lVK8ffSWZ5bnky6ZRB
hHcVOl+gE4R7qkz9lpinL0jh5so2tzlUE671wxlNY+w5Lzs2D7ARqbu6ehLbdmX6lGWERSWES7m5
DZsFBnquQZ0LXh+ZRK0KJI6DufZlElBuMfaLM160XsnRrqb+w69B3qvpNkAmz1mIFdcYst/jBQ6c
u1mlXg7pntW2pm/Eptq5fQU8ko7usLADJjl8MEidxiHbM5eifxP72/u7uM9ucBE4sHmLjNl9C+Sh
Xf2f5M4nK/8IAty6nZvV7fxQuAafRKF0uPbfX5uvc/T0fJokinqxT5gBKk5Wqg+FoF3jFw1kvEdz
SzeFH60kGNX+A2335+Y2HSLii1kEfQaIGZOdWBUYy8X8akLSMRhCWlm/B246jWEw+KDBMLus615L
U74GNDfh9MRvYsUDutblu0EidntJ3Rx5PW2YJVAqqxXMJNnbiaY1a2Q0vYnwKGRB3a5QliudwxVh
gP2CkGzD+YC6gGAbzpCskY4RixNOAOOsQNW9pggTvbTD//6Nn+odsWOZ1I89seh6KzFsXDEQZHmV
DNhnFadOaBdXe6EW5FAPIijC3HC0KSSLISY34LuAAgPIWfzb4n2GcE67g/zfHjta3sRyoLJBNSI9
slK8catsSBzX0mT5l76yhJSq+F0sD9u5FyMluNKAejvShys/j1QViaIq7bmPlt4gcJMuf1DhmIEe
B2pq8iuXF9mcngUTUgPWyPwlbYTI/cJCaHFE8mxaXuMNeFdCEnkLGRdghaRN2HBGLqImziyvEzC2
DSVIolulAH04cAfCeHjmStJt5Jhb/Sqlqghr9SjZnCmml71k1f37puvKAO7lY3gADdCQ/4vCtDMQ
46JTsblVnCTX6f9PdTJ2cNokOQLf2o21Ip0yYRytDy0c2wQe1KBe5lCXn6tf2XlomGQUNxdscbpi
ak8p0aaJIorMhdPeZksKUVybmP+GogKFFpkAIl0/Y+8MbJw3cKJ0nvXYheHTMYP9oo60i1j4S+Vl
kVfJZFpSrtY0epw/5sIrJ3C1i5UFVOWt+Vpi+Kx1YzlaO3eCKsPTVe6b5JPjj7dp9sWYCLfLRl+s
LWLFrtNox9O5FcByNNbBzx61nSD2aiH4tb1wlAJNKTUr/bEVTfIBtgKHKuw/pV/UB10hipqZGQ0w
3wZOCOMdHuoA9Tyhzuu9zMPW49faoW9D2lvv6mB9tDrTjZGqA/T+rYtw0uJehhqhr1qXleJ8KzmK
5t3q0ebwxd6WO9fCkFbrOT9q3G45vjLq5Y5Be3Lv3wq/L2+hSoCyU+CNeIiKuvO4X6uzN7YkVOvs
mGQgGL69Vt1/F2I30KfFk50FUZ8SYscA2JD5N5+lmYwAUIgtP/rlYlb3yWB88mpWZDulqUJpd7NR
GZT8MK985HXFn+gNlJjZUDYnoSGbstPnRXTVfqsUnNY3PAtELIX2BYHMsDlowgm4lML43sDumVcq
t8adIG9sLN2R7QaFoBULHv7oNO+DDBjsUREZ9dvtvapKQxCr9BM4PTaVQPucF4WDA8hXufEcmPz+
hL4874GcDADk5eeA/zOgh3PSuVtNrZxaRMYWSBCLusiL7kPK7BPIYY+9Zy6zaH2oFusuTksb19wy
xD+yb+tzsVGm2mNmuy6HPIUD/UEOQVVeUn8GHO2/8b6VM6qLtnGxb7XFiY9G5EKcwfkVEaLXBBUd
xA8KXjCN1DDUqT/v+OpWsH4wAO33+1YAijEe7Z/cA54TIYq45N9GJg0pCg/Q9EOUaiqUZNNVuOv2
7W5QtHKy+GuPLBN0xtBYTto2gq9G33gu6BHbPIayadBpgjVTXfpzvSlWsVkE9rDU99jmkJSGvR26
E1JIBwk62QZz655ItIBSdBbIXfVOjVfODgK5vViFYG72nJCbS28j9AyamPsIYRowpmsD1CF1y4Iw
2NxjQ23ZB0yNcZkQOum2xKS3mx0HAWIcZn7wSSUjOqMdHCrS9gxwUzvgZeAar5bH7310ZzUYwhT6
kDcDxBOezQo2IwfUkQ9x5fVhfWSkBZTLjieBtZcQ+jISx6C94erPmarh+6kFfl+s9DNKq/a4cV9Y
NRQZVQuHjJa0a9bIwu0W1bHhD500RtjYFL+MD/lISare4P5zgaJaN+CwqAcuKj30+1YU58Xju80G
xdP8brx/e5KbknTHlZ6cBwvU/1cyVZIiXTij/foUQyQM8n1KEReBrGHxDqeWT7odszij4bkdqXxL
chc318B52q394vghbromqLs0XB2GOgUooLoJwK+rlfPDm0Ulj19daL4jICmiotT7r/0qIVK0ww3Q
YqShbtduLE3U4ADWErDGpGwtReDmRVUUruTvLL2/DKPxBmFNKHvmWxJlteikIfBzFnU8r9+c9NXh
siWw7jvGURObKcfueIYCHoye9ldXzbUWxRkva7E3uU/8IVMZyM1T6Ug4u8hS4eiFsmWirTXqNbsa
qF5fz7g+wWw+kBYtLicXCq+vVk4kFFSSPOme5kcK32aDqysl56+BinNsbnIOsza52rJeFQ38TkMK
KAh43Z/HsMa0hO+Eio0gxI2R5I78eVb+J0I0nQNXYx5Zv3iYSP7Beu5EedTbhwXjy2yaZ1FuNU+i
PE7libULWUUgbDFZCQpug1I1vB2WBWcadTZAkeVBPi33AelspOzOoBYpxdleCQyPpzPkkxiisuAr
6jyghWfaeDulcVqOArWPmcRZiqMNYmN3436eF99yfxosCmr/VP+sjUlN1duYa5OCmBXo19uEYNNE
8ufWtnBjJ1HwSIsfrUwJbW2bvAdW/cujQilZfJvKx0nRjVnmHcA6vtoEj/25h6L3ESV/dGA3/s6U
Grz8qBkpqi5AzQoSDqBI8j3isGUw1QuFPVKfOqpZZ9f8dJ/iJNcQODRP8mYQvwJTdIqcZ9MJGJfC
nqyROn13kwsbE1rO6Nm/iwNp6f6cQEXIfjIWJaF48GKOT+3I2ekxzdv2hlAcLNZyYEiPMuzuEUgj
9W6NN9tSS/IeDg3yIeqQe9Mf97/VmoFXySAX93b3oKi1sPV8OgCAbwmlqf9ucotd+PYgSbiWKfTK
Zpoc4Ub0bcYARexptxjJbbasGbBT6Am9IumpQKZaNm3tLPt8LSoc6upeYU8czHC/9s1HWWNw1rmf
K5GjDHhRhetL5sUZW68E/X5GldfL99LZum731RROLk2exAlg+gVzxsS3eqFwtZwWqgRp8o22X3NW
Ofl4lLuZ6WVIAvSMbq6A3VL+sqvs5KhftP2RTUsPGEX6vH9OmPRhfzKhfOyd8ufth2W8E0NVmie/
SAw0nhPW7tgiWacFrRDvSu91+emY465ig2lzOC8cBpRAtLHF6LDVsq/ppoqVbha4wz0zxJkXFRfc
oot+BTzhxrKhJZQ2a3UYwdngheHXzEwheQGwsOnpX2oaKv41fJIlRyOcQhASzEEFTFIsbYi3fV9X
mJ3/5YxQVvZGeGaF9zdQoWjRGh2S6awv6p+E6p87VY8puvGcfMKoPm1q/38UgvZQ34GdFtbZiSEy
3oQ5MB8BnZweCAwyiU87pEUvt75qYi3rz2M1EIwAx0hgHQ1oMqMLWG2p/zwWWux7lLo/07F8SPM2
52A101By/2eb0r4IFBvBNeeaDcYjjlPcWVs+GT5gUG8pwybEAakogCC3j5oapnvrdgmVUOj2Qns0
yZORWqgr0nvCOxAl0b9pLULJeY42a6gpuYliXpUiaR/Arb/POtANsrvVY1XrLLOUHfS7S39d6W5Z
FtTvQqO6IxnzsznW90DzqF9TuZzyNQ2nlE+RwksIgCJ8uBCRbugfUsIffzrh+kCD44V5nx6NAvsP
6DBr6NKAi/E/YuCVntuJL2VjhQy2NRyIIdrUEUYXoMAhTo08XGhn6l1DbReX3h0bDGUp/H2YMpP/
fIPgftVynYrVBKLKTMF2E0P8qavNk0ABJ2redUMSPSxmjcQi7wwwZr2H3rZY4+vFNTxaDR2E4CB5
71OcOvRyShqzZ5a7tvn2zSna5tm/fvM18dA0GWN4OM5/1vC43sZ/m+RyRxpvWB6x/bLcutELtXV6
fz+4JcqKGfuLLDsEsaCaLcQe0MQ4UlFiyUeBDjkyBa/jt1c/CpB6aIGgVMiLWjxUSGuVNxrwY4Ff
5zpIdVTojmS4yi9G5oIPHwzIZJYTGQk4WU4r0+g15BmZ8+o7r7SKQixY1KrPJqz7pA5X8h682IWO
Ys31sWgqegiu/Fukwe6Ut3mPRXwAEqWv/B6epE48fshq22IxfsonaQeX66GWcrUo0CUyWplZPFxb
C4nj/NWKgui0evZSbIYmgUijqoorUELLswz6JVnONT1WXariOU8yV2YdyJRvg7ypGTaalz2zEXmH
2+kSGuJ2ZN+a9qRF7UNylEplVzR1fwD+FCza+q/DfVNUl52y7NpnbOG6Tzko08DReBXFQ8bWm9/s
8RAOcjkH8kkpb7lEfC80DtcPHxBI0HwsDla83vSRBiUsGrJ/GGIUhvsURMjtT+Pe5jzZmvhV83zw
no+Fj9heT8mNKU5f0JrJw6yh6s0YqRdolbSYXKXH7JaM7A6xSugOcYsZpSzbFMD6J6VHFdVlBm6V
oQCADNnxZxn3OYhI0t4totgVnSEX53w3hoRJ0tYZ4FUPxRGDxB9DKe2w4dW0Mz+yGqQn1LuRiH4k
yzbQta5hq+bECf0KEWskm8JCgqqxznvTtH9VP5Bms22uEsAFFdQXpuzM+qIiy0ghT7l9eCJWt3Dy
2mKkyzcaf9f3hTvGewqWLhKgKf8cCBCHnUkBjGapELeM3jexgcFTyFoeG4tnovI6GKVq57mw0e3Z
TNwexlnTu3BSO9lft4F+4D/SU209m6ZXJHoZOVyO6Hqr8FDEMzxj7ihJJe197b68T7X+nQhsYST0
rua7qvPNXYrgQvJvA21yGR1zhFfk08cMJjGOTz8niFlMIWhEIAH0PPbYFeM4XmQcRsSnYQJ4X0Fr
H4JQJrAES5q+aZHNOcQZo769/k/2R5v5n9snQHtqk4TcfsLJZooc2NFXFZp1h/hL+xjQ1hPDdz9P
o8bHj8ixYWoPes15wkcqYuhA1srlJBkNPnfSOu2uIRTccOO7sLUhXCZGyaoeiecsfNiLdW+I2PvB
jGn89hgNxyHxNaVvjBwkz9nhjT4Eiw3dLIv6uxkC4U4V7BY9KRZLeg0Z3khz83fpbZY6z9Liut8S
6oG3XEQsw+P68Nqdqqhd3O/laxMFdqNcLp/rGHui8UJhv7DCJEmhWXgKyiK/+CHybh7aHA2Xe0Nm
S608dz178a/SUY9kmW0Caep2T0vUJ6D7a7KnzwAyNLn5JnbJNB/VZ4WESB0Oh/PAgm8CagR/9nqn
XjQGiqWY+NkBICX7Y+jyTeqgHf/97uItr2J181eT3ksxHor22z3QJFIaXYfPUym/EwtGkP2CCCh9
dHZxccb6dWkKYwteLjM+AjOQB7i4051DZNdaC7CcnCbIgIoOLqzJS5MuRcENULFDZ9TwvjGDIuPY
n77W4q/dWD5Ie2m/0aozDg4sLHz2YlqhbsK+Q/OTtSplF8yM5ERW3skK2LeE04HPHqWJkHnq13C8
9pNLTyNGHZ9XhpZLrnI5KKqOJE+h0dKFGUC+rKBR2p+zCKwgRDnPBGgEsRrwA8GoCY7ktFVL0Ile
+VY+Bq/esfN+eemOAZGnLWDrH7DpTc/7ICzKX2QkRWKLJZqsZmDHJ/iTxKln5GT12K+3/v6Hhgy9
q9BdhNzgzY4rh2RZ/SDLAppYI9zwE3iOs9ZAmDws//LLLGaISZBYDVFNpBmYgmPH6mvcdh2je0WB
twOQCyHQPA5RnaVcJVbpjaHZgFKJCXC5bL1AfCv87oE58OCracjeNB7HNOxCBOksEYzNYSwRVN6B
3bj5d//jmbnHrRlzEKNSiTQPbN6NM2OnpA0tFWjFKl6j6xBnQn9l8IxauEWXxu5OxbB8P5w8ZkSJ
uXnNouIgwF+xVXF3QEq1sWgorOR1E80ibhUj/bYOj2OMOhhjnOGUpCPNPsL5g36a6NOBjwoUYnfu
IH4EiCJmG0NO8WTh0uCH4EgaR2EGDxZP5S/4uxjznLJge+NlzK+PcyPcb3GYS1sgZFlo9j6hP53t
sCAAMo3CVFbaUcTiOuwvOufPKY6AFo17oLvoTrgfV1daT2Y6CvXG1WC0rnx4CjFj0lzzv9mrsGb0
Mb8LW2yVddC00e22/LJazEnXNcCQ0npn53+vxscIJMwxmQ90cMl88Zgc0/jpZFkU8gzo1kacBRGs
YSnthF5AmO9tUcYt7TT0BB4fCMW6saL4vMO2AHKvbNEsAc8arYYJG34/vfEKPQAET4ZP04Q5pPz7
v1Z6+mEhT6GhtV56pIcVb9Im4p1VPkS3Qb92kYWebjqE3yVp7L+xqWpGlpiyDnKgxfvVHQu/99VI
8qtjLnbQnZB23YbvruQ4/ZTnGU8GWKzowKZkP/Airrg67sl2stWVEkZndQWbogdhlGmKgYyBFF5f
7urrjkmLEyoo0CuR3hbnwVVqTUu/eGYKxJmEJjLmOzeCVGegx19qg21yunwOh1cz3MVnfl7sLCIl
6SLtExvkrxxZRuQJg1W5Z07TG+ZaxU3TEKoUpQGuXO4pADKaAO8Q6pOJL3Ud/LF8K3oOt4pTZ8T+
61QQ/4d/ZLz+xuAvubN2lucuBBJs5DjjFamt0kGyfnzghBoLoDoYjh0xyANkQ8wFR55Pvbv0HrBo
SkWCOihrqrZK6C8pTgvLV/8e80BoN/Q5Fqu+zdRWb31vo5QEi3FUwWbZYPE2xrjaxzdXOH0RCMb9
eRVByI90U+UqdsvLLzOvNz0V3kAoNRrwCragH4AuY+Y7AoqnRaU+BJt93Y6hS+DVC4SIQn+NJGwE
MDNKT1fp/4kKVDtVapzxJfhoqeNTNC8okCxHQE6xFbF8cZkSVfLBSAGtQ9yXW+xgP6jlhnL4eml+
pGu5rd2y/t5HIcylrpOWS4LVX/tw4QFAkDysvFJMH1gpY6btYf3CeSrH5bNhw+M3DDCMJma62Fa3
GeKwrn5uJ1lzeDKjaf/3xMjaWF6c81KGuWoenOkz8SPpPpriUOBVrOFUhIj2rX5IuYf7Aq/V65wl
XuvxxgHCRiKRaNZ79ShwzJDWshRJ5pwgmTmELgR6/RvuJzBhtdVHcGauE03R7AjPVLRDwoudiKI0
7DmSHCgIY1Ljy/K+OJG82i6s2qOfR9VCsBSeFYSxCM/FezA+5hsuNAJ4ZhH/M/WZs/d8Bkr1cbX9
OIg4sRYZDL2RESlkmJf3sFGpDy3IRnn6xZvu6IOJM8sNTpok/yHuxktPbhR4TKPhWjXfIMBcPq8B
Q0NxYAQGFNVA70ktqUScGkDXEQRjV6noTMtusczxJw1acCb0XEWAKznyySSQu4/lrqrl4KcSSVD7
bCKVJWA1SlmYstWivs3nRtrGIUqpmh22V8A4TkNgCDCAbHOTGJx4FD42dmu/iM54oK0exhDUlHJs
hMvL/tsD31kKrozNRADl5XFICGnnJOYuYxvbbYSpEVHBu2p9EG/PPO2haKGt4uzU/Qgd3kOKXfJQ
VWL7EUthGIqMa50G6IpxlKwwjUMGXm1UfhnZjkVq9H5mjhLZko6aNq8iYTk1lOfBlQqafIAzNH0v
92FWjk2YMAqw/eOB1H9RzNf4B7ND5Jv0hGowLdLfi3XnuJ38blCrv/ogKO/owFDKY48RRFZIUdw7
W+GmDgrADTuvHFCB3F10rU2nF6sKuYtzGhkETba9mzATM2VjLuBLwpveebfNQvs5e6wp2+13hIn8
DtAuqdCwiY2Sq5YOD3tSFIVJLGycWu0maIHGc+HFBvfJQ36iTBCDXHwywwXYApyPYmUtISKnEXtN
VySrrdm5Z//15UisPjjEF7iNhRZkafPxfSrMw5k1EnLEORODtTzRYYcC8vzEnHHN74DAbq97Md9L
q4ELbPSvH4+Uk8xg4gbLC0GjQRaXqM9AxDm5ZFZc5KnTGrFpRm+J7v9SgLQvVDYTsGhOcKqDdWcG
bOJ/cXsvoNq7tl/KEyc+fG3uimqVLArPfuXU0oTRbqZtYDnxLWJJaYZKPwpc6YhHSMAvIGwBx4nv
juHgOI/961a13RPC4QGSZSK29tTB0zs3M1v3zPIQhP1HNylInkTe4CFGkoOYZbicEQ5hdJl8oDy8
BJZ1SfZSbS7/Zy9VzCkuiQ5quSTVqA5OG3mjQpd9h1hR+We+r2EOV50y0J5mmCC5TRjxxK4W1//w
1bKyjtPDC7LS42Kxvkv4pbO0bYhE7YY/yBqRkn+V/HBQjVPlu6kGNWFUM+zheYZkrEkCcKhUbegE
+8t8Q/IfgyakJDFH5m39FPURScwCd579u3AjsuRk2fBz7ykW5wsUaBxH3dqVl20wRC4Aq/Q4bTXF
N/+UseCngbzXgtq8Tn2e+WnxLm8JfQF5zOqS4hJvCcBtM+C++wG1y52HbkOcn1c7OmV5B4fbfig/
9WLFvQYw6NjXgNPmWnKX+QcnvhPfr+NiEZOkoB+pDFkAMIiZP55Z1JbE5bdRWM1sEW5l1oVB1uwQ
T0DeQ7cGVL4COplqddXRfi/nJpSTX2zyP8Va9YXgm8wRMuuqoegZUajPnXoD2quznTthehhFgIAY
sxyx8k29WBEdfIhSJtnwQi9kYAVg5Oe4X7EDaEc4YuxLSMgp/YANtPYaDG1Z5ACGicxNc6dJcSCe
nyHac4XUtMxnx/Z0n4kM9AcnUPv2ocNNyl1BO//ClKmxJSaPSvXsOpcm4sI7THwP7xO4+L4LHcJu
1bHcoPUxwjDWEHo/qbMxGIIYTyuPSY2CcHlHt8/K5WWzfCVSkSUPdB+psiB3ZclD6oENlPr2gXph
at9fMvRk0sZWiX3tgv61uI164E2jnJbl8bQKFzyI1TdEBdiGGJt1sJ4D5YOb0nAIU4xsITFZYxxL
Hp3Djqwqv6+GpX/0nSHZUd+YPvdpRGGGVLdni021W5eBf75QJ14jS3t56S3aSrdLZp0H2UP3qIeC
XWeBuNaBliPW4VaUXrAIneOgwif9+56kU9AfcBM3w1Twaq82FOkxkdvNSW6YJJ/aVM5olJBp3TBw
j8SpVPCqVoBfpcw4wEBk09aFJ16qHw7SrifoWWk/bmX0CpqSKdAnvB3MLgYyICcFyxQZxIk+uTzJ
xqz7CSY+uQzkwsqqqZ2wm6gtFqAtrgyHZWxCFQW9V+gdX81NkPpFhuJ5fSAaH3DvjjVFyVgxklEv
zImHy+py5Ru0ClqoCEuvok8dKHMYk95FX9cWRT8mXfNajL7Ahr59FtAZ5bvPUYS8WnSjPKR2fMcH
K+x0R9qdc7oOfPO5uaeTsNrG8fSPsfGZyxEL515co6xppHeysN26m2kSlsboMFMrxs0JU4xpBAiN
sPEE72AG7EvlkIRcEGV0LiaZmKSPydRHwE5D6sjGouHDAfn0VxNYk5tlrkV28GVuFnlPSSFcJr0W
G/NnVShVtDID+6gkp6dVdFOHDYwM2+VrQPJhaw+QWBG8K8oljcpAl6JSnG2yf8RR+d6CqbwweNc5
xy2CPaCXBeSOImpSvZ5LNv5zcih4iAHlLHXikOwvEZ5RAK8xOGPd5AX6jvDltLwerLzAUMQ8pimA
SOPSv8Gw/3mMU0sik+ypyoRS+HX9wCiOvj5Grtn2AqJD99VmNAjudPG2ihzJW5V81tyk6ejyyHyA
rH4aZNHi+LSMuxfCXMNW9ytvZcVXr4oljOqY0FWpi9sRCrvbbif8uGZJ5eyvj9iFs7NJvB0VkNzK
WupDYO2W+Q5gIRN23hHbXb/kKmp0KHmbKGFzj3/cWjMoVVBykzBmvvqwph8JemoZPuxl6HhQARxH
yNlg5pgjlU4n6qxiLn7202JU52Ptv6WFAqo6P+vbmgQ2HqcQu6gtROpyQX35kt9BmzsN6rTd7LRy
MV1kNpJidrtIFJYsaYrvl84cKJebst8F4TJlfx08jzivjcisn4tUSKq7O6cQBvwEQGqK1LnWawVY
JgjmCJTcN5MpukbjJkLZOHT7F5Apk8qBJOh6Vi81QJlAWQIEAYtepWnAZ+Q8KI45MwZJNnWDIaTw
BLrbsMlvqqSjMJe74LO/voCLxWroizaCszStzYPXOXMAwckB8hTllOP7VXzomklyp5HaOeU7o2z2
iEDTP6A6MmbpiU7NrT1miKiIbL/NoDIP9C095A2Qa03YVYeKk1yhoXJSoNVUq7FY4SYwNxelx43d
blsFskTeJIcWAVHiiohO8GBwx6NYiZ3+21JVLBAokTdYpQmPXWgqPUmXK54Vt8RUXGPsOSjVejo+
0L6b1bR8dy9kGQ+Xuz1Kjr8iRURfDb2eP5H4HRvjSqZJwRl28ys6OYCDGVWjiMk3/rSbwPRbUprF
on3Jy52kbYgw7m48D0pqCJTDnB5pruxfmttGG8CXK75ZRjIuqJDwY5dJ584liQaOfdGOglwv8dwb
g27y3Gs1hTwGCnWBdJeFIl5jsAiIPVujwjiOvSn4g+aeFufEjFpeBvCtpKCoKyGa2B/yEpNo7BoX
kv8H+glbi+xf/5QPIO0Tv5bJ8sVHjnWeS+2fxws+Rwe/jqqpy5CuTIpJ24OkoXdh6ZAfU+xreEz0
nFkFo+CPvGUvC9Wi1S94RZaiqLWxVSz+/TqKhSv1eXA0njcNH1OQtb82C8h6iNLUZZoyjqdKSw6I
y4vdtHK2I58SKot5HEpbUIr3ZRLiocT0WtDybBj705tnkpiq1c6J0A5b9NfYbzlqqM5C8ki8kCRT
p7rCeP7GfXA+h3xViVyLYhShy7AS7mjPB1EoxfTL4NoU0Y2A6F/eVLvkKwCpnsctiXLdxarg1gal
sGQyCRafAwqXcv7BPiERimxdBY/+a932RNOSdKpRpLbYYuabwwEVR6Q3FEywbqiYr+t29dP8bVmg
efeVY3rrKFGX+VnBnujmqictvKtyKIK3Y4yFbv1juOEvZ/Xtrnd1JAqxjGkgY7xJm4bP0EUa6wOr
WlYHlz1c8wPF23YsiPv1MJTAhTSQbnH/D0FNCO6j8lFQmhxUJmekZIj69cdjF3ztp+w1s/j/EhbW
gxyi6j2gcbnJBuwND9/3CbxuTqBJ59DZSCDQsVgKK9iGUUu+4QmXZlm/x2MWWdTTL4AvvkxVVAC9
iqdlgbWe4r06GGYbtcBPtfiYDzS8v9659nwJaQHv1oyTHKYDG0XMZvFNqDCSwgS7Wsg6VvnYSXBw
but5F9zd+80EUgJdtLkzzchkVwZfpnv47tWjQJJhII50Iw+R7tJ+OGMazuyqGnYWK1NRtKq4EFOd
Cbq7gCVBj/IdM8Yw/QHSGTFhLQJZFpepRE0qq68b7LrQvybF2Yw9aOM3GG4ptVsJ1JrmbWGqvMFL
eIIB8fuGea1wRtw0tHS1wXqYSGjfg0W3/h0kZEeN0ryGU01/MVh7VlHV/9s9UVCnhVBVNDCKLfCC
iTaV1QuWsLl6XJNzd3oHwrVRFDJdS+yR3oVomX0qxapo2ija8LbfzBGJnyRNp88QT6+O6UfjLCSp
5LKdYc5EHcxAYJ/exuDJSYHHtFKF5gH326n+b1qTxf7wXkPU4e5YphTqegFLtP6uOoLv7qtTtwPC
rR6zOTeVKmSank/ZHlSyj1lmFn14/Glx+FroNpeNTGqaS8zL5YcqSAyCdWYTqkFDvCDoTTgmovRj
RZPBAjOBGs5h1iupMNPU9jn4G+b6lThGHZmME3oW/ro5VuGJ7HtaQZaLioTeDwdVbGBFo/7l5ueh
eyDx2QtDPMjV6waZ+yyVZPo1llL2bCAsrwbKOYUkxMjR5/N65zhY04Dn+pF1ENaoD+ofarkAIsky
VlkiGt7d9tHu1iQgUgci10FVkqpk8FNgN207MDHZRBssdTPbnvJgocMoLatPXPzuhEsXbz/RVx7p
jizcaNG8E8VdgFBlodVqM23jV8DLT1FQZt239HfodHnAgmRfUB9NT3foYYvNQSBrw83IYuaGYYg8
I0lNJ7zteS7jcRzoce/Il612pN/jfU4+3UvypWM9gaDV2jRF7xBVG4kvAd6MgJnryOrnhlVRh+X5
NK3C5XSlfOaWnVjDzW+OS5WgKJcxmN6yOTGOKsBparb1McEOgQM1tr1UjTR2HflZm6uDSBhoeG4N
CUfLAmUpybToIg8looQrhKTZFhgQEGu528aFx7aUPIqzy/9RZw77mCL6lVgU7DzEUbmljX+hEymG
D6fGvNRi199y9bUUqvnIqhuUq220UWRtnHXGTCsNYGANCcoK3iiT+SXYA9jHxRct1zW5SrklFNWM
yBIW9lLTWxnulqD4FxJtQRvHbzFQqTmaCj2aJyflSwt32LVu1uH6IdYFUS0RJHp8HfAJ6BCLDU3r
3aZfsHGqTHiREbQATgf16ezJE/T1K0xMLy4FhY8WIkBNKbxiCrCNJPPXkg0R5GVFpWd9C+SUc85Q
Z9HVpXio0KFhw3CuqqAboySi10GeARKlt5SfbpbJM5AXmXPnpW2jIR+aW11xjTLHFOXB/WX/Ureh
ru/aFFriJSxuU8l5lwbC2XgO5eorvaI0N4xQz5Etx77Q4UEeCgx+IyPqy/o5hQuk47GSrr5qr9YZ
MNjxrgpCW867+A33INurJnIBOtOrbNu7LrhzyWPiILhqTBZhGiz/IRQK3t3W0ITM44441mXGNpjm
fiJ0iCGHZhOsC1JeYVI/ogv9SVczvDf2LbRFhureJd/3c4BmktXd6maSaj6ylNn+FP4B3zVCT2Bg
REQuP86AIh5pmg+BjPTMjC/sKQTfd/g5ybWNg238qxoEQZmc/d0R1TSGpDSyvjkeYBKAe+Aqb1K1
uONrkIDKhJo3s89l4RCxkplAn86yCqgJdazVsIwhsxo2HOfffI5hKbL9gfGHR+6Lp3SrZqbP3pch
LWlNiQkw3WgrzcYjXk3/AKvq3gy7zo4sZqTw+IAVynYsTRexjZ+/a8HDAcyc/air5b+ompNX+5Ym
XH/MTcBi/7xXcnJNXPXcw6R93tWRguSOzNenRBGglKxuCMmajzwTVh9MSihnItnlU8GtmW5eqLib
/AN6Whge7kRJem/y2o2rgaUgq4/pPkeU+IM++L6Yvq5t1BT+meY3h1Ay3WWYFnz3O56pvxt3qjmt
iucf1SePcaVSL/0erQn840a9bVb542G6FvYTN4huytwQ3lg+MFqe7ucdfnxfVUIH1OjAQ/yCvYp1
hilBMBUhl+X93fA1X8zAxpHtTQ6ikKdqK99y3J56Le3vtJxd5PpKiQHH2YtDWTuizZbI+PQyKG9z
X+QCg0YutsQ/RjLO5iPjfRF2KbbF0qbX/qPUJHvQ2Ch2VDuxpn2ScU8SC2oFzNAM0i79Ph3D9HWv
v1zXN/pPwSLgs2zPomJGKRoF45gRUTz9pbfULYpNQ4aN5SUMwbDUZEwT3Pb6LSWu6jedYYBeaBOg
VzAdIITEJP9T9USX/rJNhqY76nAhfwdpbOUzpHKO+w3WNwoaVD0AIP/JIsNzjf5HgrMrY9fSdH+d
UoiURLIob456UzVvMbsPG9FHRUgH6FAmjzkeHMCYWNrgC9Cb3+LPtnftfZPQcbTkjYaBHBwr7Wyh
9KadHk0p5uSWNrAg7jOOArLdzJnNx9a69oEHt19sMPQ4NYeeqss9+fg3P/r81mEcv2XRY7O/yHe+
zDbUtPKObkz5Skzd0W/ei35wDoC4gfkAFL0jApYGsr6l814hjjkq0V1neGfijuKMor2SE4cLnUjD
lJV48WkvI11I1G3f7AzlF5YQipgc+DiOQi2qBMRo275dGW5xCZH5yOFsQxKUocndHikeVfeAclpG
zhka9WDDhn6N78e9yAldl0HdTQoLhZbicLvVuebu5iTmPklSsTJOyUgXnLgbKBqye9gNOHfGLA0I
bnbNJCKKCILyU9TODrof4Qvn3yNpRa0wtus/6jklZxJ/xDWYItw7ssAYBIsIfNx0+EBafFLrUYhY
PxNzcreM0dLkL8+CsQvvtXy472SDsGswSp/ZNf4GI4AXqXE1MLVvzVkE5EFfHWEsvg6KpKoVr0Og
4bgIBlH+0+BAmSk9bRWP7krDAx+tSU3lok6WDe2GRXtHPEvLNiyW40R2jgdNBJxH2TjCJQqSfjHs
TjzojKGciQHC1JWXHm0BPY5g44nPGAHkYQIgxRy9fPfLn7f/27sxfT/kvXFq08i2KJSGhDxYenBg
fSjy+S9h49dLGS9bb+fSe4do/gbWOqcJygjIefHL0fNJ4ClXsuHeBUsk2//xn2r3eiWohuO92ZaL
pSr3ZEeUTyvDUKDd8Q0bnERP/bpM+L/wxkNzdabpc29w2539F55WXaUrV5b83CJaK53JSEMfcuyE
yFPU7pkLztS/zt1lkC6DMNGyTSLDTkyjCa4wThC3zvEVypkCXSwlNnTkpMzGaLFpy7LvpNTu+sLl
T5fG+SeOdvKhyY8dG2n68g8zIbYUtonr0mCnaKhQSubbhUN19GhS/LTwLgV0x/pKVAuWghEmCHSq
XNWhk1WG3lJoxk54n6ca4dmMsiFcX28Zp+gutclO2hJ1zs8pK1MpISWqcNGJBVZCdhv4XXV2xx/E
6ZBec0qHYM8eE8+hTwGRAL5292/2a76WCcPMVjLH/t4dS3L9e9iJDY4aaKuf0rSn5CsivOyiXkIB
FhDOpcgOfAUl580QpqxwxAJoYKzFypyqEl3RiGv7gW9+QqMCL23KsmSMMUGznjiuAmCve06k5pmy
+30NA7tsMcG/sQ6jRFDyQErTB/yOYPE5mauMb4N+ZDD4ON9rmA/vdFybKU/wZAkJ434uWmYGLh7K
eBv8YgVso5EdXtAsLTdNioa1M6VyZyUJ8KDIIu4/vSuz327jQRfNiL8XUB140z527hn+RHX4HEem
RG+x7gXc39P85U6TOPqh7r7A9CMEkUaJhMyK5gLANiKoTuNj3rLvDtIPDaM59gusM4+35ge4HuPh
D/x7cCS+06jlWcZ02YP71da8egk8YXAAeMcX+sPtqiY9w7d4nJ9inU9lUIrhGIHx3UaJQgQmOliF
GDl1BoHyudbrLx11Aa/xPv7M35fzzSK/W7gzU34JUKSplfxMpXy9tYUcqDv3HOl9Itdj7+ChdQF5
FrZ4zjfiOvKsF6ZanZfIuwl+cWGyejOqMmJNjBV9NdKLJeNqW8uX10I09rVcXlHiCBnLbt0Yv/UJ
eatsuCKTl9XD74Hr4ijedy6Av2NbDtwmr/7oDi/OdC6ej3qktwYk9Y8CRtpQLcgSMRlPrTrmzunM
3kAdfikmZOMHVckM0MepOoHRnUel4YYc9dp8DXt/tC34cKuNfQhIeW2Iu5cWz+Brc5KqQ5QVkFDq
cDOhRzf7SeKg+hXdxM3dY8Su1Ytv4reqhoYUQW99rnEVPYfhKDhlXevSLC5abMDHDki6L86Rk9dh
9yggF5PFp2EqwZOyeYPACZeY1jZUxD+wJY6ZA6ZDkLFv4O8e/gl2kYkz6YFMWDMso7lzVx0IWPbh
uaq4mDb3JWyn84HXP870Vqf6FK9r7Yov5BtKdC4S2iwaC1MpjtgdnzwQCdJgilGzC0oSXzAzBj0l
2uXv+LnbOmfIhGL02gGqFKTwwEMs1uIuf+lI3gH8GlSeP9L1b99DhclVyCCqe/Y42ZDOmuxva7zQ
DeQQbQ3a3z4z0m6/ICEs+y4XrGFfJUjfSigpDTG7+uQ2xdCtbKPFk/M8TXZCZHNNZ6JhtfABaTvI
qL4PsOAbKggQ90i4WEVvHNCWMPEthWClyhsFgboPRuUMZst+EvzIoDnJj/ZQ0l1rmyIFkNl+wK1O
G6m0M1F8BltUNPBCegPE6xngKVm++SSaPrFtqfATKS4T8/dd4Zv/PLyDJoLqBV5KKlqLCl8Nt9cL
zXu+KW+AAYiHjHttIzAxtAlFUHAIiB/6m3ffSwqFoK/G9sjJAdcjRMwVdqrvo2x8bLfDK2hCzdQL
O4qy/TPOOOKBuLpQvCbC7rqqYUkA6LZwujUdmsTPs6Of95bq0HShA5TLq+cVqJ+0SWNsrrp3sf1z
Zf4PA7dQ9izaYAK3YsX62uO5nAKaXUqOeW0Oq6tmQMCth2EaBP2bWGAVDTCioSLDWjGtGCXI5wQ9
4f9m4l+7gsmXsJO7sEZ98kWPcqWun53oSSfex3HHT+d0L7cV+SsijD+SFVV+hFEntJyaidPjUkHo
QeW9c0tVPOwOMszp65tqUbVc1eLSEdSITTWWtSwt9tDnA4zBJgLfpOPypscqHt7JF9dMas6u5QWH
MKajPNTljEpbPvJtd19bWfqzHyVHo2boiFqIJG0O6FN+aF1X2WEKYBjMf+OMOdY+IEUqndbk/JsJ
icJ1owq4yqJhNQuLNR+6HJCABxawp1D9OVgc/dUzghQRXEQQtVa0cfd3raNtRhT/lpQZgMWtqZE5
urwoXyMtLq46bt6VlsyHcoLrya6984XrzhTjTvCG46e6Uyo6qnLehNbxYbasaIZcfgJbKiK568Be
pQpSjPNHFIWETemrd1SnUmICZ5HwKQ6M5NZ2dviSZfZxW3NiTj6pV07U8lFw0O6OMMEvikJWoEke
AfWg9xNTDM+sU4HJcveQq1DVmRNC0ySQamHcwZaORrurGs0djmetVyZu3F87TuB8Y3KDE7tNNSiG
hx0HIG8OaowWaxnv8rj+HOjUriK0rOaQuFADgRCl63PFA0+C6fB3lOtvok/raBYgjafSjJASt94v
9UsLKHJdEjmCUcfKioRyJLqP9/ObCLi6ANudbI1w6IaDSZtuftgdJCg6ziUdICacuccYpHxNm2vF
TCb+ZGG9hfb58K2AS5TujaoMTduWi8Fa/hK6pPP/O+PTxI7dQFmvmvpaTkSozjxCrSH7ceQBir+7
I/NF1n4IzdDHI7gIKevAa31JJ+tNLQZB1HZ42n8VOJuSlxjwMZvJf8HWtVbZ3ayJRqJkwY1oiyXC
vEX9uq7j33cRUgFvLyBA0+3jFQQ/6m/la+ggqfdhSFG1bd5lFyBxNsQyTKT+fcQPYkJEGSHEOSIX
ZYLmMdpYcku+TWzTMC7/gXsz/Xodpws7+YwqA19OUeY7Ez0UO1Gnm4jStRl2dmu5F/ACyMmRSkt7
Avz5RBMXA2sdUA112lO/1M7nTPPVp+VuY+Fbb1eNIiTOzoF9uz0C41lbZHlIIEu0nd+fiscMI09V
I5yp0I0xFCd9iyvAy/BGqtXsZ+wzFVVD1gqJ3zS1SkbkJjTMPZH3nL2vfyJ/XCb3H7cDy+yeuWwn
Dy8ES7IOvT4yhUyXtqXLl0CCCuxClf03cOGg1KDd4RQIn/kbMUbZyVpqIQPcPgQsG1amVZ16f94b
XCwQjb/uJvDtNkfW69cxJEDyVwddO3LgPDBEK/KvbcF1M87459a1WPJym6hMtTy/1uc9Mg3+Lv2p
jtjzAmwPUk/83WgcOygP99JIkdbwz+laTzeL96Q/C2HIEbeCTd8w8M6OzUN3K4HA2eHEytnEtvJB
orw5Av+ugKO9hAe5/8+O/WfvyjhFucfxfBoqQwvfJN7rxry+O304QhPCVM4OgDmvQF1D6CtAU1mk
RqTBJh93bnBqQJcljbs4t8k0ERGmVi1lr9cEvu798tUd2EJKk+Vx4kknSeeZxeACVTsi/s0152pc
M5EahH94mTU8VIdIpMdoEerxlquyKQGafQ/SAfNRLl640SendkTeCpV2jNw6wZVjrVMZ1yAn/h7m
LpLNGlS3Pkdn1XO7+By87B2mK/yMTeQVgfuPDxKhZad0nx2iLJHhsvVgbANE+HQSJYQk1AAAdiNO
OaAHpekWTmNZS16Ud/gkzRyQQuFek0scYLfV9djW6nUWVjfNr/ToLbZ4W9nhfUyLS8Fsk/BDPk8j
EbZgJAtJqaaicU2JXZZrigtliOX+cF9bozbR35xXtTKLgq/4RMlBbw3SNb3CGUZNhkFaDK8RotSL
8ricszHA2M/N8eDOThsDBmGB2Pwc+dw9OurNSJC5TAIU4OtTKrj172lzKxMfy6Q7yJAHgIqI9kgh
sP48KL05melgUv0TPl90QucdryTFyxdv3GS47J8ioEe+V/Vkd+Wt+uHc1QpWG9hQU/JAXOMSjFaR
5oAvP1e2o7wHDCe32j94Tf4W0BiVgDZ4c/YNcJj2tuCFjc8x8XkjoLEWueZDhPQ2cp8/joaGfogE
vrbSLOqzI26boega2ajZs0CYAEEhV1LbHD16lRAGXN2bU/zAJbbXlzQwOntyJu9CaxHR81vnpUUI
mDVArsHW9CtvNm9/hy8S+wR4KeJxvLToKA6kcQ0DT2P5/1N63WZk7b0UTaTD5ROCN+2OZd5jErzT
zd2DZ6RN9qd8viik5bYwlI35dUiZ9KcGeueIc/MWuwlyhGZPWo+g4SZEO7v2C/JB8mkLnp7E7BZW
MASvX6yfJkTPsCFaiCLIQ46KqtaoN8wq8GR1TkR4iAmiMkPUq89Wiz7RhzjUZj1z/fiG30cZEziF
fGuVQduFPsVXjjjVUuinLTb3XSjQTaCEadWp+8YIpNeu7AunDVBZENvV5VJSkomF3SVhttRLL9ea
3jcirm7WlJz8tl++pmbZCDqnkdbtKk3b3lYqLIcKJuisCIgkN2LmtvjTTm6XxOmJou4NPXci5Mdo
lpLLc3rpWNalrCzSzM/Rqkn9YQCh//l5250bwhvFsYz9sYyY4ZcOdDW2OQYs+mlcedj1oJ340RtI
GdQYhtOFlcmO1xapAkVkQtn9yB/hfEMFKj3002ne6mGXQhpe8MQ0HHSf6KRqnnubn7yT+ArKCmh0
DTNn6qpRDVeevBinovMzNx8TDPe/HMz5f7DvTsj8QuaNle+K6vTTeBEnYDDXWx8Gc+LNHU/8nj19
7Nm7OVPMWt+wyEW/K77w/4+hY29KyiVRRfMG7MlfEG3G8XP5qD51hpWZ+AymKASb5lDcS95bb8Vx
Rgg5K/ae0rQPhXGxbOlXpV7EuvsbCYXj6jda9AXXciRGbPqGdndg9ZDOZ8BgHEhOk6rmpkqpqK3i
0qELHQfxh56VWJXzo6e1ET6sdh22YOyEe/WI8bJJ57vKa1N1erigXOYnvAN/gPUlHbq0o0VU1nlS
fyTwetU28aRDkKGSuoYvrqAr9/H7vatywT5+zuBc+une1bThnls9SrIFeFSPouhgwwlATj24tIKi
8X0Fj9irIZurXrOoBn5HOSGkVtfbD6+EUtnhDToQlfbk46HbUtImXHMXwdPKln60gKHvoyXc6Mc8
6nCyFSSza6CVkgCPJUQ8tlwjGW8hVd+xZGiSltWpt0nJcNR7hGC6mOTU8cpAfTfZOQ4SL2y9C8ss
qhNFkmFIIJDwdoKODrrLhC1CIXjPdvsKPgzcejUn5xXEwAjZhiKD+OwJqNr3OVGYIvhw/OMsJzLj
JhQkcG/RHH4nBklubxpeIMDfi4vMo0yjiRe4+4T1dQsyTX2wSI6foexH2fk/7Q0bA593A5g+5SXB
+953td6nYve8zPkm9vl0omCU4FtG8qhivjDhuYFTdgsilxRU3R8gCmB9lyJMqCr3l/wvIQlWTO/J
NkcGW61uklWmqEROEM27e0l5CKbJsHxkzLOh1PtlwfGt2VZ1zgDCgRbT2+w7sjhqHIyVJUGFE3k8
j7yv7nDhEYTv2OFWNZmoH/QMo1udJVPMw3d0y9IiETa4ggt8ZETOwALbIrISk40S2QrVacbdg/ZR
jCxKEf1dqNAuNrSNJaTOWF3pasaBhailLXlVJ8ZwMOezvcAritwv/kIQ6lM/JgLd6o8SoyKuZd1M
if3spzo9i4mLUG5EQO8i3QhAzDOYHx+icagOYJrrJMUeTTkMG4lJ5sw/OLlGVj3xNmY20MQsLE6+
+zcJwh8jJIRJhC8aRLbrXzSb7OPtLDcW0FF/Nd1pXKigtNWkbTYod176G3pa4J+qf3uOh0q+oJwa
FCcb74espZlbxxO4SYiyuque4331WAiPdyk3l/CLdoNqXBhHkPxbTyq5tn9to36x6VxULC7T5zwt
lKzmhgzLzvXZF3Uf0kk0308MmsatMnxb2NJEsO7Er9gaZQN5jpQDKu/wc1ZNcPJ5pEdyz7lM02Lx
2Dqwb7VObL5ZxB9sg/SHefp5uqWhhjsk/woC8soRg54AM3zWWGOMH3f0Fr2gWOfmlZN/901sM2gN
i4o+UnN0WCaCOiwhZttK83g33quCnkSm0EfUNd4ohZUxN99hxjQ4RBAknmZ2llfK2OmTEByRwuqD
YNhdFh4akLnYTMFwVrf1saXOR5oZlcVgDdB/4knl0+4dg6iyoJ+rLyNNVxVBigE87zgN12ISuzNy
DK8d+kzRbOucCKRbT//Yrxn+qXOYJM5aCz7ShTObI5DzbRUx3PVViu/BzgPCyL39t2X6yOnCx+nD
k1LQ3XaTJ6ChqFT0kUy/DjA7nldoIhp6KRPemP8OAtcYTTX5xB0unaCve1LinqQWZZ5wS9PWo+Za
i0QU9uOehK1E/zORBH6107HzuodUyqQAbQn7KZtdVRNnMRohEX/7lAQkPRXWjR9vaQ4MgGVFyYHj
PzBVkwH7J+Wb+E2kF+jYkh78lbjQ079Es1fExQXNSM4FFFvs0W85pCJslbB7XoKXiSKn4rBnm2/w
GGid5g4E27iEUUUgMfzw+4bCrGaT9dwHXNLbhiXzOYXXHBkvy58tWt9XrnT6IGrTE3+U1NCwyzRD
hKsJr8s3MtGF1Fvqni0oGyyrdUz6tSZjOBgnH0xDgL+Dq1dda2DgCl3ceg2LXVY+vz1prXx/o6q4
HsuHFWWiLmJF4WeqEoB08bL4NQHHGXkb6TORQ72SpDGqO4tz4U0Y9OjruQkeDnQ2wnAK+8u/L0ss
MsTgkCYYxiBrBssuSou8nU15LUEo859Dh5laEesu8ihAaYCi8J/8i+1C+SWR8IAg3H2vKvb5kpgy
ctwI27iVCpiFxnJ6rcYo1saEgcHADbLUpPmI5Ipch8h+vr8YX/40vsFyZPtcbYoL3hgCEf3lSA6h
hjnXgaJAtHJsLfR+d9TIGL0xq6TJL8FW5XUR80bKRMnYqZ/DvOvh6ZhEWtwETFS2x7luBDTyGxxP
/q+jBTu5LS/etfznlZ0Yqz5i3woGxMCeNum3EP+TAkBZm/6ZvomuLl0wGavtm1qpW2tjLGgSSCXh
2BI5SGreqNdo0ZZC9CLNTckv28Wdr+u/jbsnuNIC90RAp4+/sC/RgrLm1hlFk9rO0/gZe0T9FNdJ
rZYE5qA1Y9Oxzlqu4DPfAIlYtnKwolFtGo/YMEBCG8R3JYaStCcoLsx727y2GUTQdjzUkhfvnaUm
aN2P73CACS9dHOdZTYuDwARiD8CgUmVol8x3V2IkqcWDu9xZjVw1yGX7lj5cDKSfGl9IKMGz4oaa
6/AzTFdDQfuOwYxulh6Z0oUE0UZSAfyX7VQRouKFwPLkr0n1ZrZN39nlN5nAJVuvzF2rNleAgv9q
d2xbx3hLLjAKw0C8SwGIDv1d0mguCh8lhaAxqaVvy6wFtfV+cXqA797uytSH7HQhZwMT9DBamWqT
aU7Y86YFVX3Gvr2yYHBs2sm3Cbns4Jaf0UYfpyqhot5pCRyaSMx2kF79XfMTlTcylEDTXhaW2Apx
K4uys+b32DgIfF6iFFto3OXshtopimxJR2//TAG0XX1phcpa305ON+x96h4yrbWQjhJ3Db7HLhd8
4DdK6FTrUgv679jUqfQsxUNMhwr42ZWW7zdCtnFVOlMcBjWbbOf62KQ6k/om1+JN+Or/m8Gqi3or
swTtCcLdwHHJQEquClR4oDoAzuvdJqiEa8eLcaEr9VzQH6IB5/c+iUhfFnwTCvpYp//Cyp8NoOCw
QSr1abxYO1xf8S1h7S3vFSuCSVRtBLE6xsN4Y10vxwwXWT7oTqwHdc9lBzkWzJ3C9S76AE8h1xBc
90NHirIDIJJF9ZNdWXcVBnX7m6m6T1VRqT8XfFphYGHHBvuGP7p1D7apEZXr8nIGiR1zTYS1njH9
ZCmsvU56e2b+uPf4iVBgHDJJYrf28Yw/8e91vYg6qeY5R+mDsMZfyI+wlLSlvywA8GLMJLH7uK6o
yQSV3+I7Y82eKfmwEVV1y3XVG8601i87nB4VdWtYqe7RDW78GGIsIP2KFTSdRPNmdVxpdi3uIkKV
vYHqfMb4i2p4HGt0uRtWap+237VwyoiE+qyuxpYXRA7U7hilLW6CwU0RYNlr32QUw47kcbO2D37e
GPKLbj3YHhPCOtQIB98/YejCrlIe3sI5lzHQLKMBA5OBhnkDYwSXUZeARD/Z81qXjW/lRACcs0Vw
IPHaeVx8y55U7E13CQAgCtkQBr4WWWyv4mX12GYZR5svSui6didkIcf73hfZ2AtOUGbWZFHsa3iU
puWs/p/U7MQMoppGNLvlR97mhmvtCRkcAxYlgSLUU/V3PeDzO3vLd9UYLyMI/REWOf7/HyLO8OLo
8HTJxS3Xef0nEdc8PeszM3zlEiK+jrFMW9mq3l9y2ZlPj9FEhnd0L1W3CW3WU4qr+JJMWfqsrq6o
0EEvpMjYqB2ryzdCZJbbylZ2x0IvCjQb7DugzfEac0DXGVA60oW35cIKBH/PiCbEm39J81DWK1lF
fXlQT4ZDnaR4Bwaxn2Sk8IVDcUoLXL35jLSgdr/L6UWkZZnS1FnoPxgkMYir4qEl8/6E+6e1XwtJ
VeGZUr5NoTgm1UbgLTJBADzf9np6L3Nhhpy3zP+Vy+z1L5c7npp5JGeH/Yu6t/BrXIX6jj0o3JG9
ZJDqsuSN80HtQjteVsXwadF5yE1J442wql2N9T38LFYqdfv5+mLl5SvVXdreM5QY83pU6QSoJHIW
r1QT9Gtk/mm/ylMMIr1tYHT7cWPa7F5BX1nCWymNAo8fJ5Gj8fVVmUj30MYd0j0GKs0zSuJq4Sig
XjTwE0w8HelDBJBJvbfWOvSwx9MaRgELz7tSP4ExOa5jL0BaJEofZd2h1YDhqKNrvYRq6lpIoT56
0mFE7ewwtS02VyFTQot9mNay9qjQDJmcX6CXq4vfiIwVN0jK9doCIKf9HJOcUt3A0z1AHm+kTB0l
c8qZeS3wgPuhveh5+wjpt5dj4V9agyUCtqFZvjhbKM4NMGYkt+hK97qs1vR3qLNtXlax6zgXbn2w
Y9RZ0x2R3DXLAd+nlT7FxpkZtt+1C8x9aZpDUmTuV4vYG/EWl+q9tCCYA+0CX0ngc1GI8PQiuGlB
7Qd7UKvC/xEPMZwxHRDQACiT048ZwwyRrdIKz158JKt1nr0NllunB9RUBzeHGUpgu+FhplSi7Zqe
Mg+ho3nIfvBBUGAiW2aOwVY3+IbNpapc/U4G97Mst8FxRAmyDn6MzSLZwhxvTf4zIcEFIQRhy6IP
kkg0QOBglJNSlZM4s+okr9iIX0V9zpibuuWbEzvhk1oVj1N5iRM65pp6xeLScEJFGIj64S2LDLFk
OabBAl+nRJa+jOsjXdKp63JjYYw263ys4KJumX3nL51SuVg+ZmEib0V+ffBetqIwbhi2ob/Ni9lK
ax8hpevQ4mLcO7DeDbsM+MATE37i0ICrRRInI3EZUq54NMl34dg1hsTleA8dzy6J3li+x90tmlTU
EP4ForIFjVLOGR4jKuKhUI4c150h22zzl2Mr7O72xLW/jhMlCNbm8fZpep2JKlqQD3KdLVxFuQMd
Rl5P9TPgzQlVWHgnvvipOU3Pxv7o6C5304wtOfDH56NSAq2qGiDIDQ4VRHYJRlI1MnheI0oHBTTW
AFpNa3v2ef6dcsydMAfOi5yGmJzGK2GUCvDHnnP+rcOV2AA2dojoNZg2lutqF+T/aI5dooEuIISi
k7oPmPipX4yAvBlu4fuECaeWwQL+U2pG7TkoRTWh4EwNW6hUbET5lXgnUKnaQZ2G4Ld4kgH/GQxw
r0mVa3kUwlTiKLM7DW7obATpvIFs35QptW4bNn5jAmVYJNs28hD+92Y6huLRUShhVUmodxJBKYvL
xtx/B/y6SvDoW31tmwqe39vLw+84PiFiuS/xy9OzfgtxNJDLU0lbNAdGjGAwMP0ElRDucIQuzXjY
hro7emgCsR/L426sMKBpQi3QwHuFvkVYdkDfL1jbjrTe1PqYKpMtdiJ+NeoqcPUpkcZK2B1l+BnL
tJDylkCli//XaL74PLdNdBrPYYziWuXbo5fgkmq0sFKGXM1UZ8H3n0b+ZptnpOsbPDEt7ApdT3r9
eCUiGpln3nbcr/53b9DWIPML8YAQ1YwzXkamCLmmGzPlEUij2xf7/HMdrlLwxd9/tmBfVpqTWxy0
IXuGOvOKotjaVcMFn/CMqFRpAV/2BZB4E99QaRwR5A0vddyX3SsDEwlwrd/cXLyDRI+2W7nFoano
/4lvNryPi7+6brM+z/TeC4bAfnjxYTSgIhp92yKBKfKAJqKDOx9GOmTxMXsst73SVSkapy0EvE8s
01LiARYhQ0UFyW6ewb1lfQpq//QcaL5lZiJuMKbpIAhrYpYSG0VEberbtpHX16IA1C3x+GiudrH5
ijCdld69i3ltA6NICE8KYeHgmyaTHZxm55urtXHLPXCBpjt60tx31I9PKqAcp0932XYiRpf1VZ7X
Kf7zDrESG9vttgxbeZASBpAZfFsUqeb7qzOBPYCmKoOf3mvYuRpmPtz0C9qbRhkPE+8+KiSvWwoY
hqjr0iUF/47K3rS0sam3ptP1f4eUuce/piSMAfx9/UIsf6OTVTNtZMZ12LiBsJ4DHyHp2W/N0Lvt
D4xHWHbsjbPegS51coJniwi943LhnXW9REJdoPD0OpHSsLI6CLyaoB7IKJeOTGXJgDeTdzOdoTXk
1VgsIFcPVuuOqqAkfe39ijELLWE2ZANvR4Rt5duKsjv9FKdxz3uduV+mPU4iEHeKPGP/sdwKN/XZ
r1X4UK7165FWD+NlkGYZofbrUJ1ZQmw5OvVPN7Ex+QG0NBhehIdpxHFowndl5lIL19Jj6bRH4jv+
3TeV2QDv+PCJOyKgl9Z/WMFvF3pv5J8UoPEvrh0D3KA8BgAeqQzCeDZv7Dal2ioVf5Cr8y86LKGe
hW0p+RTe0JPNiKdTThUYPx8xLMyT7EvqHh4v+K3WpozcRooW6j1x31KyTp07FXDogAqHwoC50FIN
1t8mGKkzQKQ+BU1vgL6biE9wHqZ557ANg+DKTfxo6bV7whupx2PkpYIC97btw2fXAaLtwzOT2u9a
ZFGMp1K44zoEFDhePAxLGSE8QOP7n/HRvwMbXri26d/InuUL0VRW0fFsgbwAnRRqO36KLwLBg/PO
XpiW8/cd9HnasT5Yte4vfg79cno3ZGiSxIirjEMGCoE00Kgl7x5KQyOEbUfIcN0ZGzDJwLDfZFvo
J/UW6g/CEN8+7DIxO0BVDpY4nJ4AfE9EOJKGQKW6DqwFA35+XI/remfxH7xmyLjgAoQzFdEsrKSW
T5LMAQDBiLE6HUV+wp1lQriVG0Fvtv3CLpx05FID8WkhWyNins/6ZbZYZ5v8MbB/36FPURsnO8II
r9cm0DNywcZUrJWBRslLDBKu1O63QBgfX5cAiJ8daEONA0C178xFqJSsu/0JEohpspxYm+8rUyFQ
H5+MUHIBbbAg0qZxucAhQ0WMBegg/Z3pSOOIic/7rRn29wVSNn0vXpSMmFJWI6oBJkjIOKzYuBIs
vRk8ZyISLm8ZfSbsx/hf69i3OAY9nKMmpDkF7lt5sIg6XfT/gaFO2BpJ9K/ErHqRchWlpjXN7zOu
EWFoak3bJ2BZIMhnbdfn2U/B+ALVKn7djyfwxhSfUbJ98W1NJxtg+BnEKF+Gw0L79dOMf+MRcTzl
kWONsAiRM5Qpwi2HgBA8lc61SB8tdmGZSU8KWS4jBAjshBIybwR9DVEscjzKBs9YP5aVV+SrAssf
sQz8mflBP/utz6copm6CSDy13X8OD+gkscZ9WT7v/iBjsHgMxI5uQrSluLzQ0PEXicjKM7IdXDIV
xnKXj675KFor1bWUu8t3CmuIdJuu8cRhR47P2q4BKNgD+8Ua0Q/gjNxlUsu11NYDWjhI2gRBrIG2
790PPicegjCE/kodBTuaq1TZqBN2zxr4oaC8fwdTqyxKwHEflBsc6f1f3JqfPxlekOm+pC8HW6os
a4V+Vza9u7GfDFgZtKe23oAJvJHr0XRA2Ae3myCq1X3aMU6AZtpKAEHWNr9zWqKnI74BTjxziyNB
IJve05kgcHe5uJDQvzaf6KEhC30APQTizOyE1BSKgIZBUdqxbufKzfqfgsw+qn79Z3skDUqI6Tn+
LmMiXIKyUXX6Ji18pwoLp1ZmwYrHcfQYF99Yh4Z2PUnh+DNE0RCfkExvYDDySUa5HbW0cxQP3d6E
soYeXUGxPCB7kRwM4Fjl/qE7yZuNCYY7AHBNDHCDezD3+A0n//3ZoNflHO6+riuPZtHTckN0tEtt
+zr5Z3v9wUMxrNfcnWfwc+8vkD197YQ0VtTGqSPOvLEhD8OmllqnKdwNFKZXXpdDR0m2Ed8VLrzB
tziSWFtrkBAUwJKpBu+oEdNAJ7kgj5KqBytxCS2I7hc9rzXBw4w/Tcsy4GudsfevYTaZRyTJfM/5
rnoc06uQPwjAyso94As5LqJjQ8dZ8V4ty2hbL7/aHLxdS6GMqB5uQEvCGU1ZxzQKj5PaZk1DL4z4
g6g8L96y1qFWUvTwLg0qbi5bPn2im9BNrJ84vlyNNrFTIEYyAmaBFF+I1NK5Tlj81qX+dF6zzyEt
sd9ru8OZqask7PwSwbWQs/kJElCdvi0JPuQrL+MvvN6+fxlJTt3iNvRQXA3zxkVT9NsAPTA+zhLa
riAOeilrE4t8OUl+f6ugnwvtZowXDNsDAssdtAaLb7elCJc7GgSEUOYopR/JrBY9II/2WQWq01MM
706KP1reoUV1w1nzxPYuo0w6e47oCVetfLDiL+Gk5jGwPxsNINvcocM+YIUr+eE0bkaYAWDz2wbV
EPl3GfYMxQqtHFK81vRzXy1j6PCSDnok82PbOAHM5m94YksjWjyaIeoohmS1QPj79PbULr9YLILn
NTn0vI6fBY6IZNhjU5JZpQr10uM/jc77Mozm7zs7+9S4iFrNXpZcnfRToCn5qBElHXC4kKzN12pX
dYyjFoqvZIB1caQDTov4gJzyHYKeyXZyjeAKlWbRekhH7e6UMcWPpMUvmxVW1oYu91nPHKrrSdCi
a2vubUQ0R5AH1CfHYRBB8rwdVeP8pFbSZzzIn+8Dtp0Oyr7D+eMbBW0U0Yn6fi7/4gQmvDyZpL6T
dOdDxd4ndhdGQ0beSSZSpwgUqnWe6sWEA5UM88/wYiELcBTSjrsWrdpZqJEEY1FRtgYn4cqDSbkO
3aGocFEj5B9G1fksHiER2bQqyMl11kgguzaVmZos3lokQshoXaSWXGBPeh/Ou80ecrRdAnixJL5H
QQPfQ46xb8rKvGWj+XXj+1fgcy79RDiwoMursEV+ZX7/BG0DQ96NVRFZy6z4DA3HH/mK1WZSCL1j
TO4Ma67+AiX0c+dY78kbVSxRpFgIP0NF9JDD8WJ4T1+VYy8BuFPEIuoQ2J0rPU2/rGu5chtC+lC6
NhYc5o1n1O1Jfh98zeN90cYhmbkq2SCu9Ge53q4t9STfDDM0mmPDsXF/Quw/ToisWZ8U6gwR8344
ZTiEuBhh1JN6FKVFMfgnsvo+yrNNzRSiFPNxDUTdeoZMGW4nf/leCTtC+bXYm9TNg1wWaxAe4BJ1
0uuB+8DNWwnnQ8oEgY911uzOrrxXK3tjEdZFXb70Ya0HbB7wzkENKs0FvLixO24rcxeD6Qj3wL2j
dKaISfFKNWGIfHg4kGNTOazEntZ4Xz5kcnsscBMFNqphtnXjtGv5B+54tQVnqNS6kpxVqBJkb/f9
+fEyghoofN1GrRwoNr4RD9iscv6elBTnjNSOI0AQ+0i7+NVAY2gMzLsY3tno2ZrNnsdCRJmS+AI3
LTkYO+JFgRhBLlB6tmqVepuL1CzfbivxDYYnQIMopIocWn2oHANZ3r41Z/nKSovt+ZvqT65cfOPx
Jss78qNmIGjbaJfzrDFjYI+gZ+jWOwLVOmYgjlx7IuYa7CzugS1LRnaLC9L+zJUH9OZHLrWC5/Xs
wjHmVvvwbZmnL+3dUqzKWp5ZffMwJq9UZQuIAQkCdEACsxwyd73zfgCz6kilbWYamSZxssQgB2c/
FmMNIWxb0VXKGKBfhdizBq2WfMqrWt+Y5cmjihn1XKxrPrOPBCrACL37m6zZ7XSogTLBSr1b62hn
b9fKD1a3XOnqmQcNx1WN/fTr0gd43nJ8fuDcOu+Rtq8enIEUE2Fb8rxROCBSWFLZvU4My/coOz+2
5+XvNWLykIQ0VV/PXpNrSRr+ldAtoJRM7TrRiXGqkzECYXsFrU3vSd6T6Ol2Q/24ob4ZqDzGVG1U
zcYctn4UDtLVMwEEqjKifVNH/bgY7JA73ZxOtOanI1ZprxS6ix24sZoHB36wnAjk2mcYDIiJqBjW
Q2VOJ7gCm5w4KrckRd0Cf81JxnHx/38pfIK7GkEE08DvdsiFiJ0FQ6LB4rmcBiKN2lH6RK1GHBfj
xpx2r7ok9PvkxqK1YH9SHMHuA4rIzHeX8ejfTffX4aeG01o5HZOE6jEnCPR5cg/iZZN1PUewS0tO
GCnt0xHC0owp4ta9XKGh5aHDgsKBcj+cHkdZo28O46AuvoajL9evT6snRmHs2XuEYRpAclGwZ8s3
h1zRQS1zL8JonwQUsHb84bCAqyhyscGNyWRGkp89cyZHSlf7yVPE/1+nw9J2Bs4kqinyGgXkZhc4
zlGukB5W91GK+T6PtxEfYi7Dnzmt8Trw/AzD1pYLvkoaYZoJZJDqWvg2iXrukSY4+dN/hfQVrs4i
tCmBc7ly7JaHdKztyPnlBd+ruRUrRbzRTS8jYsYJAdNPw+fl0+DzVhZQeEPKJZI2CHsjdow8wvBr
SwwJyDhAXJqvMPRe4MbX6Zc2CGPoit5w1C6H8qkC6PrrxuQ0i7GB23ThcLlb+G6gS0NsNOZdo5i1
2Zz65G2yJYZA6qAByho9eWZ4kYmtb/7JTeLiaBLXUo+oyIAGHe2NcaK5sxSEHVMpRZvngsg51A0P
IR7eYjt1IfPyTfkk5uMY9AP73acu4kFwORHS5ihqVLnn7b5wNGPumHQJIiiMjaHFb9kgIEp5jb2P
TRUhIIWwK8cVywKzz3CVq1WGlyEa36a/5OBy7snNCBeeEkqpSlbH3w7OlqL0aHYBbtmrNt4Uq6O0
Zd1UX3oryo5SXcAtXx0yV+3nAe7dnUQdyXnBJO4OtoIxMBoAN+v0yiTzZFjLOW3FB7+kv1hWpGxb
JIES/pgPQUUXHcQUvzn+MVmoPxlgBV4ciFauPf0HyA5uba8cCG5p5gEzeVXjtYa01oE4rYTEYE1D
Rn1R5Xai/4mr+qUnLwLdkUPpQpq1rsv+yVJMPkuaeatX+YHKCivJ93z41Q5BFgv/tafo+2E6Gw2j
+1CjOD0llWz5My8mCIi+R024HwPpXDA1Gx5NgZELXTMXelXRhdvbw5hd58P7M/u+SopSNROITlJr
95NmsdVz/PsUkUbGKR1yBE4bFc3kGAS9S1qJx8V/4jyjFjBmIfjTnM9VAbgPL0zIjxBI/IVKSoic
k08O5PwarVG2nIXPuSiCQaFsQNC8XkrSWQbRxqwkcbVBoa5vgOLITe8H+XjKnPRzYsiMZqZIn+X1
sY8MChlMmLQ9J/yTbxSjlpnwIY+7VU76Xz0nMHUu5xyxASM1i4m17Gh72G4N47fCNRGIk0rglx5p
vAi1Ou4aJXVYSM2h+8jMa45eqC6/BXtmXiSjjzv6HRhmmOtXDc6pZavzPUbrWhqOuXWZAO4AE717
c2vzh5cuKyadioxGA0QpjzpDM9zLtc+mWl721czlrvep3U661lRdgUK3I9yzqE/7dSeik6upNyjL
OKw8d/Jf0M0Li/bNi2Pqmz43ZDPLQIoTEjT877onzCsYxQAmW0bS7xANlN7YNSAnJKgHcOq+l1fr
E7zl8ePMINYTW66rUQDANuxWKi9SsmoXhI9eCc64tVUDtKKJTleoosvLwZGoWRt+ng+FYOpsmarG
0nHnE371vD9ySZHh1odMwZC9HuK4eUe7QFxg3vk4LZZV62JgT3MwOpD0ybDJdMzd9Ue4uKfSSvPP
J7LNH7rhIPI8Z6pFVLRoBeouAm7UDh8Czp7LOZaBmelTVmGI8v0cZovbDZzodS7jJVACG4lTNhAa
I2mRRwatYS9bFeeedluO7tCpRbgYe3AZR9qjd7TFLZuUijZOa30n95pSCl6y0MRBWd4J105pySqk
gVd3sqeOrYKJXswmWv9A0rWyDGtUuuIIjM49jOHXNdDRbFKukPp9xryaGoFz+5MhnasNiRwnyzKa
GhbWkZZUaWRI+w5Bjf+f7TnzOT/BJvSc0yjrgg5qaPiwGOC/aR30bosEf9NSZPAgl9Ctmo5+o6K3
XcadbINp8GXh3FVQXsEB6NXkAUR6z7cfj0+e1Cpik08ycPeLTkrmq0c/+IuniBQ7NS7QY26vqH5/
eTqpigBrm9hCIslZEg5mYqFGZx0SUjBzDweNkhlFWbhy8wCVb+9SKQDm88MHEFOIFBudPh1n6hBb
Zh4JkXh/YkKGRI40kEtu+aF93gDieMB7u0YeNcPxd/jn5c9o2xhjIDy3VIMQkGcPH9PaaaQpkckM
rU4915HLNDnOkvNn7oPNwC1BbaBL6mO9yDpAk5mFJ9B8reK/TFmAwS5U1asrTXh+75D3D8RmH/Ao
hX8A5hm94HEpnePIDypOD0BLAE2Q9z4XI7MmqErChY60qCm4y/M3m72qNUIsr0QLLfJWYiSqDAeR
EinNnr51wgm04GMkgdVi357f31goBF+zLCWRzSuV721RVsrT89AChulB2EfynCfXYc6xC82PTsTm
zNjYYLTJ9h4X4mGiG/MNQ9CGxWrlS16yPFRT6dHsWV6NV/lxbxTTTG70nRbRAZmsfbsuaML7W89e
7t4M7eGhoKF6xn2Zh1Eggc3iWPwrujL6mthN/jU8S4swvuGN9KaGIUOzGtDGNKZ+8tM2THLKYBLc
RyW1dlpAGWLKk29nDYSYyq9iR8lq8cmd0qinfWT5UZXyJCbZpRW12HZT+4k/tICQhvWdlfiAfT0w
Z0wrbSCWbytWpNPkKwA2olELD3EiF1bjkNeCCgfnFvfAalp5MvOt+kAvQI7m4YRphmxwv7bPeLUJ
iOcNMXw5OppXjgkurxHjm76NQxxOyaC+1/dizYHo77ACcuzNgnV4ifk0Y/tAq6USnBEAMJ9ja+4X
KfJwFJf6kqsDnYTa/5bRpV0YZaU5Qc3XBu+EGgsZ/owsL/6O/fHXiL80rsktbGYMNtOYnInWORD8
sjFCTmzTnNAQ8OdtMD+U34GGSX53OXRXrDrUbTwz73ISC7dDkegMW1TYLzxoHncdVHmDISgxMxFV
tOO0AB0V5hySnhRU37n07WxnKhF2TRPhPKKF+Fg3uObFXPo2uLZnoDqzlG2/R/P/8/dfsD7ybIul
SQMcuTXyvm3lcmAm1WWZFo2ckQma9hWPoJI3LmBu9UqJZ1lVkncwCSuXJ5pP2QJlWoU17KKZ/GR4
esUyNdOUEsuyh2Okrur7MzA23nkPKsJs7xCz2LVFRcBYcGOyhxFllxH0fFeKnbtNpxJOModXJlp/
Yqfr2gpEZsyVuw/E/fVzZVYf9jT26MJXSCV+V3ZGNWN1gAsugyKAFMZqQq959Kv7jtlccHJB7euY
KgyiSPx4okvnacspw5UOXBZkhNFctcvnv0oezQaQXn+pLYei6LEgHA5oMYwW02ZgBweHwyC41QqE
luCtrImHGCDqX012pZZjhHACfg+74Z0v1Weth+w50DYOJ3VeXgUgzXJ+x3J3wkHcXFzmRGwbyLPv
gWL2favVZ00ew/UcB6z24t5XZm0D2qh3vkfrggfgds1OEgiqsBTKiKAM6VMChuhDKlBiSlOKK/wy
GanI4zxjBbKLOOYYpPba7fENzzYTqcpjX1x9bwQXuf3wkzWu+x50t2vfFKmE+1jPT/qHlRNeFfC8
IOtMXbsXVCpDzBUWEVcIRj+4Cc9eFaCFz59Sc5q5x/TbDyiraQBBJlpnaH2VwoboQqo4HGn+9uht
yB5byQcKpE15tuagBXZz/ynWx9Sbt56EWENufNm0cWWCGOuEbIyQ2+2tBwn1DNs0shu2NDZg5zyu
fIgTIEr5t8p8Y6Bpl/g9RLAhi6Ygh1w1QkVkRui2GbXyZ4EiilVVLv1AVk9U+/LfhUE3SGIu8FUt
WhaG3I7qVN1FWKRGpbSxa8PdKl/SlvB9FCTNYo4QLAOVEOGv5Ru+UUVkU65acO6nhg9yjcRP9xzj
xmbhAGx0uTc6jQn0t5SXL2d7efcRueJTK4gYYZdlgVDOstCy3jM7Untyq32PDDfEtg3wqzHe3a1y
Sl6zz8zcaXgzFpVEAcIesE9CQiGj9ow/0kSBmWVvJJxB2L2MSh3boWjhid4yar194zuWMm8QCqCI
Jqs6a4rsreFfMJlCoQEmLVP7ZpzP0fAB9YlGStq3peoLKDNrvtM0gSgWQgT71lnlDQp2iPihS4wW
5yzvTPwGewYIH5x4mpdbXOE6qcUq0kpi/QUfS5KzXCqmPr9JiZip5NDi/uDOs+6EccwI/sxcY4q6
gtPydSopg7SbfPZDpffxoq4lcDQ672SdnsiJ0GYjleNaf7L9/7nSTGXxgN/Orj0t0/cdAAKfKm2V
OWLenTY0pkDpuI2xGk11B/zXJulwYsVYFG25/jK3zM51Z6NjKzYgNN2xX951daOzm1nDbxkpNzJq
US+PAwmoRTv3t3Yek8dJK9/enptEp8io/hfRk2D3qFH1QHtuSokpDS7V9WPT3DP73f/9Rlx0mBgg
kehM1qRBASDP7Pn0hXXuxVP3a/DIFhYFyooCdcyrupaLpquqzCNSygW9sFeWUYzbj00Se91z37pb
Lk2Oyi4Nm9fkjiDokffsc018gHUKMX+3PJgzhZo2WYOzCUrrtJOnm5nGmct0OmfsLQa9z34bfx/I
HVNiUTUaziqpCYEOHGsO4PUEMCtc9ovpsrtTnt7jejte/qiEHeN+8StF+/HyuN1CCkOibPTBfhUp
PA2kuHvSlpr0pldHQPqCKBGoGAFHbjoWpAjMydOag4eK5a21/4ZVNabfLcsc9z6V8kfyeGsiXd07
ihohvuDqGSCxZMPKNn5UjqcsL+APHlX1ngPEkysrI1ecCcGeitGQ+ZsRMgoLH43sntjhmPl2dISx
v0fa4Cea7doAUUwZrjlFtR+lNr51YufNbKQ6NOM4F8zzSl300VGPq15jryGuQ8LmTQwCfgbtdCx/
v5UfSxOvLP7jXawgZdp1YIdAO/5FIEbp6mfE7HP11Wfj3WpTnbiOdWHyw//rPA6/92ozthjAk3rs
xfDC4/JYh96r07EXs8T1gKPov1YD/vqslk3hk/o6EgZQZy0MjlKgyJ0CoVArv6ufVcdKc/dVsHOP
1IxXB7yjnoVxdoXgBzmQ9BRdr3wZ+MDoR8LDfocOkZQOJAvDOMgOVLG6h4FSHNnirJ22kQgJBnMf
UaDdZGjTXQmibkw+A1jpk6xCuZ/aw+BYtz3eQoJ3z+tQSaS2McQtTvyWUj6opN9LxP9AlpYhy5BI
NV3FfKVyhPyO9y2e9ds/yAMhB4NE480cOxy1PesiLAnNMNuwihjxA+leM4ZCAWyuDbTwWaaDQCjC
nfryP+qTNcf5EmuseEqXkdl5Fjm3nnnH7CzYAR9XTAdo4S+f97nduSla9BF+qtKpERneT1p0qNVF
tliqrDiDSFpHA+0H6t1IZ5+JmlfHI3/4zF3PsdXVLpAcEWpR8DRcbtagpG3EyhQR3WRFTHsxWtCn
2p8h1yOcgTfzf3F3MJ9PplXpz2hVxH7nqMg8ft7xKgPHRzvjTn22NpnK0RhTDV0zEu3uJWcw+7h3
hJJda46pOOmhrgNAN7WJcbTTX+aKBqnfl8EmNJ4nJrt/e54ASep4c/L5f5vQ7IF00CtoUW24QH8K
G527OHE3DGCAezHnFU0yyVIRixJYo9H16NJyqxuj2sGu4dBzis/b2i+0pyFmflE7ItXfY5J8RA71
3T2t3Wr+Wvtcnf99jF0hrai7MPjXVtMQK8a5lveStXBTce5TWXyl0o7qEPpgiLvbLGefkuSTnsQ0
hDJhS1E2ZOvS31v2GIoml31U28HEsDTmQQuNnr12BY61lcZsRX/nxYoQryg2WvWNpUPLXBd4JQ4t
eKDkuna2fj+K0LvpKDIiem28j3wAJ8ceF8qS7wtr4UxDBg7bFK//r7VHrolg3ap8HTUZhfab9eB0
g4kBP5WUDQZPl7UN/MsnHmoIFWD0Ll9O1oRwGWjlikOQZ0Zjt0teskDNA5+iTjqQJivKIejsyqx+
1Wn8emDfJzkuj5XMTvdaFtRRMK9kMdliew9/q/fOwrZdumRACW471SLtq6/X27d8nzMVtwRfhOb7
es7n9KO0jKLIJj6LOUnYHX3xeawBrb/EBh3wLvADfQAM4EnpXB2nhIlUZElQs4G3h/uonGHT31iQ
6ro+T/p5xigfdNedR77Un7En12/zyyCFHZcN4+2WaGC/I2y6l8ErrL5MIquIkdGA6BzEY6ttdg8o
KVVLJrqE1B2PBdaNuovBx12dr92znds9NLq4PnlCKC7KiIg4mzWmF93x5UYhAOdNyVpFJdkAv6dY
T2QGQGStSKZq9chE8Z1QIOz1DyAKiRkZsEkgOO04LmLIN56lQimn33v0gQrvC5kRfFQpePtUMWVM
OE5mxj2mleDDVOs69AzfAL6ehZ+/ISiCAHG0Kzx7yG8o9hNzOGycNSCp/uwEW1w0LbcZbE030VEF
1Ajl6qS3GW5cpnWjrqsQmYuTRPp7dR8VWY+Xt1+J1/SzZi8g0EofRxf2B4Q34v/rScSgiCAWOyju
o5ixe5/QeP9cTNj1nLYnIXT2s/CiILQPxyGnNyEJzMmevfvbkfBu7Q/zEd9Nc/r4k9qFqPTz/nqL
ceSKHX7Esx+1xJ7JvA+XYTwjzp7ixyJtq05aTCpEFFahxKakIhRxRGAfz+y9aqrHsrN6gOwWQFEj
Wl77oTPNCrltNnHyadDnQ93liafrf+mR0YAm6i9xc+d6JI5gXjq9idTjEU8bWTgLLyzCRPtZHnz2
FfYADRjSR4JpmKdj/Gdc4PvdK8O4wjW9dGMsDYxvahlkCtDH+y5XHs48L5FIWbFBq1aJlqkNLnRY
Zwwn7QGSLKXne1ECicj3Q6qndkPmxmyZqict+UVs4Ba4bH87bYgvqukkruQywOIqdV9ZSwbq8YIa
unCQi8AxakBMh7gk0/KhUohjCztUjIAp39katsOqwdVEb7HWMXGAdubD07cwZt52a+L1+QXleiuw
edifYN+lCiMtgJ5FlPp6p6dySpDi+jjApeshUoTRMXE0T2yCNaDI5pVRhzMQCA89qFMStqBqMEa6
EaEnG4Ks2r21Pm9wFdKWlHXiPa8d5HRhdUtWDx024/Snw1OQrgB3TTGE7xEI5PL9sa3InORw/bu7
YRPHUr9FN6XGm64HE7IOnxvMf1+H7gmQ8Do4S0c6PL0YHF2pYgGDE0eUuXSmoPL8uw0Naw7LXHUB
nHINUC/Qun7vwGSKB09cjUNLFGrNZBAq7TMRJVvHdrAXTTz7Nxdog/iYk4FR2O1fCOVRsHNdbu8g
3/hfhVu9W93hrHCJiyIIqm1f6fiDwhLDFa0pSSXNOdVTL7QJDpbvEmtTJV7oBR+KCRSNyMzoeE1d
LO/2TwlbK40UH4dNOaNiQ/6vCCgzYVqkFfvWbZ05+C62TfS/EvTBAqpwgayGz0g9X4NqIBlEJPnI
T/d6W7dvv2gH/O3octVUqxz3MvTt4cwsyikhnH+WPyxNQCjlY3rDLRpP1lDMfFlYKrpxfLcl/K8B
0wwgfrmW95yKoyLaZ6l0iM3BqpuZoAzJfWs8PcryYNvQ1fzoPz4lsnu+AahHlCIKbQCXFyMwWRrk
lAYSb3ooUsskWBLeC1uXpxWvvf+y2l6edn9DmFjBgIcG+weamFbPigGwdioP4Pg7bAUuu9HQ3njU
AJ0bqZkr4QIZpYF+ZUA7WwzYioO23TbtrGe2NEkYeM3ogBGLq8/fhGE2aiydAwfl5vxBmkH5/06N
wdULON8+Sg9k+R4iAlyTHYpVuFh4EFZROs9yYzkydWYVZRd899bOsh83rGY3cNVYV7h92E6/Yupc
TAOJZV9vvRMqSZfDP/qSFgWcjcUuK0tCdC1vZdemEirMGlwWKy2C+n9qLBBEbeJS5E/b77fOoM8F
G3rP/u6zhcA/NHHRPjJeoiPYyEc2mBHLfHxh00VgD0rQ335whsyyixdVv5gH7gG6aYogej/QAuBo
963wuqxjRyr+Rba6L6vfAh7SuDe+iryx95vKnCNX7wliJ2RqkuCfYV5jHzQB+z9+8zyWgmkf2A9K
kb2t0Q4pqoz0iHdf9mRbGCw/tfiq0xLcUjbuT3WOSqDrPzYi5oE1mVmIp6U+N4mBfOXWncbCNnFE
FseWGw1VK0KHDasgzIAIwGZG1QmdmeO1qE6txpE/r6UIUxvM6PCBBXh8fmgEDRNINPGEHAxEEMJu
gFxjh5d865qv9G0R0g68RhbcENlGZItBJcseHVaLjLXa8mo85jbzcFl40X8vq1pq38iQqRA+/5Yv
N2L5XsCuc0wpZslrv6Bz/kwPjtwciP7w58yoOvHFiVoyEhfcDBo4ewspu0qfYXaTTqy7BTOiFr4T
IISL3H1/8JuHPZXZeWOzPdhMvld+ZsX2GdlgYuzKNiwnzshCpDulg0UEsl/5Tt8/RwognCyTR2nI
eVRKu7gS0GszNUdjn4NUrIz1aEFzwuookBY/UYfDv/1L171z5dpMowHDcCBTKxuehetuyoGS1MaK
DcM70Bl9LUTbrdMJZkhQSCMnJ+ig4GjDUKVStlR4klc24ZsXnWdaLl4JhLSpyX6hYoKvyp6Q4+In
XH3CxD5tvf1YGRDaWqnr59Q+JecgKvuoV0r72zKIQ5ln2fCH5VEjTcM/0HcCKCwNsZOjcmUhMiJi
kXYhNx+Mo0/l0v4OXsmaORI7KiFEa8gxjuhkHanlZL3/eJO1qTuXIrRNCZRWnhYbp6soGwOcKUbA
1i+qI3NHPujsgmi/t3Yd6LNnTQyCxfILjedlqGBDdPKCN+IlNBHrikimkQ+S6CsqTjQVF/9bFU3v
U4A1az+JsrLsnOZOfn9RW9F8gTOsDLy6XoUpTfSvlWkFF9rmsCODaZInl7OZA/xtFi2I/QAN5K/4
NTk9iWLLVASF+e1zrMBOXggikWXmLUkFcOQP1etMUde0naVrgLL4uTh5V4vpPSOkXn0RPsB+gM6M
kuFBFlfQmpcDjxEezx/uSdDRAU5pn/pbT0emZG7WjpnRhuK8aatrMxZCJPTCCO10wMNhgKOx0Nea
Yqk0B8N+2IrnBzlQvztkem6iFVaKvs+m3y4kvv1bKPvRXfO5/t4Ji7TstyYsQvXzqb5FaJw6NBiO
ZghXP4dl1kPTj6ade3igvioTXFXjtsjloq+PwOaWI7aVmvADKJofBOHGkXt8ta8fwsWzfq5nEPeN
AgFl/NSmHXlpUC/njegNMNIy/HtMUVcjNBi1H3k3IbtIGpb731H8LO7URfvvXB753hg8taimNDrW
6rf1zMC5XVLKpjAOl4nXyn0cETNt2CzDZa0uDqrJyBGsTiebG8YjPoGDMPKt6LT+9yw8vZPVJ7vQ
KTX/2HnDDj1hZ9fwmfBr9dw1k7kfLqLcnSCKabzrXjHxFJSH0PdPCOWCZkedO5h5uX41a10UBb8p
KqdltbdLaMOYyvAMdu5fTs6MGxhvl3U5/TWSyTEBlyoEWWBUfaQK4fJNogWlPQMidPjLeppDSo7u
fBbjIjId7x/YQFqOZjWePEcPGBtqXbJ0WzUfAoCDOZjz4jwxHKHlcCdk6sIkh8GxlMT2tEEM40WN
+qDktecEwY5Pp3Z65vt4gBuARc8rQ1uAIuit3y1LGohfe8dw7XnAJH0wTECApsd+jY/GOUkjyvFv
ImoWK/ErZEh3BJPMfwAgjJoJhiAWVec0j9Bp7lY7VIkBw8CET3BC3qaLs5tDOlpUk5YV9JGghiCX
oOXG5P/jgBw3TYIMFKob5Zhwld0vo8aRNjXvXqSfvxXs6SOUAeiEABueMnBh9aqcZq4A9656Q4kk
Ml63fm4Zmm2pao9VLeZjLzVTSnbC/LviEYEKhN7zn0Fu6t4tAy9JjLDb/2p9UffViLz/Itur7V0o
sX6ce60y4IoIdJEnaAGfXz0N0kOd+T20RSitBugLu+V/M+kWux1lQ4Kc0BK+3SL0A/SXV1vkp2Hp
KdARNuH9YK53I0Z2Q6D/Bu0pv9HLEt32qwauY8Ujcn0DvG7CTaDsE1i1nnwnP9ORwkXJhtsyaoGq
1EIRYdgDW6fr3fUL6pPlGB9QTWh6T/oFiYTMWI7o7H4cJ5zuiu0dKilAjiIS5T2iyTHzenRkUpOw
BmOXf2NtBmUq16mfGMYvumf41z/6OBxbjgyOpLxhDmEsNJDZA7VBfAbs+n25nnwNuZgUNdXabv2m
7s9rqjfu4ClSTNNWAVz+/smCPrzFTeBrVkpzWHg+N7HdMuQSCfo7cx/vH57OPFHWb8dWC7xAxuNm
UeEtSUMZAbWhdVr5tSN63giGYXhH0v6WASZ8RvRHHAMk3qlBJWmy73VMuy5I21KX01NHRkSWnpZu
Z3hZFW8F08QV/CP93UUjdWr4x1QqQFJy7DaOFcKdwsYxZjGVjD0OF2atcijoQArT7LYNbu78oldG
j2z0ypmmgWNJq0i+YWOazJIHzyn8CWeqxV/YeaDTL6LEiQ+/lH75f9JRZrtTvn2+9iSWW5sC1SO8
VBfVjj75d8grbSRRWO9k8STK7qv24p1eydV6etz4aTw0eX2OGZRiw6pkr/WfvpCt7dHl71XRHiFJ
pVhm3FaWsWAUhnEcRSmnKBF2OYQc4RWz4rAI637ukxETQEenq5cpA5sjyaShHR99oPRbSc/2n35V
Ybq32ScB2fPyHCJIJ15pSsM6n4kKpvrLSsjRXl/7rWlAawKnFZXpeBq2w6myY8gF58vBapd/sZIL
cuiNjI8NQrqKDsXddtbTm9VsgdZlqr9jiUgCVpeLVYDk/jNIuOgUndWNzcSxsCmppi5MAOq50vIs
/+oLdsuRYS1SqPKxLg9UNLWvKleegAzPfOlmWn6iwqR+8weTGQajJ8+kxKcMP/xQKV0UJ/YbN/wC
/e4AY84U9iQHGqhFKtkhJVYAtbj5HZZx5vAdGI8EPfJ1GAQdi2rNVfK1tjHfz71Nn7RVaiSJ5LT1
65xZFE9m4JCr2+B3wnX1pgFatI2UGRUotW0x735WlfurVs4CYPhd7auxMULvO9tevBdh+aQwaGR7
dyZ0qdtR9TObq+DuDsJBqtQ1s+MIjk6oi+NQqqpxRmd1NRs96+XXH3c85saQ9ox3v2kEoqVVk+tX
Czpp+FDckeOoOV9WlKqMFXmPBcve3wkX8RQxFTxCKAG57aaZNGgtvmF96GbPbrv8FOPjH+vq8v2y
2WZScIhyFa/kRWtyWuPASsFvBmYblYnXJWXAsb+AB2VOHuW4o4g4EnWtUxqdCiwQ/UIRItNEi1C7
cZZBJBDVgJgXTxAsdCAuonUFkSQ6Tm7gdcT9aCyG3an+PhhU2ET06KCPUUbyTl5G3usC5N8coMwg
k7X0OIGvJ5jh9ebJ9Jb0QXYZog4Xvtw0PmUL4kfUU2dni6urfW5Xpb/vsPcZTRUpuLFDGeiQnmQT
Yd7GCnvCVB+LKs074T3RhXpF+Dm7D78OnYsIXpNuXiWSpf5PcfN6COeyqPwJv0Zp/0u/pOPXrhBF
64CpFY8a8GvmAZIow9/CODT4qfhA5sYZRPdRMTATCZQsctqJQY77tXgoTFIxJBUOOlPP4zbZIwN6
LqMZrgaA200EehAGGqLXUol/4iLzttHMQ2iDp8hSc/Fiuap3Tr9IdlnVkMYKWmNOuBIloqOcv/DY
qyCAdjhrasditSA1Ar/0vfkjAHLewwGcNmr/kfAkzx8d59QqLvF6ItLuujA3KucBAao8SQsJB/1D
4ZterjpCEbZJh0uBJJu92YyrYCqysSU6pNcqgQnB1yBWCcFjgqZYx+SH/PLqjIy6K9vIh2He1jj/
z2Kr3e2rBsnJ2k8yfSHv+sD0ycg4PS+p+1XH7tk8D+PglHobMOsOJxoZR44oCICpAS8Rux7uLXzt
TTG+hIg0ym500uzyB1zIvbB848qOfJTUkExp8uCeGoGD/NPwZgHIPLKUW9/p5LesUnqCojjVh18o
t45NPqXZglWrZ+PB7B4IjNi1Eo7SEGmZUDq4p2qDm01Bhf0WUyMB3eDe2fxig1ALTnCaqYiNQTrX
NpN6rXB08nr3WcyZHnT9guYMBlT+++eBFxAeSKWotm/xL8AKF3QxMXGBc8QN8T6e5NYsVrY3zvie
Y2SJ0vPruWW6jbUTqEy0S8h9MaeXNpaTfQQ+F7jEwqrjH41H46hVTvIP58nxB/DdJCr5lcwiBQsF
g7/LtHhUJfL26+VymZsRih6wDJ/96oTPw4tsQBobRoPMLDjlIgpWrBPrpk3E6u1H7cyVWmQIv5wP
oF37rhFNhwXsaR/6mxrCSvCeNdCn18qHDP8q1qFybvfT4F8UI0LXHjw0ZFoW4oGpAv2UXBmMOU0U
UCc4W4LnoprZHdfVekKeaGVpLLCvNjkxd8EUpwprzxFyddNCHtEk557jipIbWvaRKHeC4H+F33pF
hwuyf4b7J2cQEIy8whBdlLhlbaEwI0134L5zkH+l+fRO91KXqM7cyEjUf0mPn19v+L6yOekm7go5
vL2SqNPd87V2jIT9gS5savqkxGMjG4oslUtnp3hZQRswDBbbDUITKHbp4za5iSVZ7IQTWiWblGKj
DNedUlUy+fWbePnCfRXzZplcvwT/PoUVmbxdwaxKIPNl50C8vZ11iXz9VwAi4z/b84wPE7RvBc2l
kZumgQQ0UZnaW+3NKM3SsfMAJfPPZLO3eb7gqEnwFSSzfM9S5g37+VUMbnv8PxMUs9WVA19dFLng
2EyIeciGsmeQdZA51YURWBVnvjycMLB3NO1rVOKxi0itmegF4yRtCFmgoBBK2uEMpssmiDUOyFvT
O9mZ1PjAgUoO0JrMhEKoqz5CGFULKKqrBcha6mHBWV1LSGt0odGQm5uNg+H0cnEuwJyS7cfNtkKH
eRu4p2s5bAj8O5KEJzfkKkiwHrh8ppx+yKd6MaZL0km0d5OCR2B/1sE5kDqR276G/tL49NN27gGY
v6wtNHQptHJ/syu0F2+7426rgP12zxQ1vnUTvKC/dOuNJdVQE0I3400dOlxlcxdMsVCjer5o/Yf7
l7XDzMWgSKoKzXDrh8GWnu/FfP1OeAe6Jh4q1bLFEytftx/fu4jsP2tofR36WX16WJpLSrRrIMwG
XHj/EAFVWEvqW9HQKZNz+ikWm9qV75L5NQfPT049kg8ao6k/Jclpe+ouVI+PLk63Cw8i/5iZsHlK
k1u6SlEaM7XRSl+Of270SJch3dpIfZ2XAJPp7VuHyuPd5643iW8hsGAFvAtu44QZgrH8vsC+ufjm
0uWeDWUNaZ2azL7wNmHFnS58ANz+PJ6zogepOAaxg80rv2dYr0I3WRqURrtY+d2w9uRSQfaB7QuD
eNBt8pwy4prSkM+rxLp0yPS6vNZsFP2fT5Bgs2FRxD9PgC2s2J8bgEXjfrGpjOG2ucX6PmEC4xtw
4qA/9MDmn1PmdziK9hrCO4S2zGYwcncmagVrqOGWBftf+e2SiIqRIh97v6JUf7wF6NLMDG0S/cnD
VCV2D8TeUcOuBI2w9Xr4W4ECaygK/MO3Ot5DRhVaHQ2/9iLE2qyqCd7EfDaKtdBaSU247sZlRXE9
rHK9MMdYC9K8JA3mKxwkdLSdLt6CpxdOVjV1obzu9hoEEBZ7aVQFms7rCU0tzKt8HEiELMR8UVXH
V2Qn/mHrvhbDpKuQpLYzVfMnDZTrvVrBFgh9rgBl9Hqq1fLeMcEluUj1ewnjbNABTkC50ivBvGHt
eTqSScy1UJEGLfvTWIl9mK0mlCBOFP1dGy5Pbr4A/2znfrqbVmowiUWsiIz60OvIHNa/4rjY1mHl
U3LN2f1MOaXbhejEw2294N50TYVy6I5yKm0OBFDDdtGO9g/gE3gUwe6nyLyX72klz7ocFzncaaXD
v16zq3Hr35SdN3KfUVccNIdpMA8uu9s3aotUkaogZO+eRp5EKpa6mTnubzlX3pVLaTNLg5ozsl0x
af6A40ok26i3XF4Jsv3eGw230y+iiAdkf6LEXinf5ANI0JKyniX67f3pR246ALZA3cCIg8wgKwGk
uZClhyvalWezlOf/86a6j6jl2MZ/egH98Jzn429C148Rus7/nQGG7pWONaLPFxGKQMGt5NV9tTsh
eWJJ1VCc4mdVyk6slfY9s5ScgV6qODKPnwdNAvJNILu0BcQyOpQ8HWJvNG6PyTCfPoS4ApX4om52
QapNhW8JzSO+/O0keCxkbP1Bf5fxr1E7ONeCq/EP+YD6ibob2L1aO6biZx0ZepDmyYrtsdHc5Lmc
IlCeN1qjT3A19VmLqfKZ7kPwwgwu/+j5yMi7tF045Y8YLGMQXiGbjDJ8VtfZKLLfFCyDBtsmLXkN
heUhCAoH6ePqLTeF93VPqYUKhRFbgiUhp1QDK53hv8zCHNspXCHGWJmHdGEppdU+BCdOZAd257ZF
Grycc6bjj1CkVh8CxIJpQeYynk2kEi6f+QwWdi0nhV6eX8R/YcZ4/AdHq8wQx9d6UwahLX64aEZJ
LJCxoeOmIbEf4yBGrf6sIWXYdlbIPakfbuEXMThr4b20WVvFqdlHkqJ3hK+Nv1iOLpMXHokyWUue
iCkB0z6di/ubWh66htV/YQaNJHNZVgjar4UuPfb0Vg1gLbbinugyTH909EXJVC7RGU0lDbBmxkaB
ovm6/tlWTpPW700g7PIqU08ha4ViAYlkLtvAds12uYwJRrrZFxbqmhSmJCGOm9yBg6Kbfh4D43+W
eZ/6PM0xqWjLzLQVbd69yGAzTmnXeMBhvgSj0pAKJsZ3a3AL8v4f5vTPLvzWRDcqnNKng+Sw2N8g
DV4yb1h1eSMXyAiEc5F4ki59srZhvf3fqIhn/danUvGy+1yDQB1ON5Rw8UEHZEyuvUjpElkdMxLi
IDqG5/NttJGcDG5f7137o/1Tv8e6dQv6hrhR6J/zZnoNUkTf18pxZ7CPD9vx5aTSCDDePNVUYx2e
WeUZvbRYPVbamFml+MQeC0DFBqGBr2MUZXpGEs4lfVFEQbFOFOp2yLuQvoxwDB/rZiwXAoMJAL8g
hpbGagNZ12qw8mMLUZwv2qoRXz3g1doKZYGjTxmAU6OlryVi0vDf+T64Sma7eVJo4+wYeF2btbS2
4i+CCdVCSvTz41vKSbPnt07l+WrYhGgfgDrIuFj8ToJXo9uhE0x68ec89YWCQmVVTelKkAygZceZ
ZnSmjqQrM50xdpklx/eUgihvEVMuU4Dw7XlQ/mu/gzoH1M2oxYb8GlqlRJ1obU6bym3Hh/SYEL/w
OHa1du7ca65gqmx9ZXRVz8jwPio8o9IoB+5WBmyLOqcRr9doSpcMbCvwYEHmSgaBkGtt+UYbmmX2
vh+O6q+i21mKzgbZJrxGtSNy4YgYZm1mC2d3Cc/2bCFi1y0N4/wxINBYC3tb6rRaedrdCPKTPP7i
Ghvju5UpDLrZrPCRDp5MXYBv/01FqQawfO/olR9G3691veBgTLDEr7iwcwt2mKB9AGNiXkde1nZI
g1USJ4TAebJiWEgKDDBEfhjauqNZTtQRRcRd0tWbYno9TLNd+dHYdPclw3chFkMvNE9ea8wKhXMv
uFv6pBIf1tGMuGMF1VOOul8PpltSG+jNe78fRBAtCtlJ6WHsG3SQeTmPnX6aS03yn//vcdbiMUgS
v+MtuMXLJpZ0+BqiED9r0cDXv2MrDhtYfeubYbm2BGMTThg6ATyGL2yS1lEDz3AecZ3ZjDmUiEJV
xVTxRsO2ewXmbtP9kUex00MN9ZYQo3D2OQeeB2vtKaMlIS96gptRcKW/Dbg7e6tH/oy6S4cP3OaL
HKw8wjNiLCB70Ffj8t0r1RJAKEVOiLl1QxLxBX14G73I8+tfShbLaHdVapDO5DkGFkZcHx7HOBhi
qQjYAZbDbPsElmkGw4P+9wTNtZThq3ANkVIucOmhW+uQASi4b1Gez30NoD6w6cdedbCAOZgD5vP/
ZSIl8iro5vi8vCHgnCKa53nUUibM1kWGxbofhm3Ydt9M2HPYzt9h9Er43ipmxhSJTCGyP4Gf+0fy
2Hg8TsBwsicTVXq2rDPpNU3WVtM1Vzx7hkpZ+XuiI9dJPMggWw78Axqrpt1heJud004KIBKPuf81
PoVhnG+s5vgMkj5IzHIKgiD95Boya1IzcuQ/X9NvWXqsQWG2tcV2r/GjqyHcJNy03XNVpsHFKoDg
9/JCyDPZHp/I1sMQ30fjoy1FAaC5K/szc8pstkjJuBtPG+Kt3E588cKs96l2fyc3y5fH7JuFp5VX
jJRQqe64wTkhgVLMf/k79Eog51CP7J+q8vr6QYlrXusRR0/+FLA0p3jjDol7fu6qQ0UQUCl9fZhl
qsMakHZOoO/lJlX89C4b1TCTmJYI21Ka2xB7VwZpvlN/Q44QVQOoI6IAF1+3CsmZxfEF2lVb7XbA
X0P43IBlcCqk4vbsd9Do+tKKXc0wJc1EKK/0qyovaELFgVSOCYq9xPGBewkrURg/gq7yNQ9kZebT
1ZiLTHUsjC91X2ySOWfyWK56KuV9dROWJeqSqi7czCGfbGVb570ekpaLQ3Kfx5eN9j/Ib+ZQ8Ncn
lqH+s8HKo9wK6yh13uM6F8weF5GjceUy07L6ao4A/dgnMj7VzK2o/iw1pNLGbXSiK8J0UXah+zl9
ICwZuvhwEa4ax9BQG8eE8Qr/5kNOacLKl9W2R9w4Hzd/SE5z0Sdy0DWxfdSs3HUgCnqCagDkynqU
YpQ0Kdw+kQ+GM2Y5DBeZIjPG6utQooQIKgb8qyuL2HxiZlmYfKFZP4pwjnk2sFqOO0MI/WpVIkFU
zUZiJh9N7lgSYFdyc61nX7x9sFYu1UN2q5UtXh8qgg5adPXsohYugBDX04kg0SybkMfock+3u5d9
DTedy7GvPr/eESgfLhYhMjJk/UcAn5w4HGdlZ/JOogL65a0K7Qkji3QK/HiAumOOop0fYx3lGoaB
wxHfHgH+MWPDzqTnNFHAZsdjFG5SP+NTdPdzQ6Xfg/2xyyn7eAWY1fk011qGX/2kujaz5p02uQUp
s9gmwshYYUufw5s6C50vxwtiZn7PREh8tzrtqpQzTe7P1Pc6gZd+UyKck1s1J+ePeMT5YhzjYvOX
YplAau9SAq0Brgbd5qAhlKGj1vbFU1zv/ysTwrGxaV76bEn4wzGPcKu/uLZO/s8LAVxvFFjoFNO3
K+y6KtE2/KyNydMqmVZ0t57CCYbfe1qQd3XAB0MDJVj2kpMv4Ze34lK+c4YEXk8LU7C8QWFzNKiX
DbihpkE/u7Mqq0TzNDbSCyVhqdNQ6RArdEqRBEYrcn7nrHN3Cl1SCd94kZtD7k/OFylMAdrcFI9o
4oqc7+e+az/DQLwvo+gYOuVIs7oewXOyc6ojcOf71xpATMulgxEtoSwbLY4kc7ftfx8TSLhTHRfY
QRJHevKt+bcH0jh1Wod0X1uOgUSo9OFEItjZDdAtJxftRL6/cC4nXRyj5DJJ0/ncv4XUX/ml05tX
2IsUqf7AHg2C5kGsWazXK5HWrysp1JRMWDWiOy3D1opl/HpO3ftvGJ4Nu66MFamD+9tm+0CyfRp0
BPmOSlEIgLaxMuGRsWwF22709yq71ur09xaXQRWBwib3Wa4ACFwcLP/0cXfzuadksnZw2ftLDZEj
MI4glQX/z7BCjyNV+ROs5bpAELNK1jiNOUEIeFJ4ItVSbgPo8D7W7VzVp+tHD/nVT0lVop78lEM5
P+Zs8zHrrD+vPiFc/ZhCMlH/2KJ6UfIsyZ5cuLM95i3P1Gf2xxssQCDiGb2Fh2xLHNZs25zFM7d9
/UUY6/gyEiV6J0Nzo0NRKCqlIO3bQJt3LJ3jMBaQkWGcBH3kdLFdhPx75APUPiG9l95wppJBXpzx
8hlpqB+s6/sQtwrJsHOirvfuTH8AOjpDEPs0cC5ibGPFTK9z9jNAHNRE09vl+alJ2B9rf3NOyEvH
iuHleWCAZ17h+vDSMntQgJOKw9b8+cvKriTbIHVtrivyrMbxkSqdiDWchZMKlKEP80hF7BbKjMqm
w9ZDn+DXsbx2bypj4UQzQSx0xov0vAityhCI8w2bSvMtJD/clWr+czwG84O6Dzb+fFLoV1mYNRD9
tNdsQOuurMMnb104mvs2tfQGBAMlC6FUxrMYOdbgQnqdg4AgmBHs51Rr7+zmo5MNtqMBuEdya61q
FdSaw6nziCuuSK33V01XHEkDHvxGPiaH4mF4PbMDb4+sB0H/3D/88b2QdAaF93AD0DbdkGNRXhIb
id1eNiJRK+n6BSlqGAU5EcLTydDHskcS2icdxAW3SAjCGx15MHpGfvwJKHVLVU2JcWLQ4/ZXFIO6
k9or3uSzZdouNbi8MBd+VQRRjjO8lXH2NxwUN0hGAWMGBdQpt0klqVP8Mfa0vr8km0XHcq/c2Xf2
tzhNrN2m+vaDBYWTaNiU5jtxp3yMdT0TsmLWBzhWNYIA6Uc0q8ArMZUOLC029KADY2P7ymxxhPTL
xa21DEbr4XOecBgQMHGh+ztzt+CayJaBIFbznaZmtkUqxdYb24WwwXDUFNlt7BC8kTStJbOzzbE7
iBPbEE6WmnitzPd+HtZ7imt4c70J2DVSDGvaeeQU70GtQ9jjxjonPCxf9za+c/rUkPPTFTbUWLuZ
Qw4J79NKhdjwnGtEk7FDJp/lDfNbRtRO44K8SR+mcn78o2h1eeykx18wHXJxIYYLC77Urhw34uNr
6NgmoMzwPoEl8iRMY8E1IKmTFFRA/Bjq5BIZQBYxxX2Q/uRHMfVT1kDwYmUYJQSdvM+g1FZia5z+
P0MILQxXrhAnQROUeU/uGQwkq0xUie+vHU6A9kbt6pNtCSYK3Yf7Zo3hBuUQo2/0HkqrbcapgG6C
ZmsNX4w+yBggKruAjXJYvqQqSkk5C1SKmxV6rkAFHGo8uR9HX4Zo7JKYjiihgjjo62V594aP1GAZ
fiMzakjUee0a1jY/flxRQbucbh2KYHdWtoBHUT0+PS+RJv5lXPC9ppH2eGzISjArnDFpsX24VHcr
SN25Y8rJsYIuroTo86is8zU8peBNWskbtEehAHMQNjM+Ly2PrisgA1tqoLnNDGchyCiyyAvTKTgX
9Z23Gz0wHUFeq8XvWoZIei9rN2cvnjxX9s9hSlT0bY+oq+eGzDYXdP9N7sGeHJg/U9HfsvhA08gz
jFZb0dIq6did/tPL/doLb+i3Y2kzGfBsT8duolXxXaBV8ScGAvGY6l7kFvz23FGk1DBNNtQasMGB
9/2lMxb3XgtwZl0dJfYvtK3O8aJAd4vffWxDmlPY4vgazFJzHMouopFzu9kNRqoMoialIOfwUFCR
2ajC3dSJZ1zrZoNFhW9dhQfgxw38+Bkh0uRDb8MAdRvCV+JIV2+A9x56R06hLRtasBEnwi15mulF
7oD4aSweNrKCb6JUUS2BrtLeMLSYNnJmZc3hNiYI0ShjR+6e+6imOyLyt/O4CYZth09lmM+LXkBq
zczoDEbOFCyvYhkH2GtGWaEK7knD3CCvklfmWBLUOh7Ze37GhubDUCZRpqkebN4sRNLILL3SM/Z9
sZZZtKYqXiDHshH5jNDf02Sw3kGPo8fYdOq0FiOuIaMdC2kKrXnrRW7jzAVCB48L+z+wjw1P+Svs
LsHzBYNB1E9O0e7qH94WmaHiCSkVrlROy3iXDLYO+H4RM5MRzUYoA9CbIb8YxlQHmI6LC2Jc9BBq
eO09NMH9zTIisydybuPml9ZOO1GqujRfEwaWNQmqY9ssmcbN4igQSpnKEMfUf97rLoj574EJCKNK
MS4mSGOix9sX0lI0HYhuDCWX9esnhUWP7vDyUjVO8XMjbMIvO51QKDr4YtdJtMpQpMN1t60/pDoV
XRQRfhsrP1l/bfcU9tC7W70ukUTEs5Smk4AmLMEs4ccXGr3qIIfZfazf/SFZiBPilcWBVgB1nKLC
1Oh+h3wakM8knkGbmB5iN/Stu/THykmbYcQpEHK+t6DbS8pAdEHPwz+RZ5dD67tJjYRPfKoWSdi+
QooNWLkwdSHgWsk3+ni0nMMEdrDExrbFATvQU1moyylZwtpyNMo4Y8i2kMWRHRtVtw3FjS+0Cf4z
9veAodZBRVca1PJxExSsKXO0iz/5xKaT6GgXMvePmqQJVkD3OCgRqR8czwOp9rpXYsK4DmB7G/cM
jBlyNeGDQ08UGtkA3iOGkWywor8hfVBQ90X371UOg9ubHrmm0AtxjRQb5oo0rcQPKJBt8WxOQEvS
gmXT/ws40HTHJf6Aa4w9HB+lXJq+VPBwbShnKLFUabM31Btm15cuKVcMc1qbNT1j62Qn+8cB7tH+
t9EkJ2/o4fsW53iKNS4aMhY65UiyGn2vUfw2wb4WErTBt8zBROE/Msodcx19xAV7dTZiw7XcwuvP
CiJ2viFjp28dz60/s31G5idnIQ1NDp4DLxZGtxuEL8OaaSmhcW/T8ybEirLVihfxs5oESuN2sLSF
aGRrC9DHL3u7Dis9v6bwXTKC0uftBzob+YlreleKHaE1IJHRqazoHTN1I3+TN+w7ainKOE+Jkoob
d1567uC9u2RHIQ9jmcnxIf4S8ZmBJZcPPQ4vikRhn8bXoaUpsceeLjDbZxi3gYI7DPVzANkqBf4h
38S9V7HM5VEkeqa5aRDGRwEdeMlBbQkxg+k0mc/dSYRz2TRi3iB/BA0jamX+IANk2JkfnRZu1i0o
ejTzK04c1mBwl/6qoeG2/BGiZZOl96q4IQVsjPqpKaaMDrUZYB7bWzpnvOax/GmWeNyWOpi4eL9V
3UvMevWbGZNpSUNnDL+1E9bMsqWKwlpuW3/2+ZJMq6CHTcGmmolxqE+yjyqRv5rLyKyyNHtXXSJK
7TfBlI3kAVVp9j5pukq6LJgTFcUwJkrzbVFaRy0P+Kw9V85zpQjmjiAxoePXNPVE4+i26yNtQCF/
0F4wKpJCyZyVa5UgasyEOc1AYbGr3It8VmkwqE+cbksh+GNOj3Qlaox72dYBDxrNFxh4eDOsx9g7
Ve4YoPZROCQTRLYU6+MfZ8Sh1ifN9AQ9W0nZmPx3OrX3RThMXDWKuiTDbj77PMZIiqd+FtJPS7Uh
NMi+F0kBBaz0Tu5aTSTFNugcxgCLaPbIsoR13TgvibrnGg284RwWxPBW9ZVs2fqwidW/DzGXVbyQ
gHbaQNLLqwzhy/4IawY6Iq6aR26x/eJ8CeuDLTXw5ily4DOAr/a6jAybBdU0D7nuUqhk6D1WX/wU
TWUNe2VIWTyqkxaaABBEwHLUWiytyPNGKF7gWR0Cc/N8eB4JqdjS4wndqCLK90U9w6htRNkrJ+JL
iwsrBsnyDXWoW8eE3W+A+Xcb0JBliK7+jjI81lMtm6XbW2OZJLcCP7vbrNH9D4OLSl2YY5dlzYlk
GW1H56UBDa5UQ/ltwAODeXLByuWleorUEAls9/yZLiU/rVayXb4pK/0uPSmX3nMvUes10Mqs8Un4
Qi9A3XYBPAzONfPcq1FlShFzMvHLwsXy3cliNIs7ZwiaP3HSQC28crBYxz5OfY+P0quyVN5RBSez
9N6OLmDjkI5Nvzyx98TmQygQOi70ay+bBIFWdo62TtlibGMJc1jyGDfY4e9AMsidDx1KMfPaz9rk
3KqCFVWbyt3DS1hkqVtUlr6KKk44bblXiTB/AAi6CakXM60YimFYaJUpnALj7ifYsM/ihTe802AW
rJfYW9d7Ll0uck3SkJg26ljjNa4TTe5wHKhWgLPuOBOX7TVHO7O1eB5Pz1epL8icXte3esUdgbR6
/B8t9dSnD+JsCYwxLWD/vgbQXIdnbnk3Tal0n7h/IFRvMyUwWIVsx7uAFcYmcHHoJslp1wBeslHd
rgr8/oeBjGNxykSJOSfR//Oxny0xDfykgIPHbCVkbSqDzHhvUiKwg5Fk3/trHHruXS2vIKPDOX5i
PzfDCzEORdGGAd8fjb2Y5ZpIoFCkFnJA1WV29SWQK86Clggo3zZkDiqM1WLlcEhLg+ZP81cJ3tci
7OHMlZuQ/6x5Z1JDbhp/giimGJ3I4Noo4AV/sTHYPQaPCQYFUvtLuhRDCtrObmo8yAVM8Um3ez+5
bbU/G6ARW+68F9vn53O0EW+V/8K+qOvF9MhgVnth180LlcN6bOakVWv1wTTgPbVmfjYxO+J7xg4o
c/aZu6d6DFeoPa4MoX3/GgLJY0WyAkeb4p/oLiIe2LcFBwgUU1Q+IJllkNkeB5CZaapapXTTlud5
+28AxrGfl8ItR3FreHWmAf5qJWMwG3+4CU3rpp3lWo4K28vSfXSkGp9FR8jZvCmfVgQIBVprwEOk
ZKG/0Nfgc/Tk8oxzo2NoWt20ajBdlFIVclGSlLyX9g+xJkpDQIKebol7By9VKk2PiB41Wg35fL1D
2cRaafcpS0wfMtlkfwQ+zzIBzDzRQQXQnS06VtTU5pkTOCyJB+hpXfl4T/9Zd8B50LGEgwjzzcM8
kLV1aOMWa104dUSt44paKesd4dO4dIRDKbl68GmjsQyxsTQm0/6UK6K/IjbYiQ05anQUcxF+CEyo
BCNfaIQjNc80pGa7TlqTq58MDHZ33bjYOoFaR8WmHCz/9z5rq/bGhKHoBFfmEM8cQN2KrYj040I7
XJiIcZnYm2hieIs7BvSN6ImfmHYTJCdCSJmUTHhAMy6+u2SfbqF2aV6dFi/Dta0ohroHlzeYvZkG
MTCNYic2zrTAgPCy6vxHJbRnG7PS2Nj14caryW4UqzJrlNwH448WMRybneUu3JZazVt8VxHN3uKa
Yqju1MfgkMrtN1p1T03JZ+7egFTmfkYeZFlYfquBT9BkQziYKm6I7o0wn5sfWCmzEv/dmNEYdbsN
qMsWunPsJ+VKBTB5m/OjDd3s0pM1ermOLD++pFxH8vwed7IhIU0RbAolH0yigo3dgD5caKBNmoPf
eOFaGJvROfzpnRWLvjplRkeLwAAvvvwccRewBJi3wm9+vKV73fiy7qr/c+IsqcGVZBH1woHc/95n
2kSnhgBuHvvJSX6qY4zWIUH8Jz2oRTE/gYRiZhm3o3JGivzDOtZMdk17j6v3NSFmhJCrppol2Tqo
fVkzTf1sJb+jYBH1FkkAd7yu+1w3mpET4V6Mc59JxXrQgAaAKr5zWB+GJq7HgfTQRXrFj3nFuSFw
MXn2O/KKq6mlJRWuaS1sPs2UKgPEewoF0EhfarasXQLutGCBpWmLu9MZ6QTG45Kklg5JK/eOhuwZ
eJGzblgnYE5ZZOP4koWGdVn6YBIAwx8ge5DDBmnGv6PDzz5KzFpyAzcjZZf72TaK/AumxkX09pC5
xu78PSIkKFOo5YC9drAwr39b7UES6D9vXUKmPasFSCK1hmszYwvYRfXLEZ+L1Ck/NLyFap84ZAfW
p6JjmY4TrQZuQwKt6F57/tZptG/c5DHTkKIzhBs2zIcbBjhtiRoJPu32TP35L/i0295SCnRFEcox
sfHff3x4Bz95TowNLaKo/HdSfzCZ++6xACP3Ozkp7D2C37O7jmrDsF/DdCKYdtGYGE0qKxlMiLjr
7qNTXTRafR0b/OjbeoO2+SiytI4ZPOru0j/hCimRma2ME29tcWV+MmUaITUMknz2mJHxzf2MOaNM
ulmoUm4f+EB6eWU8TXoUWdK2+/KypOeuB3GPwB2Jdzkrk4kaB+6eaLeeZi4qGcfqd6inTJzPKVnq
mCxnC350QdHDIxCVARBU+Oxi524qnALXpNXQLvb1qDeK18dHrWhvMqx0BYUQCgBrX+2PbjrN1Ix0
KXGIDHhG9za/zfU7/ENJs7+tY9j4l+NJNfluJQwhQZFAsTAPUjtVr8G+52cHrQJccgcLQsuCuHMl
I3fzmWzVrIV1Dn8iebI/3oQMVobpeCutT1uecxW+JmHwkIOON6hANb6Wi5bu+QQZVdrTOdvvlazB
pb0X6zpA9TP5FrHZ69DLEszUjfy+IM65wAFSbyug9uva9kt0XRZJU578LJsMPHGW7IEFpKCQ3Kpw
7e3EuADA15TtQV7dvXmO2CjJ1HIJRDpipNPV5QDTXLaoeg3mh6K+ALsbA+yD5XRyvaEmqjihn5tj
KzPWv2K4As+3y2CKi1tmVjfn7HBWHnqus6fkf22LOwUTcP0hbsCV1VNdaSW60Q0JZgl3UQ4p0OTO
uW/9dTynq8agXw1ygNRk+huugb0BkJqCKR8cfbSSfDswf5kmToiV/20GnfDMvWBQEpzrbrOfuBF1
aYzJrXVedZPPL8LbTc/U1O3gStaTRGWWsvojxKHYaoiTNB+oER9GP9R4gSkFw+k0dxSIsVmeq3y/
PW2+u46NscOgsXY4fdfFy/tZz3ysbrU+ntHezD78lMBNEzCMzp6WO3QOlaLCiZq5kBiUC4UL2FgX
rrlAvejKCG8thJjnAJr1mobIze6nGTVO6+jlb+tlwWNKyN7RUSFx2oYGeNWUCCq/hgHlIDaQVSnb
Sku4J0UiF6pDV5uektU+D+zdKssIdtGEBF1TCSIDD1eFaXrD4KwJoithQ8EwdEmq8kQ+DTRrcxfF
w7+hYk5HBeDa+l2tXryegygh64vUdAzP8lDWdP7aQGAnAW64uPtsV1CH4SlB5NMS6elxI1OCxRzF
MdjcetI18U8mCgoJlQMfXoJzBVKkDy5aFagli4CE7ewYr6OXDRxt6inBXjxAo2MPbZGHSTjH+QU4
0kGR2E1NZGcYW5g//vkv1t2Orvz5AZZJmrHdj+hS+q+Eige87T6HFU6LzdDkowg59qhFpXPul0iK
ap7mqyma0JMb3X+L68NRoOQGZW5/mnmifLUuB9z/9MnoyuXDhSFDrcc3uj625JdyZTmyHQ82zZ00
Q5Mw5JItL8q81K2JE/lAg6lQz/sbWPv66birG6ds42hcC3NPcMJooyHYVd3yW9pAXPDZBxnl1qTs
KtFbvsHaJj9JW5lVGRIRiR2yZhbhPyfZfUyKxNkqMh2GED/Mnd8kSEjOr1eX8sjfxRACGIeny6Hd
70xF2CCiI9pLwd7HitxUhpu9BgwNn0PRanxMeYDJGmUxyDWvpuT1BGUd7aDVD+1pIMCp5IJtY3VA
TCOYCz/MN0fZ+plWW7Yb8T6Q2brf+T65LGXiFLB8YstCskQpum2Ntv/i5Ix2rbMhg6ocnQ4fIQQw
LXYAfyP7XBedvuizLOb00b2Gkr089OrTML3uDJzCr6JJ30Q8hd2NWx4V9YEDRhGFuYOB266ntHuj
yZPc7Bev80tlIMDj5g7ugFXEZHj4mB6t6C0XM4FgiY2z6Keo8sNSXxQWp+UlSii20sxqLlR93q6S
BDyl/REwiq6rOW5tVd4uEzPUfRriPsnFsAvkPdMqN6Ui6VEuOkW/iKMV8ZKo3HEWtLvqR4zgEBsl
2qaawi9SYp1P+CD+wTwk15Gm8GJKlDSeCQ2rxgmgCNX9mwrRW6I734ps8CrsOOFLo3gWOuZLFNsM
VnLVrYF5CN/hB2S7xNucstTRaV08j1aNTXU1EVwz8ISj+OQIhZDE+0E+qr/AGXGL3CbZXA2m/WkW
Akzg9/hE3po9d+hL+9/TUfK+CEWUsBsyssbj8YCkvc0+SguOU67hiqIH2qD+nQbBIAB1ob9TXtG2
AVg7KR0QC5Gn+MkQGbd3qt8x2/Bv70s31RBkPm9l31dfjhu/fGAQOy1QNoDI5OD2OnraSYYroz2S
PgIqY6+UT6ocYuezDsjZixYNlY1Qbyxvmuf/aUk5F4mq/Ip6Fx6sLiTggyJ+ZIKf0aeezC39B8Cx
kz4Pa4bGzl3lztRBY4BE5tgtKl75Wf1ypOw2IV4GjzuwNT110pCUmCCz96gyD5TVEc6CqnDuEfXh
C1avY8S/dTHnMhBuglakxo9x4CiHSxtfRcrkx+dyCRIa83MS8uYco27qbcf9/S0d3y5TGYQDJ2M6
QQ+1h36nRIWUyQV/uRlsRv49ssJCJSkjGAR9aAI06KYEKpDWkVdQkGrHlm/1ByW4NOFLiJ+q4Eci
9ErVDMNlH/s05ZxfT2V/xEWkRXlpggG1FDBahhS3kov/JMS51tLeqUMm9QtDneDPAm0h6t7wOjrn
IJRDDKVIWZY0z9Gc6nab2HyRirkd8dZqhsDMLhX1ieriAODCC42s8/Klrsr4Yz7Pk9BfJH5okXvO
yTcfJU+x8gPLWWPP/ZACAELSkGuhgmPcHCD90dTUI61Ff4EJgMRxsksPsb5uZabFnNixGmUBHXZn
5R2TUvv2DAhnooVxcAC6ybh0hDNZLyjTHVCT9ktJmRwMBYPGGSyC8gOxMXBU6forVYWbL1/Yd599
Gw0RufINKd/IjkU65xZk2Xs7nw50EzGRgkQ6guzsIuegZXrbn2xwJb2JYu71wVMPmDurBnDckvji
fxO4i7RpYUZHAc4sU3ZRZZh6KWzPS7z7pqrMuakUgRhwC1gucsp4+TMK7zWbmZWObOjUUYN/FlzQ
lwy+PeptjNZGF8KmKLvyof6cuAe/7MmhqqbtTzRP2VRXsUGaLTk/JvihG55lHF+kJQakbut/c7fh
2k3lbTcQVP0K9JuKMhoNGpPC7ax4GaG/VzxgaomQ8LS050M3rMN+WEHSBjIyLMbVhbnYfqP6+tiJ
+ot9yOxlYfnTLstxNZZBZxebJee9R+MPxsbqhYDwO8SZ2YENVMukfKiaQn5dUUc8K2pS3Bx6DQtb
za7W1FX2eZiia2dGZE+GkVAXN/8yMjQRBv03QcIaTUIYDyjOiuBpNR/spOwup7r8WbyIfjx5DtHE
e3r/K/kBo3Mes8J8VTfoj+Qnf8YP5yrg9nsA8RyUEdrJw0SqPNnvV6oCBmwTsZu3hjUpjVHiiuOG
jFoqeySxcmy5Tf9zeUk4MBH2NGaHgXYIirTMiaV8CZoUyu0vtE6Asmwtw4py11Q+tj8QBgcHPUb+
hAMj4w4UYz133JEAKnmWjKTmhnL//SF6wemElmzApNnnBpmVLJxEO2VUAXK0g6L7MgisLeB1wh52
eCFmnRe36EKTI8KDIAUpSifMY73AZU26lQ/TKLMV51IPAmD4/xFZwsdxJbST3Nm+DgzFMz4TCTLN
/6hEG8YHelkhPSjunoddkspnlfzYWq8N180C0fIr7LK1CwnEFpK/SydG1ylJvDPiVk3DMflI9B87
LB5N+GEQndPoXZyM1cmI3Jtw/UFqPGzUifdgzQZ91xeHY/ncinc1f//Y6Yu7L1BEml2lLXqyygY9
SqzaVlilpiCOJFvmEMyyZlUOAiGGsxPowWtlCQa9c44i+9gropCOeRxt4yx7uxo+LT866tk0MyD1
UICs6g8HtLVuEmLolB8ZRpiEzkk1Vq8fWNniaO6+8IgTeCeoyk9/QDHckCD+Rlw8otRo2jlfrXhy
lBGagMQQI5CRIZR8/AwVUkCjfVYiNv7e7Y++BcMWHd6pXUNQZZdssIT69d+6zZ107kIC0dEruOu4
CSOWQj2vBs9GSBkEh6DLkU5e4uGWlRiTDXu6FuirVJ536kK72q8Y+E+H/024Ypn16f4125U2WMIT
AAdUG8lPT/DczN7tawPSWRJvFzJXc6zMqsFQWTCzuWHt68awGkf454HDcC9LSOw0Q2LOfqb6b6oY
ik76fwfHliHsvSx0hfaCBpBpOLugZySH7zHsZ6JxyufiB187+5qGiAh7f/Azw5hOaY7PNrgSjYDq
c7s4B2p5CYeJiuDz88o44McVYv3hXrojxaCoyJUpXzyFtEN/oDgaVhpaLLCUvUkdaNGfhhWY/t3z
STR833Hei16pVuvUL4YGWsnJrIkgNvWjzcjGCVVvc4uodSYtnW44+NqIuNLy+eEKid7YvB0XOkvo
cNG6JTfRLQy854U0iScAEsiDfgAf+p0XXLrcXJaaGVX9oCTMhxwx2wMpvhKNHCOhNfBIBnXSW5pb
kF08PV+UWDEFpfx5W2UKBX5epVsBUf6owvhhMIj+E2auAh7C1DnC7g41L5+EiOd+P9JRj1DmiG3F
2Qw+Q/OCX986czIwFtDOjw8/JEcC7F86VDL2M5iXzVO6BXfUiYfJPAh4BQQClrJlVUMb5aFOvrzK
VocUbsxTK+LrGH5oHypqLifeVxdmqrp8nfZ64wogZBDbK0Ecx0wk0NnosrWDWvF1psRP7XCxyzTD
o9PE1CL2SgHgc4W2nyFnagEuzd2UbW626i2uszHf4y2swSH57aAvfHegqdCwXm6epjbWxg83bQeO
krJQjC5lGUxr7dXe6WPbXIblrsrsAp4N/7m2NTP682Di2bdMhlCjklqK/2spcDcdAqmpnCZDfy86
U63lx/0wBYHuDJIfjf28+PVV1b48LcFsUI8W+jI5uW2JDFwlXxjRduT9wtSQpn5SJkZLTatvX8Sv
aTrVUoygzv9edaSx+nAA1RfU174QpG7r1d/Zn93v+eiXF2CJTUPhDtzQGWxXEpqNBpJ2T9mHwi0c
LK6QWP8mSuzvig5pe2UlVPncL3hgA9jYacrg5/rng2AodYGYze5Lk8gIToT2aahqYuO4ezazrY8N
glVKabyZ7LMRIc/Vh9D4AWz03H4TH5NjfJmtS3m1+IhSsCN2h/8vhNZ5z3jK02SVCGQ/PxB/22PM
oxSCH7mTMRLy+ibcDIzjLsU/y5Lorexiu5HAKl83nchHl93CG9SYzlJWaVeiZKlqasSAH5Vvg8XA
dS/Jah/iW2kOKwQseB8NEClo/bwc/3puIMJ4wBDOMM4yGa5NP9gavhAouoQeAPBtuga0BDY6Xee1
tTzDmb9fNLLv4Hhuj6cBAHN2Nc/BYTXQGZWRtfJyimio8uc9oh+XtPM8k3Os4M9zDFywxoIunrlP
ygfBjntbTBElluZA4X44znj/uMdx4dd/s2cnozDsK3VeQ3U1/vYhQoFlXpTpi97aM/NSZDeqAUsT
Q6WYDMLWONk8zvXD0vdMoMIX1VMZUKVYr2ugUy5MHrz3waq79Au0NaC2hzc1crPnfQW0YcEh06g0
P/AjDTHZnTDRmns7kiNoxIoRUyq+VjuUvdKSSPWvP0lRkq+CcousGFSkOzbg2ExuiF1YbAYYPLyT
d+eZ+HOdxgqCfQJnds+Wlhx/yDnwTwNwC00GPwZ4f2+S+VdeYG9qHXqISJDMZZyXaFym9/CEkYLE
DXsk3//5lIymGJt+BVlxHnWw5KN6cYnySEDjGaiKWj68Z065r9jBYlRvGk0rNJkU/G/SsCPceTVg
MCb+pHrq9rvmRY7Ahfjt1Rikh9zZAkV9jrcmdYJm6mrdNGpcQ45qu3j+GJe8+BvliBAr3Y3smkN+
3poD+q0ejH85yKmaRa4YEeQp6D7blsXYNkjE1zI7UtlMmZHXg2zYYSF6RSDqsendJuEzY87XpO7S
F5q1lXPWR5jdJbO0bSkPIyeuGyenajID0frRiIc/pVspUAaCaXyfIhm3RcJQuOSNmwaMyRE/HSxL
PpOyAHVUc6al+iZ6cf92yuF3UmI6osi8rvbcyBYbVySHuLvIAqgOo6w9+aijUfe+yn+8hEcswPZE
wor7AA7RO4y6ZalKeFqVHCt+54PROpvwNFQ6LQbXugRHpQbFUzL7gl7TWgPcl2/X9/QWTDYexxLD
GmhEcl0deBhxOe9dosvK2q3cL1PUjheNyRCgwtXD8LCVdxkufi8G1mn6Q3AKialro8MMtKkqaXL2
7GtOsdoLCTsoOREzFYjzYpV8RdgtbrCAsH30ZVDXU5igWbkJNZ0+5GmPgojkPTS1NGjMhqhMH2AI
7gcbt6UpHlYrB/YxRZIdhIYYkXaNtO6BDHM1IfmLow59C/mj2WGcxtlO5GKdSD7abyAridE4eA7+
mtvtt53KydM7zRT7ex5s+6mZ/sKywroXVRvOIGgyX6KnLU2KIIJ+cjpVLACJi8k4z46KpncbgwxB
fdZwIR6ekZ4noIvG7ItrlSo8zppIysA/+CehtRbf4fUmPL8d1OXUXgbXZdkLudonVwEwHoGleXlL
NuSavckVc2y4q+eh2s5OMlGBDz6uTvBvQmYNPdddt2PdM95SNIS3xlSUPpVLPTGuVM//uF5JnYU+
vbx/+G41ID7cPaRk2xjGaDmT5fR/6kC9CMpdDbJcnIar5zZ8TPlFOgoPWtx8+0lDaFqECTl3o5kP
RBFG1EtBqXnJz0pQzqcc0PhfmmsWU87SDyat7BoQgvdQ5JTEFAnqmvAtugLWtVutueNFKpCdYMsz
fZONpDboR7n868IqDjpDwTWKQeZQQgNcka/C7TfTcRaKGhjTq4hU5tK7ha7LJ8T1H97BF4FPB8oS
RlKw5/qE1MK7mz9j5nP499Hjf+37Ickr/AfTiC9kOsnjXDaBrtqgKOPZteK8sKGufo9UwZTZYvie
9LUOyDD4fmYDzmlzVUrbn7jrfoj3c0p4TDvWqnXyh0xDXhu35P1dcOgm+zH4ZbMyi81hr/18Ln6I
Lqb4sdJVpW4j8QDNiSnajVucu7R+H+Co+3afBpQSeY8eG2Fnssly/zn54n0/yycOLTxuCvblm8IN
GHMnBve5TAigVymtNLtm7ugdlI4vj5MODCn0zyZaczPKoUarj1EnTZMlSzJrHMj9l77hhdhUOejD
RpgNylRjKSeTnR38FYEEPlkDMASMTl/CQ8Li10SnF0itBNd5gPflbpQXUduohc3nPFbHArq6tqJx
+7Q08q/rMQgr70zrGoFu4NuWkyluR8Oi7z5xM2IMmT8wpN1im8Ualql3wtofwrSCmuxnx2Tw+pGH
4v7FWwGw03KXPC6a7JCOUP+ClkSGDbYyG+hwtv/YpokI9wR2qqLOYMN4NwGCuAIv2hGhxlKAfUdi
w+GsmW+rAHEyV+aEZGHBwbe2K7LCdx7ZBcqm4dEY4EjhYeY2D2b3nnsBP7VfbGMwdzKy99TmEX/x
c0I9pVLt3pbfbBM6d5id53TIky//b7WBaLHuHMPKFkm55S7LUlWZ2MinsVx1PkOVvlOj2FvWPbFp
gPaZWlPAdN0u7rbTfgbimLZJTOG/BTSF1KNH3wFzXs7KjnzOQt6zc6BWXl1xXkGAAHfp7IW+2ogB
2qFlWU1saORFBuaw/07NK4OWCYN6gM2AVr5V9vH5QADrx3iLngzKk7jA0CCHw5SC/sJWt0xqxFea
LDJkxhzxdPbVZEw7c8MqcJz+9X9V6JHxy1PcdL/xFlh0oZfL93gBDGgNy/5Mzx0gO/Y4ryUf3eET
T9kciGd4nAgjvK2vr4iE4S/GQIw8yuFGahdi24bHMAghDrqDDRnTqrRNn6bnhEAnrczItBgGbO3c
7ajgR6DX2jiO32JbP5RDUUULsjNW99+jBOh2+kwV9xpHgUVjV8pqcD33rpCkJkvrz17hXyf8xwS2
L5jmPeomHpltBn44ZhqtQBhG5KcrkAAC5IG3HEV32laa12PUaE8thWn/227zvo3uHqkr1C8uVlr0
w6nKU8V5ZeqC5JgOqakHpA63ThaZlBeif35M7ZEr1ZcgWGwyCSKt/xTezDpwN59WdeqoB8VKIJ9b
rQj1NarckGiezm2PHfIi2fLRB9PNnBVoLZKUqIYJrdE7NlTxs43b8PV53ERJIDAf7P/BU7fzER7K
S5XjWmSwUiRHH1176/5C45EJpDWmCIjR7A/oJ2/5CBKWmq/JSOTw7pP4p+KFYJNHRPhR27T3K8Gt
mw8eu5EKnxU+adIYVLo4/gJEWAevjmLEvAmcd0Pyesu0lNR9g/dO1V2v0+5RdH8hOzp24zxFpiq9
x1zo0nmqY+xykzi551+ADHcuAREPxg3Qnpl7/f2R3LTys7x3XUSEBoB9lPFeiQHN/QOkqenzRlRN
SfKEBYbZHN0cP/udRsH319NqYS/iUZgRXKaxYrB5nasQ5itWlDV16Jt1o7hckAwr30jAgBMTY6vg
DjnU8FeoMeNbda9IaxEM5xRXGp8YxmYdhjjDz49Z8uARqYEQPw3uNAKGrrJiAr/jwnDGgTHI/cCX
GXGPJjGFz2qIfcElaAs03TT298xioCGnP0lS/4zC5u4zkGyrE8+Bv1czLT80MUUD0WXKfejaOJdu
srVGWxGxNFWhnXWim/66+jp9w4ytloHHIplqf35Wp4aA713velzzpsj5pa181BHzAJqAoiCY5MHK
9pfzF375J/+9Xjv1h6JxEOG333boz+jBqlWYCHR/ZszgMA2ouMQxqGrST1/c+FWGD+jzFCfrcGis
MELrq9M9VH/Bcv3Dcg0TYKFO/gaH9TWzDcYF+HHVHpJa8UQ59zzGTAM0WXiJGstpWAbutWSplcqo
RryAz6HmYuxkKG9O0ZqdlfAgwy81VOq3wsm7WEiLqdW/Mv7tD7IFpa4aV5l40RXoyUMH8VDIdgcZ
dqI/TNDZDMLfasAI2NePJ8+u8DaY5jJw7JBM3xKyG1DRtypwSGgan7wZEakc+mGm6WeO+SqDGwgw
FTTJxOHNkbPwxAb2pYr6nz1rr+M7ftIsoCo3imQ6KzbkUfonhkF3ni3aCCHxsdKdcRuPZ1QRCP5J
okv4q4lEWmNzJMkFwcq1G3MDMJhLUE+O7K6T0FVIxDm1PE6IBf4qz3/HRD7vV3M82cKM91Bmd+hI
7JaL6xsne87zXXJ/3GbIsIWXfqUYnKFOXAWEgI07w6tkZ5dLQKS1yMC6OqkHXiZnaqMn7gCSYoDr
THJinYUR/5Uggbs5C/PZ5Pywf86x49l/51WSLYZgSScdvbLaLy7mxR67ke8FuyknEYCKRstMvUBJ
sncGtohU3Zp0CLK+NiAYN558KXQ50wQF03ahSI6QFzzIGcOdHI0KGn/YJZOHvDOBjAc/IM70SEJK
RZ0oUdDk/bVLwLwF5NwwtiSdi4wUZIXXdPOjg+qX8ZRxwfrsDKYyInkOasEFFkottDbdoKFDfS03
h9PrrBy1/u906qAfUEqXLeiYfAB40XTpxFwPYFoYVdP0R4v7StvRYE0yD9LSHUEQ+BunC0mNWKCE
OrdRVim4Ij1t2NFQYARgZBkwGc3FVChYRAYh4oc/CdkF6+NRZqE09HKAWRcV+OY30qEULIM81hxG
iCJx2bEEH/XMzPoTz8AXN42D33uDgzTZ/1k49kgnWxTKGA6xOOirOj3u/dZ70R0l5eRY5gR/rHTu
sePUlo52lefomePkHzVbGtMQvaLNfJ8vhNMpNLE003LYK2rDeSPrYFL7Wb7DzIPw8Zfo1rExQyKS
EFmwonmKz0tnb9nW32XrsFfQmRIWvVIDu6jJK4Ne7w4AAYuJXCD9aNiy2wmGCTZ1Cc3JkzWkuFzt
P3rHBSErndOMlubUkKktwNdRROplZNN/iN6MxWv9RFrOYjIze3igIAM2VpIv4VRoOb6fxCmMJyrI
dZkgby7N9ID9BVxA8XBVrVmE9ttQuvgSWZhbY7MwyxYalhkRJPM9IgZOp0ydpDGdaB2lb/fTp9hO
ToTSwA4s6mFkbI8/g7kY1zSGV+6RsVOMu14W8aunWTPWEb6ObxQnwCRhuBOD6O51gZrB8Kbfx8wo
c4iIH9xF+yfYjby6MEWZ07eZE3CKEtQTKtmP6d0/isIPnBthRue1TCRjkLBcDUt/GXs70JnUY8th
+jvEFBjdVERcQN2FRnvLw6ApcdbbL5GYPD4ygCwopj53cWTgl027h0KvlMH5CmEz4IEmtpMR/Zn8
8WSdOYXneo89s5N9uDtrZZVWUNBoNkP4Vd+pv9ZrGd2461VV3Hd0J6ku9Ve7plwVde3U/1I02o11
7UAYOZnszgAgE4mNAMkoBwlwrYhLOusZP19Bi7hO76HSkoFtLZDd+E9T9+JGyufqbYOzeTJw8GnF
JpkLCLZ5ldfotJ/7NcbOGvazHyrcxT82aAto4/NLLT6NtrpfUYJ3+PPIYZiSe1liU9PRCaF17ThB
0KQL2Dt4CsfxQmeyPJo2/PA2xrcE7FaWdfc1meNyH1ILR/b5Fx8zpYJVmiygT7kS4URoaZRFNwiL
k2eUvoNyzFfpGd+jDkIN3kKucnrJZgy9TUfHuRQvfdfz2pd0Q2rsZxJidCOFFQU/JyaLh9DO5OaY
uzPyglrrRYr0RPMrl7x54GvqD9RNGV/qOgR+uIPG1M1dfRV3QWX2bY6VdNWxLCKqjnmhhoARArGC
KXNIi0LleQtBQOMTDQTXFyGpcVZsU4EAMI8fFUxT0ZxMJXwhytegO6LnhNZERpNI2J6bF8TkDSVp
N90ZcEF/vS8tNUUsnuPupPgZ3fUyjZ6wx8TlKrPqDixw1zjyyo2bByoPkGaQnLhmLr1XdK1nO22q
JGi54Bta9a3RDUS9meQWm84iNJRRR8a+xzhseL0N2VOsixUUJ8gnzfwufyW+vAGNEDPT6uEZ87KJ
EXmOMwJeW5iM12t6i7bEK9GA++uZD8kKivlobhdVL4pD3hmnFRtTlAApVZt5L2lSLcdyf4F74Uw6
4o3Lt1SKEP1W8iZMuP/S5DhzWMCL1/lhlt5/9PgLdaxox6SOwJau5sZWTv/PPEnHNil5A6fDnXBi
fjs/wghQrAnM+SuDGCnh7ncoFyz8hElew4SbZpM+XVi95tnxiW1HP/2pS2MmWGt7O2i/yp/HXnec
V0wqALZroJJVG0K/QxoOY6b0u7LX2FiPZtp95uKzPGzWjz/FgWEnoUsz8UBTW5iYguwx18goTLdW
wTqSUUxxD+ZTIX77jp4SH9wPaTD2eDj2Yi5r/0Lm/u7Nd1AGMTBZX5Vfig+X9w/Y9zeT8le1j3x7
ozN8pAWkVUhBS8BD6lI6oLktlIkHk4TLDUosxcaY/mykpUW31mMeSog+KiSdlcD50Lcjm04tAH+w
pM9E5bK8wls1xzz9AiWImXzRBIp6byjcb5wnu3j3iZ1mIhQOcopJBdjInDgTpT8kGi38hSAbrXul
+wwVNW/nCzvGhbNVTreKq3bos9/sVpIC/SM5urxGNqIXm7xHZoMT4mGCjUq516swQ+OrDbAYGcEh
y2nidKdn9Z+PPsqjvHCBpDoIxXrqwEcm2Fnn5+SRoJ2RMahgh9pA8tlnO/5XYpKcjPc2eDsCbW1q
MDwHgUCIWTLUoy837pzEuHCk7JlIoBnpDZq+EGpR85x6ALDHWleq2PVfx5nw/myQOW7gJbeoYaue
nXYgqNMqiZO4wQDy5nK6uhazuqD6Q0df+WQBDsVWrkGoHLqqLaZ9H2Su4bPfuouq2t41ooPH6nmG
GbY8iYu4ZvkEJ7VUvw4JODRR+PPi7nP7yj/0BX/pWLscjX8M+35mInt46uRLoNLbn/6nKMpdaQ6H
qANctom6lQUasi+STAflYXlObIduim/ABnKWWLOSLLC+lNDE/lDrVvQ1SOBeUVBmJhIvPzPUWIei
36YzyDVic/Z0uNgwy+PlD1m+AxZzSPB7sUPHHxJXO/C/dZfc33qNY7fN0nRPd03RpNyFdIocvvq4
oV8XFYiPB9LukK5Zj5RQuXq8ZVOy0UXUrtgxJReViTgPfC5Huq4E+yI44JKCeWOnZd0dCqwhOU+l
SnUN+PVlyt99Sk2Jcu6q4Ogajpv08uO6Uta2tny3wHS9HPuEyOtiv6fT9RDN7+F0vEXRQI5ya4aq
r6YnrID6k4tw75Fggieow5AG5crbmAkL8fXWJjI9EpunrMmpms0+bS9LY+ZhIODBchbuFsLeK5xh
1Bn8NSWre1/luSFzmER+gW8uiHwwReoKaTxzbkR15mCvllUtzVYCGJI6aHna/4nV9+S9xGqi20O9
YuZJCurW2rYoCzhUgGs++vNyOD9L9A5TG5fzSX6xBYFzh2lW9LFIctDHLjpgGj4hm0paW/CXMnxd
ewplQAieJRC+Fatxr3S1kknR0hdwF4VsqPjhcAFlLHdwWB4ClaE5o9UfQmufu64AuAJ5OXAkd+eX
NUWd1nODB1Sz2G3vyVhs1IhruqH2E1I1G4NksRhZkzejyae+61DpeQRdiPr81v8dagEgOXW1fs6H
XBfKXkS12C2C5YenfVbL9GJfYPbzplmjRNj0lHB8/U2qpceGN88UduwZTnQlVmaMUVcrLeAdIAfN
TsKsvNbDhfRPE2qb2DIebkmtZeZLomag9RcO0df0y0oaU8eAIaaOHgZchP5j3FNr1FGkIwdUvgcR
SvgKYEMIGuX8Xdw3qjTs1M9UGmDhktsOd0riQgi56Q/TcOiDDKEKksGY4bo/MKr0po/3VPtJOIX/
FGyjJUKxC2qzSoUinU6BWHnfZv2dbihUTPM7F5KmVAhTCRZbZqAxW6dDd4kVrpYtWhJefpCUPnfl
NUlLCnf00CfCq3OjhyXaBV+G0xMIVjhTgL2QL/lQBwI2C0Oyy3sWUnqbcdZF2VQVJQupuphAVQOD
jkTjvW3++lpuvrMZ8XoVJN+Zv8gPFu5j+mQ3yUN+trHpJpincLbwia8yPFbnQbGYDTrNROogVl+G
zPLNkYYoKFja1Oz5GvqEIFU0Iv/YGqoqUS2K9QGCjB/SMGTiX5plaE8J3DvT8meJfTdi8y7EaSwE
iFQSrUx7JuYvaQQA+XLITjcYcFcsZ2gCWwpoDMmWPs1MkZhcymcX2w3COESS8D4ZwIhI5TsSXGhh
nLO7AE8eLcydxlGCjBcnq9zDRH27NOjdQxhGToSj1uyWEINPuccqsAlXfZDGfy37ZPCStekhbNbv
nbuWil9WY83piPpgcT0tic3d3kM6oVvBzJT8H8NB3Cp1Dy/zMPfp1toPpeCL5QQFtKwbskyWreM1
v2pRhxf6LAHNSIGMlfZtvLyKspngSDIRDwexHuhLOuxNW+lOlbbdFudFR6IGEjkt6obSZ5uj7BBk
pu8vfQCuqpwGrpIJ/eTHmuvteFXLEWzUZbdifhd0v6eKegoFiFLqkKtcTj6VM+enBtK/mZbfOrin
gBvKEacz7gGaCxd5YtC/AulznzP1hwqy2Q3kHdc+9Hw9aGeIhpA9leyxAyvItcsXy9WZc0I1l6ML
AUUdP0r3VyJqcngwh71W0kT+4wK6JJH1gKzAuM8gUNUuEIojsuYPcg0FBMY084uoJmD9SmRpHDvB
djRZGrsspwdwWkd6pCri9FSWvdYvAkjy9EAwXDJArs3cO42gziZjcvHp2SPl9qziL6+srdt3Bebk
5iwUxwW0D+FDxkO0eOOPsIoOjZc2WtdxsiERx238/8Bov1BYW6tBqoBefQn1OgA4UtuNct++2Q9Y
LbHVtlqyFXT6tgCUAVLJoDQRNVznnbcam8BzbygXvWmR5YDyJv+HcylYw9+9Fyy0DnxE67Oo1qg3
CYRhWIwxlMcTeKjMceMFr77/1cQJEAAzioY89cS5/JtEry3nZLSF2zXXgWrALquF5VvrCkfeflJi
MtrLA7hYoaQ+I7s9OYcDwM4ssYi8JDSZeKLqOrnqS1MCzl2YQv3OprhwaVT4ppvuh+mL01GSwrO+
WSb1Gbx9g/kMku+8aQyXmIMGywgZQjgwKXbtd7xhbOQhDxb1aVGoFNeYzTZwq74V/kqit+LjU9WH
pumruDd9/l/Jh+nVVtFcRw7tZbCilqUa1GMOV3g83wQR7ASq35faVtUfkm9w/r4rDKq9hx1Q7jhD
Z0qVCLIVM5tScMuCZwcjoF3tG7XZ8y1outVnGwPKmZ/3RPcRonj8LKIk5uRs0wcZrlVUoys7y4b7
H9xVoONzpN5bgyip51cz+hKK/4PER8YbyP5kYsGW7omXRv8WIw/E1Qnuz6HPeUmbmTeib96+qfyi
IqDcgwPziiIcV/JIOn1UJaKxEuXDom2j2LPZRGrR2kjKYP6IJS+eT+67/UjZ9DQ92LucbgM6jfM1
GLR+tXGhzKwc/cuVGeLpe4dMc0aMnKNYUnfG2A5XuNh3wG8tUU9ZPe27l37LONmUb6YHE6jQossd
0k6Pnz7UvxCAovP6UVF6CpPkQnOnvECG6cGU2MiiZ1X97BBNAVYOqIkz9GozdSeKqObs3drUJm2m
tE6rmM0K+S4Qe6Ofjjammfxc5UYtFKbg4hz+AqyeV5YNdEsF1YnUVTs7X7zg248HmxchISSTo7dV
oQiYDDGnONjRSvkx+i43AnJLZESSug7Grhtk6mjiqox4ChA04EFH8Ha+GoFmRJjkN5OVx+jQuGWI
NPCtCCIihUJOvvEeZ53MzFTJC1AIntaEVCZ9KKndkAkFYnO786SnwN4VvwUD8pwUZ1ATtXJ+cxSp
7P0ubFfmy8lmtI7sawiIozLe9SLTniegiBLeLeGjGspBVQr7UsXUpFyR3KJr0VG39arQVYHOyj2b
g7i051wZezNaDolx9J1fXxyBwyf8JpwC1hxtWATC/qxdmqVGD2NOeYWVzqdaBBLdHAGs8XhsIqwV
TSI6GKMTfT0D99/8blYIsKoc0KvLh3SH6EIrFyrKoY/PRlTn+86DTJ1FjpEVzfabDnUAKsG+rFrY
QWS91zGViEdhuusqlbUZ2aRB10VVyCcirNqPFWGEKWH3YtGxvtHtTEY/vTC+1NxTff0SYwtR/PLX
/qCQKlr2bKGvCN7kJRjjhcFtMWJ99O8Gp0HRhIsNiCwGwJvljy8VbrxwbFZwTpfpArRlM3hMIsYv
iiUZnvhHM8TYeRDFCaVuisi3KcaMYDIlOKgklke/JrTcQnNfcp0TCf4bJIYkwUF67PDgPTN4vLrA
c1lHPHPrgAy52ULST2FaJsZrS+Iy5D4r4Rixm97/XosmHYk1YzceLZJpN6SqMI3diQ7pLoMyKTPp
DtXLeefKOrDYQSK2KVj+n5HPchbYUobHdVG6IPXPrVYGW64qieol71HClVOI9qB9PFG9xaVF1OOz
JaxxiDCY6tBbjCNsbUTLbijdUFDT+oAwb6S4RebMInoC0zhymzDilzf2M+bT7vTNtrkYdFQxMNM0
zan+x/Fnqz7jQ40lOO1qzUaCDDGdslUQk+/IFmoKmkPywPIU1oizXu4KZS8oPBd93bYlnyrlWEzs
avIU9c/74wwOeIpW1wNqpk0WAFCJXcv6jzmr1n1LKSM0AnEFeyIUfyEL9vktgL1vCrkv9jDXO57G
883Xjlf8Xjg1uDZEX1j//PAQyebM3fPAZZgBl3RZTJluVbBcuUq3MvO+Luktr0juSYy5GzRBnFL7
EezHyCAi3nycFEqexP52qVKCkKedh3hCH7dnTJWh9vHJ1ZmxM8IKFdAWHEZFq4rJTmkjsqew4YEI
l9EyqHWkqHRE9SjhXgSvKZiW1Z7/YFkZpvL9dU8voSEtkRvRjsgah6iuWmgnPIURYUxPjJ4w8X9F
tghn2FkRzu+LGPxEmJu+y5ApUK6CwCvdB1LMQ7WDJaNQvYiddsZI9Ugvrlz3k2NEsFLVooTLalFn
Cl89dTB/ctxrLFBqfgTw5dEnfTE7NCaqsgHxoPObuQxlDTj0UvsB8vjGspw2UjCp+fL9ARyy2BrV
aG4wCF4/j6nCcwUx8bmF/9G8qOSg+05ymm/IeJPRER06qKDPhSvNjqs9S5i8JbxKa/UxD1f/nwwR
qfcqfU0fhtbm1fW6/8D8r7bQXE32bLj0wmjOUEP+S46PH9b5rxAG1l3uhege8Vg5XHURltxODwQ/
ogAEymx1LTHyDLyHrnXyhIt9Ciit73Kp5rtJq3qq0DafG7rFd9XcBgoQgn50GQBZWtlxPCf65MFd
GCJKi4vP/REwoWaUY4Z3bmXR1nO484rbZ4PNXhE4CAKKq4Mo7pDtedlFroaStF2HzuMf79bizP8z
UdmbYPKHXI9Sn62u23wk/SyOZxRLRgpSgI9ubLNX3G3NqB9yCF6jZst+ebKihGCLVvCOwKBGNQNc
RQ5MBKF8poEjwypxzg7RB35SDe2d1QL5u9YfmavGYbWGuMgis3ciB1zF0pI/qxjuK+r/kV4KrRuo
4j4T+2ER/JMoL9x9iM376izeui/3kQ1T1jn+ynmAopcMRr0N2Vl8ymTdORXazjnJaPccdkFnG8v9
frEpCjLe1wUf8zD7MrUapaluzvJgVFO/vXDpz9hOkBWTxwNtRBk/Brt9RTPC4dQy0SwYD3cH8+MV
zBcaswQHZW0ixjQF6BJOA0TdYXagvX3ji7jd5VS00Nxy4Fn1HN/7wOWmjg3Is3afOT+vDTR9NlYc
BePxV3832kl0qD+hb216PTlWZYciCh3X83qO0atL1BeWgGjfv5LXGrw3y2vTeA0VNHGlqGhs1yZT
wWTMVDJJIpSYrJyTAWq+zDO2Uc0F3vee+272vh0wwejCRqdBkwSuyTd/x/lAd7qm7bk9acFAMZwF
tYU1bGyHVpAGngKCDVGFkD4oX4JsIcmQOFh+NULDbRzIbtYvwiKGWvHlVeQcpApOiWYBjpunAlSr
I+re1ditvTIMeXzL/xVsDpFv8dV3n6xIer9A9MCFoX5SGQyFYNLkrEC4JNuImbYJeK1tLn6zzx2I
Rui+0eU+EfU1lTdkNsYCljsbYQ3z7Oy9kGtsZBt1InDkGG3FvOcIn19jP7QCfgVYLKuhXVaE4LMP
Vdb6CD2cJCO2GZ6VOnba6wUGpokp2gkZLyvXJ0myhl5SFPD141JdlnEWMgpNUnblOjrS0uG15YNs
wcQmlOpz5YPprO74kXFGtuPKyen9plnWEK+lRsrkFFDhjJLAxbFkpmKJSwTU+x80Ab1VtNQcfG/H
kY1tk8N36TCVMla2StrX9hZyGr3WDyV7pynlcyHJCIvBdetU5hjvMC86PEOceD+NxLsbJKr04rKL
LmslnNaId8RajgcZxr67+6Ai2ybK5HFIppiVkqWazKguGVOXdb/AvlxOABGgoFWjlW2fmAnQsO8f
7vAV8b4mHd0VsvXMYL129YjnMmO5rI51gYPuXeTznuxgTCpzMndATEXr2GKuFB9dO9hIavJgK1yU
m33lWHouKft5E0wAuyskpsUFi+tDNdjomxj+WrG1yM1CsXdmqhZ8s+vMF7+9ah/Lv258OABK9jRJ
Rgm+pjJ7tYDyj8KlNTS5jbXfi1t6VDNCuGOUMRcDi94/MBbJT/uhPS+cl9cmMfjw60WEqbxeA1tX
dRm4MaNysAS96A1zbdL4o9cBf/zh1Yob+F2eQo6GA605lZfyR2sSk8TWixhEO1vPibFzVImOe7xh
f2ZWXFZ8gfRzD3WdZ9NV6Xmq0u5UpwIvOWCgyOoWOkH27+m/tEXT6ao7rgowcUKAEx41kwRIlfDe
RUd4HTVg8f+1vJgVUrqHrFl3gzXJ/ysqNTIgtjmkr9NsApk/w6l309tYS742z4vQCvX58ayFgEA6
MM7LboNMdB7LYVjxDSIXk1sgnYAoe086lxNu56dFerWwVOwLFrYhF0DdZ0iqeXpTHaaZhfxDs5tM
3RBUGP7AGBSmobZoTFyWwFpQcagQKtaEuyRdPa2MnbFgiLBHpe48Mtc/GnSU4ib3YURjiX97beKX
JvYQvx/hHk+RiIqG/sv8zBskBpBLiZXj2zsXC6SJ0A74SuZNT6ljpNWxBbTIjKPZt5lfkvvMp4ZE
ydYSOC8xyU0KaI7otGypRrcJvs6HdCzP0z4XAZIiAq/xFR6tk7xv85XrRUE+Ll0kQ5RGbHN16Bfv
0Slzg42s8lbWoG7ty1IQPz2UblLHp1DPcmT25U6qdlOCJACRjdDbiTgofesMpJNmKXYT6yDa+c23
elfBrraTrH0wS9ERwTu8Ast1BFGwSgjYj7VZaEiDo1vDBdilL83Lu4fpMf2p2fLA6fHowaPRHG5z
+GxMc8coFu9fGj1yiymVokAWXqCSBiogkqvLmeqAHTGwE41ndvb3nX1MitNs+Ni4Dmzsk8zcU0uI
6m42THNX28clRQMlgqmUWbuTxOlqxoAWmsyVUWo3hg+lHQl6h/jgyTdeNmdVCWpm/FsBLyvyrSqR
54y9aoepdWs1XqLIHDVEknclEy8BaVYUwvMvmWAqyBMt/nEsVJw0oyFAutB28XzuPOdSrvXsPiVv
9AkHs+2pNUieCfC1vZRKgrxogEvj0vv+qX36lJSzsEwKfv6ey1aR4DXfmSXpgUBFk0z/IjBBuCcX
Hs4okI/j3Qp2hucKSnEHAeDktQaN+8qKquwj14zX8EjLSbkVRE+A2BPUmgt+JQg7FMJTKmswHo78
SDuZ1c2kouh6FVNwSctLW+zqt5Eia+q3+l3INsW44xVUjzYfY5wQW7aK70HHrHeGTDX3GnsxESjZ
uwxVMav80vNVBFbpYV+u1Rjt7Rgj3m1iQBgUaHYIJX6UM7YHIbFNGaRpNPldcKpdbhD/3sB4sqxw
ILWdN9cgOHF6Dkh0TX/HPfxkech/hBHzZ72R3wA+1f0XKK5ZDRJZYGk4cGFEk58rkSh7Fpd4vtSJ
bAk+oPIu9O8wWSsGirxnYlUF+r+iqzFF9If6r4D2WZnz2UsQGBBKWVykuqLCb0WooZ2NIs0BUBw0
2fDHbPAXKXq6TeIAJJ3vyY/vVuD/XUreJ0n/rC+IAEq09STcZIjYz1h5AG/nUdutfCKRzp3devWK
Y2pvOVnzPaqcfW4Fk2DbWP54+uvPE1w7KRq6XMGSE04p2sklnvHuFtwzmE0WYFpZS4St4utn+Iu8
9rKIA14knNuMCqXS4xPibnV1dDlkMO/1V0d/EWQZwimzcKWqYywz8qwV11lxDgXSSh1ZNd2TZc0I
5LCNDS0YwHQBEL5P9qavENrEHBcm775Ly+tomM29Spm9hV12Oa7p4bjciCBLoQNolCEp0baTFS+X
R6iPV4QGb3swDTgdpgYOOrhCLmRE+JzQnryNgC4Xr98MJ65Zqz6j79lw25WqVYgleJ7h8mSVviDe
lkZONGwMRS/33fRLc5R3lD/k0r9C3rFI/v0hoSCR6rU0zq3s3mM2bgiKmgOPPRg7oUObYW5S2ABi
Qh8FtoPkLC2xjybLVrfH8noz7EZZCxa9EncnKGnDj028K6c/at3Rm82CovL+tYOWB8k3JHeqI/y1
dI+lFc9zhtJL0kejk9VoqVmqGe7dkEwjC7TOt3DA0kWn41jDLVl//0eqDaOehBsOIwgb1An5vMhm
OP6broSddWqqCp0EUQ4ERdO12lrZsHaJVbPk9ZnJvKWroGDcf4GvmYGdKW+PYEdOFmMdJX9noBMo
y/qvg+C5xAveyEFWOlznse38bcS8n51Agrtn2YfAIxp4J370rPfewPbWC7iKjI44jYEK19CAtdYP
20Rwg8s+xo8nUcGHC6vLEmiBJHkWDsY9DxM6x/9moAkXzZpsNL5iTlHh4mCDFTr0EZ48xllDuK0a
pYJcM3nnw2AaCLIRUeIIUPo+u0lru7ib1pgiCxjlhCT3RzsShNxvCdLgqeq+NV8LGhuB42oXsN+Y
ly0H66VExCCPlFkKEpAs7FuRbumuhSqO/QajZ0s1si+ncXKSw+x060b8BqtZQEO/JjrGGoMWYln7
fjHCcht/x9E6U75jQ1oPbNqPXM9Ai0NcY1Sz+Atv7TcNItcP+6qOfmQ0eE+Swf/9E9YqMb5Dbg+Y
h/7P/5P+aoZEnlzhkTjJgbnotpIsirfelqrBV4lUhHxzpTrtM59iAHPNb4XiL9DU699RKD2Sm/w9
+AFiqdx6am0aL3AjSEO/x5UiWXVFh578KHM+1FH6RQZ/NKMOx6kMby52G2VAimjRM7UNWIn2tp4p
guXFnWluzAdBpD5vqZllLZ0yU6a5OsybG7KsooLejg77CL+xVxfE3VlUI9r95j0u+bxaz/ypecXZ
9/x5SVtzdCIjTDBjZ7cofUb4Gltegfez5WKRlEeVo97jQaaoNklKC60OJB7SbAARkYu4x+KVTGB4
wjv1rO9ZoGmzq2VGabayDFcU2ypMSENHCgz3OB5MT3iwmSdsY/Mfu7FPEq3XdlDDpNtz/7JF/nJf
71OsLV1keyHrHmlvZ+bmrE1si0Az4oHGtu05q9P8/LT4hl6lGhzZgL7Uv7JlP3FCF7EzaHUpGCjr
kbneTXKSCWLSQOOrtM+B5OP33gKYHglJcYH3FM5oHGPMLXJhb9yCpAnXlNqIMegfbMXQAUq3do3r
9h0+zN5nV/WRe91eviiRYMSi7SJ8wNfihhxslU2b4mho6fT0pvLzTg+0PUVKUUJjXuqfruNp4Ok2
A7THVCiFL23hNyiMThHt9EgpuLvTPUVCsZnmdHjFdLKousLGenKjFqc/L2AiVtbZixPQwHdg6h9Y
Lq4zbz1vu1zsxUJN15LhJHqjDohCniKuC5LOwEkFVjfMqCT3Is4jE5fjVuKmz42odWrp2Z8AuFWJ
xFbPlY256Y02iooxGyG+5/Kml93nzp4eXm3EhDKbDU7AhVmPId1RufxKz/FhXgylIJhVAD4v7vmw
LdkrcXFmlbBP12STRTZFivvZBER9D7TM9HQ5wj1MCUlF1+k4m/8H279zMIiey1eQGCLMFC1qdiQ9
1YcygUFmIwJVbv+8pOol7fzyO9FCmWWjSf07nCpVxZ5TXh0Q2dgW/YjrgH1oD6Z/eoSLmFf4bRP6
EjwwcjJPavc3aR/pJCQKHuF2rIlMIhwBo1sz99L47OrZnERAPg2BXhl8JBMdirgf6kpj2SXwmPHX
e+1VBEjQfb1tZZ5GXuqbswlk/r559fTp018jzX4VsgcwA77CeulKYQ11hFTPrHpxA+BV7pIggsrZ
cHCBB5DWPpkCYnt5qyboyJRxOz146e7zehWXwuJI8Y1iEezBEvD8IT3BtJAhVnNkENmt+DjXxl8I
m9u0U0iX/bDroUoSRBdvNz3L8c8KTUMfZ6egnGmf5ZDyM0OcM/RBqjcaAvbt0SgGrnyXgXJ/6eyJ
pchGs32qHu3UvGRwHthUEKzQjxvZDsdnWNCFIdPie3z/NANW9/9TxafaYjurEJ+Qd8VYbJxbRfDu
lu2l/3JDusPIen8eMp5zT+OTanLL/xiHX77rRY0dYkVbrBocan7RB+YebUJFGQ/cxi59ep4+xMTo
I7pkjgyiiyR0s2k6DcJkm3dtYli6w6q4UWLwFjQjua+w8eoQAuQV2baLl3iXRlkXskOrVthfWHSz
udR6QETG0CJj4i0KIqLIgWUcgf6sMWp0z+7sO5mxVEfMgGRXndEXFV00QAIWmAebscFETkJU7Gf8
dFCNYihGC0lwrlW4Z43AtjjVz72FlEHkDyf3P41Dl0xnFxSiFKh0NXCD5yZdl1EXEAqpQCcqh2qe
cgfH0XFHXwHoAPIhzKR4p8KCSXgHIhziTbda6BkiF0/rYBplp7jB7x5XFnUHV0UBKbLkCSZ/5fXe
qiV3jLg20PnObY2AQiyD5eqx9RDEi3aKkQ9QJTBdElcPkM1vV76AhZsGkyrlOjvs4+JJsj5J/aaV
0exu/mePyd7f2Dlom25fOsKp/hszxE83bTdwJphU0CkC7Le9VjRRQu7tDQgGPgUYVSSVWU7PI7u3
EXEuOEHwL/Ut1pn3q9xKKwzczSGNQmJvD/8H9G1GFq7C9pv3vfBZpwcaPxhPmh7Z0+gw6wEr2mTP
r3oga4zeo18GauOx/7pmORIuhi/n1pV/lobqYE7nrWz6fSkMYH0b9QI7KnRc/hU7LevrzeLZe2i4
I0DcL4wSlqdnLMIrYaX4xhy5YVw9hzJnCEh8j7pjlNvZgYSOeP85E0K+QvxM3NyaGLtC9evuTKos
3mhKqE24m7icVdy30ciMREjSr50W8Ikvwfm3IuREoK2e/LIOHqnV59rsG6TVuxsu54WytJ2NAqdA
iGzKXZWa1eDPcz7OvgLgLIjZvXDfGIslmA5fEiSS42JgkET19ViXk6AGVY/PUvCh+6lX6s4zkCYA
gdXrIV6aks4VswZenf+/IRAJqLokDuhiCA9MxA0lEu7wSX+HpPcy2DEvVT9QQyw3YDi5r2IGgUar
LEbQTLTlGB3AjN3ysgtmyu6EaD5kYUdMZj5SAYv+bx8QZvuNMk4U5Ow52dCbJrC0ixLRs06ddQTU
jJPugRPanoCUIFTyGDseGFyC7KahPv8iyxgjF/PUV48dWvLGLP9wstEnXzzC+r7UcAm9v2lT6Pse
nDjh/w6wBSJUzbj/HTJFcNwLZ7Ohinp+GusuwaHoFu62JEAqVPTlhWq/G5BnKteYPfPq9xPJErVY
6gNvjBniU7C1K2mW4Nu5Ic5BFgjVx8dS90Z3hUGxFbc1rp944tE4KnRTDAZ3ptrCW5MDtYIEwxfX
tP6ebwuwvvutDpXGjiAPC3XYj3HlPVZutFARdrHriAhIPSL4KOrtN0OrKqvWKTVQfkXI1VRCpl7M
4oUkP4XnANCN1IRY250n6dJSw4EAnHnZWi/LT7PeqkH0+e1/NodydZNlivQwW/tGVn3BzNA+gSWV
xoIzpmXDjfbQq9ypN61f9cEo5qyW7N4hkuPXNXLncBKRFZVmGc0zVabgmSIuHPgql7RqI7n8JPjS
lRPkRiiA1N/9VShPEpkhweew292gUDih4gdhJFQzrFFJ4LL1g+4SWnrxd9zzHq0VdHK7NZSOMFIO
6knB2H7RqJMEIWFvYiHmUKBizh0nQcTC/0CW5+jVQdobJab4CcaIQfaTgeKZC+eHg4Za8SY+kqCi
9+SLSlIa19VgVqNL1r+yjbflTwrI8CbIDykgYGP5IKrYlSV+27ZBPCsIoOBNfssO+e5jFsbnNXxH
l5r+fDi41WNe7S67b5NUAM3XjQP3LC1OY8x9k/yw7wWJ7nj4oYx0984YmRLpbWGbx+c/A4Q4zNHg
vQz9FO6GjrCIM7H9297Q3w07s3rW2FRDf2oYPsVIvxaGcg5ucha3K7/hHGnwmvNV0e2stLkO4iW+
vWANWjBGGdhypuSdvmZXc6OikYQCURbeoA7BT2+UYsCybdRqoGfbqrbFSxEELI5q3hK90AiozpdR
LJ85lvnWjYEC+EWRzVeVgRYnouCW3w15JmNfIdjI4Lf0qhcfh3svu7RPzsXGQLi1CSfNE7Lvh26N
wgzEQGMErXk61b9jJix24pC9Jvzg/dG+r598okN8ngpt9EbdtIT6DnqEiLZaLcNtpx44svsP0r9t
f4pGWco9pKU4ODUWkPdq33znZJv0ZP8QBtMh/EZZA3IaNYcs7w0c59qDcpGqksqE3oeLkYIi2/iA
mrDWaXKvwtC04bJwx23++8ZGGL6bL0LcS3zK9wtSFfHTMcY3CsNjxiTfkTiaWWY4YQIi75Pb+lYd
9Ys54Kx0Fk7mtks1MjtTpXJGwHKxFZOTYR/hkocePG4QrpCA2ZLC3WbKqxZd9Q/C85SPWg9B6feR
5yvrvViqKVhPt9sCRmvBlhRglGiKZEkWNhmQX3KqyoWHZ5NiFw6FQ1lvIoeCBGH7rYTSS51+YvhL
nrHP94uRZeoeEOTcHFTjr+TSLKs2En+hBmXsKiX39sV5t3Nh98wtBT0feZQJp4XJVCAhugEjkcge
OwMg8DixYFVPUrqrPEvPlfG0OgiEORoUKAYSCvFKePYgKghVBy5Ku4PcK/CNMJ8iu0ERSGCJC7nv
ktOsS5OCQjVXxi4Afepg4q7/xurJ3HTQNZj10ZUBEFbMvQcJbgtL/w31ctNCmw+g/ly1YoazT55+
9PSeXOEKVRJBGB/CPPYNxY6PniEkb5k3gI/qtSwOuC4T2CaSv1IK6oYVcd30HFtJXwJ776/y/elA
sBhqqBssNnfPXsOlanHlME63bQfTxZ7HQkgkwq2mPj3d432uBOvUgLzHyVEowGHkWwVFPweAfleK
kLSmpCTJhraI0C+2TqrZe1F1y7hBJwTF6HRtIu9wyPICboqbX/exZnuXZYq38hub6Clyi/L7IVUb
JaPdhsSczsJA81I8FABZwTKTMDrHSO/p6ZK50EFXz+Kp+xhCUQuJPNLXD2KipCuVgS93KD4cH1F1
sOyvoYhrcuRwOyy4246oCu4mA59MDiUuRWqjEBZTsXdptRDzqV89Ce/vPVKkuKO9sUxj/YtT9qXA
qXzpKTmWt/yehHYyeEjuZvTfIxool4kavExjFiFhnV69+trfABLpnJ6jnAmQbWhdywwpQbWwZj0+
h3feJLcqkDkzCUNLwNIwWqQeBP1KTGeFrQZXTfngug/Z6QCuLmL7HHdcQAvgc0e36Nx25B5dg/hW
59qXlbldiEdtb0whynA9e5JxEPr7PdWVvHbqJMmGBhI4cLdH9Xw0OJ/jkHljJbxTwts0odiU2NPA
n9WTHwsH7j1blGQulRhsiGf20GrRyMdt+tVgY/pnhNfa7F1cI8unWuOa2r2L9lWqNEHeNLT+/HSe
NnV5KssBovqyqiOMMEb87rwb5lR0ntbKBMEpU2gUZJlhqq9RiDfCmM2TOxgP8hXMxXIPrKqZlAeV
+ciMN1aKwvC9h/OruoFaTCDufYphU/Ir0ZiyIUk3sGe4w108fWNJB4H9i0MkERCuwyS0MzP2jo1G
EHYDLl3Z030J4161A0N4qGYLs5EiNEwtXIRWmeLkcT/wUIEbg3RtIF/YPN1LgOhRvMXZSmher+TH
xDlg3Rzj0fxSFS8EdIqZuK5DzvPUHgd6ef2SBnj/ZW+qhoEWwicaLzF+SV1mNa7RjIzDxuKj+Aw+
bFCfOBWvcNrpg1EQtxkM31HnbU4X8K1TNW3vRMGleNVVJ0LcrhenKla52SVmxznS3fmMU4KkmDce
xyzd0eKV3i11tO+av11icb5RvsGBve9SXieV0AYP1NYcgiQoMTcxNeTZFtvMJ6v9CPfYVuDowBaJ
rNbAq9Eo9y5b2Q8WkeW8NOUqhljQZV3176ZlopLx9hSTuB/CGjZlnOBvUXF0BKNoBmoTaeHw8/jt
Gbmhcxkdbeo3KV+fPRB/ivAYmkwl9V5RkCaf+URhtqJu3EbpDip0+Ji0DVEsD1KQsecwcEF7Puss
qvYTFVyhBRboyam5g76CJrA/QxuuUeL/zYLbWp88+g1MhzFm/ItlNjSdbdiBoT/Y83ZbgltOY5Pr
0uqLs5ZfytJ7zqidn6Op+VUeQ5qTl6ARbp4I2VRs8pJVK+/MadBgtJOV0yVon4zxBKC6ep0/qBS0
6udgCnBKjpXy5McaS7s1wSCMRffvxeAb2jvMj2fQ4LoYeErFuFeAvFjTsfYFDB6In9sVTzP/jlik
SbWiSk66k8JKnc64qtBnTCyP2GVXGWpwzIIwvkq96fvEYHYBA8NBkSCBUBYbKpViuDUEbUDv6roC
1xZp8RG3U1b5k3bqulwWC3kl6QSvt8uRltzmwxnBi5gIdXHax4BJ/KN3U7reMG75FF2pyYZp4FDS
FqwEbLRE6glT9z5WUftym0cKPxwLiYGFDjxM64vIQDeYszJN6k/zFjtuPLpD7aacS6cZrkW2Y1Lu
Y3NzrgyClqQY7oTj5aWuczoHIudbkM75sliwhyPe/amNBZQJpG2UvnduRGu8cAsQ3DoMDxOQg8MU
JPkisJo+SHl3iwk3Tj4CSz/j54iuPT2By5ASq7BXfKxA37NISqF5vaCJ7Z2nVfTCjkRy6EjtOsGG
Gx31sb0+6PmoGa80dt+EVVnCR7c5AhTExJ91Vp3/Ko0BUJfI3uTkFdv+FwomsgmGd5sYJXwp91X4
Oi0YyzTR/aaWxT+AhfBQ2gzVPZU/78HC2avZijXE4lm2cK9eTb7cw3CfluPDQmCxbxaLdp8RaTMg
bGN9zeRY79OXlgLx18jilOkg/OdumBet4ETqRTNZJ9kyf7yg+92FKKWMSTF4dGslu9RweLCsU1th
JKLW+IDPBNvzXxCWq7etqQQtZhM6d+tcaZCjsW0o/tDmX5vYnZdmhCVZrMrNlPv55x/qAWVrEkIp
zM0bZsSgdK+hD6bpBFrqitBJftyfZr2lcinn1HXNLAojegjGuQr1SUaavMpOi2tK3rW/zECGYePd
C1Neqh11xLhmJjZdvHhqdn2Vl+aq7/nmBpO5WKHDHqAamhE3KgHSJo4AUczG34xa6IX9Y29gpVSz
khEXeZTpTcxFwVrAxYmaGFGIO7E75n/msf1O7Ak1j0Wrrv+Fng1OyEhIhrwJgNrCNCatNYqbuK8h
rJiuiDxQZeXlyt6XBo1YqwodUSXnFK7r6DAdtGX9DWY4mwoRaN+dkjhg0tehXZ63jbAgrzWHW0eH
SYceSZcJ9JcQXRrdAqogJKNyy0F77MHkcDcbl3gplgHBWe2ubJecbPCw4wXKx33OT2hI1JkyQ/8z
pSs49QdF68HQNl4dbJefDnFwMYsnoDPhqEXqjkQlBYh5o+o0TRcqYYch3Gqduy7A61mi30SWzReN
a99ljrrEOW/o2VL8a1SbBFlAeb7FySfln1XYAxVCBjhCBektzpPeEigMFOjGlGiFKuGtNj5zfBSJ
CChY5XYdqftvO9jrYEzIX7ioeFOA9tKWipq6wUZiQ2JUBNlVdMRQsY/tHAY5QjHwAO0dX0Hmgzul
t4mR64uIcaDL14lEsI15XcUC5353GpXa1rJxceyICwZiHR7MQG30rnGIW1z4BlYOlg1BPIEUp+Jb
9vjPvd/LGMMPG5jILZs1KUIn/Dg/KIO6JIUwQ4TAYbJt/CVGqZZRBo29rgskxYILdghuG0iShYOs
untbTDj/uydbvkqmbmtG2OEaFAQNOZr9kDJAHcBNbjfBG3g/NF5pPqr80bGCp1c4jI8rlh6TUV5v
7SKpknyoHAhFNaOR38/sYM+u/4Rp8YZdnVcyR85TmcXq6mik2gWiE0Bu8JuFp2+OrDX2KXslYI07
UJoL0rX+tpn173S+PcycyTvAj8MPo49diIi9s01a7l8oFy+gOoNafrE1V0dCiQapSHDw3Sry4VwG
odVhBeO8iguAGPa49ZU5Lif3pf6y61lLeyyWI2vMEkdlHCDIkdiT3UePImgrfuygvAKa1JZrVZcT
91MfkiurUT6nBTAk9if2MKJPn0aO+Vf+1oqUaaMeSAachhol62EfRlvBLTvWgLs8GkzvW3VBh8c8
7h7N/OqVQ8j3pLLCRcZtEQFf64ZwapG0VeeCRiAPbAnXZBZ84LoT4co2TA0zmv787h4FrVmgPF36
JCeabk+aIMNNvaw0zcNc1HTrTcZGsgpb+jP1Zj93Q9++f5EaLz13M4wthTZ7wTCqqiJT7RBFD8co
nQztwENbq6lcXsGAUDXHa+7pG7ImEk+2HUESGJeqWhh78jT9uiV1C7kuC0hba0w44/eauYy7XcDk
hxJoN1HxHkzKMHOwsiyLiBYIFYHibU8YGRdk38rB4TzuNoOOQ1nngEuTF96mz4WJ1x3qCibxJM6M
UM95Z2YbBgSil1sB+0tx8m2gHzArWzan5eVl57U8Ig6OcrtB0/vHfOPlBfLVx9dV1upYZR6swMKO
J9MWDiG9w3XGjIWXu+u2O7bg7eBQyefryc29ARXIqKCk0yObLXi5V/HFkVgG6oEpqHMstU1Kwt7i
oJbtddOYxix297pWjnQuHGiipKGFNn1tJJqPE8+1vIXmXnRxaCySy0lb8lpC3K6YJO88xZajN41A
6H59WzyefSeqlDIDk5dbPsdP/jtN9u3rY/avk5nr6w0C2yUloqQBjZzQvIJoJEODhRRiXBCEwFLx
QZKI0IxNGp5KW+jmPTIIKca4UyQb23jG0sUDoZ30FVKXoDNG8zTiSECLLLW/j4RMM3eQArYFt1X1
TjpcrvVaYYScOFBPjaxdyxT3W4hbd1CkAI/wlgo1QkwzMa4xGFYHGu9PLpjkIMRFKmt6Ir0k2kw7
HM7a5a/17w0h18E/+xnjula7Dzp9zAwK3lczxyVU9ch3prcd0uuO0ofExNnVWMMX3WxHWbCyS0Ge
p2nuIAf8ncYui/Ou6PRYfopXoQg0QBKuyRt3QoeABlfuj9oWr12Urqgha3b54JItM6f9D+0TWEee
iZSwj0xZ2iqY8lRWMB08Jw8K2cZyV958a4C+2RmUhkHxbxAoiL4NwtSF33O4RxLk56st1daV/ymM
KznhJBwUgZUv4/z4mF1XLITorvdtlsCO2iVyjqKR/DJuxJUkri6VwNzH5NkNQXzmuO0/rQO4ix0r
eOy8tpbwecx7hTjf90OOWKRaqQdCC/CLDwXxP6kXIY14y3IEESg/GwgQY8gn8JtMPHyz+cvcfv3a
g+ODvs/7WYGrvr9b20hSu6Mgw1iN0oi0xYN1aRl58guHs7LWIEuQFs9IsxxeumthbKcedzaMcFyH
rVLOgRJG+XILyKLdMlvdz2a10xr3BHa0S3cZRgvuJfFvMhruRcr+gUVg0ZEQVXntF1cLHezI+Sc2
fH+Dt/BLUJ1RsbkpR/BkfTY8NdGoO4zZ1PmZURMyZxNd+OWcel268oaHBY24klcPqZGOtGxUD1xa
KoPI5O5m2q/kDKu5cGxRTeaDasnhNpC4iClBtT9HOt4/d443UqyZCuJYr3OwASjBFCZmGNU8HBcs
kMgknU/86IIoB1ev6JRDMXrIhJ1wZPrnQeDmdBnYNz3HI0rKmEt2YeWuHBUfMwmf0f3VEa8ApQ9O
l1nBZb44Zd3QJRtEEq8ke8niWGRDBKCdzegf9m1HLtOEV8PZnbp13gwXr+4kw9pyAtYXfVbtUq4J
TyuHu0iYe1AZt3kum6MpTRQLxAzXDMUTqLs/xFvi8EEd4OgTMPY75IrdzUgwY/9WTlCApTmlRVxw
4eWkRXLgfJJzHJJQnj8xDLOAKXpHZvB/QkOW0CkuNnjPwbNaXbuUazZpsE7d+HaZzPyZ7XtnZky6
lW+9A57gGyWK8slmVACsEciXbES7/IcldNVhbkPF9NCn4W/vSl511tANH5NP7XjIwcsZgsfMjdry
Kwjl+FEMIbioSOPo9nkVhrnN3C9SWLYqp2P8K8sFwW83hsdNhQiMPVRu5CnlQYF9XhOhG9fPbTtz
/4rhXq5mMBDA6d/uBLOJaYXeOnumCc11obHm5UUMzNrEo/k7y8NtqBTqUZJK1IPfPOm3YUx+1oa0
4+o05uf59UPBx9bPyPpwmSGWqwiy9WSRr9so9SAaUQe2DrKAedB2BP1HdS2DkzHAMY3xtC/lx1su
Nm0Rl0MEYzjT+blRJm8Pgxrsvgogqt2WjY0US0KTNYCU6e7KNPXNCqubzZ+koHkzNs8Q5Fqfa6D9
+ylfSyKrLP7+8iFKdu3R82bxwawftkTVjKSMpJjPg16gYyBOtrfG99DzEdFCSqpWI7/nkiz6YLO1
fahIEr8+Juhy4+Js8z+SLXAgPcN/mPiJEj4E545e/mes76yuX8DitHu9I4UmBOSVS9dqsU9i2pfW
kKOMFB80X1g2LKNxjDwDsvFR/CDLLWZYv6oSLiG4OfhzJKmM2/7ANJFoqa9AruOBeg+Ul95Y/4yw
SjF01qaRUdRoJQP3hmJquUyIw5Ri/zGKJfQ8jobq4Z+RODb5ENC5e/iCJyAUB8xg5XDbfxm1OZh+
cLCLKNBS9YReL2HL6wjnb4DdAyyhWFrbIWTzNkVaI32/iMUWJuTQOOu5FtFF6/WHGyLRgEfeRZ+W
aG0Kd/KDvBRLuLVuVmOdavpWlD6avRT+vZ+4EjtPM7cLZQEeXlP4VrR3F4GPlsca8a5uWrmhb2K1
VxVaBqlkPqd1iX2e4YDRVkoEwYULvbj1gp0DbiF+JbORUeKT5b/aOiZ/QSdba1opnY2DaGSxvL4y
JEEefGAYgB0OZFDY4fnmj9+peVcE6qKHRm82zquoAeFEYoBHn6DxnIryIdc2xj8zfgc6G8XRNufw
7M2iwybFXt8YLD9q9WYKOTHAs/Vdks5ycClrHE3+2boJsG439GTYExiuhpigGH4MziySy0I4f7qw
+dj2LIAD2x5SsBFW4nFhMwXYWL2hS4qOung77VttgPsb8YCR3EHlOcQTui9hU2Dj9UyDcch5RaHt
11gZIdujhAPKDgqrdsXpBE907ZIuTEBUv9Kf95TH9Ef7vy/aXa0oLj19hREoNsHEvsetIqwlZzBt
wijQ2OL4MZtZKS66Y4jooF9tJ9Cd/7h0EO3taGVmQqjQTu55UJjZ68p7Pp0x+zgTJsbqzMff9gN6
/iYGHpIVANiRcegaheuy5xvgEa02DvjQKIsektzyE8Gu3ISL1+j4N7FJ2BzwrWqvtH9TygTykM9N
p+9gYAZKAr/HY1JOdXIHnvw2lC+JmYRqtV5UPMBHWZ0cgE1HClH6iAJql6g85Dd6SOlZExWCrUhM
Q0ly+k6CdY9TfDYb0XKmdjAimSdbR6eEGCmidmv1Ljtjo4bvTdXfRfb1+MsDVb3aQTwEVF3Ij+8h
xKrRAOK9OXfe+2RmcOckSrH23Kl+giL67LNT1W+i6SbyluAwImi1HNSievkjXo+ZceFbgFTCu3Sg
sHVQi2CHa99yNtW9cjUNhY+SixCiks+7+V6dVhaQbZnetzX9c8MgrNmq3ROTey/b2G9O6hMn80ao
6uzOjgY4tvK+yJ9BfAstmfIHkP8EO7/me658rKkiRcFbEakgIuf+ExiHuNks5XoDdi+dmKJHVzaV
4JVlKPkBpenihK5EKVFkRs8R/KIDYUK/7Hcq6xdQ0hqoZdCnSExM+uE/GWY1JWpUD9dvp9VGQf0Z
4N0PalRXf7WNjiQ4dMlVIcMGDp8dC0qNWbkx71R+cenrj2AY4Zo/Vr2Nwbqnrg/i3zqyP7FsFRUH
hL2tLLOu9+GRzZL4w8wPRYFJBHdPXm4DR6fEUoDxeUZO3lwK0JtiKIGeFrQD/AK/flGzPw5QI0I4
tb9x4Ios8x/M8UIbqdRbEUcz+MctMHRKfNshykjLmR7JnzLV9sLmezjVTCKdl/0KVYk3OiahohAe
tn8F/LnN/OlW/NyWKnaJufRWIodzJJRTjCVPrdfCCdKTAQu1lU2aF+z+MT9FJo1xxg+ynPtrX7IN
DLR0z6VsX5yROUIZ+bCaFYLOjsBD5E/KfIddTYo4++FoqfhIJGsBFoLh3iasuOTEbOolL/IZY66c
PbN2WPPwmGB+MOKYwMdZWcMQRzqIcbR5/FyN5xtYOaAEQb5i8C75+tW/ZhZ1SwLjjLZECf3zH5Lj
w8dogX5YLLKSg1x9YuIWWiFmJ0GUNu5kO7AH0bTknmf1ejbt7rEMxXsl3YtDbFjDx+JP+UQ90K2O
c5NZWHjX4x8HegSe+fyN+Jfvo2cNfjF5jEcEAxLHa1I1y5ZdTip0F/cnaxC7nlUa6zKckOl+X8tg
xsez24GcLCMZZR3NiqLmU8693A5xhuurzafJqzs7Ey/EQPIAbH3565TX0npOUr54M5nbIoqzjF9Z
Ig+f7Q3f8HPqb+0QnZchTxTqQpTsf0Q2H/0CwEzlpaOYQbLMuEYD6OpOIKvGmSo4K+FqX9bPUqo8
BKVRELklDAqvHY/ggCwzcmVZsEzQmZVZ0XZBL+X4M/WNqzRFVOv2OrJx9ruktcgJwNYdg9qpx3t+
HiXztvR8QH41Ab8/PcYHyJ6tatRdX9Ho0lH5Reo56+ld3I18VDFRQOg3vfPr5QQD5NvU2cplwumu
rUDyySvQBJKvYpInoXUVrZJDpg3SGcOF+9ZBQvmS8AbtAvZ3KjjqPYqbmsTlS9QG3b6iY9wWHlL2
DjoI4rQkVBLyckqqmT9yBXAZgQcSNB1kXbCQPCZzPta9crNZpKkcA0ljMDb7na6vgotCsZHnKPNb
kZy8SG1H3P9LAtmXkhJSb90YLQBAZYSAQ6uBBw2whGYLkU+1NLuI0848ALeyeLs90hgI2HsFcYAg
yA0nrxe6m4EcuvZ/scgbAlMFQpKRHDIRktp0x3nLtfDkK9zO6VdxcWZpWVOJnkhKszc+nkV5Nt5A
esD40FquJL+4B+RaYG4ULaaH5sSm0qVeqUf+kTjN2WZkVk9XVA7xcTcTw4rsmVAAMmfGyopEYyza
Ba+EVU036qu07D1ieO8k3cczrkd5I7KHO+jAtdhh/If1qBjvznVNrbTxvNTEOVsLmBDRfrC6dBim
4SYXj9GmpuFLtWvCK4nxkPcjDXgORZT9ADyY9kNwJO485Eq1/A4ytROhtMtT0yfa0dmHDfV7MbmZ
+V0FY8dLHOgxu8Kz3s0sKKilvaoQ+Hqpt/oIVCPjdam/tQI54R2jcwllM56pR/H7gsuh+w8196If
v8r34YVRJpP7VXUuJkC4F6Em0cozU8mf+2jSNEOj6+qYzvbt8QMYxkiFgy1YqwCfvXxXUNjbjDqi
MffJbm1lj6SQoh6aq/BiNuIrgdMx92hsohzzjQlpG4OK5PPADd2y2vdGjpdRpqBf687vtdR0w+TU
7pxBu/bufeRDTGcHhVzgvPa0OPZUj28p5N+REsAnSG+dkZhRffHikUKUhvUFyocxMCAaSIPQvmSs
HpvoiLFl4VAjnMr3PcS3+D8k9KKcFDHYPUDM6jOIs/Shs8Cjbpv2AXWOkbOHwOZ/YBvOrztL7bXk
w/aaK/oy3khpU3CRU3Lpx/n7KfVThuXmcM5soxMCvti/dmAA74lbbf9TPgh+mZRZ985pwqSroGy6
Qt5tWuglmC104vK24EM0gehPNvvFdnORWwbmIVsFIt6n9O6aby7HDvfkDhD2btuj3tDg6Fs6Ks34
ObWhEFTI8huqSCVwC0ITxeyQ8s5hwEo9g3ZWHVVroLCfSEY5mOOq2sQaXpdS6WLEudmi2VNrlviC
RM/sDYLq2KXG2vgk22Pn3XQgzhnRqq0HIECGivqet+3gDca8oO7bHd+1z2R7mJGZo8aHQm/qLMbb
4lMXU5XJS13Pm06yPuf6X1fkvuLUkrtZpZf1ePoVQRBP6jRSv3ZX75mdueGTEP6YcpU8EeSFCfj/
FEEI7zj5WUQnUi19bzfzxcWatBDc3Tig/JKfNfg2CXx3fFTrfdDQIDEj7Xw0ZKltWTQgBqjtgbPn
jamffyU4M+WvyKAinRvvN02JUeLApeL63p3FPMW6y4GekGq34gIS6SPeO/oBdgXq7ay3+FhnV9ia
36oQfLxr2B91HnCKDLnZgsvcrKJsoVv8NJpfssqIIGGOgt3dpXP9ui3x4L+KpdVDTc63YG/aF6md
XnLi+LlPQZMgijSMD9w1+kEPB4A6Ffrs/uPU/DJ4mo0aevCS7tFV1E3ndcXdrewX/vG280zxTbuJ
Fyw4HYSzMDiesKaJ+t3bbBqurJHhacHxUq4DO+QK1WR5If0Gzo2FkdsrbkQRGCtvDVkaYQhoj21C
XEIHvbCFa1iY1RGOaZDGA3p5NiWcbCBbzCf/i/9DF6RRGUghpe/vv2NDDXrSblHvpiH4ElnMvbbF
+vdu3gHbojJ8k4kmn+pPk2eBAa+JkOZrYkw/yojdXoMEQ+6d4F79eWb5Z8hkc60Fta9s5/Vf2BQR
x96u3ejm9a2dfrtLZ/zmve6KLOsbhkuBw+LGkPoIzgiK+udZUnhrCtOBD/R0J8aF9n3uR1teE0Nv
wHfzusUJ61jFKcF56fnmVY1/RvRvzNixGprdtfW4Ot9ps3XcSUJDfJblpF+cvKtmkB8TuSYvTqWS
L0x/pF3eLMTxTGBmZxYvT/rHm+plFIWNdDThpfs1LQl/7nXcWUPqr1ibZ8RdZzviclfKTwFQtNdK
A32zvwBtQfUf8+h3Yt68amXK3DV56C/cAgCXfbwcPbrAqy7cOjIxRCKXlFP8MEQdtgKgGrBrRpcX
FCvk2XzittxQnxvMLlcjJ9zaME9uWnPzKAXMJ86rNW/MLKnjvOinDCXKrGhj1X4FY74lzPRN/cVA
zXwIj2342x4gBhNyZTtHP9FapB0FnF8m+kiTbY9WajFm63S9Lup99zyKVkLT/MzQjJY6QCfep1Jv
jEafT/e2Jg+Qz+QWgHo4o3dp1lEJ738Jt+GO5ZaDnFCtdyM3/24ENCObqqxt0XEkffwQrevmq8F+
wRlnTRaZLmYw6uNacaU5s13AAQ36t8i7rD6/eYeARXRXP8KFjne2MORHT13tzA8rvaQrqvJNrHlV
5E/qEGY2DmWhy+cQ70YsdfY/jfbNmSX9ISVeZRPLo+CIxo11AdGO0+QblPG3ob38NCsWOopKGOEb
TlxVJvWZixUrQaCR3NLU/0j+TWWxRxqDv3gMkZEoZyLByXSoSUI4FHfJJgCL3LZ/64lmtmIn39Mh
Q8kg/JqC1QddH09QKdrMO76kPaou4yMh4xrEI/vKBtnDx6fnJ2hLUtdHQFvd4hj0GIWzrvQoXv+5
CGgC+9hcBlALShJAGWJggmeclsXwQCxkyRxlef54e3dhdnI1J50IfqFeYNMiGZBUqv4dvt5TTcRV
Pru7cF7d+zHGXp1wMXjeR8Ga+8LD3gA6yDGN6SgoCka2BTptxk/ro/IJjez5tyPTkfKr1KxWmOT7
xCCZKP+U4ms6Pa6Q62Mt5w/xubavIOZP29jfVZzKtzjxyAs517c7NOWvrf9NOV/Ea4nTFKVyzW7T
ybS1bM+5QegntLudF+25BNCZIdQ6lI7I4PM1C3nweOwJ9TwZJ3K69DfpjMZj0Q2dfULH7hW7NjJ1
iP8rg8P5mbZJPNn/GDxx3MH22WhSLWfc9XiQuRAS3QYKGvqVGCoelYSvRU3FiGfAmJCTr+s2RgND
0oiSP6dHmpK3d7sMd4yMK5GTNHmAK1ZBVHoBxd3t1ARtK9Az2iy+KcK9hSJWQaQDWohosyrMeEZI
8NGE5KpT1u7SOFoKkCSARnu/PsERmOwdzHWNN+WBkVawzP09CGgM0vdpHMAdcjfIliiEntCORL+q
3fRvG0N0WN1xBkQZcttQkwJ3Nel6d8d5ANyoQKomqahudKi31bdKYbkx1fxfzHE5JYJ0mh+95sDV
Yio1UR33n3bYkDMmnf+OOLIgpRgz0PUmz/pI70r1UwCAKeQtBaBKSqKPlwdLQufyDkHSqCbbZ1VG
KhS+1biYuoj9BJ25sir/13f3jm7NpWAtIKy7+Bt6TpivUHcEARxxKK9WJcEW+X8oOtL00lsyYFdq
eGTUYGD5Oqdw9klbVtuofBN3zbu9PPXQDNOZ3S30LNR7FLpCHQjkFDCRlsmVAdtyUqXHf1XOMPDm
/qIZvMPJ01KP+5GBFm4oE8DqrHM3Hg5MmBruOCInH3/ABVtWzr/JZuoddWeIwZrQIgWygf+3T3Y5
vJYt/UB7SZdB2t1Qg2Tvl+JQcEkCNd/RuhJEaMsHJUVyjCansAyx7z8sljDJyEKRXQNsm+kMYkBv
xl1eSH/hy9E+H14AO8Vj8qMjeVo4l+EDnR6KUwUsgtDSX8JIW/iE/aFl3IuA/mKsFlZPio3HSTwb
zzlqgz0gqB2G0JG14BAjOvDZXw4g6xF1l43MdtMQJHgahhmLVNPVfT5GRcwM1RIRr+lV5jUF75Vw
pfy9VSanZ6jQaidZJQGbas7E5JlkH6kAq0dnFpaFmXVkJAyiPN20uSVEyRFnquhtcMyexdNCe3Cb
AOy5RxxtD1r2fNr0CafECPohJhtWMLbkfIlf1eE9U9l11/06sC5WUyULUBnygqrD0O8wZZLuHYiT
BeSxAhEof684z/o/oSTBBZB3v22XOXz9fMuKurDfcDbeNGOYuRp0JyuYM4aI7chNXRhINLTAyY0g
02sydlfapl1XRX9udv0gg/cpM3TASgAjTkJNEdrJxLwEUtvtJQtifWr7IYM6pdMRCvSE4+FOSmaV
6dBmMGBhWHBbuL2ocn+x33Ie4KndMhDOA88jUReA8fVuo2SgzcsTfb07lwI9sz2ABqMTZdd3Pp5i
+oJ+zKVS2T2R3qOYSqZJPo1GkrtBV9V8gCVbTA0OIAxjU47uCAS8QCS3OQVljDmX47LJUdWAQq4B
9hI3uFByuOLMQrDeIYtcsH4LgDwUR95aiyEyp+ufjjKsQw7w7Q5PFNAOSda5vzEZ/OtWI47J0Lxy
tNE1v1eOSJ53vI1koU02wy74Nh9EMZA2YXURgNv6BMwNTmkLbbPgMbeapnaEJ6epLKlMFm1harCu
Z7nlloUxrXcipEUjwXXWe5m6+qcxTK4DiipkgwwBuWBiJUlMnW3vvtcISrRatuRRIWxWFH3cx2eP
EJnk7QaVQFVbQUpjmxTExQ2Pcy6MFUCQXZ7mPORhXqM5y9ftodwZOoRZ7R14tJv5S2A3+kS/3rYX
5l9O/+YPriSDAd4TuERe+yXSJL1emHp2BHExRNOcgtLSvAHr0XXVyG4YAqWNAyDpOpRDRlFK2Emo
uWL2gRuRBqWNcggp8BsX4oapLDiFSS7m+j9gusU9SfJ6D8tkNcHENDvUfjwHAz4qjAsKGBLHZlAc
Qfa+xxOuJLYWTPUdc5xAFydbpnNdgiZm/r6UiRNyb1pTX4qOQpPdmgxfhDLdK+zHHIO2aHIX92X4
9kK9+rzvgUtd57fDDMx4VRZJhRJFzEfk+IzIertHa6z+h2Ri5ZKMSirOOTEh5ADNf/Iyz3g0pxJk
mt4BqCp7rGAH5/7+YY4zf6iEPKOn6XRNnAGJHJI7f+2L0+zeU1otYrkLSZsuuU7wcUJUurAwQ/0E
cAxhdODYST5duXy+ZIX1pnq5NghvJS+uCeHEufPoiZ2YKH0vS7cX08dRhOENUKrNjOQUW15kFNxx
17VYkIGbuBg/67IVUnW4IHq5BA419/6W9hjUnks+mhPL8H90T5WHmTjpC4NcZazHZR32lwjQLpc9
pLCaulTilAsE5xadfYV+H6TUSzSbNfE+AxbY6Zt3SAa3NczSmMB7uAM6wam42fHiWtz6auTnjStm
sKqHpldpegllt84AuUHSko3Ghtp+g+hReyXX500SqySL/VufmrrYVJdEg74z5k0PbUG5tIqZBc1A
gTUscErP1MXPxP07CmZ6Nbis6pfsZ7Kr/OnnNmfhk8lBy8sJlIjSh95WFWbZ2tMxO0g2+IIAvZHx
N+9Cnp81L5d4mYbZL6bNQEAg9FEyQipBE4JrzEZGp3m3QNQpF4q2fDoyIEzCH4GRyjLkIRo77v00
F6tJ9qXDBdSd6MvuTjRcsTTPzBpZP0iHVu7KnNPrpmkSN9GjFJ1ko59SWGfIFkFF+TyeBiy9xFj7
wiNcbeoJLr0kKNOeiWyjstbyqwRGU1nnroBHPs1KehxZF/ooeB/kGp8Igfmd9sS0947f59qpiied
puZiHwImZKAI6+CEGv1KSi5/7oq/E62IGcJiACwAgmrk6RvRU3r9N2hsfUyphp+nxytUY+Qx+N5K
H1oCZ49mWNYTXS9QzdCavL4DBZ1LiDweAwZ/FX4yA0KTjp+TNIRX5NcBohZ/A9fyGWBJ3dmlZ+Ic
0Q3/oHM+ggNBv2H2NcF/ltr4d1LIyM2l9ooCD8PjDXecnQLMqlzdyk53rLBpvo29cjHtAoJlYZ55
/4oIvWyrjeNGWQ8awghh5OiGm7DKWkjeqp7PhXjuAN0SLv6720aWDe9zepMll3/gLmXyiUgzDiGK
7SiGhVQ2UqPUWB2PwfWC/+VFla3K5/iOKNDqCe8kOF/QIe+w7Mo5yL1FtWpNFjCTJVtAIgKqRQ1X
GfDGKGinXG6HiW5O/tccnJJV/msmwkrSpkG40yZw42RIWlZqH0rbUMczxnseKDjNnLp2I09K71Mx
PKyOlG/UZxz5zljlHjVZwT7dL7n3l1uyGzABO4/HLu9gae/K/6vgWTc3BbeQS8ZlxM8s8MHWfAxN
5vrqNU1xHQlyF2F27A2F3DAdhEIQO8VmrPDPjXR0UMGzOHtVXeckFlRciVulnA6gxo4TpGG9BJIa
3tv/amXCr5jsCTZSXerj0Cf/NUgC7p/vJeZOX5C1GUNHsF3sw18i509n85bA/yYc2cX7zBabtzJK
HJDdNazQSL0iWWFokeTJKn61hAwjcKUBFhacwYFd0WgSsrT4RUL+tm3gfX+muFOlzSYz8dgxVo7c
vbScqtatwGBN/rOi3D+g857kWHbGkeCeInOF+UgN62DjEFcqKgVRXIjoeGagJ3JAJDmWY/9y/BMx
BUKuSX3KEnjTwYNbMmfWCO1RTT9yc8CVpxqSNnEaFyqH62zjwkB2YnmIkUerOUaupUrYufREdWWl
2e0gSopKVwrtS51zU3urz1s8b8pQ9/kae/MedyGUbZ2RymnHFddQmOcnIe3pZIIzA4fMl84djUEi
a5CzI66M/RIclCfqnWZ4o9QX764HPBQRbpLfOAJdZzAhlfs5TFPBfBOLsslhu/DIi6oIwL+a6TNz
V5ihO9UIeYHlFSH6FPQmSHhBrF6n5pTQoOaoaR67EPL4tyEJJyKLbuFpoGmhgeyDlP6/0Tg3hfqE
bmdSXfACAgQ4TUIVEG0cd33kC7+WNImT8CErsUPyFlim2y0a9WNSiK+KmHFI5aEJfb6U72B5FU7B
MtHdbIarK/tHTb85tbAjl2ZqOZaSrhNRyN95j+1DfnkvtvNrRznhwjTMlifPX0Abjuo84LCUZpKe
ZC5tIEfkOrKikHb++aU7vL5hCnviWZ3/UO+xzfHefQdMb2VA/l90+RzOwUdQGq2vbLUrBEg1OLKg
djnaTRc98dCtzp+mSXwRhlbq3Obz2ekRawaSpjiYnBRSdhEVHPL+cChd5BGjVNeVDobdbc4Lzi7a
NnsPsMQDcHIkjacZphB3pc/ixiLGk43WUz/oTjbecGwsznmmp89nG0fNsuW3SkyNtSH+Kk/8gb8i
v9DuEsDqprMTHubDJESJ0C5ozmJCbtc55n4jMeaf2ADuGDmRhx9UzTQ298vkIGvs4G9TLR7TbFpC
eaT3l5BxsOkD9s4SNdkeQ4hiMivJapQKQVDySv8qq9y9qZwZ5D1qiGaVEClvhSP9IuZY59+7NXyO
a+rvYcNB5EQaITUjV6y4vymqEe7a5Qn87FqVcNHmwuPY7nc+UTCFjuFA+HBCqT9CDDwiC6ncmr1F
M3vdf6yMUrz9DADfrFN3b2fsSYkx70ZR2w94TZnaSv5Nqmm08rFGccimPwuXurIAyAX2ZLY6+OsC
w30KOUsiuBjZkuEzP+5HnvRnYf5RiAW4nM3FHMvIrYmqMw1NaK6pbbiojcbkNxZuu5kWTjPQ92jV
mFZF39l5fHhuJv7nttVi6Ihp3nQVVsPIKQDaWcpowHqRw3UrkQQOIN5vMjT5wzk54Tn/aIYwxEoQ
9D2sWL/x7Qr6vBR3srKsFEGWtaBzLtsxyQqAluLlptzhTCcGmg1XChSrceAz0wevgQLD1zrrvS+k
bsUut5lyXQVpFUS10KFM9r1ti9d/4EGR3JB4ADcjA9TZv9ruDVAqlhFzhbnScU3akhnwv8+oG40e
4x9x0AZqSOcLURijQ6mydeCu2NKwSxqFew+SbI2T50ZqrUlMcImsIjfXHWTZBE2865RMz3HMv1uy
M1+88fkpN/2TSYWgM4idEh55B2LrpKE2SrIfkTYQYKmCMA9H0FZGMgNM6DpnzR50JA1h2RHLnMNq
nH0+qn9HKO7tJyFRmU+XgA3C5SuJVO/FnNKnut8Qul/hI2UJiXfyWmI2sxDiax2NjSZkG4YOwOD6
3/zlaGwzrcWe0yETRjDew60XXu/XZ1ONYFWAU36oBeIS+NzAdK9vxs0olk7f+iQi6OAhrxNQzv0S
Qb3wxiHIFSzngIzlRbflcYwX5Bfg60W22oQ1d/E8Nm8nLAEP89PxeWsi4wIAy3FBhK3rsapB3B5j
EEPHElQCH38IxatnIXuPxTizgYdPHpLNjvyfv/lDHPsgJdjcY6o52chAe3ISXyP/qecuUlaGgRoD
OW1KMPVo0ETy3GwUrkq2711FxcilFtTjiX+7lybOR1nRSDUero1W580FgFAPZ5XRW5a464UrOazO
jrFWnLtRk02bl4eqjG3bTVbF8SBUhWqTbhoc7ICf90FsktNHKPjuNcLfLnwsS7XvM6RsudVnQ4DN
i6zuAzx2YyboSR31FDwEq9GGc25+PPpzveLq5+EfcBWGELKzKgA3QHu577XLb48oMoLwrdaT0IFz
jOcQUge8rqBPtggn9S9gzy2O03EeM5uyog9/e/AKi3riIbGM+NR0cb8T8BN0oZjhPXBpH55YYtP9
UT4kJsWXxWan+uiJiM931KhHzyZYoQGXb1OZTncaVdiNUyA3tp9X0cBIF++hDEbpsEgNX28+qHi5
Tw3mEOaRw3FtxT3+ZYOvj73/Tpig9iUL8jQn9b97U2jlPRCScjEuPOeY9TaAVQHSCVIVaQlE3PYx
O80IS9egDKER/sdX/c1UVZNBeXYP6TCsEKLrWhM0/q9yOQYX/7TWrLPN0DbLknfBmzNNlXM9+Gn+
D0T0TXgMLEwKEYVd6I/Fmomh+mwOITvDOztrhy1gQy7z5CUKsMWAkNU/Ej9znB3USfA4leR1V+9J
D0JxdyJM0QRWUZtetw7ggCnYo7LTT/NXXUIc0EynqN5SU6BqS8r2+YJnl1xFB3IkBY9Asr80//9V
y955SCbj8FPQHtcUyuv7vG9xpSH8oyCb0SpzXyMC8hawnn4Q97zjXeLhTF0v5hzqGghCztxyy6v6
rUvZxJHqMX8yONJlE7oI2QHNZlthonPzyK7O3hzbXmLNuq53tich3sJX7nkuCFAGyFhDKsQHczzf
hQ3jWa+kZ+lt034byshjEOWXLI5VbDdEBbRJLnBLsScjqnNWWKCvbTxqbt3m4FRw/rz9CLTU3lLS
hIgK71WlToIFwzfv+ynpQshslYkhuGZvbxgpVR37J1eS5wTRXSKI54c2tM7D5ew2A8N3uy43DzMW
QJTWx0Z527dpbgKRMXfH2bJhccU6Sr49tQTjFLW9GzD/Eu8w3TfqAMB+i7STzZUZNSDP4ZOTf72z
XWXGtNogxGFk/wss6V2R3sUaddM8etafCW24vivNyWSQHHMb29RM65V6aXWiQvcnMlxHxWqT0vU7
q77Y1FsIlOrmSy8ZiImm5yyAg+3I4JH4N9iJ0CoNI3p7ixYAJtDDlwPMZMgTj1MJv5GmCDtAp1Xi
koDcARF5oQoarhs73sxfVFVJWlD4WBfV6NVgrAi+IfdaiDEERw+TnQwH1CXKH389ENf+fMObH061
IAe6W2ehGUVdt1ONoMZgrzyhpZLLBODxnEH/sbBPi3YaAibX6oXmiKl0BC6taWqhUN6Crm5ckJBH
AGd6TzBITy06k0ST7mSmLc9j6UT7N4St7A7yxxkTphGJ5FhRTaDAvtGENYIYUYjgQW2fImvNwOY7
xTU6+mpchIsHBPjUNm7Pok02UdadGPf3LE8fS2x4NFeRHl12hkcyKRecMFfPQ/yfHb/qUuRmH8sX
wmUdEgJimqj2sAP5u+QErT4g46AdljggqufbZj+hx4d0NLVn82WKVzrj2gaZLuL1/8fFGP4gsf/e
xSVRrzN8H4R1/pb70C9JfXa/KJxUjhx2UlVe2FaHM27DOkcKZqstVTUWYXt1s9o9rTqvPFIiHQQP
qqtS/5xw3USANhoSgS3JCLD3xWH8lS9kuiEjI/9QZViScA3QO/yojZMoK5CpyOwYjudXceg1s7sx
q3gEfU5ga6t8T7lVP9X20EXUVhMTcNetHe1yJ8mPOZXUoR1pHvjnRueM0m2+qfoplncV/fPJtpg+
sfIs4e9yzI8a6SaD0Y/d6/Qe5UZynqtktyDx69/EVNUAHYR5fsn9qlIM3trwzPAqq9wsFxPCwBkk
Vv7rjsAAed/ifOLjKYsjOjJHKXg1VFa3s/aARfEosK+IAUgLw/+UOQxbc+VBitNh1987tg+cuGIi
WZhgAqvDVxTa5FFYQ+gpkKdz/YEMwzzBXFvn+vnJpdaZK/Cj1DCEC/lwd+kL7VBJtrioaQjoD8zJ
2pdGMjNDthqj9NwOs+yIBo+n7bCyJKPPqBwy8xD6toJTDPcLGWyi99SG4mfbzsLo+BKut92Jl2Uw
qjfb8l8oA2eqGQOBPhsx0foeewpmAkEVwK8fYYBvSPg048fOwKl5aaW26lG28ay792f4IKqtEDI+
Y2b4ZV+mY2lbAuu4AKwkum0td5K11g4QRJVDdxMXo6lnt2fkvTb2xd+O7TFwo31vfVyBXvpxecyE
WlrVN/aa/3zZf7Ndh6HiN7HGQeTznwMD1aWLquZ6ZlrT0YbuNkNDeLArm8S6ypwrwmobKz1GruLX
l3PiUS2ogm4fWP7YNLmN+ItId3s/oKI/1gvACX1Wxr90q9h6QjEfXQrkS5O/YJjAWavl40C9dzYX
kC/1smSi6POO5fmztQw/6B2BdrAW+U3ZDUn+DavmYN9R59sbqpUSlrTdZS86oWqpTLeSxnYCxwDM
AL/07hB3owjzTNH3wD9CLfAQbHSFV8sr+LmNmZPvB+K3KO0XSgUIfDglqaqpD5bU3aWTpLOBgUIG
4HigBQnSG1VG5MiAybJOVgghV2iLVIlKqstTY7cyZBTNitKj0xGgK9i37H0Vw4BHwkc4UcUn3vyB
i7gBV0yEU+SPb1N1PMI+AY8Nwo8Y0GrNaxLhikwCLF03ftXcoorZ6c0NM4nBS3KOINLGJQeEJNDC
nLrPRt0ItbFZFSdJt8FmyuS0rjb3N/XpYwn7KV9mA1jTUXB4UHpB/9t0lh4HlV//8MA9WKF30JHh
D0acwyv5HiUfFX1nuANsMvx6iL34+sqqO7bKQ1PPTOqeye30yBmo2rjJ3zQPeUW0H28DECZSS2QD
urk+7W3flqGHXvJSHm9/W/u537Q1Xnn0BjsUBHpBG5YcK3HEcXSEa/+hJsHP/UMaXRpks5tU3k/5
ZMGFDeYXM0ZafToFbC7G+BbaZAl31p/d8mQKJWCOfgCMbFMQ6+4qNmyVSJDHvdpbV5ctjsPu+32p
Tn3OCXsGG0qJ94ETpWoUe8qPwwPeemddmXwgjS+tEsjCNPwylcG1Yl7sqTQgSctysEtIt4Ajeb6e
45xXBfauYW3JxW5I/i7pU8rgLZ+d3dpfE5a8fvzj6AXhu5n0t1NgqCwJNzj5R5fgiWhrr6gdVgrX
GLTiBENdcFtlBduzw4fkoDSfUBYwaQ0Vq4aI4LGI15EwoD97OHEjZPO0iwzsx3qRWgpYP6dGmn0I
LbE3HBjyXlKdJPUE1aZpPM1usjkzrxkwJ81BbNDd6o5pIANTLkzZ1WETf47v9fGUvr1jyZSItWeU
lnzLM1KxpcTcGQYfapbZoLeKtxCdM11ZDcgiJrd1qi7qckWE1up2yjPUFXR/04A92vYBbcTIXkkx
epIU7CWLiRLW7JnvX77G1PjPtwX9GjRr7tavI3hHnwe2aIUZR3QiLklyea1gS3Kgecw4pvUTgRcZ
txJwI60gZoXaMA8QygK1EQBKpUwfizaTKG1S1JdKJHVXBNUTKxA0tlYG/PodzKWhp7NCYnipD8Sw
aAbayIDrXG1g196r2EWu9T9xvq8Q6sh9VzN4eGWlVQ+WVoIc9Auzq3fQCs4PZM3evL3LnSBpw5tX
xeKU0RJNSJkDtVVE9yORiFE+IoPrFpGEGVdJaLYO6xXZO27mcKtDJ6+MwAZeB13n2I+os7Sj26cL
sSR3HpYmnLJvPHzxez+5L7hGhw+iZBQUvmWj3GMB3sgO7Wl1tmGjy4KU6F0xWQOZkuuLjhgnDwl2
ulZD4Kn+TbJvY0WHZXjvVRUxneobMC8yysJKr0GQx9CP1lbHDt07TC/U5Gw2n9SYRGfsfyst+IAZ
wD9X9Jdn6AWAju0O1RYGFx0xLkPVOXPgbm6ghANEHuvOoN3u41Pjn1LUs5DcOfisT0UFJcQBxj1E
C/iL48pA2PJb5sDsrkfDsvSdlq0FllD2894tgHNds4ZgFDyXs8BFrSMTAlXnMv37so42BnEG0QoT
CV7QDZKkQNspVMWFyJweoO9aW2Q+71NwaaCyPbALB1eaDwt8vtXsPmpCx+i/O547jnj/YhvZQwSs
tEOgoqpFAXmTX6A8bo4JAlcTmc5vtmZhJ6VQbjPIRautqyff/bmjw9aUc53EioEcdHK7ZQa8J6SV
+3tyIPD2Etvgq1LeKzGUEFwsYUqpV0YTLSk5PaEj7npzP6gTfcEULC2vTQpQHvijOqiq6shIuoMo
JQu0Ixy8U9ZqFBjJE+gjtxo7/iDHHDNtAXNTwq5BXL6KMsJ4z42u8dWgyi++H4GkoxdlrZOZ6DDV
58tBksxfo4C/OSv2DAad6DRwup5R65PQ+p4DFOnMcuDtCLaSOKEoc2pGIEkxHXnYY7vqk2rEXawp
17L+LEHF340W/UwEssu2CwsPGh1/a8sjHSc3cQiwwmdMiz5HDVAZJFwB21Neu3xRj59VpMGEh2Yj
dZ8saArZk3BJZoFflDi352fWGSkdhXPbQsi4B4J9lFVtVCYjypcgLdKVHI68W6PQcm9HS2NnHxxE
yIdGaedufaI8gq6hO+neQn8q+x9sjJSo9JPvBnyh9BJM+c1PWYmAlnWtsxlkd5z0TPizgPqAfSBL
kP8Bdgm/8Bs/VGw93n9WgVHzhb+fFw634gR6cR+aI729/QGv3H3jPl02b+3fB/jbFd+wNI4jvdAS
LW8ixq/UzcHQUj3pjbzWRzUb2jKdrlrp9TlFaOZc5Hi92JVS9HPf7I7/Y5P0EYR0CszAStxrSMFF
Bp8UAgqnTMnJD8xpaytgUYTPMQE9wdCec6uM4smShsWa6+xs9JgvxsYX1tLZ2/VeAt6hNPQV2we8
YuXh6/4Q3B5jkAL/n+inaq4H9r42dsuA5aj8v6kUDZQWBRU/sTYThW9BA1350kjkgKyRE/c6+rMo
f4Ga6plMC6ztFqnumwFywnoBXqCG8wIDoNel77vTcJjzFSiuHlcphc6gOF/T+fF2hZ/bVHOlSdua
ll9JZ1ydoKqMKX7kENiZsvXfT5UJp8QyVqz8Q1RGJZFWyZ1KCfyiu/F9o//i5tGRQG59DUuKQW9y
FvyHaxfVtGWQprxSCDBi8Gpu3S/d51vK5+kdeDEHwoA76PFUKBi+SA6NzI1ktwnNMY0/EntflJC7
kHjOW2+cXi0oEu96tXNAo1XX2e8Je+30aiCS66ZKpi8nHPdq3Fp9S0Z5VivFT7bGmlMyuSKKBZnE
OBzQJgRQsxWLzASNebr5KUNTQBM9Ar8OznAI0ka9R/atyGDHNqPP6g5bztnex0fpQ8CMO6uo1j5e
E244v0IUsYb5xkhTcK6IdGMGSDee4eR9P1f2UCzh70b2og7FeRxNBpevDR4qviK6OyAh4JvB56ph
1CWq8lxka37iQCtoLMTf4QyroPHASo4NdVY+4Q2x3/2eZ0zzJwxgg/5JYTCP53/MI1NJlj6XwX5y
l0kB3JHbdDxA2Din1Y70eMAK0g4CqkeJ6UhL2jfbJD17cGM4ptaSQDixlYwUCSOkbQaDFdb4n2EL
0d5j07RsGYBT+Uycx8gCyw6klxIlVp5Vj6RYvsZ5kK7YQSUl/asUIUNGYXKqItnx9HZYDjUJRBrR
mW27jVdj9Ur9BjqOgCwmzKOJ4ai6Rg430BIljH0tGWKy99NmHKWpoJdUuahmlp89q1djdt0EfOsH
p+oLgd4MQuZnibg2gOoweH2LDEm0zAy4NE1aCtwroME3PEGaIz7Q3hG/zCcwgkHtvC3mRMQ1XsPv
we9VzFrXT9rwdCloE9SCt1CTbU/h18BoKxhmg/DAvHZ59wKn/jkDr7kca9X05K2YsDdTsQGYSTLT
h/wPiJnP4bs3KLuDJW1BYeu20UWmtN0/BMqwUBe/uYIDFbDLEnueiQr96R2+CVFymRnRWSFzJD+B
kd+5YGpHtCs/1fxoPa/zv88nxoRJMxcEi2TDGV+OQ+Duqf3kOHvpQOLyaYvP86ydmq554Fvmz1HB
joj2xyr8etvV5atrpWiDM5E+epLN6ELBip2qbXAobBLcs6Fn9mYr7AU4f1iUZ89K0V5SDekxDT5o
2qklvo50zeDNLNFE+ssFUpOmoo/TL7Rc+zYD5OAg7Lz7o2FvkCoZA/Y4EktyHYgJrwHH8fz2tt/5
KMVgHQej8s7p/o5Ze2V+YuhH+kP8XdmVCtNXqMVj/Z1i5jNoLNIES25Pi4NQ9RUJSnSoM8lGcYNm
epH0aMlGIlF/DB6Z2aTa2vXuOAkV4KGryLDwnbr6ctuBQYOEf12eAJkQZQOd2CpHYF5z+cdrW6R0
ueOL9uDmTFnnsNZref1WcKbxWl7Jr/40Y5Rwtex81Pp656G5ogl6qF05CuN/DyfbIFEjjLrru6Ol
1RZy/2wEs4onxt9J5C/Ly/gSUhPRw/R0hRG99R0HKKCkab6XpMmVgeMIcNxK7SYgWAeKZ4h0otJx
6+g83OXpE7ad/u2eBLPAlAIAz2NGw3TBokxxA5KVKvrGfm+nemYjNDGp/FxOOg3osVQmfUgYTwsJ
qX5pcsTKaqA6dEoo5ZHTUzZnmC4QK/c8RqlaOfMzl1sBavK0rMswMomAeur1T8MSYbSNjyLmlGo+
CmSndpior4BRNCFzjF/HI+Nhz+Ac3gqQFkrNhMATW9e5psJpzWHumKc/5DHCEWGE2mAPClJ1lVxL
ZLH/JXHiiziZIsFb3NhpOXeihDTKIOz+p2higWSgMQpLlSQgVDOuFq94Hde2WC/GJsNrplwPVuuH
0DW/Kewx4tP26IXgS9kmdDd3AlMbJz5npdIu2fICPiq4QOCaaNXFlGSrmOMigpDWSj2x+cnH/j68
xGd6ty5IWrMDFOrTWl9VgYBpAIaE5NEMr3K3mh7ZgdhbLRIznDEbcfGDUIVVUKuGuhCIjADj8nS7
y5Rqoo1kpX0jpeSOgQ2Q2l7B0GTCff6noJSgbUsGm3eaFB+lcHoFcge98pBeSeIAjtBTUHRBqwm6
1fLT48R4w8PjNeDonxrct56aMy3zk7a0IbXxB3fscuXBgs815A60bEfDfc7rguHVY5re7m0EcV+6
CUo6DEb7TCoX9F77lg5hwoc/SvjlNz4YE0eV+5CgE/8j839/2RGCD+0u+e+QnmRVV0sz99yo9TB/
9e5Cm1tn5qKoCUevEO3zQKluP9jgIHExK3a9c2UPxpxZzRWYisx2IRUL0LjoFANlxEd3fNKOHSq3
DUKDjZXwVQsA1W7XT+gfg4+YHupcEDLJkal5SxlFvuemC+4eSREhVc5b4r2RbnxooChI0L0gNce1
k6e7E6JkyUUsqQujsfIi1A8VGJu0fMi2gvIO/mSImZJ8uUck23T1/WyYPKuWbd1NtIbCEQ/uhlzj
FVw7dBeRyPk5pYsPDq4OfMQJlca1ka/tEOAnGfvu3WSd7cjLKDnbvkxuMkOmux7hpEE3B8d8Rp/W
4xNGBsPzBUJpuqp2fU0386M4PqMsE1AWz2bZaniKDmSWyrWBMihK4IWhECHKYwr4y1r87tZP+VUY
qbMd9ea4cTbS1PuPO4BqYnMEESYBdvOj/NYFIZGAvpwt9gao0RJB1lDyqq+l8XZJqVxT+OnSTFXv
3DSh1NxZ0SyVODU0EeH1WP0D9WUzqZC7QOCOZlCzO7v3Vi93VpkplIyXYrRaXHtNYO1V6Mm9VPae
+Yes7yb4VLC2qLZ3qAzlPojahCL9XK5tz0onUCld8VgynT0lQHKF0EX2Guten+eAxJB7vrZLKEEe
VusbqSJxXppdekIqpexZ2C/enbSw8YEuN/FWtRzrLbdQ0iJ9emuOWWou3IK+T6ysT0+IIO+AoLIo
pLLlqs1varE0ZjTwhVUkNlY8n4bOZefTdnh9UPmsanjd65DXqQLQdv458OviLFqk9WnOM874r2YS
i3HZEIpmmOUmNPH9DLnCIzWTo+0oyxfPnq+1Z7BMK73cPwycxaeDcwKjf8krSehu69yAxQjzvfDl
wfBA2qeViD+ZR6AC49e7VyRP9mIM3ZCCFPxsC948aIgv5us7asio2ukZA7LpfXNnEIBZWEEGVRRu
Ff+vsq9BkMuSHZDRYxlkVjEaqV5kaNTo+x49Pxblw72IR7/vLMcP2o2cemCLpiWHwsHcyouV4pzm
one3Cs9yzkyWC5QEGsOJAeiorsgFfkN4czvMpTNOmUlLFvOHd5yDorIBl0o9/2JNSSZu5xlSP6Ic
/5YH1hZlEvfvMROVKrtPhfpzQLFStf7noYZ4Ny8Wz32a4lb3g81MM36Pg3v7hpBdFVxG2TYmG0Xk
NELlBCZsUpwOruuLBsBerkjx5bjWnjjf2RkoR60pJZb9afO++iivkhkUywrtsyoki8UYPjGBXJPE
9K242ltNzH2du0OOOlSPWEONQ4wM9602Jb/VsFigJn92AxKWtf4uqVtfOlJHPhtkiBQRxvEAq2E4
M9q9swkEJEF6BVRCvY7L0ykhZcBgJmNnePD5Exg/dSyFzLtLIn8tcdeCdpOCo5np7DuKqB94mIP/
RDeR25oR0xGj/MWj7fNkNXkjC81+/KXtpdQCdHL7ONFJa7tFTbDiOTBOS2HA8DkgRr/v1mzbEirx
5JPtBPuPbiJHQceq5wO5TlpMl/T3HTWhm0eTHwtXRNw/1JDVcrHzoaFeGYx3gMVjj6CgrG09FsrJ
TSLxyenXxx+jh8X3lx8BQ3sJ+ZHlQceLak5i1xeZVMXoo6P6Y6Acb9WV9SdHM2cS/UKQFhwB2UHi
pjid4rBRhtfiq/g7JDkYk2+yvQbxW2//fvVxWS865i/yIhEmnfJtg1i0T+98O9c4x4vn/y61QrYc
DcHpdph/f85d5/xPlHfHSTOuXcTLdq8hO5ZgSKxhUF+oFIQPEMLyixMiwuo/mrZ6QvL+JwsEhu01
p6keEVxjkFeeS+K+Ccj/Wnj6lnRiR2gC5Dqp9LA+z4SWWcw+y45XrIcBJLq84y8XRGCQOC4J16rM
Bafbx5FFQGD6K9gJZCDr+Tpk/ePUN6ovtmTe5SV3GnDgCM9k3QG96K8PxZphAGgVRol/ir0a/btk
xxZ0cq2LlinwHtu5N56bieQOkXqP0jE2Ob6+Zm5u2qY0eVxz4oNGLHsJ1HjNfgctEgBnKXle6iNv
9ATSa47mV9wZLBNjZ3BNPqM/ej6JYaXicALIVsPWxIehPqOSI1DIpRRPgtBiguX+LEGvFS8UnLja
d71PM7WyGVgM+h+PR6Rgkg8cKYcQJIcI5w0ifctdaTFHSpg+hPO92byN2xQS8Q1o74eVc5WK9WP5
ZkIyx6CQmaPL566mVy0Jv6McF7pzBtU1ws47u6Hsxwj9sMrZTTf2/M0+hLNtlHbVgqAtktV2rj6T
q0uQ7c881nMhMuLNSQiUWoIWFxiNBtS6f/3OgCINX0n7MOSy4+7nVhDUNpZTeRDj0eZKPXzQSrTF
QJbtat7R+r3DmRQSLC92Q2Ztn1qgGMg3SMGM9EglxVBDx9n6WjubqqWa95JXG2EiztVbnpjNLDAV
4btZG4Qh8dNF+9YgAjsQfU/HzGUyS7gXZsrp2xgxdEytEcVoYmJdJllf0LCzQFBNmqmhNwyiAJVj
xXVmGPLX4PZgSqxtsoz86w49hilwd27ZzHbZlTJOZ/+AM2E+K70cmXL5jDUCAcgBIhZu381CxPSw
kdzlutA6o0i76u3/eR7Ec1asNpv669x8dYcXhBIVzdA7mWsbrcmRruLOhayCLF2/aGVRvzVUa6V6
rGYoxLnegsS50Aax2BEBUciPTh83jPe2NHuldQvgWxw29flwyZCZp/sqlzWZdtEHO8pLlIE9t8ne
MZr6CCx7pZFqkdkLQlhascRIlu3H5OWjKq4jktexbclM2XPvApMG7Jg+ZoOYyGxZl2V5Mg3fj2MA
4IJbDadud80DeYcMjfxAbohZUO9EE0KGxLWt+NoZRidyGS2BYFKoiFXvfpilknnTYrahHTIwZ0Hu
EWyoID7CIxbAhHaKPFq8z0mFOvCj1l0CKZ/wGuWtGPMI7p0d/aWjS0c8yKWsSUeNA2+ZFvrZCSZx
cwaIEXy5lAM6Fhh5y3xBn+YglTzfQCVqRexX4w53U0+f150HZbLAdngrsojAaZYprUg8RUdrPCxq
+KpAPyif35u1YZ60mJUHEKXjt7d/ULY5jOGZ7dIYyR42xqDqeMhslSNLlkxgoV3Lw16wLThvwS8O
8VTLBqqSFnZbnLruQwPjjaktnT4K2VbapYKlms/iAA8sdZG3mcZZkdtF1eoWyAOB9UqFLAghvnQQ
B3BSQXqXosIX+shyTVlx7UOX6VEOcjeJyLPf8nnvLYoLiHUi9WQtJiLcDWl3EsQTzrVPKsC/S/Ym
ekMK2lqqKnHcFyl2UDoHQCUue87dYIGBHhK6UZcr8i+HXxRQ3HDyDKUjAwxZYG4QaLIefCJ94x1Y
v2DAWSh3mDwxSO7JVa5FPD4X76riNtRLJzYPzQuY7Nj0eVUesSthdAUbdNWRwSVclPOwHMynJVlf
Wd8tMu/gAJnjZztGvekTc5p/SorZtslJvzCMW4G4HR41RkDJvTTPEzHALdsncLJB7gK187iqfFqR
nnLeNa7vWZjbeTL1XnOp9ABf4OIF1/uVGkd/c2BY8H2EekMgHPDeY+AxX0saMxt1GTjYfFvdjBUm
WY++Y6PInwrnGd5MkONRlLcfKrZ1rmaOZ4O8sxMtlLR+gRIkosuNHFtlhwdjuIQmf3zRJEzjyWgA
nsYQmSwwFlc0Z8+YORhi9xKxndOz3Mw5gg9S6KJqbpEg+Glho7goROt0mtnQIp0S3/ewEbFOxXir
HsfOgZvQDb9HY1aQUM0LxAkJa6xNkgTFQMVC2vN0CwtT14bQa1L0jQCH2GdK4LOVvZiqo5haf4t2
GETccEkYYMJFLbH2ZWdwsp6pxK9cibr3HZhpW8mv6+EY+CGnMvm3VjnILFY+gJw2LfD45yeWvsE5
tXi+hTOvEZ2P6RC5eVVms9XEh0PdAo3dDEHiyWrnXiWay4jkj485w3rA38IChgtSvnjlPsZLHCvh
/BiLh39fxR64h9rGwqqeI8Fi6e0RGBXcDOHROtjDHNZfRNpeONr8c3Lb+dTWNams4bW0k9J+uOsd
BlahDFf1WVcYCdDCA/dzBcDe6lmKj96D7D14T7rrNGCHlDptXvv0/eF3mwZW/CD0dI21MjWxsfbs
1/Np5tD63qhBQmuDvlPcM9x7XROPQWqvteiIh9+hw7b7laqzrsmTVmAkcNyyreCN1xDO2lb2aTH7
ca07xRxUFIQpvaHC6OZ34Ib6UOAcMh9CGqbUWSD/OFYYZGmXy97b96s4uC5IsSJgc3C6KUwTni7d
8yHqKDshmqRv9ePnnSPQjV5d12UfJa2PSs0b4ZAw2siU/Fpce3+fAM2dfjkRs2qlvOWJ+X5sV++5
fk7NmpMS8kNxVpfGu7l0W9efOHFWOrAaJhiukVZg52vle4YrKP5DTuvIda4aoLmwiIIEAGxZZ7aZ
2tkgmi+urcUqdDIqP3W4Y15u5AX1oq1oSjLsLIxKdgS91n5EyeY22UfdL5xd1ORLbjxXQ35obCtO
oEWoWZfAZISHAfzdX3wqd3TdjIDd4EzQneigpeOTkX6EtLh5fKLCN3gr/BU/23Bb/TtUWZa4qRbx
sRDIFO1ftG2HVGl2J9jcdXIkQK1BPZo+nn98kxAhxvyBKVbGSHy+LiG3xyFtJAII+MFV2zP0UGOz
NCNiYIWjbQurunUlzYNmwDApax2KJRU7V1as3M7vB2OW8sP9TWY9bMPDJpZ3b7ra5HpBEVmLktJe
2qykS0wQO9Y74cn8j+TksYbm/NkMOF9uAiwtBPyVOC82vREML7eUbJ8L0ZJBqDYkUHMkYMUd4Wgf
uXW4Z+9ReyUOTymyuqeWQvBN1KEUDdgt116MUSqby3XHb0McKeE0rVVjJMnS1ODohbCwz/hEIpbH
oQrXNX1RdIYfJY3FEz57XpleG6Efgj2LbNX7HwuCR90J+OlrCT8YNgh+TesnOrt4LR9fsdXd9Uog
JseNenvzw7Tl+hpCziVe2l0gIcAATO7NpvUOyxp99Fbhgpce9g7wmlP5vhQ7/4TJCdKWl8+SRWam
WGK/RYYVbEi0IZCIro2y9kNYD6z6HBpH/jVKKy6pWnToleKtb/d/h0KOPTRkhR6DWLAVNtfxADHo
YPbDzSoWmW/041Bv0uGT4gUZdj5QZU6gdQEZ02TSyeXKWXREweYSEu5Yr0mfotX6r6qzlpyBE+iK
bB1KJEAVLOFt8JmSFUkeUuB1bNU2X84gNZXu5gQG8RVY0k2X5aLHV9qOU20N/NfnEQaNtB07HP4P
rrDPzp75TutsTBI0y53nL66EOxzwWBOi7lMlgRmXxboLUIZyC0/MMO2dvfnYSbvfguolcUddlGgW
pafziMOkbklTh8sDSw4waMuZs7/FVGacRTrBjci23DVWchIPunD83Gptt0b1JnAgte9GwaeiBmR+
rDsO/80lyhjc6Qu0a3JHaC4ao9ofTlmq0GPqVXZJi7ACEU2f6zTGjqqx757zROd4PjwYtw+ABSYi
fm3zF39HCZSzBd3yDVydWkpxUPYVDahU1rpA/qYlaS9YFrAAsO7V3rvQgVLKhwucBoTB7Qx6sUUj
HGMAEzUTMS0KmNDykIp/wXCqMgcJstSxVuZEPS9fsp/aRiZ4AMJrk3pQi8q2pGyoOg/ghRy5NW30
p3SGihayau1Yb+9AuBt6LM/815r0ul68AvqfwlQ8WxR53v4El2Dujqcbx97+2O1+zjpZ3XGutD4D
RGwzKPRxkAS+P/XnYBBCWmTKRBZDd2z311l0YfkupMtB7juNSdJvmauYX4rMimOks+gj/3TKBXv9
YSnymOYVY+ahBKxHmQma4SUokCqVgGfpoTETmr+FvkTwqF64PeNbvOGiVtJ+jcW7yx7lRfZruKvj
AFF2Ijsxc+gf2mq1GIZTaEzRbU31ykuxIbVxjK63E1TILjRPTdA5G3PpaSSXmIzucWDUhDK8KPJv
Hnz+iZGf7lysWbjUDTOoPjZuAE0QQPQU0ql11mEIJt9x/XlomlXcUXrSP9REefSruuUq2SwAvfwL
vtTGt73SPTirxZrHFi6vguRPfGUwYYu+7cbWW04CazbpaOnXev+BLrMqG16NDd7iTgammzWTniN+
L62cGCHSzsHnw/3UrQhaZq803D0D80Hp9bZpeHbMFiTapz9iSGCbfkPlwOd2yjtAZmbY2RablhKN
5PAS8SbueJAbVEwdmLbddtpcJzdVG0hMn38uHPrpulmQuSgKDVmnQ9NTARMH+NzUiOdj7ALBK+JK
/oOJZmRFE+ncQsk9e4astrW4QdGCAHGbYFaAl0B8MdLEIAZeTQJ+JVX7PZ33WzI8Ncvsaf0AgBrB
JNZxaZvvVO+Q1UBpIFI+b+nMee+FFa/fAMHS9JFEaTQE+U74HOm6msjDwNAPHxvd2loFdtXKANgP
iksYt9Z0mLqnll51TGjhXb0BKuFSzQi6g0DYu8MpC28qPk6TryjbbMuZPrA2wxszy577Jk1FUVI1
ukEk5oFExZZ/+O0IIGtg1pYW7cxd+0wLwzCnK7T3+9pfRZegcbCRUXJtSoFBevsdVjOe1FtFTxdu
1dQ7R1a7eeMGeYhdRP+yE18cn/f7pYkcNaO3pw4dur+6vQLLH4pXnypF0XTbNKBKct8cFDDZqQlj
r/ZB8o3guGjPOmSMecIdZu5cSJOQbgoUK14e4kIKfYLNwm7LvyXX3XKEhJO6SAk+3+pOg89rp861
S9GovLyGXYGTRNcxf0Ury3OHBcAV1eU5oa2kYm0+GUKAGZqBuCfvabKydwYxIA6wEU3/7oBr/yw4
diYTqt8CtgMd9r8CH2Xz5/YgcAAGCX44YsRjpWLPLzcjDE2GdUYOWoLd/aLfIU92nAO/V9qhzACL
JN8bYSZ1qUkYrGRZlJQpYdxCtL/zmdhwobStPaoM35spvHDeuWsXCvOdzQeDmf5MVjuhMdph+4MN
ONJadoDsIJuKTZUBOUs0dHNNH3F4yfNCGQCQpW6ABkB146eumsIIKgw0nAYkAY0IQfCe6WOphApi
iTP8GQfG5SWMOj2npnVfcmG71B67FY22VJU6uU8tgXmkb6R7KhiDWypyxkEi+gV9SfaLa7p0IYZT
2zysN7o/ToVxetmomYi28rBuRzJwPcGQTuqKcxuqV6JKxCyKpHZoFmCVreqjdBEibWMV8kDEGiq4
lHXSHZrD+g+w07iCMvDdUN1nADWH7xYCZQv8e4fAv0pnzqSCemt/boFS6J65/89ENsyfVSAFSyak
TeSl+Vuub52ZLMuNcqZYrYevvlmk8eOl/SPDvvr6xFWnmoKhavfQmoFKWsSZcOnhB64gdZlwHgbz
Qu3ArtGHluC56DF6yjhuyHcr53R0rsVnh3R2i9aemFkNygU0qID6TD84LnZ+JQUjZkjqJ0J7G1rE
smpVQj0CpHxvVH2/fjvVNTBqdo/uBuWyVMYqeiWKqJyz73v3+5xmbNq5jLOy+dgMeB7hvex7ZpKR
3XNwSx5awutLeBdiPd35pUK1ZOBk+kxao4XDOOfwGaTVQaaMPkooJEbYEaPtW08dY6ZKyynTNqpJ
9sQs+pDqVyv9IsJEAZjuIRGYCfr9IvnPONgv5UxLAF76rmxzudoPFk0ZoLnjD9Yy9o8uL00ZUMhq
Yxl6J5DCKnkwZBP9IjWmyutzlC7KIEHelyuvT74pzMzT2sFGoxb9b1TYJ3BWUqtQJfWtEWJ7O2xb
P3Hb5tee80rMN6sdlCV82WdKcW4ZDjf0uDHR4DD9A40AKAEcJChmY5mkaFA371cl0xQQdBCYGxhA
ImF9ju1HkIJCwDJ/E05r5viCsmmris2YRPgzmZlF2Q2SMGwqfCtpGnxflkaFoRXHPxuSxKzXTDlu
nXpAcEQznQ4axQlkQtIC8PhpKu4FFzio6hMMROWqDxJrVcg6jkGqYXZmXEiC57ku/4I+kOXWSU8a
LmQ9EfvZwfqhGUYma6cfq8eZJoyKXMq7nhw0++OJlLC1+6eCP+BRU+tPnI1iqMuIIQhwcg8asP64
o32hhXPneD+/rK9EqsXLiYTm6wku632qHlbgZ93rsHZt1n4BH9Q+7ZKxJb/xKRdYnTv8uIELd5aE
wzXMcVpDU9GXSv9UiY/mL7ajaaalTyZXueOSvixcYNe2lKfFlqN6/Wl8ON1Ldosw3CFRyOd8CPvQ
FYUUNsAvwtaihQEWsflwBRIOS4oGwSoyKlmbRjbikYlCO1Ry4TR42/z1IBRrtUmmOsKLbEVeVaKj
Dy5vNv78ACxFj6byzP+Q4QZ0rhBI0j+j3de2ml2v/br2V253tKVrutireuX/sDRiF1gLIYJpIJPQ
GrkvBXi2xyaN0J67tlBKsjFWrnnO2wu2LcYKgyX3XoTw9xOMlXGBMAbUwVSBI2Bnd5YLIx5X5wTF
ANBuwEIJLDmH0OHgesnwrruoNMBhNy3lyiZ3nc7ECub/qdz2YEVibr02fHaDzJqGyh80uX5bSBX8
462hxP5QHMhS7rlSoJoN23dkzwmgZb0NAMglbycSU54D0+UFqwA48ty8LjlePrKHk7dXqP4UNeIY
llxkJ+qVnBjYc1NCuAR5ZfeueGNN8mJJshgdZ73OtJgo3ip5MOzVu6+L4GVbxZ43w9dm9zWDuhA4
DnOf7v5WTk4Mal76WqxJVJxAKfi3M1AoV3fdCB89bFBDxdsYKpRbfMmaWoyXl7JkX8MXdL2e2MmB
bpOr2ke7NQoS12ENvNKsAizwAAvTKCSzFC/mRnJND6cJFwu8wkFPN0n5Cj0emwXZa6QRrRDOtUUJ
9dHi50l/NKtp79Px30krDr4tFH8ovgaALQkHcfU3i+fWq8FMQ1JGp3F5iNg7XDEsRcXoNJyLw35i
poiuzPU2/PEtW3wFgPmwmgYWeYrs//j5OmElq15qetz9RubYjnzR7bNdAlWhIOFYHxBbc4BMjX1v
Xw3Zzl093/ZAgsBnTB1jzoFg6aPhbxUoP0fRXlTpuW1uZcuzPZXkKq+ubNDzi1J5MEa/iAny44Mz
dmKhyzhoU6ItnFw5iMf2SpqLWLSY4aiYCLFySS0JwDBM610BFTQ0sf1Bm2VMOwTUXr2Ac5dk75PE
U1sN4yv3aoRWDsV9XtI+18zO+lqyC1g4WI8ri4TbKEoiQYLt/EQFj2xyOEUfeb8TStsvqH0ylTs2
chgk3qxf1L99px3waaoyp++dMvofuxfelpyZ7bx17qpWmQv1vS2VT1eKJSscRMjs+HbZJ07oklhV
7+r1DZyXXCbazXtKPoWRpiUnA/GyooQBcsIQWW1JDzN4KbTu0zv6rYwXkPvccKODJl9WgLM9R/UB
uxkVK9FhE6+LA8Tz6545kM/SPMkadZeyoA5Xq4RONOK6zI2XdHqGK24JsyK3FuwNj8SG+taB3eeB
nKgRpS1LBzSDySuRK3zs4GPfZHn+0U2QbD31ZAsjdyZdY41cYHlM4z+obU6llshFVxbu9UZ5vQmI
17sDANWpkXj7PVsHsFrhmvQcsphJNcsYWmaCpFJdP+tg3on9T5ZgaZbQWjpuC0G6iPaPKeKK1s2+
tLVbQUqG/XyoS4ONQkIkUK0D/af+br7C3bgshzfD6ebZRgxYxOyN+35xL1jCBSjm9vcwvDWS5V3o
IdhQtIvmWvbpZOhNSebOaiKOHQG5E8KUadhjtpLyORgGLjVeI8D7d66yk1pUiuorQ0H08opP8/FT
IwfI0dyXoG+ZiirOwrudyDkE6p149c6Q1NVrY5emif//FRcneLUcQVvoBKKqw7EGd+Z9In0jrSE7
Mjgi+odTCO5YNY3GzyfHHJ4Mveh0P1VWbjTT5FLzLdm0qRi8IJGrjLcQw67pDI55vyXLuC+02ax5
gF4TcF8j1XHFbGhkIByxIsEm3N7LwlN7GfssK3m/8vS3XxfbLD8H8gTiGehiI0OFq4MtgYxYO264
ZMvQRtpYzezBV+tMRWVzA+cgs4skujb0t6+X2Xuww6CzvLUwm6cCYH6CfAU2zzRpy6HMf3J/6UJY
1kTy73WuV6mDAqSSkhat3DAAXfZyqDBqMWirggZTJmhDWagn689COl4uXAgEVzzfL2/Xyh2u/YA+
M6bWe7JsHIBPq9Dr6NQlkTUwSwHGdX8RRJFbI39YxFszx+rTM5NexjfpzW3DnBDK5bQxphR7Sun1
s0MVqyOgcj/K/e/Ur1qP/VCESjW3VWDbjIp8nk/PPRQmBrRL9HZ4zxPpw9ZsLJvh0qzYZQSEUhdO
qC9p1stGeNNA5JrZWLa6yaH744x+PHZJ8aw5VGQ/emhmCZFp6CXV0vgCBuLlO5lEt9/etXWDwNhF
vyc/SGw2i8s419WAScXO0Aj7q3XC+cWH9okTSzytbtTysvFQSxT6rUAA9o4j0Vz3I7hvW2SefpuD
c5K4F0VrcF3IsAbQuZCDwHBBK0XNZIMzHz4BU9jFrRDnsKcE6UcvUq9yU3yH/HKgJMln9CNy5LNq
QWmzwFTBklhxYuKusIR8oVjcBCzzWq/HGhYZzpGJA2tpSpAQLoMssnRZFZSF/7X2M+QzSmv1kHRZ
Js8L/7qJlFgMg7/M2GbJdtoPaKO2ulGCxuSsFDUjW8E7w8l3a3sKI30ss9zk9yabpDxcfUFXet+1
/t6B45xj5qp9EBXX6oxBI7F5H0QsDZ6f5ATmf/Nin3JpHP0k63dles/Kbd5xblwXBMfxEJ83K6vO
OHKBOx+YWcyUn8htZywW5xHTrPuYxVYcyBsJJnBZ2VDLGH9HPiPwtLM8SqkiMKcrhYJwcVUijPu4
vRBmcvQDGQmv+cP9DtK0VgYA9vm/CIkrXkAa9xMv+rpoP/9jQCCguWrVetxULVSwsVxDckmP0dRQ
MZ8BRnQnK4/BfstEiQO4Ki5dmQIp0tgs3kBnk5tBqXi3Or5CoY0J0YQshwbgLkdm8MEa3QuSEObI
oSiWRrPnnHZDsVUsGiOTZJ6FiE/XwTCF0zt2SiF0xFKpNsFPwbEqRBdaO33yAGRKBZsB/oKO16Rb
DOf6LqX398mRyBnYdzV6T3ShOVa8W0YKOxZiczh7ees3kKFz9bpK87SicYnRn9QVMx9ZdaaG3zQm
yxCJzHLLpYFciCnJypcEgBKNPI2HljyEWum6Z9LS32NfAGzHtGvVLOQ8cKAnIrF5Y1HdZQYwz/LD
Bedg+bpFVcqVFBDEUB9S3w6EdSjbHMlKWfOf7Puy9c7L6GbdQ0X9hCpxSulZIN5SYJ1SQDDj71IJ
wwLU7wgtw6W3H5Mc1CkPrkUfj5vESTjGzjHDnknGb3Wf7s1FXdUJjD8ach48fWMFYLZSF+kl9H20
pphS9QGGeL4M+6L8oqp/1aznkFyZSNJQJoYv1DFP2AbO1b7pjddS4+C36ySHg6og+AFhyIx9e5J0
KMWFaKvx9UaybV3lkQ6YgcLCPSlQIYgVR9B6gxqJhsm9vkJfpgaXDxqSOkyHpbq0iqfF18u8xi7U
d65KZHish5HDKxImnZIlQnIHlU9f/OvG33Z0sjmZX579uqCRqIjFw8jsDMe9xpaF/QjP3asSpilD
iZuKXIbsDG6v5np4jYe2OskLl50ZCGxco2QJbcqdJW/umcaXlq2USsvGGnS8oNlVmqidAHX1kqE8
wFZZPIjmJeYLLMUE0aFBWfz1PVYAvbJ8wAXpRyGRhhauH/NbPrrtBVBxpTrU+iDC6jIsOmt4qXjz
24KqmapTjpY5TbHpLKU97yKTGRzbX3Sws0LiFkAzDud4kx2wWR5MFoY3flAIiv5g5ZJn8WgFJkDT
xms4ym+FVlXkvW/Zz2BlYUWF6E3Hnjsvca7dRW4AA/fvs8vkcWGXUz36GR/nDltpLyiPJo881Zzd
gg2AJnp1cUh5UE0Ok7YCa6niGwicUjIyiLvY/+mzJzXBGmxwdzrbTmKfkcYXSArzMsgxWTffRgjD
MyEsYjsSlVgNV1x7PoxV8SQpwnuhdZ2bgz72QBR0gzYadoLBolG/K/zqRtcGCeC6qGzwrTguxKCC
C1UHMfNzymgCEmtR9qd5IezqKAjgNPvDIxor8a8FqQR/V7awN+ckDYyT/Ekyx+TS91cx7uCT/BIj
uPhZ1YvI61QLHjMGqJCz+hyJ/04FHz9l8aEQ4VEDX4Bp8vOmy8VYAUJom4YZRkBFXAR626nBfCDN
V5sqWX+/DrzQ2xgFX1EEo4nLzCNvP9PJRUhm1woBNtOrja5wxmR5L6VG7G+klYDG9WVTg9Pigzsf
8noRoN0TZnA4Se+gEu9jSaQfkMXPhQBwLKn6Zk7EpKrtJ2IA5HrQOIMx7KhPqTDvbE6xLiC2RyZo
JLaB2JqL5Ix+cy7mTLumwtqNujVLVTca/+GL4ZJ8y2C1nf+Bjb5uFebqZrX4V/VYCmnudojS1GC3
6/l7tzI18if+U9TDVg+6nP1+A4yqBtwS+GK7szX5GSFF/qz2P9MLKNjSERxFPzuoL+tSSCUkJFPH
/+Tx30dRiBInb8IDhrNm5FLSeWk8IGSXDw2xGe5/GAkLDSmGATKz3H1Mktx8tmuS5mTHj2/xe5nd
1uUwIRKQaS4UKdq1APbpZjR/hH5gnZ7cYf76MLnYw/lkgUMblHGs+/8I5QiPjFxjNjmhj79vjG6I
u9vOwMfXanJ2DL753tgn/l7Ump5+MPfIzFAKywYyWTw24HPwQAVlnqbcNW7sr6lW6Byy86o9FF8A
+vwaVZiuJ4GZ4v7zypkcTf54u3QxZh4TCfxf1gPM/S5Htwc/sOpINg5I1H2iZAecX3Sz36/EK1HC
MQfJY+L5AprzHT2MbEA6YufogXWB0wDKKv/yfoGherr+loJsyDXV2V3zPKcfJ6QldTRzlS0XdQqn
a9dB/hb6AGv92mzICcjOYnoxlVFDPCKA7i2/e2d9/VS2wQfSF1TTgKwy38JiwAwgoZL1kisBlRB/
EQRDtqe4lIw3alBEz3zDrSgeiZIQ/V/+JTgknnGDCnXdjSX9jI8syPlLDLOhfQK28yRjQlP9FVmG
m8Ve+8XGufzGwHIH4+KpII3Q+uT8CmM1XKRXzgZVq1erT7TbfPFjbNgtYx1fuVrIXToRSyVgQu5/
wIauMUNlfrWOyJEeRb+XTQrBF2EM4759UJ7LrcV2YiraQ3balyw3UDrbcnovrXyakohViSYJS/3X
IIIW0vzzSxWijzefDFGxe/chmDw1bYnAXZyqQAY7SDDFk+xxl834uVruQqCLjaElTuPNzU57UEPX
BrfuMXwB1JJxuv6sUG/et6s0tvXzbePDHi23c1JAgFwN6UW1bGDOqIyOwaJqTLRSQxqNpMa+kdQi
/d38zS8PvqFNYb6u0ivzAOczT4NcNfMOtNX1H/NhU5dNem/f8vWpuXC2GU0Azf5ljDJ2sAwBQIDK
kBEkVw7HpBDqV9yvZAhqljKM/5p4CJR925UqcbIwYxdhy0mjifT1D/HA7riwvmh34kImH5uhBGTc
ZBKghfx/3aaZbcMqpt0gnbjfupDrwlahlLYpE6qBr/HeKOwd1fapADThn/Yc6Krmve+fpItJ1kbb
O22XZ+qWUBV1fhOuGeIAmKX5InKboZ+UVlNsJ5Ly8F7R0m8Bh8XlKQrEzzXneiz2kNEn1nt1FULo
LU82oOgmHAIUUSVcXs9H84HanFuHPfNJnSWHiuV2DcVBu3XwMrmxdC1EGFu7SSzbkWbw1vVGBXwu
tGNvpDJ4kt7lKysvc+KVhI8t3076R+mmf5Rfo34m2+TXQyvwh9lCRCtjc3nRZOh1K3FhmYaL96kA
UN3+4cBKFJGuqibWLBUpKtx5xUJkhrBZTNqanJmkKLxS2QOncHcgBVNKE0Wb8gyBlyJ6cgn0y7oQ
UD8FZkoBM50K9M2NsooD19ueUXu4LKfOfv5R352mnP1BvzEgDxzNhul2qgOxtxAg2Yt1y1IVV7l4
vuXWrqH2SwkMa72xOZNS21fn7weqLkT8O/lf8jiV5uV7E1xp+VEw8AcgCalqAKcyTyWRueEFgu+a
IL8iHk6O6twy3O7katMqYPjuWPdWuJG3cRM0+Ae5sxhXH5b8K/wkphXhVNdxFjvZk7z9TRXPphCq
cklpEyoCxlfu7BK4NjflqNQGMQ9i0OOQflFAb5XwX39i0kGh2jSKjTGEEWJIM0p5pc5IRCMqnJ1H
ht4r/VgMWJwGqLEvUCdjuQEmLZ0XwtPHZdO5rI1vWTXIW/lByuZp8rN6E0N4GAk9qWTex+TVkOTl
eMLipICQ+mVefeudzbG2eMn8T/rSn6VGsOd1/sQ0WzQ2W1myUzYOR3SmjGisvRRVJK/efJikwY12
h2iGi9xvsaeBrvt64RRzY882K1sy9rvwOtYhwJKuxYcNvRy/OyB0hw4gAaK5ayQ1qv4e5rNrzlyR
4Gt44ybRyip4I/wBJlprCKjIDoIgnpgf8xB02a+giLAPVoSQKuc6h5bxzz558hs4h/F5+fWffKwf
raNJpgmLVKtL9niw/sNjlRD5tbhq8gFa1UT/EsX4VgBohdPPtvdKTyoPtvPHatWO3rqYo+p1+jLO
xxGnVV0Wl97Fi6RM+o7crn4tIaiMZOQlWywznJa1RG323Ph6Yd0JzQARwSeg6fdpQMqv5GvVLlU4
lzIk+WsdXTy4yupVMDL3XVnKMiG7xRXfMzf4fhDSrVqXt0hmCMdvfxxwQADXkEWK2Ac+i+x3MPeX
Z5H2gbmJ+giFpnekPSsS9zfewwPo4JpQJTJ3iEygAvhUhVkn2tOSj/STpJni5c0bl6sg0lCOYOYW
+sVOAP1/PFo6IwaF7vt3849c9ThR41BWsjHqmG72VBTRimUmOEPXPmETjxb2SZ3b8wNDkbTKpP+5
aCKlNEw2wkRCkvwji/SzXtXi6waZ7iWUpLyfEQFT/ZMnLfvx+IGDV025TbNixSu3390rgQQS9gsV
UX93tHVuKHioQyNgix2Xt8riK2L+P4hkMRuUwMx+dU/VaEJt4jhJaxvFwXpiJpkEdGZWRKEz+lCg
ym8PJNVCzmuyJX7Xyj5PjmJ/vsKVc2iFW+Cmz0vMfGDTIe8eqORPj4rCLE56uCwUZzkPrxF6e/EF
8V83RuMVPUlyhcZ206pwqW76NU0h6RcYZtp15sRMq+dP2fjSp7zqAgTKlFlKnnuC200R2ASOClPz
iltxm7IwXyvTfC5GSMCll3U9Giu+Ut4/mESe3xUGczQrFy74DVXc72esc2+Sc5mfe3eh2pfCzBWQ
AhNBYtcxdg5/9kKxEwhzuUxO7dNLhwCOFAhm7zVTQO3e1N17WgfMFxjYYlk6SZCeFuQ7jf9riaeB
wDnADrtJ8uTHCx3BUZ3doNfi0fo4pI58S7u8/NRXTT1D205Xer18usUIoOSjEGFy9ffU6l7nFzsQ
pYcu8mzwrS/NET7KXzwLWlRiXjlLT8c6K5wVLA5pMBNhqibsVvREbfmqBadOVYM6gKEcsEvwWBYr
MC9g8Vxi5o9B4QgKXrQw8E3jvPPnce6Z9WlogTOhKZUwh+IrQL58IhsbYIVT1E1OCqtxO9ZnDjrf
+9VvBwTb9awWR/ImNg3StO51Xcr/Umhni+sLE1qQ2v9o5zmlkSAU7hQjewJ/UTkXVF4oNEtZH6uc
EFAvjesx6KFInPx5mxQL4mcnHl8lMuDcDforXeHx4Z/p4cZE3+HOJ5XLSOZb8BXU4O8kLUhhI+2m
zW6QyBwuuGI/KFzH2qdq/z/MSwZIvP7Ggh02jqTDlq0+4MaTmIhehn+RrdNoAAzH8hlN+QZU9c6U
WIvTZFGruZFwoJpOX+gnklQLd530HNOst446Z7zmWwK+8wYFFtFxeNoc0o4WAdUAKDKxMGjCHNb3
EEh8aHZC9SzySdh5txllQz6o8r4QA+CQnFCBiYm9UujKcC/0eeAcEh+RPfBwjApsi4PyaiFBhjcH
dUa5mQxUyJ7C8AhwG9qoW+2qJBu2BxKjew2WZ+6JC0eGIj4gNi4lCycg6J/iOY08wzVtPxCw9e8W
jo7m+RR9zqipIZvwD7c0SjWp9+SQCJNawuhujLzT6POekg09KM8brVLohjpiXHoPMS+MH6R9HDT/
qIdFnbKy3yk/tuTzzgv3nrIVNwnBETta+ZcAqryemZwOj35dKLz9UnxQTtCjwdoCXh12190oO8T2
2mouGPXdphkSCBheX5137EHUVgfQINoFA9ynxl6aAKlNHpp4X5gIz+mNeib0hwywOvSmAmg387i+
8GF5RqgsqysUaKHj2Iqb7DNE3ae6d7yDV1kpXqHGCgnR85n7Veic8LIwweCAE2M1i+csHp/j9Fv+
8l6v3bQ/bawxM4EsXP+TkI0bkCvQRhMZ1rUbDRn4TVRYbE8pMX17rh7P393z6q9UeT0nlRPhnhW8
Rn+SXNJOnVM7Gny29+F0GhNMHekCBGNdanb81CyXjeN9xHeigMsIxvGk06cdUqy/55RX82Mw82u6
h9QRAOWujyccJbhqIsCFNMA2eCFK4LyCZ2Qpj5pNldAnC4Pc5rcDUg5zLJ55KZPGPmTX5DnaO99K
Eew1+cNbKjARyWO/hLXuruOYoo4aFG8cj8XJoMeU1jYn0uCQ1LGeyLBfpl/YVqwnkhLo1ZDpRCuo
8erPoeg3ItvYSBFQewH7HLN0m5YougQ+sfnOJcDSjev+U6Gdq2FTENPnnyLYJm+bdfFd1pQq028S
Nyezg4leKON9aTeOQp92oJNL2olp67/9Gvbvoc1bpN5cTcK+ihe5fFSjwsHCZQqwFzje5EDr44hU
xbaloDy2YX16klgJQ1cmDlXrzpnNm6ajUVsdxTxjRc0qnl1cflgKnW6x1emmgppt2yGAJL33bbbS
sUjcsSkuhX4UGSO2vrtMl/DrjwqeJUPNN1knxGQkwOIygvnBdDtEBq2Ig8AEWIkP1oSFnVZlDmv0
0gxMkktTKwDJn+YWxQOIcZMEHpN4yl9iK23d3Q9E+5f4PjPoFNmzJSMSGq9fbK8Cx4QA2h4hBjQR
Ha002H93NEcfpHngsZrUEoDC6LPGOgIoDrCD/uq6NASfSJ3OpmrObTDIGr8zzacW3TvnQvC/Rsvw
v78/SAW6FfILll/b8RM7YYc5Sl3g2OqoxVQie/pvu9cTgBj4B8w/7LEUr2EiwVCvv5SDsT81ctpX
O6bjXbIetHYxUt/XE/XVd3mZHgpuwVt56SCy1fyhpH4wkjjrR+ciKtxG9kTULsBgzZmdhO5GbP84
FivD58niYEbYjenYIXcRBy0CTFHfSb06aKrskMUEhUdrfXPvBTF28v4BmCOBXV0d7eRMZAyrWxqv
10QPVSt6pRL11yMpvTdK3cgNoBBZfaSQp94YFmHXwARFMRZ5xDcEOClr9zwzmXe2Tdv61t5JAgo3
Ov8bYF+oXnewTac2kpEhiF3Q40cPTK/rwnqwH8zzylEJmXIxUTVyp0V0CM4o/TvWlp5oPDfntldl
+DxEe/q8/HsQ6cQJswJ04/mPrqnAnRBUteVCzaDXqEzYzL6Bm/KWU9U9hT+uwRqMxcyXfKN2aoGb
Cfz+npNmsDPG9N1crHWvFY+TIOmGCORFJI/fDQpQWnfBXxNMccY/HDgh9Av0ZbsUs1nmoyeRbOvi
J7pp+Un1KPZ5ry03MTIXcUVYlxeoyNgk0OVrclU0Z+LQuY3Mgyosklb3AAZBf2psCzqT6x2biMmG
k3Ri5bdUZAgKhTObIqAmIbQny0LfcWjLkb48O+v+Ao6eLAdneiiFM8G8hm9etRzXHK5ZH3DzGuPn
56hGQnWJA5vsWHNeJyiz/xrM6K7jZ32Jmz0ROZBUPVAknjXGR0oqCsoP+vJ1pi5fQxwvluM3i05R
FTOTizXM9BHXBP3usOHS9HQR5Cw02y0rx9qPLnvk29B5pue81V1dbLGenrh7lxplFQrNeqR/zUOu
EeGo/mEPTOqkSNapUunahwo9Scqq6OwTUVZ8CrSc6tIRUvEhmprh/fhUdv/6KesvIUPMvW7rxwlU
Ckn4H5ATkGt6WqwPb8xBYAs/tI2+SpEpYnXdQAO3z9KkVWGTJg+wvasw4pfVpWOvUspc/vy13Hlo
dP9B4RSZy2jvQkZyUZSIBZucWL8ZusihfsoP4IowIRXliGKby+QEx6r59YIrX06zEEDeRIHPk0SF
2PeDqdxzhp5s2QF0lRxtpmorhFY4tLW94BV+tDGU+/pnGr3+B3WJXhJCrx7uUkbQX4zOh82gbK+5
1i1UTkpzHnDKNuopO7+6wzLX0cgsNL9KWWzzmh5ETkhEHZOd0rKRBYtdQDcvJUH0VTdTwCw9MZsd
BEC6ljy6cwpJFexW2muEvQ1HT1Qp9Or+mVmExmPtBjGuov6iDNHoNOmSwuCa2bEb34uH5UJwqR2+
ro0Nl0PAbW5tHwDrhiiDmcNEUDYAS47pCOCJgFzcHhjx0gzeiEaKNCWkd5GQ0fiJ1XBLB+/Pb56P
O7+b7Ool3Gh4FhSQ3Zwasgqmb6BYlVAWaVwmx8y7Zql27bCWE9oGq79IRjnNRn9G/kxsFFp+n/mz
4uzWiLrxDg9vffUBuwVvOBzGE1j7pb+LD2pxb0qdxMaM34KwPe/XXF2OvvUUo+WM19W1e8JaV2Ik
5vCN9Pj/I+dtOs0NQ8DRP0uFZ3HBeGjMRum1dfWrAAc4kjkQxc/WB4R0YiO2HeACRwPwv635qGvQ
9pMQeLOEVnjiuSI8b1BS7Q1TXKdj/Vj0OUP2eOCxS+ZiwhMJ+bK8oWXfWM60D/8cNM2Yzdf4JNCJ
lou/gP/aI7GyvRm4Vq37Ga610fJ+qUmLNQJu9f1B7BmhYoh6ci4hJj1WhaXfN617Fcj7Ot932/4Z
1aOFS4YE6+Dv3psRP8PMU80segTCbWFQhfg/sP/tj5RocCns7HAUdaOhBa1iTmQjGbozO41+M6da
JwY+BJH6mEEaBudNa1o2E+BvIf0tJ/glx9JzBF2Mahw1i2VEoMDyC70F4DlEFChKaY+ZLMIqMCDx
5ehBEQORkyt7lqLwfDoIdcigIhfkHkoiOSezFy0403PNL26eoSDbnvC8tqPdlW69KKFyNzvoo8Hh
fjYgt0d2Z0J4vBdwKZ63WCehnOWEMB2lQrPMXRo+r14gm6xERIwfixzRzebdTVFawIjCPSN6aaye
grEdYPZMZycQYU26IYCLgTooHdIKZegBTZip+2jpHzKzKsg9aeG51q1ePoOPRKUquxEfSxcGHLrL
kV243FUAJxPBFUXZW4gvCwLyp441kaa7hiXSxpehztPtUN/8PXB098m0yLhgfXVea7rrTADUmY2d
6mHpTmhNzpuD+cteCRJdBkQb6gPre0Vmuv0KEj5LJX3rnx8ZhomDHU35lKkB4zlkTDS8VStBOfKz
2/O5sMhoky06joDDWNVInLxLT8skx0YgQkwcwJcSI7uSLV1YMnmcDy8JOUwzVYbWJO7/5Sc6U2Pf
q375LQ2s2mXVBq/JPB2ZBRu4tHhl6M5ZMlcMB1FigaBwRgzhn/Wa3X+I8XbGv1otsfMS5KHmp2UZ
VjnMSkyfZTErrQHmLDEy4ew4K7iPAjMeamQvlli08DA5gx7N5q5H7LmrPEXjcAnSfdkHxV7rToPk
YGOSgaSF2hMB9uBMHxU3qMhjCvozGJoEHy2qPsIEflwgp+FZMpvGfbFewSANNKaFv6QtBLEytf+O
3/mM/uxrrTj6V8H0KeEXBzNgKPKwhMaZGtwHvISIP084iSSvaYbNI2McZJaSvEgJAan9MgmN+H5U
qUyS+pOJJ/eyOXDI//KwZ6yfoFaNvd9hebR2ZshbvbpIWau5Q+Bo6d62usOw9OAqOD4LGxu+pGKZ
7dQQVwm2fhvxzPtGu8WZFqXtzJoRaxXW8NSrsgZaqMwwPdPmPoIF4dYijiYILj+GVR3n+yumxRht
eRCSeWs7HtJffLX83Uo20NWraVPaAh1MUqYVqbywUf8mX23muPUelgDDoiG4oTrbHZIvmOT4dQnQ
PsxFivZBFj6Z+j3N8HhaRcMtrwQvt4KB8KOYEPPoxxWpZ9Pup5Yoe0Le3bwKSJyJnJQUx+GQMZ6D
bpEGZzXDVGihSBDZ57ImFjviLa/AjAsba8evMATcosohYtyDrbC+9Ee/vL4uosK9YbaApZBI2q8W
DBSLhpChvc07pgvDeyuBGsYIMPzeZjqoSBuLsKIbgSX7/N/ME+LqgPeAX7J2XlUJvkQ73x66YWOz
BroSZvhzNSi8PrZwfW5bRz8fzNYuvDgpF1s8+ZclxvrCQtz6EKK8dN8A7I2/q4FoDyY9ddmQOJ9b
h1NZEIsr82EDb6ndZdg5GUOcOlfT34sp/FiQfKw3fTtGsw+Nj6nkf360FxiT/nO5P/cfsZ3wzwq3
4f5GxqRkgwHLERklFk27MCTm0uAUjzlIjZDCf5Pl4cyTTtqzA8154LfwH3dMnqJmh/DAfSKpU4jk
zzuVJR4uf0ZBYcLgayIUo/bbTt8B6wC/ziAmM2XInFgqPGE9XgFRBxvYE12lYagBJRWoRlQ34/1B
lpgPixGY4EQ2aUjfMIEadXvfUtpTTvzThwbXOriPEdTiNpvRbZfnBwwkpZof0j+UkU9NR/C/4O4+
zPXDWUQyjz2Ct33AENd+rwbctcOShyJSkOs9nTh/QpUWP0Trp1lXmPFhGHURJwB38PhUtXDTkaka
b7ZGOsSrHZBCBaDxNjKNWYaOXtv467ct1bkYMa9UtG2Roi0XLibYS0wTOn4uA29IWAXnKT7iwSxO
+osOvgaA7uqzt6iiLzYzy0qps85tFTt2TtzcYeOWV0B4d1KgXljBfYtXBsuRL8T+soKnzRbNjLDO
YJ+zcaYfnAzc7d2vS4Su6s+s5Gomz5nP7KEQ+nDh9DVTGmDq39pwi/fMokCS0Om9qqFff5Ph++7h
j1G/Ckpqnt68CvbUROTcih8YKTh2vsV1TP3+Wmwm3FRcSsT/dLfjf1H9BFeCBavZD6s5IWMyRBil
FWyFcSrzWYVtJduJ5YNhQK5WUlRZZGuEBbYTT35qR9iC2BVOvFZWNCmnkItoBFFDTxWUUmTf8NXB
yE8PE58hz+PvsHLoKCnDEY/kA9iNS6UIbmQcXVWtJHqNaGzSv75yW/66UHOyti84SyTywjp7B82b
buAi96CNgzUZEMIJmYq+p58kjGKX/DtUfts3gxOklwLobEvo/MWt8llk+Mwqitx6LTs57NMC+nXl
TGf0Iilnjx/n860ujzfr4zXwEhE9PJiEZWwT1QPtpAQuTu+YDN8q3WSVP29aS57ClYzYXIRSVBzB
lO6mW+/9nTATkbR49QmrEw+salJf+AFWLZkGFnqS366ps7ZD/N/fYkplvAl78VrQDY+avoJ1QFMq
rmjdMGYAcQ3MndC4CQm8zegxO+MbnL/DivQnPsV5jK1hGqdj8xacWi2LGwKAkApS1hExWQ4u8YLQ
Y30p++fuok+TF0qAltvFiMCm4ZwZ2nogVPYDGYt01rmDcQIHFs4GoNWuRiMILGxvJK5pQH2VNz30
hzpl4nxkr1lfjSdUTfgPbCMEDU6vuu4ZBKkL3Nb+g3F931G8K5f7+gXc4tY2q1/ho1/07cBMTpOL
yM9MhX429DF7EX2yxmD6obDfALp36pblr9ftcJUFl8paHp1WewcpU8JrqRcvrAYCzLXnz4VLHstD
E9WI4rsXEFg1B9V7fYSQV3KRA/cPkZWTCbjfkoPDPkTgko/9qyvkSkhp3Gbw9o9MCUjXPEnWbNcl
Vpqfc2pp477ugGcGy3yARgxfu9M96Hb0sgBoY+V7ZwAQY2GGX8fuZtzvc4VPARdyiOzigb7ue9/q
ULJ9rSanMF8KH4+6+7NWQ7xREM86KE7WHWhcO69G6lSZFC9HxPRd8+kDqw7VljqI54OQy0HtNmHw
WPz7bX1itqUjiHZTSgN8/UnVCTvKzvo2YfzAmBMwwCjOgNOFeaOic2tEwlOiknCahiXG0sVYdzB+
606nkmYNEKFPvX7ABonq1vviDtrMfzWtG/WSfDP9DsTGYYHCIWABzrQeYAgKaQXuDAA8GS0ZPp+L
BhdpTgRJwR+0YPvgBAcffaeqnrWN8344Y0MP5oQNeORN9FIfcxxys9jKmJDVZ3bIfTwkBDALfnKa
VCjZvoV0A3q9voMm+HtL9AzJRyBWad/xsBCWoR+w+ieaXaxE/vC8FJ4MYU1hICDG9ylGUfdEHqyS
sIlUn8TOAK8y/hCMprsg95BQ0R7Qf5G43bTQi/LCVYMwYFi1AVJIouUXwrXMGxeI5184Pb7oBdAN
QzEpdGvZDOiKpczYuuc9dysfdX4q2FFwug7Y02/H10VTso5jtWO2aENtfNhm14NhVVuMCjhbGwfd
qDyWP+MGeMBbcF8x8F0HTKgz3UYWJ8GCtlO1LR+YcN2sFCwzM4JoeJ2Tu9TX+9lWXUdi31QdCpVv
Na7SpU9uTk0NIobPEMpyU891MXdVjOwWprdla9evlrQxQrz9D2CwYnPi7vZMUPDpascWuFyekFD/
kt/FlegDv3PqTEfJXScVL6NIkzLQnzKRqhqrFCSI5+vIxEoMPl8tiX1SV4b+airer7RkJQF9vVeq
GjPol0po6sQrSof7KdP0RRNOMBnnU248oMfP6kRpLXxVuzqYBN+PE9auq4IA/QGlzQK3ezI4IyQL
y3C6ttPeK5N5htNrZXlHLCF12FwXS2rojkzYaYIaJVO5TDdGtlzBlh3R26r4C7Xy+4D60ZvsE7oe
fgYLxKX9a6Dc6tmy9a9to//F1Qxgj9v18OBPBzRYgFAhNSR5HxaQvRtyPbUeLjrFjbY3WSQ4jAHW
sgPCcrLlbGSjH2d15Wakc2FwUypXYU/NoaoHjWkW9W/gV9P/K2pJEfk/v1VEPHcR/LGoJbIGjD+6
DZ80VgrWe2WnhB+x3c8bUlxbaioIC0XwTaULwr5S18bHa/D0HxQZHmmaL5Lr4zTTRqS8ySDFPIcA
PSYNjfgmOhU/GWgnuvjsSpVWZEGY8Q2uz9PXJsHoHfEbgv+I+HNL2dP0CoeaAcXkp5d/GY/ktdcW
Hr7KbbUBwxj7MeTSrvVWV2zYRRrUDCMf2epKxwBqwZQP6NSn6t+jTytA0ZS+raw2W0UyZHIlL5aD
lrii4mRyRPTWt5St5w0OtEawNl1XYOlUOPi9GZ15E7cXiTmixHD6D1//z57AiThRAyAPiKWqUZ+l
DsS26cQ3M/LpAzpX59t9UyKix6aeNajhXRwGwZhVD9Rx5xL2MzWx53000hmu0CmxpWNTDHbQqKzD
jj+g9XLWMLfd2EMx+x96tFrOyjF4fwPUEDZkSHzOar9Bl2itMpLOHA/T7OlHdD1sxnhcGdl7zz1p
orVn7PFwJJ8T9Kp/ybjDKPKim0wvbgw+kN+fExa6vEPqqPY/Numn/H9QJmWBO7mFdBwih+oYijyH
ffjTd98rk/c7tG7W3dMYjswTOn7AbCfS9fEp9TcH35jr0Tbcoa6M7SbP0p1hcZZ2HsOQRA2sA3gl
HCqzVvJIAUL9wMU/ghZlawT1JDW3cFVXBSBcNbR00svfI2dXszyPTTuYH410ViNI1T6S4YGZP9nO
SaT8bMQSMmxy7rHKO+oFx2hS+vbFAJSLnWXjrHNO/V4k1WKN3SIo4vuCMKXDmnvxD/DyV5n9zerZ
+TV0++yVs4Y3bzrOeXz0rfbnXV7XkxC+yBI4gj7AYITcxtPpzldXfQKH02hWbykIJu5FObE85Imo
5RQsGmKIn/lhWuN6h/SiZz/tky9N2r1NKNz+MUrUsLVQkL/b5+Q1zEqzw/EaVQIzy+5/ELq1+zXF
dwaFM8Uu2ELqVq/h6rfr5JxMFR54TMkfBcEm05XAZ06CciMLRmfFJigSzqmcr2cGXnL8gPpOcT/A
50FhZAtpSjJ+BNbB23awjarHAl5xfeJw6IR2tXKP8Tylt7NXzavMokjjXbOioRV5OH2lT4lQT38R
8TSEWxU522N3Up33Df2whq2xmEcvE0Hdxbf2o4/B8LqrqNUNmHE9PmlRPeFcDefgoVlT0tPoC+Ck
NuYqvIw/D0P4LUKF3ZSRA+CDpvc1bc6IY2Tbid2vnuaS6jOEkzaqz5wrCOLUbP4FpnbWGGs7AQXd
kCzsSETRPOCSaDIjIAQXLBwfzOZvtEtUO9uzsbPUfxNTrBDq7mUPVzQ1MgTPKHxqBZr2HWUb/3PW
egmYJ8sknsdFbqCEXyacKOmDE9ZZXET4ZV3z0NTB3/cETAJddNHf/XU6cjuZ8loAxh+y86lir7Yg
0ViVpwi++U4NXGWQbhomr18lg3V5r+lIAizlbklbnUuY4mesH0kPt60CtBbkjLgjgVBMs9Cs+TLF
z3GuB+EcOz+phcZkPBj/csozFrGJwDMpQPnKB2NXM5SUfEWAh8HsBtsGDGVPDDjjsj1LTYYMMzdT
MYHLcVufq0dvn2sgIPk8eMFX8xiXtPIyHWxwrUqR2zwLjltuo/YPvt7JUdovXxpt932VfR00tYeQ
bhJW7BX00lfy4W6PslFlhzBMu8LICMSan7n73BVtkPG+HypOts0UC5jtgBvCiahpH0m6xYzNP01e
6ZmHIYSTq2BTPqOT+RxBVjyqPngvKZsBYjGgGWG/cZXAu7AOWAdHPRkOY6CRXRh0qZmo153uGJog
BhPj6YKc4dHDSy8uomVhlQWTt8l+TsXV2y0CANRWggwcCKizwmXY2eJ3AdTM6ANiK18EzMF/34NP
850XKnZKvJ7z2qJrrncYEq+X4PpaLlz/nPwhGeXpvq9FvkNA+wkZfLjxmGSZeM3XEhNBBpt3pIV4
V/gU0Gaz8fCe8Ea5Uwj75purd/zySo/v1S5L04sP1gPDW7FcS3oTPEJXL/5BDw94kgRAYHIFv5EY
mH9UgEfymwJEwW136qcUXSUfHRvqzzw+7Cg68TO6BoQKzxRwHA/tSItdyrBoT2KYCVAFbRWC48Ib
sU1DJcVqpFZjT8EOhxjhICi/w0kGIBvDG2XIPu3b3qSjzqodGlmbUam/STWNZ3RgShlJ12LxoumL
AgQjZqsREEImZIQXJjtecCq1Tz09WPXxqWdAmdn09G2wzyOH+/yk7uDNeUnsy7Ep+yioGggzVGpM
YsSefjMrEW8vTqaNsCPIFx9KNudMG7aUbGaZZujVwAXbehn4hupTyl+WHrPGnAo2fsSKP6RFJu7t
nEGhPX5NgPE4+nDSWgtvjWarqHMnaQvANIdDTTbyQluHQgcCn+NnNzCKyvH2mNOtVpemWoOks6W3
XJ0ec2KN8qHFgB0MPWp2HAANWtIdzlqg5D7487lsKrpuGc03oTscYovRRp4PvhWxZ0IzfLxiFzHB
wvd6elWdygNgfxlkBUBY9zK3r0za+zc+Dc+Hst03kU8fd/UZ/aEF2mEBqdurTwNOLtebGRIQmrcp
QEit1tLnuYjFNY3A6QbNo1OsroayjOFh3DOTpyZm0iJJye8qBR9UZQJnQx5YF+0KTbAtDHxJY+Ep
mydETCd+ZDBSKPoL9oy+enUaqzSI11+PiGqYv0lsREg0aGGbk9vB5/51iBWJU5KdxXuGUysctidr
B6pGILFcBHag4cNyYhgUcT+e8tU25TvtR/t0JCunrGbzI/YB3LZwdmdksH25N/srPUnOpzomQiUA
tnWy2RRFi++f4B/ITDzBCqJc1CvaJgsMMTI/G0igHqK308kBLsDfO6ThFoJUyVdVqO2JFDLLt9TL
UDhvlR6EDMUaZtckt80lgeFEDjFQfAS9tJ0v94HIVrBSr341BH6jwbb6qZ/uYpDRtkXHMC/W5Nuq
cgDoH5DgLQuA6iHeX99oa4XBjBqxrPHqjGdrbJce9EtrDuwWjvEaWXTlOUzCw3mikrnH9oda+0li
rO5ZtfANn0+5CViZ+EJPfmMoXp5z6/grdbfkjkRjBItTgj8tfeSq7/Kxx95OwAociEgN9Pzb+tRl
5H638RxlhUbMUfl+tpEBC16NpFIhahVmRk0qjHmm1ucjNJhz+ek0sRHN4WdS8CoQfvwadXCs6RlJ
OhGVeJENmTt5kQjoLRrx58aFb49io/nqvY0hEGd8+XZwDK2IGDZxqLuDsZQodxkyfazX/WqhI/sn
meagxw+etg2qpHM79ztIjK8v3rfu0bcdHGxHElWX7PN8oZAryWZcihBwm/vgJ1QpTcxAUA+P8Akf
QipYSDPvlpWfY5hfwixtP+ApjUX4Tgr/qIvRjXp3rGLOmhkMRGYO21RFXSQnJ5TBGdQZGGz0/pV/
OySZFmafU16V8iADuTSvXmf+icdbg9Z9x6yqNTsoSQqAWgjiWPkUeR7faRKbHuNfGvpf+7SqbPUB
dO4qVD6by5pz9PvydDxvS7fHFKfy4D/kotyjPbR6zqTMmECS3JtWCx5jJ9kdtn+TjE19fxUfn5Ao
4aM6vvW+ogPTeTFact0ZWWHkGjlfPHoZbP3rsR727SWcQyttu9Y3/ey+aWT3z7QB763+QkQE7/sd
Y1RIvdYmPUrogcJ/zW0PtoDZ2WIJtCZ0fORxASdZcSkOj2YsdT/jw5jJI9gHCeJ3i3xotGX262up
xw4v4bp+ddAe9EgFPagvxjWe9YkTqezttfZLJpc4p8CtHAQcXM/lfIR/6zya/tTvS4tJq8dtjF59
eGLpJyA/RaeZoDe0ulpQN2jRo/zgAh0PCbwSVfPimoxCNiBaXAmNHMC3I9kBNvx9zc8S+xrj9mer
FnxjoUn0LbKOb8KIBVdZVDPbM8Wv2StSOVjwgW1NRBgdhJND+dQ9Qq61YXS1SQZ9SKQ3VOV05BLd
dnWCsGSY+tUZlLDBvUjHoycUIq/dnm1zCRNwZ25HvgG7yJsU+w8khYRfZMPrZjgt7Fgzh7FL3cgV
TZbrqKgqtKDfGGiPWX9GM5QE2wXzXO71ebiBlCTQKQw1qNuqvVrT0AgAteExPvtudoIjNaZjUbrB
4XkMI6bVnLpiWH7Pv0jdCn4X9KpJDTpHim213JivqIM+cc3cBeRDw9X1aY/m0oJQyYRRqeJzGY8g
aN55zdfVoHxMA8gkzT5l0RL0S1GIVxhIUMygeEQcO3igxjqiJ4R09p4Ka2Ozyg3XgDEbJa+APWUs
2wtsvfWQp5WNZRgskv+nos2g8BDM2LF69hVVKMmL+NMD5gCb9CmcwCP0BlKSI+4G75ImB9efrF7N
U/peTj2+1YVh8eZyhoTREF0zw+mz+/KLXM9Dl4ubkJeb4xlmSI0wQiuuL0q5iyl+2XpHohXS4Vub
gKGWx5CGbC+J1g7f4eilJjG4lNcUaupLIN2HkNUKI7Y3lXWwVMv2cK67GKXo0i3o9BPPE+7DSHrC
658r+ljbmEcHLCxKtY+cXhS+1bPs70UqGDG9/4uChyRn4WSogATjZZikMpuSLUQjWK5LhSmHv/Vi
f7o/cecESuG3GQIwsOp/ZJ7X1c5F2nJhPdbU9vDaTPfjFvta1geuy6/NNzWRJM1r33ksx2q8MG6q
jUjpflQcim4zio/uYXNdHRcRB0ypMIh0kFL2iKi4Hc5VENfd5JcHip+hjarjo2x1RR/IpGcMPeiz
KhGCk0kljRDqOnilaQxcmkK8GUshscDHfwekqvYfKDyMU47dCiLoKafF1nn8QsSIDsz698RjDES9
JLvrFTrHy6pr2PkaxHquxfTeUhG20nFPZI+Agz3G/EWxnuovEyDHv1g+CIOV+ASDf/3GzmvYEXah
QXZeM5dTq5l3VsPRbD0cXzQaVcKqR7FJHEYu0wbG4ggMtJdsW85O1TeHRpap5jO4r3sDgxSMFYB5
5dVx6Z50PyygYO2taqdRxeiJX78AtSolVze3YXtDAjXZFge5fzwOL7PkBYBOyMcKfVPvOkQn2zQy
KGq+O58RCIkLTNk78elcUX7YDOcn39QWmHtHfcSNRv0fcNsrHmgN44OAydbVAcOoWGQHyqen6ppo
nPSTsIRXDH38T+eMdCRONGMm/behKl9mtpHfgCJ3X1y01BlliqVzrYNdvIZvaQxsHxPlb1t4uwP8
1HjcZBcqq4E4Sc+GhfExKEk4TqVOv8i4sft53v7a9iZHt2G/R9gwxQY38afnrfq2yruVECL8HD37
Z1uLfryaplmiPEGNfdejUIJQ3V8VObbDayBet6Yjzq6CCwALSzFYj09YcHStd4+zCYxaT/D5SMIf
P3qhJVIED0HQE48X+kV8n4J/u1ZCewvwfQERCk/drzOAQxT2ID3pgMUtoxmSaASLkKR7zasbAq4R
AZCbqiZygIAPBHjLstv4oZvan/UICkfO1KzEhBetFWsL4tc3wP7uAtlt2k+WDTGDqqKFASkyouAQ
jhNql0RpsTF5RXvjTZjq/NXy/4TPTeUMfsjh0Rh4tdixQvDsuWtzr5pPuIF6gtG0r66c8qu2paAN
OQX2ax+1npT3ULDlNYI0ahDmsCEfCXUjseZO3CT3MnlD1ZI4o+Y+dUp2fRP8dxoKsQBEZ7UAfaLO
pquV6vCR5oKzGdMvRMMi18fefpUgzwrQOE3IIO0ghAL64Hx9xtI0ERnay8eMXQkz2E6RdYOHfwOj
o9996Of8OA3znYLUR7WgL1Ishcf7uURbkz+vXqaJv4wR17iG77ImPt8KW2HVhA08A7c0qE0La7Bj
ktbYMQoKNs8pN9vBjDZDXydELT3yPJbB/JjMae5JrWvoDBDJgHhJxdHzsSyVzxDvIMfunl9VByG2
Zt8+TqqTniYesaBODpUOGXpATR1jExfsq/+s7jDiRME9zbAonnVttv8IZMGhKeA6zjFk4MplIoQy
weq2dui4x+sQ24q+ZNzY0n/iNam+ZXMHY38UGNPwaz0bSX7HkLEXrxIaKQziHNVMPNBuMHQnPKUF
tsLCB+u7UaFi6mvaXKwtC/QfcNJrlqOQqyMHLA4Yr+WM4g0ru6vfYQ+VJZl7uEnVhyR6LvSgAY66
EoRW17gVAlPzCU7DUCK4X5lAHLJbS0M7YbJ3ZMGHhl2yaQyAdxZyTXxvJUUzOA4lyYu8AA6+oclU
rHVC0giGC2NlrF/ketGXTt3pkcAObIa+fxvaOb38QCKYuWz2MjROZuhw2NXs2ppEL80B2IIISDCU
X/Gb7VoxCilU4+uV6kL+GFZaasJ27JW3EzgDJEagpLLiutHlJU0WM7fy8YszNjHclBwXb+5qD4v1
kUX5e335lhdSs1Vd4s5Lfx2SAPgW70d5230CdfcuQUevXkhOF+8gzShNZm0507QsbaUVqNZi6vgO
dTEUHbFssK1sObyXQ70DGqUzIX2YZ8VJmfhOx2jbC6tnDH6aNjEGh2g1d+uR6m85Y/dyDULobIIZ
t/9Z/CWHQRokgusRToeMtgDu0W9cOvRe5/0nJPvzeP2Wg3UucsEVIJ09kcmBndgaBLXLnnxIb433
UTdxn9XjpZedUw7cBX5VnNhap2NqcMP23MgX5k3BenvUlV7uBbFIxfS7t3IMV0gSkCEt5/Fwy6DY
Jh2002Mic5mEcupdTSAUBNF/wMXvP9lXRJn60sAL7wL/pNUmVSFgsnqgdN9ticl3YkhPrfTlz+Wt
e9czs3l8HcNpOhjMRbj0prH8XZVKDB7Z6eNCkIDE5hwjqFisc9z6V+/9yhFD5s4ZtKD0DoG94Fsm
th6cT9fPC6K76tTox9qP/Lhs5p8KBbmOK2bq3397jfmUNVlTRatejfoETHxmN6SbwmklAyOnu6do
7hJla2o56xHd0FI+jCs5hTpjFaWriGnb0UWUp9TtNPXLMec2RI/3WNAI0rS9AFedcIOYnyaCpYKX
AYvv+7DCgtAj0quxVFNl52RoKW5J99QmvQvi/y5o+fcWUrrkg9NZIYBK57pDXioTjovd0WysGF3q
VFyGSs5S+EpOBqbMAejSydi2ppq2jMLj1zdohBZ+EGBAfLMMWYkr2J2uNDj7yms9TdE/yD6Vf2Tw
jw/ftxlfarCpXpTLieMTl919tGvjkkdQDhSbND9MQ7I1ywwAjGi80nUesMiPqGT9LsaWqumiq6vd
3zy/dgJ2d81cnjBm+dI3q7k6pV++FtEuV2jZgZ2JNSZ7KmgfqorKvSFKMo+zPtVMAIjvI6qV/mng
u1vwEsACHBI1tWoy8YUAcYdXyDwNLKph2eKrapbgeTrAN4sLB9708C+3BdQBFDmNUwmXnxRgQ/7z
QPqMjkPxaD2afMboZlUVeXkwQlRM47T0PNxXkay/7P0XdLR1PjX8FVOz1viidpaa3DujcMmoo8A4
sIwSpXTFNu/jiHYK5slFnssFPc7Eg523s7RF/ndJqyJ6Rtfi33Hc8tse5JONr2+6JrWhg2r8JoA5
DwV8lTMoTak609NBdYtcnFayoSrSsvYkEtrUAIJLEXQxkjDl3fTVzjRZUVvieTyGu7DdA4DTXHaA
97++BLBQed4VBDUGFpqyt2t/n8oT0hq9xVOsy3FjPzPNuunsTMLKfpHeZLxKhjiegJm8MvOJkWaf
ee4sVXDzmWFZ0AdieSTqMMQEpCFaFDrkzQYZLyh47G6Ru2ok8yvyCv9DtXgUxzY/TXRMAmSJztxc
pN71bSVeFHrOokZQwUfCQ00abK8S2CwHDq+H1LhTQD632CgVQdzHfc9voWs7cw2bYVnU1T1xFbn9
sYw0oUg9hTjiFBqVuWl55aBANXCgS9sxsbYz3mEsGdKJEqi3qlVf4+mb85zvpJQwMG7CpCvH7iSW
3Zo56dh3rIQT4vgW14gnmEzowRtI+wBowmpeatKg+xvVdK2jFEXyy3iBpkd83hBO1RXaOw2DI0Mf
38tzQwiBZhr6Br/Ipi3z5jkoDj7HNqjwc4zMXPMzL/Qz19p8rFdBpl9IHXtsrEDW7QWkZ9yv0S0u
7eQfS9kXC6oBjv/ZUH6ij2laou0t8Qb69M2JOm8vu64k52iHadAsHJZscF4Y6wTroNSSaSPe970C
T+x7Tn+1lWIYShkTL/bTF3IXUaE+fAtl8UOMn4SxCRfjblxgY/EqE3vYXWcsjsTUMkyfV4DAhbIb
gG7IjTIsrGKrpVM2AwMFGDpnvYqmLxW5Kc2x+/fWGefcfAxb0MbOpGjXAP/iU88Idl+NhTyzS0Vy
1B5aLN8qZ7TcrgEmeiSWBhPraRzA71oMIP1VVUj3cAlS+5K4L0QhnlvEQS6AqVktd8HgJawr4cvt
YDeLJwNebpVpyfLzza6ArhcNZy3O4vxkx3aa5n8/b9UaY0mXUOrDYt5XVVJDgoQ9A85PrgO/2xOh
bCwu6InOaOg0XHhDXvp6cbYUdf+KZrts8YyrRMJ+lEwSG5ahvoQfyJiPDf4/eT6Uig71LjOscROQ
aAC/UHhFeIS7rG5v4VCaLvJRQyqFYTiAb9QOWB4F3EgpnUChH7tz+ECtWWaPYUbLpllf3Pepkmc1
h0tPzSTU6lLVQ++zOcb53K7eBC2LpBNXBBibo+drHcf/1wHj2jxkDqi1CPO4Y+7+iXcRmQSQiI1j
Y0N13E8qxY/Avy0l3znl++lM0Za31P7+ilGqb3hpGViN5DqvIseHRQVKK2nELJT5SrHMfafzXtVR
ukeczcDdwfg/C9kACQMqwvsjb+J8ioU7+COfZg4btzkeH6u9xws253JetuR418tz0DLphFmZuexQ
I6VE4RJPMRgCLxuc5OItcipVNu7PgMLHaAGri8TcyitbiPZTrjvCWbEtt5cj80ScqjIBNLT04Q9G
Tycfez6a8FIQTMrNlFSjtMAFNU6EUPSLG5gtX2wpKSLn0u6VJuuXrMsU+GDp24t1zmD7qWB+/P7W
q883Y10JBZFX6WIZ6f9v83vUFG8ia4/Iq4T+aFHRtkpqzdTRFIwEm+fO4/mAEBL8AVCo9IVe6ayH
Xp2V/AHSM9x0bDMjoDCNG46zeAiLOl0Rg/AJlAslxgq+Xu2Teu2EXw4qrBWJ8rDhmEUypV3Fg+pa
E46/oy/jkHrkC1Lgx12Mz8Xl1+KavpdfHrMINWrjyEPaKNQTlbZl0PFx3VuoQAc58Nfa7pcxkczR
+LqZjG/VcYsZ+Xv7lRdbLVNhM+DZTysd54uLSxRZW7bLBk44loDqV3h4bIm9IMwBalogcSacHDK3
rJ3TpL4X2zN4cNpxizHC/c13F9yN1+pTBAINVbEXmt4BRSXvRjx0H0zb82WBtkhb3nLC+CbNRccL
G8QEl3AJRXZkZUrSoB9gMjnzByEJQ8U+owm2avikhXBwe84gr7W+xyOdqi4USVKvtmpEPOEX8pYU
jPF6pop9c8bR6WP35KP9ZlUwW4OsiwxpUzOxmTKp65D1cmgL5/aPQSZ0UfCOtkxBazyXtQissX77
t3/4j1fCIiag8aA/DQR2oZV1XDtLVgsMQzOTPIDPPfh36exaVO+zZuj8pWHbUOtgzCPuByKg4vU3
9zWOt7DCImD3QR3k1i/XMAzFW5vuTYEBexo7VLLLTZ7H6PF0DCn5ul9eeh5ejfgGxVqqilVPvigW
I2FvKQAAGhusgqqf7lhefPjPwMn9g/IBt4hn50vGb0a4tcdmVAsBOfUn5kpGP2ju7YxeiuCGa2Q/
TviffvCYfcc6fSofkc/JHKYLCbRmRscGNLbfYtcrycSkCBrfCs5jGf695Q0bo8WiZkoDzuA4j9oQ
9YYsoY9j6pG+O4L2L1BaPPf/y843k+ZA8uDAT4SMEdCKueYWQf7Wim8COV8vT5KzUep3zUNI5zMj
TlZVs1RFPp5nQfiwjxs9JqungsHx/SL5Ey8PgnMnv8JO3TvWCDY7wRFBCX6tTtYbWik+69ISXNrJ
cEVCO9Rd47Nii1FAIq8IKZiCCRMvAfFQDC0u+pzsZdaBEfr6iPCy+LLTWjfGzJLfT3fopJGwgyeF
2c1bXb0ppYYgO2wc5CLO2+6eLD0kQH8aRO3un/drra/LNF4lWOskD9EvVap7p3Kwylh7nFTHoKtx
RkHGJHq3suQMOWDkcRQivKoT2Fm0oyXlB3Rh5ITkYyt1oYhwuO0Ou4gg4TpT16VXAt9NJ4QmlC8h
qyuFzcYw/TEyztJnXM/KToPuWr/JgSArf0VNIcjUzb5qIcVF0M4I7mzp/iy7wToh95uT3mjRMY+g
ZQ0dLJi2rQyfYE9xYcQ9fB86YnBfqS6ffqcr/xvBIpvcI187rmTBiagRH/S+Sm3rA9W9sNX3kf/e
tpRYFWEp+4Vwns4e2j4xNsaWERkIUaG6n95BTXlQf7DfXf2vDLWqC0AamDALjZfQJOoxwgtqGtvL
oKazcqgie8LrEWba87C0tCgfVrin9Vdf1YzZhTZf2BXfoUX64KHTyWtJb59RIaVUjh8SZsOEhnN0
55LklNsjKDDjVqbpQKLrHcPR9LYc+M4bidIYtOKvgrBOdLDY56MoOGYKA1cJEtcD6ubtJJP01t0D
eEqSfdR8x7sgGbD2jnQx49oPZv8zNpRbXgVyTyWFkV6kZ3w9xKhJVOHgPS5TsoxE+v1mx5ZQPohr
F5WJhDCS+9WA6Ml4vvP1sndirutkvXbBdUnG1HVP6Eu5fj9/NtnYFvQ5sy+E3M8ZET3Gd7OdujKt
3Axr/huAjjPQNF4KUeM/HWuVNTiCaQjPHGZDTzlSRSjGNiRoI1vSG7Y2VGmvPbMyo7N9GT7r4qPM
Pgxga769hiOyfx3TYCHdT4G/uSQ9ffZugR4Etlm+cZvRRWWgY6e8okksIKoyQ49AAN8CzVjA0e+l
/qbx0EOTID4EweFEdmDK5JEie8kIe5ExE1iWhyq706HQ9uRUyg4QvXCr/HuXKrgOdkoykMMyZRTc
MYv7llOOLk1rnobDQspCt4vwG9fixHeLDRwE4Ec6udoqlCVaw2AKZcWqKeW3jB9XcH7li/gQWYBz
QRAPCQVkX85WmgwnCdob9GKuw1BHhqncA3nVsHddLdJM/qrC7w6pKnfN057rwoYVSWeAvsmBL5K3
d245v6JeBQ7V7ptUbA3VC5CH0crIsgukTsIbLT4MUqXuhTz3WUsqBbP7OPhrALKA/Fo+of9/5gJE
ngxYx4bOVxjKkisVL2Gtb3MnTOEQyfHzovBtlLa9DIs/8+22y04w5e0jM/SHn2GyEkjMed3MCSic
icze8CCtWQcMg9FMr/YElbGfRHqu0arKBwN8lAdvr/K2d9d2ZAcTBPl7LotTvOqG7OKFIZHbIcbP
hSibFgEK4PSmF3Tk88855gBea19hKgJBD+ITsZat/7eeMS/3AmXw/jqONYNDLpPWU83Lu+v03k+0
95J2z973WxVYH6F9SV3uFRBNs9Uz5AIPEN4MIMx46PtHZVfHnep3vW7PcqSJbdKJrOolcBkIU9U5
Mv/5DIK8tn+olSleJ9u09Hie3Au+6YrZFN8ENAZE5N2Aa2GtXARpR9cRUfyFmOPCa71/Dk960x0l
+Vg5YSTU8otF2FtVzVGZbDwmoYKbiQeyB5EE7J/sCnDTcY3kTI+MhXdjKS/GX1FuItlH98fpOVwc
gE54aiwz+i2HgEm0dxsQ74REc9K4Hxqg4S9hirr4Kkm7JyCZSJoXnG9UOgb5CI4hhk9rFnj+SCwe
cdbAHFrw5e0mJ7LNWuc8Z2yAEVN7BtxChyoJDZpj9+frZJiwXDCDnbquDPwoQPHz0PVTv/tNhjhY
aSg+H5g8vA9SsXhiy8R/5TETCKnV2/7UjdxfsOauvujOTu2vKQa/wguWqNdCpc9/CJfrxKo1tQC/
5E2WJgm6cYXRGO6REbM3zbEMKUayM5LdYyDn2NkHfE6sbx/sH1DayYN2VJVr0oE9GmfU6lk+Mp1p
iLaHo+VWl577NAVGf4WOpxhU3T41ZH3rGA8U9MgbEeqfvpNmfGUio+EQZGRqlP+dusaBPv62kzaX
cZwwF92XGvHltpH/SIFcvdOGIRhjqONm920Xy7+u0bI4IZt/+nG653W4dDs7Z9zvFqoUIppVOrc7
wpjNVEe38jW2BuP5ZKeMCGNPfruS/2/TnxJGdaRbKJpK3kQi94xknpgWtAmu3NTg2PhO46xOfHmL
U7Oq/GHwYBDiYRChzluKnoDm1Y5Bd9hEvWfN4S0sSGtMUGED7qQASkmOl451srUUaySAu7pbQHnV
HsdVoTonl8vuj3F1dXIxiuGAEyWmCa0lAF23Smb8rlkm88LY3aDKKdU25VF+p458WOcGzCJhQCYM
4WujK40r0D5rl1J1vZzkD4ERzeoNNIE5Q43YRZ/Yf3e66XULY6HhX6o8j5SmbMPsik7914sTESIK
DcTW2OPnDQGqCGNEyTZu6MWQAPrRBBZO4cCsWmZwYgWtupvncQWskjQReBUCFbP4UpXWqRJ7N2wf
9id+SLlOn+WQ1iGuvPdzGJE4HA6xJU4u4dyUTyYfI1qZPcg5NSAB7xOkICig4d6qhgZ/w8C2DgJR
G14YQk9vt19t6HFsp0IKyDVGnNI94fxKz4goxl5A4LzbvEkH2lRYX+Za2uCgifvvX+jYmo7Nx7MR
4C8Hhxs1JHkk51QCTTEpPtkOFWv1ieuRoqT+1yCNkjEvpQgDy9EbnXpGGYDSGT2meXopF2GFqgBF
g58lKI1KyIQm69mWwML/iZRcJXlPSuC0ZzYu1XnkcQSDsrmmvO8lpZ1LW74Nj7+Fzl8pnDaP47hE
cPiBVk4mJ3gJPdEvAY33DSdBT6G/MLeCqnfQ9DM2UeQTpDUt0skMSpZEZlC52Z+HLxBza1JPVU4M
19++efwKWpn6cuSVpNawQ6lYk5Gm8u7+kO7NXZXQM1690I9LVOPfH3zpdhyjxq6cdl2GhYPV2KJ/
M/QC2TiPCWyKnVO1/2N6gNs8OPWfw98TBBGVbYGMCWd+2xjJ9HN7IWIJEgkr43ktkRjKaNg59Ud1
UueVIhJyPQ18KCouR12TwTw4FFFmk3zX/lkbu8ZvN/9d7B+CczGTVGq/tMGC4qLRlMr2/LVGgopF
eCRk3vKPmidIFdhiwWMqbFh2Sn0+nzE46ft+MyzehE337nq1BegLO90n3aAQjsLSM6BKG7EYFz0q
PZMb2qnu1qqb29rRSOjjITqArn7vTfqjb6pCW+hNd8oP61lBp8g05rWrbQgQGaWaT8jLUHX1OWy6
N+P3gG59f8j+n+nrmzxt9eMbMZc9xTeg663UaZ9hO5Qb2HBkOvzCIvx1gYWTS2J1EqIoBTqX37vl
cDDJVh6glI9Kls0SHEWRhfGAxsqDq8Osf28nuAep+o7qm5P4DLsXwZZh/vURbQwNwXM2A2sS/Rcl
2DFpP8BccLdiqX4FS2dE7NgL5GJON7BdH9wrC9GWpjJEd+i/eHGSlbhMQT6nyqtzbPvX6cpNR4aO
CE3nOUT8CW08NA0Osw+QuTryQ6sXaH9JMOS4EGxxiNPA06BUddbSBkLxTb0ZaQkM4qCaXM8yrTl+
fFXbNZIcm5mJwnrkciao4Zp9RuvQxin9LPz6yzg1EvY3TKlK6N5qi7LiixVHogk95xA9estAvssE
3Nbt8tI3+i6DIAxGpTFym5cJlyQG0EMpoakVXHu2Q6ydblfW60UbBh0ZWnugqT2uUVkA+gF2Vyru
lvb3pGfNtXeWoxFyANJxKlL3+MReZpcUkp8u8dCxnDpdjHsgCgAqxsCknQspZpPRvDuyavk9UYZF
SnXUTO4E5cMuJvGpqzwHfKy4Si8nXE5+JEqHKJ5vM/7Tvq/J+bLaNAM2NscjQruAsNVZ5DKiB10X
JNKRtKBS/BCkyXHc/1El9NEISxPek5Rc2mV5lgHK29Qipx7ye/tvht86Z0FvTN0IPnexLwH7AspC
RlOTDxmVJW+1fnWWpw2B8vm/0aMvjiPmSy//4Uv/RN2CPFpzBu6Ut7Ce/BlTR6XZBDhg31wtSohq
XG1iNDcpjAdyzvefwhJkGdXKTcRpY+Jv93vYxVM3vyrh69LaUOzmLqCot0FOfVKIGqcYqmifHQKm
OwjNLf2sKt3xKgl8UyvVcnu8Yp6GJFw9kT3uZYP5NEjOhGL717/KiX8PiD9fLqzAbf41FwwA+90b
su37lNDw64Z1eKqvo59BtKGVbjNO7LR0vHjflqWcbrD++nyQCKUInfQTzl+JDNCTukqy2QMcq4oc
C9ZgKWr6WvMO9HEGfDNiKBJAXAvrtlC0JowlsBrTHNK2iXx6wTZioR+Cn2u2bt/Z6WJH+c5NxSxx
iERwr4e0bPElOBvPHebN4ytDkM62P8tn/z9KPLXjpUrjgsyMqGAIl/EjyO4DPRSSxcSMDt0qUzFW
n9MSeuEjTovzJB+MxA3f9bi4bzduWj+uSpOExyYZ7JvtZPIhAPH2cgIhF3lNQevYG8ZwrfemVHZ4
1//nTDPPfcpGUxPJu3xiptbhEmokGfSjeNuca75UcS7OaL+4FHY+DAd1W5NEsWoJfTEVeFHoztGb
4Fkds3Xj/5hV4qh5D15kPXLxYUHuOPC6Y4I0JASy5yGGWCwc3j5XMLtFq0J3GTnPnTeCks102wH9
w6RPjA/68l9SiqGxfc4PLrLrKPUOAtPeeptXfvZY9FJCYU2+drpX6BQ7eBgAblCoW0OGJSKU6gTL
Lc0qY3c1MHIIEZJVOQ7Xn6SS4jU9XJBKRfZo1MDct5pHajmcmLHudvJDeYphBB7NRcNDYoKZiBJG
oxpC7hElRci+Na2yfC4r3aNjJt/KvC/A/g++Cd57J9o08Ly9jzvhtJp0X0QfY8k6CpZHSo/WVF+u
DpJM2nyj75uh7DTQIFU2AQZvKdZWzSbwYF5cQSXTrifASVq41n8Fmy5wI4ULdgveFXUD1xgNBLKG
x8qX7DMHKd0ptYFgFxvxJ9pgV2q9YQmGPq+ax6+EHWnCC6lVkQphabPPLCplWA0omhpE3DXDAHi6
MvXse+BIIfllB1IothOT8EGBeZMJc3rUVisE0f/AtJUJ/+UzdokTCMejAFm3qipbk16vWOyNEdqw
53UoOXSKSDNXobORZYYgibg5ZYIPu7oEKxeI8v+/la6HpNYxzxvOjIRZJvgM0Uax1v+A7c0fh/gJ
GcghGsNOG9qvHEgJ8SyJVpQ3EomDWcCdIHqs0FWeBn9WPLMYpRzYWMgPeSCXUTA6p6V9xWB4zDx1
tY4LbnAlQE89wjnXZAxkq5IXEG3buGIyRpMYC0bMrzf7piuMvJ0mL6GO2ZbMkdfDk6hOVgHDQrTO
zb4tzu4QJkianDPDfLb4ELw+M4A5EzWlye6ZTaSEBFuC30j2aoeUBgVCaoVAssG2NTx3UmtssLv+
jB3sEFApM4zua2BY4rf6HW0MFyOV771K5nPXKUGFbIlgjuWFNaEiD50sSW61R8oC8NxMl4qt6Clv
c1enovmxdB5EtRsQtNHFr9/iVNheNA1HcEzXmFwPqXyKOD15M2hMH5sitAh0zFAUO8ocrEfeAYU9
B7fBg52Ckat76N0eN7IYdB9kff5ll3kccNeBsFrnhn8S6ySjisSPakD1mEjtqsrsXKB6fEu9g8rq
mZVkHTR7pR8yGL+p5dIKiHC83PPW88HEp++dnbIiYx+VeWcMimvogOlmOTc7QVw3p1Mz7Uq8lVPG
cg/eoYEU7IkLhwiVjV3wBYIVCiXf+k+rrcXbBYtfSh1ONkvPUCASUVb0Bt1/DM1zQucj7fbCs8Cj
MqqyP/0v7ro3fsSSxa7pBC4mXqFp3nxCsH/x9gTY1SWYeqWqAImp97ZJJYVFEaAxVudiPyDEHiZJ
GJ/H/2CkMivG+Jk7Y+qLcZo2RHeggL1F5SepCjB0gkp26o/NnVsPvBB8MZQSuQ3n3mpsOvO+TAic
xgOxRaEHOXB3FVExNdlOb42/cJjS6SZftO3c92AKehG3hvVVVjD931pEoCkZ872vbMT32Bnun3hF
vfUU7ZUMoEbp6xEoRIk0yxTDGu6B/Vwk2S7qJEkVsVB3WgWxxjVOSy8ulucJ1qDRMHghT6ziqHC1
BMX/voPdw+Qn5LfLCeqs+BCDAih0MMs3oFVUsPkCoiHQKYHtvlO5F8hUrXE1xOSrs4tWFaoyeeBs
ss7CgbAnx3kV9oJ06PIwUwTyq0Wxm4nuZjrFDFrPYNYRCuhcAChJybQtX1M8cRe2ISv4Qa2QibKj
NJGX+gNHpVoVwNFiJ/H1S+QABvP02/tigszGqgxo2XAT3if8wvqokbOOwCM7iVGEpr/kCDhC6a37
2PQUMfF7Ry/onw6JP2v+tbLu42OK3nZ0jP3rKZajOtJgc9rLbsKhPJQahaFn9SWQGgiA+d77eFJP
/2vYmDAlS6aVhwWLCG9LWE3aB3MJvcbNfUVSbKymq2V1Ak8OkWlufs7nphmbBok4SqemSz+gb4+3
cQ0bUz4DsCAmIx1RL1iIDK6hZFqOwTNI2YgkfMWJHqBEXkJkOTSFeTJ3LJF0y1AyvRsq6j8FNx+S
/3PbwTgShwRTphNDB0SIAOzsB6iVA1rRN7ugQaPmHVnfKnytmm7jqVxNzlEA2hAvKSBaoyhDHaaT
emeOglcWicLKQXdJiTWeww38fwxI0u4+ygy3ad5KpLrYjN3UNNGp54BjMc9ur5fcdL8WBN68OF06
b1UGJOnjlN7YXeD0d+lQY1jO0c27FtsdYpYcl+ErGOH2VJTWtuuP6IWViG2YKJOI1YHFOnCTJkrz
BLSh5ySI/wO8whnv3TuGDY9c8FsC08kGpM1XPHTi8Zi9RXH2qUPdlr4HdUd0Fn4zoGgLY/YvE/LD
ixTBSJKgFduK6r39bwwo1UkdNG3g2dJHgghPjhta3LItRgQxkb0+xC5uYoVPDDC1Z94R3n1HqPKe
FvlKF0RwmFNG0zPyj6qWxnYdKsbExUMdrKsfUoYE2G2cMxWKByDahrZZ87iAHHqK9S35N7lJ4LAQ
Ukxo+qKvml15bVDsyFOKH9hYesZp00tYwZeqYMPTqGVTvcxCGnnKQoSepcGX9CpzM7qtjDxUn0RF
R+671ohwyb9GWSqb1oQL8HZZvs+aCa96B+DvHjmNbWs+j4MkbzPf1hnx0exJkIz2D0n3+byxhdqj
BLoTwvHG0izMmb12LvblcwBtwS2++Hvuw9JVnVvSBz4buOcu5O/x5CRw4lDnZVPeZZvg8f4mMuNt
I5bHGh/QAN1Eor1dOpPcwQ2zc088KO4crpc0LjZe0qehpc50YvanALTle53h1pFvBRzG7JvFT3lk
2ZyglOwcaI8mwVlHLcs+LNw/6HrvsuvX9DWvWmfcDRxteZ3ueUZKy6r3CHVT86dbzYEZC9icFEsN
/7Ddy0eiIepUEl4KH+SzaIEI2MHkG9f1YMGp43I7twPg2pe0Cm1PQ+61/TcmIf/7cpZlljDwUUtD
Fo0QGpq0IZJn3EZTLIpmyqfAFHDxF2lWh6TQw++9s7g1YQY7cEGlLb90FtPTzzYr7deQ5TBNfUys
FjI0spJOcmozOPmAwBj03LdT05imgCybXtUjKHrTRuKV2q05Z2go+UfSVD0UJnYdzVjlzs7G3QyA
nvcqWdnRr5LX9hEPevKpZCLUN7wzZQUZ3+tD+7TbDlQU31hz0UOXp1VuuPl06N+RVtF3hOuqxWak
wcs6AqVWfuaK1HUTlUV7bxk2DRb6Q47AnruBLOgJWgzQrSKSaOalz4v2lRNfy59RPouis41TrYRS
HZlLu+nicks9ogz1h8MIbm85loRshoKyYvH1fHTs2DLb+qGCI+tf+H7ULTRgZ36kf0jqSX8fr/MN
F1YhsbK+k8FB6dB53OsiXNckPAOpqXlmyH8rRCJ8xwfPLxYE/NdLoDKb7m2Yel9N2nL9rUKfW0uj
biRblFUuFX2hAVZJAeFaQLZvmyZWpIJZLcvycAy8HQnxpj08f6kVkPuLW0cCR+gT6O41pSq5sKNL
ChqoTHl8SxLlLroa7TNrYlpB6NlA7J4/tKUfFikczErHgkj88pPxHODnqhMb23a5l+uLTGzhwtC7
DbcCPGhwIgIYBia4onCuS2I7g2Ky87VMFwbP7Dgg+AP30QqtRMmA2E2+nXoAXhSz3Y5KPCd40Dr+
vuCL+PVcTlZsB02BA/TNpgMmunh/pv7CD/sOa7zCKMQAQKFpFE0DSBJ+6XiT/wDg47u/jvxh8YzJ
MK9X3L4lFFa/mdbKFtikyXYQQxctgx8GxFljlQHwxDrDEd0i+2Qiq90EL4k7kpb2/BIlUPW8NXS6
Ub6J8g36dzIlGGqGoRgOzjGGfyVxnMRDt7nJb30J7EEohkaWnnbl8Vngj8DNcc0n9Awy36qWDcBB
Br1/XsTsxWeZnBZxFBSEg1qc6WbQcyQQisxKDhDo5iJE2fXSob/KbelCaJII7I1oVCQe97jpHB1D
VAgtM5gWsmkzZNWNFQ95rjlCLPnPyfM7l1SKjZSUT0nCcjFMMIxFhoiWLurSXnV/gkpwdj8iv6HL
g3cO42NkXFSmG2akqX2Vyc60DXgcl9+vqJIy0T6QAiqSDxwKHs8zUEFKuVdZgSDI3PXHHWPAlRic
z1hZK3BtJQvrpzid5AqbVqenpBSaCCXhNcfKg42YfqnMmbj4StWvhi6Xi0T7EDoI1k8J/EXQrbsK
ZXtepPrit5JvJZy1sGYoha4X/8+B3+GxjwFCEkEvWhY+pHIjz81FCtXtbRyRX6qCH81wGjG64pYi
PWxHBQSgtceYPTsi9NJEzkv0r1xPhadYdzWM/UM2JHb98AtteNnhhLM0qGgJMPL5O2p9Z8O7z2Wh
sMQP+whpKjHAJPHmlytObCH8O+5HhGaxpvzEj64ajG//0IHHmAFk9E/2ICqyi484yhGyu/Yvo6Bt
QvuPYtsU08UT3gKfLsag6q4ANxW7qI1C3/02mSPCmQf9BTZTYgVjkhVtadVjOMz43utNY9+BiFnC
U5duBMIl/W2bMT1cxiNMmRwW0jZQthc1MPCK/XXbcSkR2zffxaB83/KpVG+tQKoQeCRv91i5Obro
/kj3vERpvc1JzXPKsAExW1FAmuR10pZg51d/RuXtfujxOTqE66SXMqlZmyNVPjSQGDEjXq/L2Tg/
+KPzv1YG8TCTTybJ18so2xmbGaFQxLdPiB9yh+0osQ/iHokO/bQ9geQvCpgDOd2jAfvw1pGEVJeO
hqLP7E2I9RaSOWr+2JRW3QUkrv5NcSa0QcXaREdp4ByarePeJDIuITErfaBDtE92ekxwUmv0lYRK
RfQsidt7SG51VoapeTdGKK5BG6f01elc1RkG2CrVPRCXnbI2tC/nh0Ux0nguljgb4RGMRnyiy5tP
U4iPd2viqPCwH7SeQuPr1lKm5OJZqf3uP6gJBWbZBX2sJySlJS5851GCPVUiz3fh88UHqF2zZltJ
d+q30lgMNBL8/RinJ2tqmBMAFbno5HOPj3SkvwsRAxRc/dQjITSAKqCkH22+lehGzoy1j1vH8D5E
KNGDXliRBXbzMGpp64EHsUC8WX+Dnf/B8gjPmxjtG5kt2jtWQHxQlqs+Wgb4JyusSuBd79fil3YU
z+CGWVOoCvdDIaRVZvgo0L2cLJPOZr+DA8LH7tydrW37LW9sCQzSD1TxxZ1FODQY5nz4bK2OE05n
x7yXywfsg0VCJhibOtnfdsE86Y7c72d0h16r63B70J3g5Lmvzj985LIMrbMJzjk1WwGbEaE3+61H
AjO0o/VqyEWBWf21boZlUHcLm8o/4d9sfUPV70W1uSleIO+jfqdIqsR4OmTM8c//ecpz6iqkh2if
Xb4KkwfgOXjR3OI+DLMfl4hWj0xF4r7sLlXjk6Lv2xnMnRLh6LfL7BPK6ClXjTaOReBp28t0fIPO
Crzgqi16+NNtpeAbiknUzc8Hkwxch2s4K6loGSOUoDSwSi+h7/QkLBBZ/ukHW6kyj0Fvc60bu22e
CGQRWchKjeQqmP2n1TIGoSiemDUThJ1QLIk4w54Yh0zTRYrSk+gq/0jqc6vw1Ei6WjI7iak7QVT0
iW8ttIipUB8e2p6ry8wN0wN1gOONOIH7x+kAXBWjOXV/JMSIOdNdOGbrK4AK+LM0tsJxOxsCNqTv
ro7mXYBgLGOwIclcSHH6fws9uKtozSACDqdhA34SSr+UT+LhxSM45w0KeIMrKLAP0XopN8juWc28
Dk6zRKP2i8OGlLMqlHcTyiT6N8LKLfCEl+pBEuQUJCY0WP6LnqxA9X5S6xxxaj6ARalPyR89wtfI
wO6trEgE+nqcS8deBlIz7HaNypUrP7WbIy7jcX8fq7E3MSSYhO0aBV5RzS40lDYTZP+wK/q1TmiP
mHZQFt+di6L+UM+5uKRHm/QVEIYzszEnYUi/0oFjNsQIVNJIK21Xtv7OaiN9PhvgT3hfiL6HgpRa
pmm8+0EQuy6mYf5wUS/b9UzTYWsUqbhlV0JsY4y42H1gslFxEgk5Osd1FOuBdcH3PYSvG3QIEWLl
AMAcuNVjnzvIZNg4Ucux40oy9h6EBM47R6zMTr8OLVhJQSiueG4XvbygljM5uHpKKjQ9esGRBJUo
w3ubvjGyhZ0P3Ejh4B0QrV+YuCMhmiAqIkwu0ala/2nTxEVBZ8plNsbkus03X+MOJENNkyiA4nS0
8iUQmND/mayNkXg6+rhTqoPAc7HpemKO3TLf/OpKSUXJcasSmoZiwunTvXMRPey0r7v85P6HUYP9
eL/chU4vuzgZg1/7PrVEWxlSBOI9rWOhgOSCPLm4b2JDDBSp5MgqcRmrNbeU6Hagw2LFJxjDtzIO
ZTToyUPWasx4SUHV9+i2Bjo+D40kJUaaeKDwDwN/ZBBWiv3blNsO8Fg0DlGZp0cCJM1y7pXQ5RTB
MxVcy8rRwMrtEajJ64uESE7yvM7p5+vFM900rY9iWEl+mi/lre3qOxb/mDp+XGwgVAw/qZT7TndQ
7QgKG9B3A+mt1SMG3ZRj7tq7JNBCfP/F8Z5B/yooHRqwE9jui0qZ+Xd+s3LI9oDDbh4A8TkTfUUk
yq1Jm+wkJnVZO+JR1lu/iHiSnypI6IJuMXL2x5JQrIM/Sk+AxPLVQCl7wcdtkBc0ofv0vb0TKW+G
uYNC0K+T4AhoBUQ1tKegdTMoRMzcDZ8YHWR89pnaJphQCYKaJZzRIFAsWNx9JeKSOVssUjgLkYbB
5/CeCsI01TFNTjOxy2HZzvYJmXtz3rFBb8GkASHjmfFym7qKgZY/a0TEWJTwNWNFinXhqZhbyVYb
ZGQSLCOLfFJjFjL7hKmV+x4R2wKX6G32YIwmH4rkLX2CugxX7CO6qSQQKGCAeuhY2MypsD281/2p
IUDXVDjfkHWjiNLcHcYQPm2DUfLMv9FGIf85Mc5csJIR8IoPH9Ookkd2dgqBpZiyRYgj1X4HhpAz
PWmzUIX/DYlYElDQ8fWdaXI+d8y0oxJRgq+38u7tA07T3qlzP24DHhNM1FPSGsNzzjXbGF1qvOUZ
PbuNPf4ZHodo5tQCkFlrTYJ+Q/PXEdFjHpzArGJ941vKxkyHC82qY55bF3N0Mw2TMnK1eqUJhRPe
gHo4U1n0MIZIv27up/UaVKXqHwBsaR8XOAXmFM4/R5/czgfOSs6BIrtXMPBx9p1UU41Qn1+TJeBt
dwV9bK91XaZRq+doJAc65Mze7pHNktNVd4+QY1VGzN2iKVgHXFMJwILsEKTzBz9LUhZCvMccmou6
7INdRfQYu/Krfgj8va6noMPx+fu/VludCxnqTbeN2f0vAdt06drJxk15vDNJzZqDXBA8JK4MvZh9
GLpGIIG8BIRcb1/q9kc2lGQ1UqGG+ioZATptFxEjb0MctaVHOO85JbNEzrsMmTdvv87UNG3l2X3O
7F6Sm0PwgsHmprYbGCH8/xr6oCwe1nSWiQ304IAAaOMdYlc2QbJWb7899ZnLtYmG7VSkqGnSLBLL
vAv1+cABieNrcMJ9u0eQbqrg/lyPMpKR0lCfQDCokBfjBYAD9abjqc1PYtS5o40q1lQ0bUEdFRWd
4nVKoDnQsQMX3GyUIzEAGMWgwsCyPLI92WIscXV7+Smf/XzzggceyCFKSHqWJQOwd6n20Da3bPic
fCo2LkHbEimZzLb/OpznXxvIZIUtCI7hyzNlRd7ZLekc69Zk3E4JrLcKS4MP9ocqCXt7rjIhljz4
sfaI+bGa0LTSZatjn3Eid9ys9B0r8iwbkOeDCSCr4BoLdv8qm9lfrVoAZpRZQ+Lwa78U0nBhaqWU
4nqEBP/1T6/hpogM4+dbHQ/NfGY2FDfM1ace32cnGTvzz1KemeP9Fd0vNEFRlfeb7T0igRIYos0+
88u9yHcDgpLc+WNvHcLF0ll5Bjm1EVbm1AsT1d0xG10pozsJbx82VTIp/bX1u22FV8k4sWCWnLjW
JFefK7nD+12TsBPrL+NEZNy21RUJ1RnZcpoww7wAtCcVsGgQNWS66NQKPYmh5Rb9yHUp/0BGp9O5
MtDp0WC92aTBuAPaoCysuAKA42SWu+1OTpChW8hwqgF7PCZ/6w6Q/QBev8BGwzgZfusF3lnHw2ak
lbdCggznDrIT3fNVbEkdrYrXLDb6HfNlR05z/T7bXsJ3Ldqk0kM5bm+hl8ofMC462M541ZhmBKtQ
jfPh0nRTnXXM/j1KT5JLiTTAbfQ3Kakww8ch2TpMvSw87qHijvGXs7lBTuMZprYaHsq0y4pHcQVM
DCBGDoX5sgpfpDN3W0NLnTLYmdMquZH5vj6UdoC/peMWkt6f4P1dEVxzZXAapxk9g54bHwi5kT8p
FgEhj8JrID8rE/wd8Te990RYFTYNVt8JHjUXUR0T1DrMIOf6PycIwHTHDrSZYpWTMreOE1vrAQo/
rSfp+TmENDpTwkvUHkshMrpoqDlokdkxeZ6b6XDgdhGCUMSqHwgf/xuRx+SQ8tn96PwSCDsmf8Kc
kFNwocZbFw8ctL5/tofA1M85oIS3vQYT1MqBN41X6zU96GYUy1nSctzg4Ea5gm/XHGctTbLqC7fJ
Zv60jqULd13oGeEyC8z1x6Ck8tZHaCgeoy4BqprE8IHXBPF2jnKDospidhusK2vB2cbd0UGy7oN1
uFFwVlGN/nFrWgUzOrhsvTzOHAftoQdikIZX+iFtUmdn/9l9e7M7aQfKjGzp5Yg1wSImHlbQgD3n
zIQp9+poeZvqsEqZFRdYlWNBs86+xeG9V4OMtL5glBOzTURt1V84VXPymX0WE/P5MzBYkkq93N0c
EFm6vxRlDXGJNiYa672LEuy/A/GE27pFyWMumXxmniZfrXao5S3oWp4fnRH/A6/lyn8W4pTaYAWe
UOuiCEAQNBN+jf/KziU2P4KKYTO61n/bFRcN9Le6I4Y+cnhYJu1nu3si3EPtrwA06bBkymRP0plj
n/gsdY7m8g7bja7O91ka7U67ox+cZbdGCpudwZS+/hGyTM8CgIaIPct1mZKdcjdRE/G1VT+8kvQ+
HNPPXmUelcHk6vAdhTNE3jrQKXnFfq3quRv6VtyuSW5h4FLhWsqwl2rnCQXnt2knd9OSISRhqeWD
ToPNoYLFPRIq8clZ4XZ0UxZM8A/4egk3Oj2fDtP/ciEgjEG9HUgWpfPswll3z6wZLYFnhIkP7qko
KvLWcMioaBBqszdEj2VJ6OMZBqnWSBb/b6zz20osSpQ0yZXYsd1KK9QrTBbGaTZY/DQHHACJxo59
QTcGofpZzxFgC2C6C1UyZwUpTc9Lk7p2WiDLTq2UrZqg2XqpkwVxHefn7j/fq7dAwahW0hqi+Hxf
uNQ9NUk0HzLHGItbpIe5ZoHtBapVUkziqhe4bGUv/jVLOTEExU9IZ657SndMZ6oQ3hykuuFSB2UV
x8w7xNoS5uQhhSm/eF9n781ZkanSexvBfO8poCZtFfqpahttmxrrtTWPhz6QuQ+REpP0zfad5WDf
TwUPQVsSgZBnZMP9i4H5YTw4iE83SYFzGKcdRnx4SA5vUfFjmUwFSfAsr0R5a4OWHxsA6eQ7yZ/p
7r8Nmb0eFGpqR1GdybEXht135disbUna5EjZXFHkSINmR1BzbO8duMy1sh3fSGfTjGH3WdaX2IFy
iSWHdKynQab8RSNxW7uNfrRIBIRobMmFLBl2maDIh/R8yMJk0hqk5i3G9Sl+/IXkamNI+I8Knp2U
9NxCYUto3luj6UZqsI/wjPxbIVCYCvg2xggQsd7bg9HjBGSpmi8oKZjQ3jhiKRErpbs+kRpyDmb5
ofDePjdiuv699K0jrwmyM+DBX2SwgEB+rlD/mODRoqkg4BS3qCxWDLq7nHAgsqu5UC8QEdKWUwnF
t5HR3+zNmvJElcm0j5WHzGZdVjJuI+x1TkjBQ51GH26vzXaQM5DRmA+fUJH+zpVhcobto+YucwPz
iPp2lmdktC1GDzWGRoFAgtpVO7MHZe9gmvBJH5KWDHeDaKy6CAwOUwvdTWJjBK2SSh2NUT1N0pkG
VhSW69zm4XizlAP6qlwhfwHaK+1M6+F1rCojNf38yRWTWfTbibyiY8u73wXvVyiezcmmN3Xl7lbM
9CXB8YUYHyAIxAg/1SGMs9AtZCaRvzJrl7PnWA2O7yAoZ5s9582RWea9vN2CzPud/S/Yd6OCX3ZL
vLsUv4ynJrNzGGAt4lWh22dH8mktf+283APoVh7YuHmzruwbE3Q5zNFg2LwjoB59jd8dBAZVJNam
BPL5UeD/OWHjDLdOzyIKHDGMSwd4NlnEK7UToz+y+4vISZEr6pdx+LJKp2043lOMEaXfRzJRGAEw
qy3TIJaa1+QDMj6OswPq8dZHImwOMXpuhd3pcTb6qkTdvr6Iok+0S/PaXi5siQbAXVIDITJuc1iH
32jm09TYp9S4nmVSo2y1xoIOkG+ukXqdDXWocK9AceyS3Pp6eLRD4et2/pbUbJ93ECi2OnuT+Hu8
1gps5NfduTNhEVfYEFIoF0YBZxMPRhhg/Bs/NAtSdOAdRbEi+zkZ728GY5K2JnwGHKILiFV79Fr4
TSIHfRHpnPxSShGhPeh1UnB5XNsqS6GD4coIozGAnrTEXdgX9SYP7P+XZ6nH1dDbEDNOQZUqKZ+Q
agXS1Gr5U82yNbcgtqgLkUIvygQOj/RaQWjmSDNu696RR0yAEINzsJJxGo8RMWxqbtvEqvvTswGg
6H/s69gTnywxxXeY6MwbfaPnTziGJcDCaglzVcztH4Smkf+QMJCZFteBUvJyoKFX+13AQoFHB9ou
W0wJA3tL8ZQOfgEZJijAxvUwnT+9cikOsOn0hzNP9NzNcaktq9QLet8J6s3/W8hwqT9G3yY5rceh
hV8vWWT75UxsX9I5BjLTGyPW/10ohdf01Lx4cBpnZSghl69+kPGsgaGVhS2NIsB1THyQZgSHNj4U
m8vGc4QOkq7nAcO/2BC4EIh3i+BeWljFIjO0EzKczIxynLmA7KpPAhZ5GYt0MJj5DdzMrqkR9B2f
mq8dqEoaFsFLDirwj/LIY6oV1yxREggwC4z7JE4qbudJNP55Azx7KvBEwdPX52BvL2CdLHISwysY
nmexr4CfvsbLsXvO5mSdfH7nC0E0NOm8sCyX05ZRCIHgxEriGYgLaLiVHzLOCTPCAGRgi9DfMX1I
laNP3TdCm1IdeG+Cj5LIzwIA/FTYhqzfi1EMYN0PCjGN/6cr+lR/kEAb/IuOrZL0Qvma43FvN7Vw
z7UP7YoNQSU3X6L/PVXWJY7jUdgAKnH6KIOaLKLkn3Y7M66cvS0ZqG/MosSEcO/2tAlMl/2Aj/Kv
mgU2QpGDVGYL+1lAM8hXnCeQQ89apkDwdzYer1Q5fYrqT86d7f2T4DxyrpzbeLXcatB3+iWFzkfK
PcKzgmzSpaBFtmZGe9FZsD7QNIg5QjULEKTOKJ+oz+4/WwLDEIAZljDhGS3dm/s79ZlOupsWZA1g
nmBFdBVvwNPtI24DTHZs2D1s3Sv9hhAvoCI+tuInnjZYLgu3u833DThAW45pj/LAWa5j2oF+0tJ4
Gs941O16/OC5QUC/ifAJnQGrh53ckUp87rEhEMFFQvkWkIaoHdG6TFb8XrS6tEwW8Obnqjb45QdQ
LA6SSv2Bonrvgm6yvWuyJrwrQAMnHiupmHKTCm/uoaAeeWzGWS3DyTvHeAFkTqlGP9ZkKbI86Cc5
Kz/B3wdIIA47YHsPwjPgtIT0Ci0HqOVKYAFhdwbjrq7benOuRLjyuO/r4cxhVfFut75DBJwdCfRd
0D2Tn61mJxgS35bXPugNQ/JLCFwSn6yCc9PpPfXHx7WXknNx91utxvzYCJkq2Vi//PDdMtw4OCNJ
pC2tQGpFWDLP1Yz0hIaUcZPalJjFyCkBc6UNx9VjDMiEeE+mn+wbblompnTw6jVH4O2he5bChGRo
IvEoZKfTTIRGvLV2yjsMmjiesgprRypNya1sbhS3YEO22N/koYpMepdVHjf9kwHuED/T+tcfYZPv
OrdfZZ5oi05Plb7aJH5Q8vulVIBPBjP9ciMo2wmTeV+WO2y8r1EWXixb0nVIfXpCkWnhdojK7LW7
Aw8ev6FcBlty+ZifMCAC2SL2HvLcW7zX3PaZ+WVqwFL+ZL+fdL7Uuy4RLWJA62Yqw0RA7hXzd3YM
b7V5B4F6iYKG55qfkOfoqokkmx0SXVq/c+qBRFc0/yyeazHQrVWx35uJoR4EGYiqpQwcZG5lD0Hi
8EZZWioDqcarQlp2ydSDrVmnqYPctsTO25wIPk8tVvIZ/j/0NYUi3kCFCWLG9rwTb/92/8XP+v2k
3Ko7SAkkOd5TrvZVSmYuYD7NStp0YtKFUjteMreurecDW6PCECQtQHYddPARWDFhBZeN26l3zjbV
/NrH9sHt0ik51elBRtoW0xMc6pRz02cmzO/2kKzShO7o85b5gQHRYhD8jaLC0I4qq5WjTCFzCMjb
1Mp9TbipIE/xmMvmGhze512kGLfLToRd87fZyv55in6fHT5d1KOWawVNxr0+Y1s2StmicyeQzv+n
2YI6Um6AUb7ucl5FqLoz7EatTJs0BIyOtCqmdnVI00QJQ/v4/WERta6Ik2qM+2Bv3yVgDkKgAQ0s
Q6H33guw8pBEHqZSU3qQR/b54zZyq1pkGrZgacbQ/yWU3e8osNccBezsWtJOw0ydqrDcBGUD78Ij
DZeqxa2BtxLGRaTNvSzgkvMLZ4AwF53KxeYfNVsaBYYZQTMMpZo5KZEsYsN/Otp/uQI1i47i2Ke0
ToMXxvOWbhquzh5XIF6JQnzkSz71GZy1Bw1mXVVOyg50gVFoNQOoZ0NB/Pa8HZcVxuw52+UPqgEb
+e5XjP8MVtD1oBiZvJgr0fV6QlFFOSP7bl8m/CT192skTCcZ3jnpZF7pf4aHOzReLUafJ6LJjgrL
gUWb0BtKwMG4WlTRAK9lPNrqpDEtbm1WGrYv3vcRrpcc5wFCcm0Qq/tch6rjKDVtF4te6two10tI
irmhQygjAVH4jTPlYOm9ByHBkIt/1PdYEVGZb7aqwdo461QopS0Bzb/Tr2VWocj1hrMJzYXBr8CY
IpjliMuyXAjU07Pyi0dwU3dpxfXVg+KaX9+LotYQJUvFJvykEYkbDhK6JHMHPigYECmZHy+0zth4
IvO1JVeujm62mLh8IYCaL+UhXPgt2QKas9lnvl0Uqm25W9veHOsiWCGhN9GqnMTwU7aUA3mLOfzH
V/y03cD5n+RaGxr+4bgR/h3B4c9vFvxaLEf8gZS2qTF4V5HOmdOkoMQrOH/pA93T7K09DS0QvcMb
6dp9KL0+iFVLfci5sILB5Sy05NKWgX3kgfh8r7axR/RTV2jG3XsvZIhAhwtg8oh/N+Ujt7WRAiWr
s63LFgVXmEJwTiouUfP/7KIjH/P1vfhdPFhVFviUnizYfCXetqSdlQTa9O99dRE953/dbrjSCO40
tNNKXhN1f/Tzl6CTBuoBXo4GjQIffegSGU3h2MfBSfkpmTIADBF4Y8yjHwB/wPD+ccD0HuZNLthy
AiAbQvp4619kB3LV9X32nYbnUP/bAAZGy3KFeS9fN6FRGEv88O/n+ICPBiSg35HVByfIvhns02Eu
LUU6TP3FDpUJMEf35k1U8DPKu6cao9J/UYZICJOjGzU/8xJeZypBzJztzzrijeqc3IWMbDdCRlke
iFWWC7+sVQWoB4uzRDv7KZZYhkhXhp+laJevl3nOgvmwNjlRLHS/V4lG1uUzKfbZxxtUsFsG6g9N
jBzup4ZH5e1OGIL0PTEHP+MpcPH4QHQw0/STGFIBefMJe1Fe+OvdW3Xd9Lf2MfMR+ARHQCCDmw/F
gj8RPHRXBACY99LbUJYtdEAi4d2Itw1DVA4ulQX27vZGXUOKX4T+cz9+BQH1AhKMaQMlvPXUq4hX
FybwVHRiUZz9f6CP8RyiPXRIn424QRxt5cpmzLxjC8eBdsCIbE4SyFFxjWtdgT2v6mtWUZt589lt
AqN1vHrseWjZHcyumQtVhfGJfxoXtZs6kRSQ8MlFDyzuu5cfNJBTeQl9SUDI17RIWnMIPmQ1rUem
Hq6OLrOPMeMu1PZ4MiQryjkCy4eDu5CqcZCHLIOUzikxAs+qzLxjbXMZDRRymzI5ecGABvlN61lq
n3zFJHQ2ul0PRNyGdAGPv5KrYWNXwNu7qwGRbvbUUdyWqMe1EMbCYCJLiwfsfDcfWRg2dtumg4GJ
OozLDfVOGbf8WHxTOflmvXKdjm0X1Jfprt06dIVZUC89CIhny93la/u4LTg4pmvqjbbHCWZ0EZAs
V0k8w5ZtqagzGEA4J/JcIiCx3lwFcDJUI1G7z+qoEDrxqqaCLreWsFqOn28amvlB77Nu18f05Xt0
Vq+1+tWC922/JiU90Bd3b0o0gHD14SmPeRR0v8EI8300+WMAMH2y6Cpsyz07viYzhB574uJxL0Is
wUUK5z4f7aHPSirPWVS2rYTWa6jSzIIX2lswFV3aftujL6mJ8RPv9grvu5T5f/i7+6VmHhEffq9n
2prg8zQfLor9ep6yt9cfSAL32kuz8F6N1PAKyIjDep2dXB2vfwRSlrGaQ0HD5VMIBpcaLiCUXn+n
WP2hc2PEEA9pbzT33/FJIC1BmGeofKYrJME4m4fnzmBzKauOAxC+ABcdYFh05sChyYEVoGLc6Jgm
iBhDAz4ZRDX+SI6Zgxhq5/76C7tFSa9Rob2dwKiwNFZZ4jT1AhaC040+FyK0M3l1/d964uq1fpqV
OAQ4SW7WrYpBo+gsgbiUBDbroTZFntSPwvJiK0zX6ie4thmuc03qdV4WoJ4IXv5Bia/tQaB1EQ7z
wwo+dyn734se22JhMX4iiSDjJGMDw68lRnhWw+VI32XdfK/1iVMUllxRfya2s4UkX996oF2WYi47
r0y0Oubxzjk0KrO0K6SY7kt3t4Zeqgj4dPlRJjx5NeNNBROB56nwUzxAJQCVpZv/b/vyPPEygLoM
4W/9D6HzAkcxNIwqPfBxXpz37bl67n2KY7x/sq1bP7tdryt02awc/EeIzx9vQWAPodtKfnbRt61b
x5UdNg/vrVCJpV698QY78Gj4AdV3HYTy4Q9yOzryzjcUmFe+WgoljNPHt5NT2u5+eLaaePZ6sDlw
v1K3KJqXKnN9A5XgJaDN96Vzt8i7Rk9MpMa/CzThXr6PI+Siv5AVnl2WcorzFPwHdciC2UJs9uM7
ZeFa3zCQCWM+YZFq+GH0lKA9ujm+lXATAGU3IvZheZt/tsRhWO9HIRVYn6Vm/lKrsuyl7lADhSsi
NdutBMN525KLzRYh/VoQT4kcqHvQ7OwP/KhMg4n9iWqwRP/PtLTR/h6d+D0PuVwP+QiprcpzKm4u
+BzDR9d0VHP/gZs2W9VWKpAZs+8lo/7NsqnJSVq/naNbpC0bMHiKPCtbi29CnlJZGKes8ekYIi3j
tQclUASP+UIsipxfKCHg0qhI+I+2Nv79e8sU7gBHL4313rqQATaoX2QBa2RFAg2S/gYqheORI0Fo
oDG/+XoyObycEtp+Ep/WeUxWfGLfkwdD1VlGSmDbRJgxTl7Z+eDRpLZQlH5gma9dDBx/rOV/2QMe
sATu/6y4PMwX9NpTY3AOCX5/JZk+1/EuiFsl46oRk6a1Oh6nduTedb9fUqeC//Zr+7XW7n1/8ISc
OThtghw0DW/YzxNwrmhrFonuoxYa5vYD6RZIJHpeyl4ZtpCCc1V2YoKrj8ikXsLvSECJKe9SdND3
3yFHXf8+D/47KxtW3jDpK6Af/orGoKgOovcf5dTXIthpSBFRDdPagSjI/vidhKe61LSqBMC+jY2w
O9h8VIv/W/u02lldVNCNUs2fDUIq4OGWFdPDkocjEQtfsJYW9RdUWJg5ThPimIUb04zv/BgdIFm3
Svk5LRcOYAj94UOwk6YYHHH/qbVUgjHIDx2O/X7xrtC3PDrsgYgYJMwV2N2P0b1cmxt/w2ngXe4/
YX24G84ItlvXTgLt2kzlKZKB4h7ne7SLez2d27047PrZTfi5TgCvxZusztYEMKH8W8oW1JhlOPGc
OCezxnF+JV5DTGkrgfyqPV54roPbWekvSEVOMa8Gj/t3MvKBpCMEMKw19QnYkejKZlw2sGA+nQhw
QvOuar2+3XiForzP71BRjvQy/6V7pudWS7oaALvZd/kaf3sdZAxixS1KlZzFKU9g4sHwmOgkPlYE
EtHrIQsII9i8J+bhDbig8LUp4QQPtmY6KhnNNyf9YXq1KPT4qF91IWc7hpnmEJYPg/WrtTocEVs/
h3TVOBaiQPykKJzHSH46d1xotCij4cFPYi3MOfyaJoirtQjSTDdwJiqeKV4e5aOfksSwlJkPJFcY
3AvVo6+qDNY0Fv4BwskaJpj3I/z2ouP+HXySXMQa/wfmeyuTBK+P5febV+se488ZfP7r7NohYOfl
+ONs5eE0svcq/JblBMhVx9OIQ0jePFUbK8iZx0nPsEysEc6YSzjKiGq1i323T1kFKmKHJ3G4hQhi
bzBQn+cSu8c9PS6J0bYqWLoUt8LjsE4O569m0xwSxEFNSOAXe4MyaW65b9g4bIVPwY1fKxhcdPF9
+SuRr8fgOV+AVNNgy/cNw/l74/LIvWSv8Km/KpIaCT0Ed19PZKxTQ6jW+oYmSfVTnKrO5f8WX/8R
WoYZOL78xz1fXmMBVy3oDkCozWBjgfHePKCVXEuRJ7L7hC9gdbLy0WzoF81AuwF4FzHMAwZSSGN8
VVF9Y0hRzQowsEvVnY90EzgegWhUFX+Uz9O7pL04x2640/UqHKHKNnamCRaxJUEQ2tVMv6gZy0sy
+vvGk1EV4s+XFABXIKiGrEs8cEW3U+jocxSwrB875AY4B+DkfFcNaK2FSzvMo7XckFYeEzo+bl5a
40PgrcpWcZE4f0MQDwMhIbvwVR+sGPTjMA4WWJCyGnIOBXoUBzCB+bbAfEsKJkziET8BlFTqUVRz
cfk29s1+UqG1NlEMWnEXK6E/bSCXstYZ7oyso3HB9N6mqr460twF1fyx8ESSzutkb/YPvtNQU3On
8Ei6LPymgH+LTS9g3ZYQYRR1PCn36BVEEOfuIJF8f5QEVSTJOwLRcyg3dTxcbKkPv3AuU01acFxK
Pgqdvm6ux9ELNHSUlMq3cd6LV/7d/gtQXQkF2/s2Q4WdbK0E5oN7iMInT64faXFapIg9DL0bqWQV
ONHe7+oidlzMfWudM6p0gg6W0ZfBINrNEVG1Hy4Nq41vlYlvKyJW9TyZnrLV/Rhoz8Z1trDSjbS+
0CF/K2QVMRhVP7W/l8hf3CdpsEHlcaoV7lNC715FoEtVww9P+3I0TzwbDsPjXIaNIsC2nqvZMxmN
J9iMVHOt5M1bBngwDWTriBHl2KQfroEyx5jdUs1QzkV/V2X8baYvWMCGC3aUI7W19iU9qK/QYmhb
phazr7/gMPGbBs3S1G4i2jAkPMzQSncLsZT51ZjbI3F4tFDT99mnk3YhKevO+Buh3Zh67d+1UXQJ
yErfC0/v6VnBmhxqxhD0/cLpS8lfsRXcOoHYOFuZoRHvqYgjQtN3VGL7TeYRvkpiNHrBWSJL91bU
RDc1WFUOes11mBscZ00Waqr3aknsrTETj5glK5id6IG5s2JsmaGvCuNCx3cXZDeI/PCmazQ8vDTE
kFaxxdwJ7Wf5cd9wqnJABLCk8+ATK/k6PhVLapfORhvf85BkI751eHlNc4P8wwwc3dLz/uqYkzne
1js8JUi6pykEciAHrSa6XJwRwb7g17XsGV6vrNa2cv0F7fkbolUkFauQA7NkRTGEs2uB6LJ5EwBV
j3yb27aLv3xoyQw9HYzJ+Mh6gKgzQu6Ksij1o7torkDs7Z0JYTukXZJBsGXM/9hKA61SVXJGaFSP
EEpEbRNCeTZS7QApBggtLVriTtXRyKG5lTJs5TR/0oBLsaynGydf+LfNms9ZcDnOtNrjJUnK0mfa
/MP02KbevatM3yEHOQsVLwCKg+3s8DMoNIJqH8uRc79TI8FPHX4WB44JaI6rwwIPYbkGqRQIZDI/
f5X0i9eCXOoPN1YLYtxk9VB5N0doVuztiH/puRaiISoBeKPNxVNNmq5PeSzp7rX0uUrcHzysLYEz
tWW1Wn/0Ol44XzTzbDEbeNCub13T7RPCyAX5dXqx5/uywRUKfz/iiukmIHnzEZkC49SF16GLdq/G
wryoByqj171RLYZMFB/fnthutFRH9yRBq8J7LOVUbXvz6V0EADTYTrUwZu46qaaHlnS+O8Iv/tA3
1YqCpEd4OvVgpahWDIHfzj1sZqDEcAnLE5XhLExBOKaz+392gnrNsZCkcd4+/GMoPelsv/BrPBan
nLik3IIVgfBGot3DgEha+Ie41dsIudv79KxnB1pQBpQa+A8pGbW+FooyjH/E3/7g1JTzG7HgSsjv
h/8AjuUQOcpFiWQN+4f9pcM1vn9tgCeUL0wTN43cURjl8xcyhdHFNzypfztRhIvvGR1k2lCnr2Tz
zna7fgMsVIxEUzuHACZJZRkKTuso/OlA/BiYGfBYoObC6XvubvsSl1WnCLbP4xPsdJa6JEUC0BA3
AwYdwrmB0ii48h54/v6dsa4fDOvXLA+oxV8vB3LM1c9iQgu9ZZ/zvVE7qcrZgH0naJeoCnGgVNSb
rKXrOM2aENXvSV4YdWjXx1476aH+7ohYQOt7RjxOLsvr9IlKOtLYAYQa1TwyGNSw9gzQ+uSMaO7H
whN5CUlejztVA5oMxbDq98LSmL2p6bpLGxN8U5DUCwDWyVnJxAx1Eu4mxS9EpnMLmYo2v4QYyIdT
g90TIyS/jme7sYzuPhO39Ny1kHvGfnFDVCjcv2Er0TG/fCH76oksLWfz0xIQY6ol5Jl5XAyuDUW1
CPltxrh3D3NW+9hCTnhjtc9jRo7T8x1CnKw0lmBXMTw0RAZ9mtsUrps+RBGL9KjdJoud0YrCPtht
ffmeqoPDspq3e5mF0I2b3QraxjLDwsKquDu1M+wiTRgf1VpPmXGLXRv5uDHd9T4D+zvgKKZtd0DJ
rMnupxirMVNnRkqwnlhfYpuzQ+ZkDoMpcQBbtrEeBBtZfJTWybX44dp6uWWj7MMBiNq9BWJuTCWV
HrCi/2NSuv0Tt87gEceSW/jcqPoov8BvybgjM1py0PPwfX425n5p5Ulx3Xc0CtVqLXksQG+cl4f2
2I++K5mKfV68dRlHRIPa/XjPTuaV6LZBwP4h5CoF8dAx6lvpBJ6+gLg0gkL3f4L4mDI3cCcShYiN
4an1HxOhCULn4rIxoqFYpZ5QUWZfsCFiov5wD7+y0eY9+5R+MDVbmSMEVf9DCdfr7VBIZYWd67QB
bNiX9m3y6Mx34iA4+gGdAUWep7+joNXiNZ97Mi38bapRkeVu2Mwx6/6rO6u9VhWW2jEa0BuIszVB
AA7SKRUTBN1DxegTBrC2Kd/OG9ns6+f9SnL7cO8cH8ang67cxMmBWIYu56wzhzy8eoHVpYYpNgEA
S8hy0PMxOLRvwZCv1W+i7C7zZHWPpxsWZ5tCXJK0tyGATfSVf0dhDxZK1Wh86RGQ8XStpmg8NWPC
rLXLyj/i4wZKkZ50kpLzXmahaug65xWnhpLxRxRjFyqvDjISm2gRxeY/oqYPWOFJL5OCqYYa5Rj1
skUA8logg4ZZJTQ5TCKkS809jMmpo2uRHKOOSn2vts77ObPDWgbrXbr18vWhPowFCeVvE2YLC0SM
Voiec5OBCaXF8pjKkWv2QsTU59NM8OY7Qf9EIlpV4qr6ehofNvJAcNh1Ca4ys97H7aodwJzlkO+6
CCY6z0q5MaraUx91eqNrfNJD/hrltpI/iEL87vTd4JNKyxpqGhrxTNNLrsBOmGR87WG2hi7tn427
IGPyNv7SdzKvJzmF93wRMiaGVNIJ8vaxyE4Gn6MTRQBmaDeZGuiVpvsNgf444al4B9P0aWaphAbm
BaVvDZpdSMmuLZJwC/HbMLUs50VWx4Wo4AHF8ytLECeC2Dln/l1ihGJnxdo38wwSz5y/oLHhmlGN
3YZqmPCtl/jeJSDun3wpTQTdTQ+n3lM4aulyu3DOHJFRrkGBg4R9EghrRBBPOpyxfJ9h4F0FqzpG
S0uLQD2z3MGzv7HWsqOigOfPGGwRHcqyk35lObhyP/NL+mDvGoOydmLXSaH6jiwFNCWtfEJGMXqT
bEhB9b6Xhb0Axuzrzb5GTMhDH5dL8LKzLDIxmtn/7zwlJauJB7w8MxXMi57Y3d23SqjTucfYeErv
LXrq937iqKUhOuIvRh12dIyZ1LNB6WQMOazc5yB5JSrNZALU6/mRnmdUyMZqeNVOag/hhIV/vnqu
YWgpvR0bj1u0eDGxuSctSS1Bej7PqMXF+BasQA0uoCYbQQNB+i951K9ALdbq8NwsgT5Q0JUZDwpQ
QABZ0UdF1OjgcBa020c821oY0UIc03QlI54tf8ZhRL5+X7tpzbwFdQTXoquKygZPiS9mbQ8g+pRF
kcmXctefc+38EARlkM42zc11ZEElF2gq5N4AQhKlVeV6NMrV8MoTB3WjVIo96f3qzRcAXRPsYx1N
uHf3THpxXkMfV5pbxa1cUzAXkIHdmBAPGnf9IHklocR/jWDmUe73GFRLHrjEj9UFU4hmbe+ofoBl
tCS7imFaEGyp/ugc4K4hEG/b4zfR5gfwUR9/pe5Tk8TLKs9SpJE4PG+hVvTrJZMfTVuGomk4tOlA
aqnbXOoWCX3EY2+bC2X9CfPu8KvAgrLeYchw3Fey0Y8oHJNTfu/0mCuDWYTB00YCReOXaE+8ZjS+
Dxzm2trGWR0qT9H+YPWk6FpwD25yWoPEnLPvyieRfkBaDCW+DOaH2gLpFJ2+CVAAnVqqpslwbzIw
bqdwqvyS/WTRE7o9LPPCIXdFLd/v6ZNR9Dyxxde+3hLZ6xhtXqAgShK+J0K5tnxTw3s70kprqVqb
3nRgS7FDNqN4tlK2/uIilwryKOa9MFXHRPSmvIX8Y80nc4Bd0uKCFWrmB1ORTVEknrvFcPwQFxmX
AHy++j2FJD//OA7jc2qolTrUBYZCWzC6RJ+d2jWOS7+i9ZUC65h0X7Gy7Mbx7ouB3yKk4O3QXmxv
khg2uJmrUg/qXMOscgmu1dzuA25Bm89R1kQGo/oFwPwtuuxX1LHhBXneXNnvBonLEtabiyXfWNgm
KkDk95ZnVAF7mYv6F89pMyxZPN/3I3hLM5K0Uq9TNjI1XzNhjJVaGFGPVIW2QT9uLDAxwlBL4l3t
jUdwnwD1Zum2OjPVykyYYaCjuXoGrZIroYA23+DYtfaUU6HLEV10wA9VOSM1h+otcNEnqp8A/8d9
7h3MASS2zdG18qXYf4B7EM0/w/ipA9PfqkH+0EpAqGxGtrnobvzArhewJ58+wfSvgVdrsFZ358yS
/F1jivqIdbKGrSTyUgmarsNzI8DVfFda/jNkk31Pkk1JraHaMPh77kwHOqkojBhwWYQqqBJi9pIt
1bL2VYlvggXXt5fUsHskjk1AQ23SPgNrdzrghdYWXONNWLnHJdHljxcLrFbUYcU+nKeo1BhjeyQL
CCZrzd/5zrrkMcY9V4U+KSs2j/zN7KUhQFIA6vzK3yX08lcRQqg9TEtuBg3NId5gmv6yLCQUyxUo
c4Jz15d2mzYOXLcrUxjTfGY+6D32kW1Ggp5pMkr5wRXVN7lA4n/EUQI/yNLJ2V/0nhmk6T5vQ0+Q
6JvuMySi6+RpJ4XkgvnB9wIPSaD+VSujzDGOiKrx6SrCjB6GTkh/jbnuEbzDoZ5QC9OqjiQNHVp6
zriQa/ejKn6CiILkQcaXXJbegHIYhQ0QGpFou/yAMMwAiqv4ptMvtotRQ9GkevP/kkiPFnLlawlB
x0BXCxwRHyzX0aXsFGdfpyhjp0IRV+RK9TpYF94P6zVokg/0EOemo8FUMYWocLRceeOjBKb6Opho
DNY5KYOCTjIwOgF7VAIewqm4jPZiMeu9q7OVazGYmeg54PQUPuy3c4b7A1wM4I3J4TUoQ+9/RuRn
w7u6neAmF7T6AGjouHi1WQTrSBSodzLuVwSLnq4gl93YxAmvG4OUvFngVMv8lZz9c+6OQcv+6mkB
FQOh5le1Z+kDiZ/nHK/TND/h7nUUrqZRXlPv/8zEvPqfXmPtTbrCi9gxYDtU0NbIw0zf9A+YhKbD
K26gquvYm//tNywtpf4NgnANuTpF5zOpYwJZBuNtbRK/ijFcFdbaJxTYSGjJHUeOGGTbK5H7oHLf
vnoXIdvJUi8z61eSHTaCQxCaiHEa9Hyqf/0kRpDn+ec7NfulcIWb4KY9pqO/tUp345G/l+ycT5il
7wpKT1vQMOSGMRC2NZ+fPIZurL6iuQfjrngK1yrfu2QvHIPKJ3nDZu7yX7OeY6CWxPwu0KK/cC8n
CB1RIuuAIybSCQYU7RvnKkOlfqhXfFSdE2z9nZl+h9Ag5kj8AHjqPURv7n18NJmALbkTnp8XgyPj
RTuNes9FpzHKY6RaEXoj6/rFdeiLWFP05SmquxIQhX0ycja9gDGdL25kIVO1wTi4bCHcVxRxEXUx
4+j1aEX1N3Z4RA7gnHv5adaQiQOQLhYviyuS6G5JA1jx2NutZfXd8Zrla8+DpwebfE32FnHeL7Rw
NNNDsDgQ6Sc9+bpojENMdgk06MprsQq6mSyG1esebo+FjKr9Cjs3zxfhZZ4kC0WdJc8E6mA4Z5pa
xXAMbO4C3xYh/EtEeQ27/LNWU0t84pKy6PHarr3wnmN5XKiaGCAgknzf3mAbyOskV36AWk0QLh65
XGmvCAZAt1LXl6AjCu8QhO9AAwR4vA+/0lhOl5OFgdKKt1bXABl44Lq4GZ8ViqLk3hORhoJCqd8U
+SgAONcKV7AFWu14cG63N6zja/q3nRYospnHqcORcpTgPogpj8FODyf0wR/YKJzdAvzvsVM4IziP
2Qc0J/T0xXhbOisW08kdsPhrOLbSAvuxWPOE9mqBi0cqf8aPsDxF9uO+qqcKWiXfdXT9e/8wUxir
p6br4RhMWhLm3Hzh+mBIavey1Lko8Cq+KPeBr9L3NUZkg2MNiN9qciv9lqDiwNAzREnPVV4Dc8qG
hEse8taeeVhDeWtqR8XyQ9zab4WzDVHmOx12b7ZSDmT9WEbe/6+e+7eLo0zWy/MGLoIrz8W7ITi8
YV8CGukA922MkP/ZshFiKmkl3yrHxguN/HKHXTFkatSC72um8ZNEE1zXrZSJAlQvZD2FxG0qAhaT
/WouZ+9ZhTB+jhyAZpNNnQ/pyQ7zL/eaOftHcGWopBljCpzKYGzWjxygkX63GXhKIVWy7uaeTDA1
RPRaHdsYLolq+hKxCiAQp+lwc26IITE10wBp3kPdu8tqF/kj1e179tPjPE6RPt/1iS6P0I+9Ja0F
Spj/CcedlCmZ0VNF9o/zTRTdAVYbIxAxExAxRRdRS/xjMGVIC9C75X5xCf/Ylaq1K24SHYPR7XOH
TthaUEoGrDFbgeoRgwNVDBnccHUJosNqMIs2F21YOKfFLXghQDHh0ltvkK0daI9lFdmRpIDJBFa2
GupkmLkt4eyz59dSoDHvJ7FOLYAYiwXtm77CU6tdFflEbgp/kU3v/ixt4RLASDKhYzd3usQCVJNv
zfghUnWn0dWHQKeMSkmtH0LQ4QDlpXvOPW8BpTah3vTmTcS+HMRxIiq57lLQ9H7OG1znYJltFFq5
DGxW7OwbcIAPizpoheP2AJN3BP7uPKACh9Ynjnq8jrq3O52ZW5l3IPblR1h5N8mHNnsJLcRNVCVD
MwVtwSSeDcFD/YFa9FFS6y9MpUo+aRDSqp8Z1ae0ooK1fcT3yzzta6xj1GLiIQPiEVbIhKXWwSoH
YXz5MIh89pDljpiZ86MhGeLoB2PSb1a5nJGqVF4TprLYSzzGYWB/6enzbIpwGAhBuGAmGrJMOTAb
ipXCfCPAJO5w76us8Sa1XuI4dVbHX3SPYnGNh2Xs/ZHZXIxaFrFXixxIt24M0pBcPLA0cvHUMgj4
5OI9doKZ5PghXH6pYl6X43dnuIUUxojw7aLlU2YrBVPJiboGWe5BRtc4JyGP4Fl1FfUBaJ/lcWDw
iN6WmIVdF3KAFF50wKRXAi+Gr6VH9g2QkOPac83kcvlw8FaaYktl0ze5xs9lE4KiIW6XF0qXVD9O
D1gfUL91JgvTVBZaSw5YsiDjsnrBjI31jRyoTx0YbwkFJ4JEWb9vTXfqyQMhHQnVR5u5RWalSmoy
kb3lgCcfuzQ4/faofrBqqtHZF+JTfSFv5vRWd6W+8T/zCtYtbc5pkK7j9iKVPvSvemdFH2PhjJNs
dOFacPOhiuxxi53km7uF+HnPSuIal9C1DEc8cPfYYHT+xFaIoPwGFmu9k9pRWemx2Kz6MZJelJrJ
FYE54FLdwzg8+HJM6xVtppBJQYPhslebDu2sk0v1HWdeqZ6cCwh5OxOgDT/IAzH4NChJfdAV/Ohz
k95UU2OVvUwWKsv7HDtYaHOWPww3n15eIe4QPbFEuL7PRLKriTRoch8Fru4sWEeRFc/Y5z1vkotW
Az/ADzMptBD9wDFGSXgP+iE8NQZI9/Qyxvhve3vBm3gLHe4IypqZJEXbauyGVtC7guRaweFrwRuN
IW1R3guLSvC73cV5hZzoaHRkwwnypgFPWOoub8TH5fspTq/XFBtoavNrG4y7ULRv6f/I0B40QgoK
QkuPQjbxYtHWnD58fmRXXcEMi29mNtd5s4mfjXCgh+mEdUCeMif5A+kUjm9LE5+7qqBe+EhH/TTy
/5+QxgjeNP9yJIU0YQAuT/qvhYqObYSPAJyiv8S3uOjH4DwCAuqGUWDlaqbeg4C/1A53B1/Xx32q
oNI3UoeEA+qTUNfDMH9Hy5Un+4/aL7WGLJzmfM9uGc62iYphWbIxJFWoHSRev3wA9hw8SX4kxPt2
DPPa4WGJkEXfS+S4K9j3kpdBgkZ0IOyEAeOlhd2UKFl3CmYK9XwY+quqOUGiV6CjE3cHNrpAbo6V
APRvLhYp8o0u6S+PK570gUYrWLfNeJpepyg90REusby9YruljXX9K2O309UiadK1+Fo/+rC6D8xc
OwpunndVWfSp3Zvq8Y4Jn0bu+HS74XJSbsSpozRO8v9AedE70V7WyZ8Z/2QRUkMsTAPCYIukObSF
ZWS/OwwhvYu146+Dmzyowmg4EtuzDJahbp+yKevccX+fxeeRTjckHAaayOoRPbejteRoUj7fU9kM
4243b4v/IW+P6kyL1Yq2yZ3Q876VtRW4YLWjsRtEa1N8b9beqpoZxOD7zflexwkBZTIjYBk7U+Dn
2210EQdgC6M0Bno0svuYzki88OONuYW6H9hTR1nqkbL0+abmpiKZMewvQlYxHUBDZjhA+nK8aRDY
/DKtkKOPZ4YAvGSV17IZrBwlwIzt2ARFyANNEksUjc4kbqpXRdZAGpVidYeQXjBWzo1w3FsKFbee
AQ44MaWekX6QfpRzYM74N+sArKT/qvM+i7awuafx1oh8Q5DyMM0F34s7NGW8cBVA2WO6iE56CQAA
eNBblBxVD0nlVoEbFYXjUE1nKMu6DByun1eHfSR+xrGg9JzqPIs58xmqxBKy5YkDrctlJpUDjNJh
TGwPXMqm2gHezXgOOukxzXRbncOrJ0Llivs+xPN0zbLillS5xqAUjKV2qhTdPKIHqYSh42rpFFtf
adu+i047NlpJrAIkgb+F2RcuAlm+8Gnaw3yBpxtiMqUYT8p7o1lZM3nXaQa4DMjnMqOEWdrn9HiS
KeQTacfhNN5P9RdR/SolwFertJ1l6uKjcX1ffJYTbMhSmJHdYadqwp0IZlS3HqYxynFhyz2rnpix
bQ6+jIWQAKMAYQsxfArCd5P1Na5OtjFQNvjEPj8JebUylWaaNqB9ej43oM+BIvI5Lh4+zTmKQZYf
YE8rujYG6sr958kMNdFwXPvMyut2Jm6Ach53/wO7EqOW9Fg03J2NJckJT+IuYORUX7Wce29a3fac
flCynbDMD5Wa6Z4EzaBsGvoqKez0wSxFAXO0XJqeWYovfyTbx7kZrlllW4mi7Y005gBK8eKzJPEr
1gEg8/dLO/vwflRw9jggbcP+bUFRwzrwB2DSYDdqztX+2JIDWcAO3H4M6kc2s8lsnOSRYo3GiImN
Epu2YiSDCEdlx6fDN48BNfMYJD2TvGLZv7oyWXsexBuPlKfOYnppgCldba8GA+YWZgwtZ/95X0//
QB4qnFg6dLJJX3OAgV3iizl4ZVtVpoxsauMIc7pFBR5OrdhcNfRS6zmSvB0+pBLO63dNwvd8u/dG
XJ64qwcClF1c53JV2Wr+r3WXjShRCkpahXBgx1gAWfnkbYnR6evsysEA0uREC44XnDS38Oyw7md3
L8VTfoFhy8NBBGJv/Hv4cRU3KQcPcSPxz9xfO+/2jPAXfr2LAeBu5R5IevNTbk4FqnF5B0Ywa6/n
1gkinb30HLMzWzHFzrpwsJwqOANKhmy92nvUrYGaBc1I0OvPBh3XG0y3YrjgcWZHAttLfqKwyCUO
6ht4oSGoqEZrGbvC4BfeMRQaTDdniWPoyxxQu1wjHE6BWIBCv4WhS7TwtNOK3tWa6x5L0SryRGF4
SuZOHJLWDr9KlhsPf8Pfl64IIGrQGsFVQwawwNszl9lmSftbRB0suzbkl7eAcACqKO5A2Pi3Pecy
ET3N/5MArgK7rB/bhHdDTU+Ru0B829AH7++H724WmCG9X7XUP3nNZJoRwxQWvOQ66VZIDP4G80CO
ujYRcrukLTygcasFs871R9ZXpygTi5J+SKu+UalJT2bYocSkpQhVzKcwbJZQBUvpRHalic2DHfxT
hWWMwR72Eo3yiIMGgUFWEuaJ7VFoZoGDA1S/ldKpWveaU+NVdj7yVDZbAUiL0jslTORflu4FUP01
8jPbT6PPyOPnxIlGBP00+QjVDjYrhrXOjLRyPmoTnK4xW5ZbVUVKGS8XFw2ZqQkogUgZDhA+q+Ts
seX6fqXBWXvTJflZX/23V9XoiQy1qcSYeuODDHixpKDiQeU9gbYd6KLssBGlJ2ROYVBhK2e8jAvn
gksK3QrL+putFpyHV/sr3g4mCNhJvrFsgWpEbrGyLtGvHvhR1SQmDu0/4yZnbxzWkAAN4IaI+aZg
A6FYJ2/5U5+QMS/eQnUH8f2KWi0x8h2JbbTtzWdeAy2jSMwPJxq6YvoirIum1VxmE0k6I6KLMbD/
D2QYVkw6DAWblMesr0lnx7bnLlW7O6YjbqJBGuyIY9dJCwM1Yz/SASJT8dCBxngeQdmGwAToGMoE
okqNqNECJUQM8oFnTwnrZ70Twl4PyMsDd1eWy18BkHuIJIksLckF6ickIlzUJkPquuZlu8IqJgfD
FVWoTKka21bpK5PlYsDR/tuOiAE/9jVz8xROGP9NGD0ZwXWBLx/sc76ElhqJcU/JAQtTa0GLW36l
73W+iNciB7PxH6EVwB7q8PC+toeND3a7XJ/N2+xtA+/BjhlDIQkj0pvzhfDdM8alZC52RSXfaIbD
kzPuND0y1aSOF/ZHYIF5XdF51ovzTgklXoRhj3xGw6lsrfcgRfTJHn665/fAVoo3tST1L/gf3UOp
MHP+AgkVKo18W7tmH2z2R/kpoYpI33a0tcmI3vP2zicn+TPQGbbV6LWdoxndfKUTq2qHNRUv7gmi
skRiSSBxtZntjjAThyhQWJw1d8Az1U/F5V2yAdcNljMYngcSIPdfcvrJzV5JMNEzxOLo1Bpceg8w
5yuJEw+5XWvPkhNW4L4sL373BflikeRc6u8GiueJUkkpvE05MjKls59J+wY/DKbMxdw9kghbY0rY
EHo1jPliK2RJ3dBSQqZ9JblCq8WOxcG+x+s7HZZ4oZvzSU8dehmD3BvjrPEHxeQxWFWu+1rRDwQM
YxmjRgS7E5yDRBcgKWcYJZWIZxJ8rEwyMAuyTQFcXddvI6QR8IXOeGnxXARJpNb4PdYxGSFqxDoQ
2CjEjGG5BVlK1mHAON0f1WcGzUIkSWiLSir3vARwnTjj1dZhe1jrSxxW1S3mhp60Z37mEY+69Bkb
XjByt9hzeIqiFyvEwlAdXaZXx/+dEXMVlgVKzhReBDeEoHKrMa1kMjrzU5OdmUQ6WUnO5lJ77tza
Z1gDRVVAdUgFpghoBSVh6ZZvL+iGbTKZ+q5ioru0u9MpmwUfZIPid39rff1Wir+9vqaK8j8z0e5F
zU1odKVeJSPyXdkxsNvNsvroF9SfyIprD7VrnP0H8AFkoW5hKCHoPlZ9UtqAKIp9GKG9KwNrAY5v
M4PJnCILKxi+a4BF/LGgwkO0nfeN7suLAaPOu1Zna9cwLbj3ZHcGijt4bHXEnytyxy/4I6WmuhMi
bgtkC84izq9D6UIIL63swqEG5Ngt+V+75n10GG+uq/8cRL74oWMEtIuLSH2QMd9eF4CZ9ZTUJmck
+4gvJx93ucXEVMRCDIoxx8U5RurhWzc6UFBDWU1E9Fqa3fOPseIux5Pb7V0mkYhOcqKQV+lCXvxJ
Ar/BeX0ZZjTlKBoUUOTwSwv2aAjJCmmHOSm3aVDE62MP16Lo6uqb3OYlnzvZGStCDsOdyPkPSiYj
FhUIj/M4aJVomHIuW7cdKu9yGZjadAug+uTaSG5NFpP+RawdTFXV43HXudjXDETvUMHUQiCT+8Kc
Rh825v4kic0y209XTk8GPXql5ZIW55oQoRXwDGrvC/HT1u4eYB221b+60TkCOuLifl/r7THXO/AV
Rd6E1kxGJ4NBmasciUYEscywI0tbYeTeGvQhke4KGVFR/Zuwt/BkBF/zHNWkOSVoFP2ljgP9mDbg
4YDEwYj+MvQLx+gpPSJnoUzY6x6UOYsLLdsActrsysL83XzthGigLPcMbMeizq3kOEcigrFO0OOp
77/Y092dLib3Tg/fkxcGBfzlell3bnkW8CFzqh8KGpmovKLYUQ3j3ZDIgdUyIBIgJPWE6iPN0/8w
xEklrxsBu1wbkCAfZimDTYf65sIwZJatqR6qu8rQtPIDBd5Ba8+dqZnJUuZv+ca2cI1EziooyhcI
QczYxWmJyZ9S/LowY9IM+Jvowjbb2H0xslpKL/7z+SCnRSVV6/hxciK1xEcWrTakxi8uZfUsHk3u
vfpPSRGv3rFQieS3QqFQMKLU0Pbhqc8uE4uRIr5bqmFH7zStMbCbtbycW0fYo8pKtGBjQZMZNHKJ
tTDTeh3IYoejr2kqHscxZDwH5YPk/RoD9YLZFS5o2B/cKzlpH+eh0/h3D6uTE3ZmTUIp0D9udRiN
5/BFlUqdQrhIJMJFqpJ7HG6U3hYtgFVnOrhr72dduBGYW9nfJ4LS7ueX6ZWodqapTaAS4ifWrrOe
jjocCDs3cblg9s82FwMmU5RCtLDfYbSWIdru6diaHQgXuZgNyCxy1LmyjtdGbIwVVZKpvXEo4Wps
ovfxRCwbI8MGX0cW48Ofiuadwi8V9c889RslHxx+EIyw75IeBvITWCws240Y8kUNUSwutKXoPPge
Nj0hL8Jg/Wy2CfiyZqN6aWwoHQ/Bg/aSvSoa2XA8ymshfE46kH01Okq13RiiGkE7GZ7/Cdb1zUPk
HigX1dByNuQcKNFN3sBVKy3aQAs0VuhknrDa5Ltoy+fLb3vGt4exDTH5dP3hnTvIz2jOymRaNwws
PJniSsold78IFQdQBKs4WwAO5cxXHCvNQxmYDAl4qKmwIUhf4CL9dEq3JKo2QjO+TFs1q5OGkVas
PtnEk1B1gqwpVZEG6mk6C7NbLOngW7StqQ7lYs3hkiD03tyriHMObmFAoUm2hCqOfLFr3qyyf+Q6
MVj5BFGF8JWgEIllzEHqb7c+OIVnAnKAHTdfXlToMMLzxgtATYgXDktaH6Kn+gReqoEcct3ZGc7W
YtbTkXaTdcCQ6OhnTKuHItWVA4+ONTV94Hmxw2200u2bM4R3sA0duqsOaGnQGOyXwyXDU+kBYuPm
UjZFseY8kGJjza+48DnrN49rrcEb/r1cSulnUXAfv9+v/eY2SwLFIi1i9hjwUhVeVLNGCEz03zjY
dIU2zfFnwjIdrYUZqrUcc7EBAAgYPL+v4LfZNLxwxmS3gTSsPSEwi+yAQiJbWmyw5vXCD28oVKv5
HdxkGIzujpvNd/8eH7E7QG/Tl5uuVrKo68Dvqto8LIdth5g79Gcw2UXjwIXQ0y4lwlwVqPEslrhy
bWGWtLfFoPNPg9rhtYVHBfbDfirv96i7P6GMOWOquIJ39wkQ1amn0vjWFmJh3wWsH2XFw0K68iiv
EDKklSdN8A+9dqOkBuIQlZ3f3BRop/2oF7JIcRXxmcEow66JaqZk/H0QEvDbivWvwg29OvgONaB0
T5n2p3JWeHciYoCW071oLW0rnlHarWrtPxOChzqsviiMUcrD1FZGQBc9/wzCnCoPj6Xve70YQhQ0
l9RFFIAfvPxb8/Gfjz3YZJgOXZXJMofqUHUaK2WmuciFue6sDu7ZwLPz5NM7aTXxNRynvBxolJzp
Ong0YHug+3wJG4ljZ5AyOgzE8U9o35e6EzM/4J3jWfAlVc/HOc8ARvcJJXM/GAlK5iMWyjyWlpFN
brCCZ2wn9c5onADgRyt4OjX/kSQ2OHQBjLLcPZtkF6QezHvff/zYMXCWZwEdX3/eg3NgNgY0Y5eg
HMPHwF+30rmINaay+TFAqXX7/zRGj+Sv4f1lfYzUFy+AlOIxQ376g9S0J8heNHSe4jELlGS3nVua
321tHnKhWBu5o6s1jAlU5DvatpfXediZJmf9Lp2KO9L3Z0zUYaBaJ5rEbfhhq77bXez8SfoWgAtQ
Qw65M4oKT7pMjrZ7QwtDaEBapWjeEtm3eUtq2VLtr1rGwpFldRwLNRH+5fQL3FEN9YUq2lV4Rc1b
galXr0uJ9VZgJw5OyO0Y5LJaIIhuGnBawU2q01Hjy9GoN5L3uvUhUt9k+T7F5qe9M55Ru8Pmd0NJ
zJTAP9XfJ4vtvwTYlF2N30maK67QRenSmw/DOIv8tprbkSeXbjU1BbXAHoc1vp3+u5wKNKP9h8f0
Y7sypjBzdVWX4QP4mCbE8FY2qjzmDcdT6HLa84vK0OpxHMneG5dW4Pi4ajAWWSwTCColSa564Zly
a50dKt9Qtu6Sret2eYL//0xGDEvaCOacT/1ZVwyHM1uzBOhY6Pwrg7Z50tTQ0DjCHD9p2CbyU9r8
kWLwzChD57TSCeWl2nHefin3F9YVWdZlY2/kOYs0jEH0FJ+aXRi+5V7lV45jnBbA9a9dvUHFl0Lo
W3Z/c50gLS8dsBsNGSsWJXPTZJp4aRUyMjY3Z1rF4SQOkuW2bRND5PJPRex16AaTGZ4SSTyO4AW0
uGpV1EXAtqTrQ/YIgPao3Ph6woe2QCrdSzTUTVO8GnkrhjVWL4sRFrGbUFlsv41HfL+aOx5oYLxl
vz/4AsHkw5ZZ4w4KtDGACMW6cfXgz8ZlFZfq8JbcXpIMJS3Lc79BMU8vOfGE+9JmYo9H92ouGPSp
EF9eU49kdnSnR9g8P/e+mKOIpy/qAH+iFQRKai5pbVtlPWclTQ9oY5a8EcDEr9eFM1i0flRf0p3T
BuT5nHEVGMWMoI4NyQ2BK3PU9jS+7JXstyZ0EGMmd4GxQCYIVqA2vmjqHJQ1YNKaOzxwspWU+p5C
72mJ04uTo8o/Sxo266kPNY+rwslou+foM5pzK/fSqxFnst8vJSrAcPQQHZbHySXfOlEuRJgCqH/r
homCbcoPeqae6x/8Xviau3s8hx8lwCdqm3otuuphSSpTMgS200kJshLaWTXfx22wzWBood3BpFhY
SlXuhFjUi5clcr2cfIsCLyhEfHTC+wat9ayImz2gIlFsXqikjCMhgu3nVwWw8XKjm/rfyTPX3yDa
YPi986VoSTK49I2xQ0CsKE9Hon6xd0ZUsnBGoeNzl0m+uK+BGSW9+phmYJVMFxTxdSzd63/C+hdA
kPLyRr3fTeDcIEGmP0wX4cdVd4OfNRphPxF1DRDOk+X6xBNvLduowRMqOtyIqO45o8znWovHQCWh
TDzPu6bu2Y01hS/dQpCGH3VMxe9pLrorr6qxUKX+W7DwbdSbIyOhzxB19zHXnSvrHNF5RUG+/YyJ
RUYK1Kt4RgUN+sGBsn5lDLgp8PGe16mgv6VbAdJZQ23MPAL0WFC6RToIouKumjw3xlp8FjzqeVjg
85iS7OtD07PXtmJSLl3EniIIODci8ggeHkurIiLmn7h8frZeXp62aOEOqy8UJ3fPGdApGZGrLKDt
jVMSXVVxmez1YuBT2vJUhH/I6AXfpoD8TTfb+kZnsNs/muKp6gOLAt/EvHcNvWM1jZ/t4mvUxg6n
YhVEmQNpdFJihk420yjmDkBpEa83v1ddpFDvzKmmWlUB+EaWlrezCCC9by6oH0R5jNitwUDVb0AD
sXwD2SloR5CDnF4F2TyVD971TFPvlpUSvjLeZMzwkxd3itiFjDgODVS71cz4EFdGVGXe3/Z2Hylh
Nmuz5Q31handpO2PBW6WtIeQNpyd1EIp6nSzCvJVjZsvAuXWlmmTZG8c7WLLOOxGhd+8xEQ7xQ5h
o5IeGTU3EfCUoIi26LGSkTA7VokNgZeS+6TSjPr1kF8bVT1sATcirSnXQO9/3XnONtStzFfW8WO7
uftg6Kr6OxE2Ats5xu8NNVosoQE4OCTRy1pq1mbDl8DB52WY/zkJDWdqaxrI0JGWhDg8GdJMpHX/
Yh8zxghRLF/uC2U2ezNkBAb3PGqs/SKn7Y3pkSul2OGkGf2qC3LPLzf2Eji5Cb1a/3RWQuy8+Enq
jWJHTfhmqCBw/11tDZeaQikSRwUVeQslxssR5TUu6if5lqQ/s63Mjhbk1M25Z7vxS8fUKsWUR9/Q
cAzy1vOkHdY4PwFvAclvdokfpHRZUHWV3OpK7gGNw3FQSOmTEao7ZPYvpQFZHYiKE8US/dzkwnUJ
ZXZTi2WdXfTxJqPC1JBvgv/D7CHMZ2s5w4SkhyWzLZ4ad6s6LKiHI0Az5lz05/wPX33/Xs+P2fk0
nv5O4+VrG2/TeedVz2t7g5YC32wQyLnmpTi9ws4RhvTDEPpbyxURhzM2Uq5y2fJtfPolGXJNd76m
TcacFAgPFTiNhypEuBtedA7dH1KCcDPaf95CFba4bSfYv/ioMCmuBfivlyLwtkpmDZpNcohUn5F8
TnzTXG6B/CEfOaTjexVYRnVZtRSddOr5s6ZsyQyhf524kIvE6fyqTRts36r9PLpTE+nxo7o5/mzn
UWcAmT/IcIuZo9ptb+iLPAlYz+TtpTNW/iMgpdkHFNcR5kUU8WUeQx85fY8gFNUp5AUuPo2p2Xgp
HHZzYH+nkOThtw8mh+9HJj7PtCnA5VO5uzTtP2vRbc1YA47z05mfxd9F/KUSNG4ZQkmSXhV2fEv1
fVgiQuS+P/NShMta3/cob5F4am/1Px5UAleo1CZppbSd45wuMOwj+KfRy9uXvcArOqlsptPoLeGI
e0LSHHsXALisPHQnMJJJM655ZwNSP5Sm7igIU3pqjEI/yIPZ0GTK5C0oMCveFd0dH0EJDg4jVUaR
ksJBbZYqzIFi1h/wBNp3C2T6iVZO2rOaTaMs6c+7oANFc9yzWnQmvwT+7zwp1Ujf+J+89u4pwqbC
ZOzQbMCfW1MPpjLTi7GAPRN4p+0GCC07t7NrKnNSs/apF1C4O/VX7kL8EMTXLLBvdQuY6EjXsGWi
SpkUnOSkYCebgzlDQePdqwHcaBCLzOTNz+EEGjTdj5N9VAAFWGqyH/hHwii7gYCBh/Ii/RLhoE1H
26g/Y7EZdqWqRbT93zGVMYFY3xRkkuyVwMQnc/dlIpUydn9BMbCrxXkVlu0R2Os/X8sqoIMKYZ6E
aDsPhxyA84kl+kFgr9Hn6RI4WhUH5qg6axhyWg9/S7SifLQbJuqMjAn3CTx9gTkp3fc68JbmGwiE
mvcSjz+R8C4SO3KN8NgmaB86nlCgEc3WHzclBassFkMOD9cZpjXQAPBzi6LTeduR2Zw2zxiEI6/M
1BIGTvUDYEAuw9WsLjEUbY6nR2RLIhcpL/W5rEpd2dTUifTK1oE3T0MtL4aNurd7c6ivQ+xM1ICb
vyPA0NWMXVt/22UCwCYiYH9ijZb5r30k4gFBGGtySflGJEgCduWuSIGJ0jG2oce/i68ZQByOf0lc
0CfR4Oa1YbOTPIOBQw8/H11/LWMA4+SWZeOvxq168/sN/ZgvSxwQUKakEDXMrSJhK2xzoeZ10yhg
M40gKCcLpFUEZ3mTssJk2dFKp2nqecBvvIwkAUWeuLcDxYZrJCrPyccJNjaAgT8TCwRc2Kmf8ZKj
f5+eDOIUU/1xmUlsHdGz32lhlM4H9pbaTmxQmJwfuw17UXzYs610K6Fn0NaH7tmRtQCPnZHKQB/r
2MRQNofEkSBk2PzOCMvXmQbTlcKU37c06oWvWK/W42syWpeM5MeD/X/WL47W64SUxvsUxuYmFsR3
7lKY8HthENx8OajKBFsWgIqzHUMRaYNuc8dGABpefwr5TO0v9crGsO4pVI3/mFVhjqHnPZn6Nsyo
zuxI3P2TpJR2Eewg+rFWlYEF5d9Hsrjdq1PzniTubDBhI+Wk5OvPSQ1ovgtWcDRdhxNSCkr9BInC
21pn6yA4dZ9gFtD19f99p6lVoCO30UIwCX7oKQ+m5EoD8lGXs6ePXm6Btu9uYYR7o3+8EiFOG3iY
p6bSg4TxXLAtVWcic9Cb+zxZuKimyXus/LDAmMhg/rk+5743+9Fs08xIlIyKbv2B43y2ooRnPykg
ocEJOkHNlRMqDFOg25jsP8A0wWymYT5nJVyDx4dD7Oup3Zh+pXzkoVlVLwiFUrgTuzuJQN2mmvxR
79L0/AmpCX+O334v8oDpnhNHVIvS1EgzNyY69bZuJXI43DTkZMw7FaJcGewX5ZPrykTUb4JvfYr8
cHEcuthlHw2cFFEQZandRd9N23Vi6nmEIlEWi0daqvGk3ET/jZGaSK3YSlZIEQZ7hmhNXjevI0Y8
ZeyEl/guP1yo3wHeTa62rSnsvxlICr820oEVPvcfuNP91cmPVqFQhJ51Oom2xpUQ9izQICOMsYVx
L59QJ3Z7plhTgbM0EJI50OmRjl915cAp/nTqQXznJuX5+9O61vEtcCKmDz0rWTCKFqHBXQ4mUi63
Styw0eg/A2Z1ZU3QnJEefjT7soXjhuWLd3JChGfkPh0P0PTZlL6bz8xtuq6FtNnsb14BZxdDAnLG
QBfXcvyz1gxtdPSuemeEw7WX+Zp4cU+2iBWnmDfcWseZeKXbSPdU/Js3HBNIVv9hOM/TFUMC98Y0
aacRQXtdF18X6k+DhaIqvn494rRzG7wlw3ydZyD2X4G//5YR8XTBhzAaep2GwsEyxWE4PbnY26mf
CBViZ3dBq+TihtIvXMN++y2jN7tjjwHD+xOopVEvSmL1Kz7M0BU2JEwagTP5Qg7tCKUB3PGKurXg
M4XIU9VJYkoNFYD4+1+xsw2BSQDcv6ujsOduCLd9yc+GFd1x8EJMxPOJWNz3LGO9fiQVD2pPo6Q5
R7ASymPL1MRvkdBfHkLjzP5LPPubBfvQ800iD55HjUm2io3dM+gNA7qHKPV3Zau5Ru/UaRQPSAlS
YWsFxEOtB9rrURc2HzLJaqSNysLrOWSqGeu7IgTlJUKqwDpdx17pttjoKq//dJjKBF7T1iUi1XgD
y3Giy+jeeY8Let+KLJjgJ4OX1qNor9E7lJ1ON9EQbsIXUmT1fHRfDUVc0pmzZE8FK1mznPSwdwFa
7uxSo5xXujqzLz7Gl8QsVkpcKLGbKB1i2kIU1QQW1Nf/qTXg5s5jzZR8/PB0hyxsYDT3UF+afl9U
0XgELyIqgD3Uyrid8YwmQYQGmqYAEwbmVwqhX6DW9ul+BrFDqgfF76HUiL7Z0vXwrlTkxawgEWy1
a+yfWOboK0FJE26jqeKdF0fZJfXetQH2waBoRt5npws0pJnRX1UZ65aR9h98A8Nidtlgx9P+t/hB
hQY35saRdFzG5ezLZrgpaSYpkQVDYh3H7/uDrTNXrkNq4evMk0CVw0jZCV/EOqFTm6mSRbj4pPGB
R5SijKmmMJ6AwXXKGvzCFTWA7WRAWupL0EvXWxsJ4C/oTyN+4Nu+kAbru4hSZNdFktQqXvsvhNFg
hxBN62fx3WmBPsD9zbTKtE6uY/RVdnuwPCfifCUa7svr1ld5BPrCx18Do32HMHOPoiX361rPcoGd
jpSqQPOHdMM2yx3XBI/nbsGN6rdAWy+WJfRrNbTQJVQ7N8aIgINv6edswhoEcIGjuyepejclZAJg
JRlOw6p04vWSmX9Np7lNeLeDklq0dsLKpoM7ocI7rhgJgFXOW7nEtfGFFneyY52K9B9SD7erS5vA
RiT7c9BBVkDZ0wgx5sqEpL7MvwiJCeKeacxsUTfdotRcpE8KEc/O/Qa/imPiX2LK7YIO2qmoUeH0
oZa2/jMcPdffTTHPpx1Gb9n0k46AFiOFueFYe6vPmtrvqm8QPrdR9l+zHHFZUTb/G8zCVZzAj/Hq
/kClXC729Mx7W+IoRor3+x6pB7JY4o+I34sSipEcPS1sTwM6uE3jSfABl+wHyouQSKoL9Xk3ZdKX
DK223fFIM0FJNHmDxnAwPfPI/GP96vyn2/k6loUc/Qt5k5q1Sjb6owAfD/WP48GZ9OlVjgZIjmur
5BjsiZgtpazLbUAbqFpsBNvLZVa1TBLZz3U3IXKc1hkxDkp+Sn4GJIWmxM5p2G/9bzMGWqcO/1MG
e9Dog4Wz0VXus00wZUOahWrTWAbcL+0Jy++HIayoHLdPvJvHN0Xz7fVPgK9VJJYRca+2Xl92G2Su
X539nxU0lEqVKkotPXJ8geP6fYzhjwwoQgGtDSCh9MBfQvK1PQFumFe19TRBlvvc8IqdJmigLN5p
d5PCMfN9SgkSIdH42agsllWc3rsExkQkTUOZbYLsqoHeHR7q9O8A292KdhsXne2TJobyV3hYEU3X
0ed+clCjtw1sEph+uIE2hZhq0KYTSQJYUJcRNMIaZDVoY01E1VnjbblYqZg296FApsOVf7Q8vVgG
cNd6JtP5JezcBKVomW9yhClLX1VIsYTc6QkVp3JsCU8YRpHTX3b77SovUJH18QIQxi2KudnIluP8
gUTRkGThOCrq2U2YJEwBb6KWGUMfd3T+iSRuBBBIaeRXNbPC7y/T8eQDwJdB7dZ7u3bFO8m+e8zF
im9avzgOSXDvZ4FLoiLdX+tnxru8hvgbeE9bLa35vMVb/1ayKXlYIwtU/VwDL6/JIjVVownJ9LPR
VqXwPll2J9VV26bAoGEso/HeQmsiajvdMCpjLvwa/s7e6xlYSqjjc6D0DZ0SkgOfVeefn7ls6fZN
L6qF2aMOEu0Azd4B452s6Py/2e5fERKOalvzrGW2TbRUaN8cGl8KPoVsrPNBVMprJDVESCe6afzR
2b6RQhh95jzfb8gaB/UZFdQuFQc57uB2jeZ74FZKKYPBdHNLmanTNM9aE9A605W7bDdjbHmoagei
kbagmuM9e2yMUlNxVWCaOTe1tXqI7rS/BcpefCjImDjlRrO0U8E39Yfj/9tUTjD+2XXSuscY3yjJ
BMgz89aINeaFU6ic2iADBEAhSqzkwfosSafwKs4IX9rqzKLXTTrbin5wIdO2zvZ4VEqOjJYpO9VV
liIlefsfU866y7ZFefqGULrDYsW7Ju6U0eyqKDdNObABQgoP7hQZuooc+AEIlxl34vKI2pWZezQA
xYTOpRDMggeYgOYn6kZ9KFGfuV1vc1QkiNuvw3S5v4Y5nI5nbeMWjoTJ+PRf5hLA1FlgNjqcCrsC
HSqpEXXK1SsgXZJQ1xkZoT4zEmSxUvhT01CxYKmRRY3mecUzHu6IVuvJ0B1pA1M4sKWkjXYaAUFN
kLdNdYF8NwEdV+/ORkxZqRydbpqpdWcc8wAtw/hkmyeTmjn6QuE/1a8Yc4PQTR+jw7F2/j+MAV1h
jtf8lFho4grEd3Ru7TaR3Cxj2YZ77UI6w3J8HNreGfYKkp6IqO5Ume70qH+Z16ZqVnzdAYgWZ4hJ
YyonmKQOX87+erNSeoPyZ8SFBnuakNoA5g3j+xMhRB64aXNdOiFh0rzJFQX/EZ01ek4yYFxQdyIa
tiZxFN7dQpN9yjGZ/7n4UBZjt/WjGdaBdxO8uRk9puqdd9CYet4n0iVEuUGRti7t9M4MVoV9Zxbe
JVeePDgRfxZOR9kfGwnXmVwftl5obV5ZYyJLlzE7/+RN3beIglB0mecMIbbPQtuEFvr9ZSFePfsC
9TaUs2XU9/tk07y/FW+iCNLjRDNctDGp/3aS0M9DgDoJtd707jfgtNFlSq7I1BqgQPEvIC3Oz6j2
lgb8RdvEUveCWe0vJO/Jf7pw9aIbbl5Z8Uj8x6DMzc6OZbVGysfFoOM0/+kf1rz8WjVIy1XS+gal
uqx7hietOebq3k4X1zYtP99OrVg0sJtlBGlSkvJstWGeEoE4hOI3Jc6TSS8wkMV6M3MyUv8yFx5t
LtTGWmRXlDqMiA1C4Z/LkemBfcMNYSIH4xKK5gUT6lqduuSa21623CsQK0RNoAwiX+y/62hWBwxs
4WoTajws+Z76cSC3j9LElQ/VRDht1o4z9QFrxOyIJ24oZ8cC/epP0wXjahNj+ahWPOSitQ5eS11t
KJToOXxDhWMG4iIJ4EQJSBYf4k9aJOOpFneUOcinidmtcbv85ynG7qJAO8Hg0vLS70xHcitp6cZA
87dK7FzNE6Kyj50SgMkSoXpH9KmgJuyjWXlZc7ZKFm+tEu8Lw/fIqPxbfkJs6Z0CGbE+WsP3sIgZ
mLl9oQk/BYyn7o4G3kdeJv1anDq9j4o7ZDF2J/p35fXza/zd8EjjmSzy0eiNkSvg7agWdGHeFtFj
LHv3p6n5Z6/czh9RVz6CfM9ETh3x+yYPXqkBaM+7EoUUczgIaeMCDYTo6Uz3Q9IafV7v+uMyT+Ct
VGD7P3rF9qCmVyPZCxCe7LlsU/B+uqL3d/rI2xzhvIPVTdE17bOZuVquhbOE+O2r91Itq9wkGoVL
h7UZYMFVsT2bC1ECTY1O7Q/lfme/DSy5MZwo0szzAD19UvI5lWYYBi920KA0UVLo2tzRIP3fnKGb
Pm/lkdyLMzZxsvmJWond/ASbk4sHTn0HCj02H6Wirtg5lwuSsihwGKCZu5f9pceCexRbkUepD8Ta
DMmpDH7ZFvLNAARHf1OD+nSVUMHp4GrWPxZh0k7vffXynoPInAqFu0BCuHB29G0ABp+Vg/xl3AAF
QV4a1qzn/mQrjvU9qQdBR0gKugyP6+9kL/y9dbeELZWU4cY1yzLq1Y7DPAyoWZBmiR4RJ6D6nNg6
mYbZxKJhRZqiRM0jaPREneMMzMAul7VDG9EJtWCzccj3D1HRC15MAbRsHSsHQowI33wRt3gLCX+x
p8P4zaGVZ2XSSWp63eHLnh8F6pDYZm88Ri9p2jEbKR+i2Mmi7M5U8vzrVEODgJS8E2fgdoAGnxJ5
1q8/T8x7WL1ilYxubHoVrcvZTUYVI+BGc5czK/OFjTs0njMgfky9gMCeH0h1X3Ce9MM7HuHgjlPt
bYRhqny3nm6fFXR+/8I7ginJPrQgdW4S84s76PAxmeTyAE4WuVDRWxY2iNAZYmkgJsAn9e/8gAJD
nPRbuuX/ew6olejvh+pwayZum5Y7HoN80fAzrEwW99cf2GQhpSqbDIEIIEChi7YO1eJDJ1q7G9jD
PhIqlcSJVc/6VFNlk2ifU2kxCHUYiarpW94jFl00A9X9CeTkwaK2Q7WBNPFU8k8JFhrDuy5rTUPp
l6AKRr4DdWOIhc5hQG4Dp8USm6Q0/rpPxwVDxEJOj442/OHBMyc4r91bw1e4Fh1HVM2O/SOv1vhk
KGTg3GRFUN2258ylYELygaus2YyNuFVdJw6A8usaliZQ8SamIhWqqOWi4urkdkCD9XlvJd2F9w2V
BajY8wKQ1okdJiDqFK9FEP41HpxfNvzY0dI16JG9UE6Cii+27huR5H1Vn8lgMyb0U1uMfOYmWwsF
7nBckgrB3hyh/9yqF3vdUeSPq5pp/0y8lpd0kbk5Ra1YoqyMAVQA/F+SSWPAXocZ/k92troXQAkj
NjYQYXLorH5gyS53C3giNMQRjl0tdtHDpapy0J6Xf7fVQxTosEcD/2uTMjjgFs59k4KHEzhWMM8M
deLDHu/htngVnlIbbejVk1/M2iAMCbZ22hGnbPtFXGaHFVFgYjjuR4F3w5abvr1Zb75gzys24AG4
OcpOgjUXBn66RlStzEIlLOvS80kuAY/EgIdYVcqCSaoiQXUGX8+EFh4T85zLqPTzawNuc/v2gRh2
nmcP4LfjlXrDSgvlDAdegaRoIAo6NEzZwa86P39LS5eADsILvImYCJXcSlsznPzODZkoEF26dfBA
gxjRKPV9LLJ5nnNWxmkqZ31rEy494RDpLZyf4Aq2IpAJLQt+uIahIGg1G89jivA9VpDvk8KJlDyu
IbwXrIuMQxrrjkqNjNOv9nmvkX9hRwjSRYSTwf17k+9N8phJBAlCfECLadRxiSspB5mZrd+CNZho
zo2NvOurDYxMhbdGSTIwsN+4hIBSDuXVQrS61tK7V7UrfvE2v+ydISRuFZyMrfXJxwDPLoT2c5qX
UaGnLqUj0EEiH+CmI5oSh33N8VhoOWxlB1ZYaLa1FbhX6mSyZmco0tDsE1k3Vcz6UVwPd5KRpeDQ
kIl/sOBuhb4+glVxOPH5ZzjUgyN9WBoCA1GODmPItywhES5WZ/1WDIzeJ2Gwa6SsWehu7IRUbzrt
vjE1ikkA5Ai6WM8kdTeG/jpm8jdMGFS9Rm3/mIXxMHBkKEAZi6G3IAceW1K+wV0HBj4MEIxL7iki
YTL7EIQWwuEJM4Ie2Q2M4s10G1DAD3V+tnX9htvipPWmlMP5sARAj6oF5y2xckG75FjqZc67U1fp
TfobM045Am5FE9XiqZCYNkJ3QDR1FqpYcOICvJG5i//dJGlipxyGPkziTsM1Qtz/rOaoBUDAp5fo
/WGk9mz4gY4w5R2yoioGdrxY2In5qHbkqwqtQlse4OWGjwu94fqHFWDzq8dWFm1NgAp2+EJvRm1M
Ro3efbcBFaajoKYqbXTBIvr8NS25Waru5fjKOg7jIypxHy1rKgQTaSIWqvZcJG2+da0L0v018w7M
43EM7HVESlkJ4yxy3VVRe4USNjP52di2At6rVf/tpEvohMkgrXLvAw1xdDW3snGTJBVmRFfuvSPI
A+8otAljoX7ZX3NcOvHAOtq0YiGKE8WEF1ncsGANV2QE8m/GmkdLWdTP8Nc9tY6KMMFuEwolpFXd
YWPGDBnJlooitK1/dIKnIxPNL8LkgkTW3/daqdM8seNh59pBCW1s5PMBWXt2guzsYjErwKLOneFl
AuTdCnszRWguklH5Gkec8IGQN0PJmku6efxg6HpRZEst6BjNxOnKSQoVa2gzWDNqZjXJbC3p/Fuo
2dQspmHnQHFmmHtphXGlogHF2Z9iFI5j1UQNK9Swm/AuJ44OUX49GBrfBeiSrpDoh3er2Wzo1G+p
Bq8LNtCTex9RJf3h6aQ7MNtrgUPOyP7ilpkHbpnSIIrBIuzKTbHwS4XKPMuY7RPdO3b5V55MOae3
FSBkuw1YxtTB4/7XlBlTjwWz/Hn1au/sOZnUOJ/b+UFpevohR626ZATPh9OMrXBXbns1qEP5OtkI
YpRNYe+ghj/awHhCsEjYp6NC1p6Wjjh+nvPns+8dtQSfh6mfXpfv5pYECVgm7eox05e5LGW5MKCG
KPQTvcMSVBQQuEQdu7yQ416nUfK4IecXKSRDVH30JKZKJUzuVLjeZDu9Z1UwGzs631iFfVUwm7Y5
hyZ1QUjSsUPNA4AIO4nnPnps8PnyIBgMPPjDW+yoYWkyoUiZXeRCGDqOBUT6sMQRQl9dPpH9Zl3C
Trmgi64kvodb2KcQycF+fkHZ3A5tyZQu/i7RzfBPC0Kk337oCxCyb1Bx03KfOJ172AlAXXFXwtL+
sgRqGWgR2fGlvyLEEga6R88XK3JMSAMhz0zSTmezhehXfiZwKXiJ5af+SFi/HN2NwMNhyT1JQa7G
f3qk7lpkqT5aMdv2JjYsX3wsxTRI7ZCQma9kpfTq2RBeQ5YDdvvqVlXqGgRgNNNr/qKeU0iX0InO
jVfOn9vMlrQXP9azPJf/2zmWAB1VWj7699kfJLnPFH5lkNIBuUW1NfF7xqYQqn2j4jDF4M/cmhpK
Yb3y/CxEIqUb0uPQRdhIyQadRJJpklt0iyYgOGzElGDdGTcCxh412Ra9V2kd4A96qDCz8XdPisdg
Mv4FuT5Z5MQz+FZqpq3gJgqg1pSHj0H203mF4LCoa9U1kDyXj7JNVWIRlKAFoUFkB2SbpoBnkrJm
UT/spIerrNCuEXytLUrje6X/qn/x1zRJcrRdzCQO7KKgW6g2yaiTx4QjYXwcT+hmwK3mxPy1XS9a
BoUrJzzr3dBSZmDrXgH+WSMKFO40sClHimafndT713OqcozPt1dbk6qQgjyAlYhSMEpftKcvKrUD
XngqLNbj90wO0kkDerei1QKDa9EpFqLUqDG1/QIAbQ6fcpV3xHp910nedJNxmSMAaGBmq5GHti6O
Hrpp3uq1FsUdp4YXMgJZSm73cbrVHe3cqwtkzHlSAToxwfwT75kEPa06joTqFI4IYlOBlPeCITnd
/HRS4WLfUe/wR4ksFHF66cYmHztB568GNB+Il/ku0511eb22YyJhI4xmRBPRRDZs6BlUPoCTEIb9
jmIM4b+46U+xtKeGc78RRUnCcaU6lBPxKlttwoBIpOGy80gvEZQ3TKnVsBlAHTNlHoFUO3ilfJPO
XRY0eCcmcHM+2ivaVkoBGOYjjYJiP/kwZtnW/E8wU1Vg5Mz9fSTcy2w5xo9uCglS0vNvoZMqBdjv
c5QlbYh5NJsRA1zvFj1nuXhR+MuPWCGE9nP02syl0QoZiNXZVrYRhzm2nWElS7UNqBTmiAGwznQf
6GtK3GcB39GEyyfDqXutdDBNPMrtxdhsqHPvaRIsFYFITVEZWxuRciPcahq7lMLq7ppTePIvvME2
mrBy7PrIaEK3+pvsmRbNEzge7YFERKUZAntOiP/iuXvSC/pT3feSghYCnl/4hHt9knXZICGteSGz
+SysBCs6lEl4yn9FALiNVeD9e4WvgqwA+NTB7OL9vVDCO7xdVy7Yhe7NNNEcil7rs6TDRKbv2o4c
NPAtWFJXB9dk94eySVuXOrMqyGw7tw8jKuOkFHLH0rTqlGiMzmgUbiNxlL9mcP4IRrhg9ATA2L3o
SJlFHEVz30jurmRkTToEWvkoM0p2djoNKz750OtLREAeSciYFkgGB3lRTyyErzhcCByB4sqfdnK/
Z7FOe0bDZOvSdzLskXLp9wg5jEKISL23zwbqtY+10Xdaeoezsij0rhDFEWx3y4DIIdqA+cY6NIMc
8MmVdCQk1vA4CXYPZ7Az+/Knib/3B4LWK9hvOKRehVNanl1uUAIsSft3zYEqSCeWmiZW0JMOca5h
qV4JNSeIiL4hmey3in7H+mUjiTViPG1X/g/SCexqAQPQhXTu3VISXQjqDj/m578xA8OvSOKokH0H
u+RYRuQ7w7jbkwD2KAjqvOk9aCgj78gpjC8CNJCE0ZK7LXOsLYAZzfEiN0hhZysUG3r0tZ+yot1O
sh8XnssrhBtm5wZ5jkLBlGL/El6h8Ww6SCsgZwIIdyIGSly0Q0B4V6VLmBOdn/5yNK4MrNSD0nQZ
NQgGfgpSGxWTazNfEIHHDYGoNhQ1dQCYMoDRTmN/SrXnjwtJN53xmCWuSdNBrjDkql5QOwVjn25A
a+af0CWy2iy9+gXW3Pe2RdQHwQ6ZC1bGRfT4Oac1Cbj2E9MvmyXQkiHBNFrPKY5JTnPMGOZmxDs0
HCwxEK+KC1o7xmGwhneGWMnSFx7D5XS3T6rw90TOA5QlwuE1iP7RogVs2khmq/b+SuY7y1FCDV17
W5Eb3Yf211D/tMFmLWc59CfpZr3+NmeteBWIWswMaQuaitwQaWI7+PCUUO0D4OyPNowGBTo0QRpO
Pq/aTh+Ff40GzjzkdeKa6HXBi4TT9mZXK1jKqFo2EGwjBlwv/9vC4xjIGF+racS57SVditwaxxxn
L1QwU+VKFcLhlDzo8sCLembv+tkexweMcUqadpmZNtuAaY9warei2go3KRrowU4lzXXEdByTLlb0
nh3kl5dp2W643/5uDh7G0Sa2l7BQQBlrOGEtICHtNLZ8FkXvtdzAg1aZBofcVZz59vN05jgrAWMF
iddKK5ZyR/jvVcPXa2iTEfI6po5jR6DvSK8oRKcRwo/dkLG8I6k53XB/KuUx1IbfEuqVm74+1o3n
P5tslh9XgpgFda6dq5Y2h0g8u08EqlaF5vWcrODNnn8/F/IvmYSBfBamTOv+t/AcryAeMd9wvJsS
OtJmektqEJ9ImRqlvZL6ovCdeQiEZ9hZaemP1YvZzWWiScJrs1ovi67/+dQsV3F87vWYXW4JOwSe
t/psv+vSiPSb7Mkrqjw8ZGW0Cx6T6i/EvfQB0/Ks2z1ZbgvAiFPYlPt97C+jGaL7CjmIJz71jcWW
RdbnN/uubY6OvYnln6aM9CbpzNVS7pdipczyHyseTj5Dn7JF3TXFIevuWPIR/K3OJTdhbtM4TZ92
lRsyDJu6Q1in6UmI1FCJZwHjyHzVVKf+AuEm6WS8W+zXyjd/q72Yiabr15p6xKazM+funn8XtwGI
MA30mTSE/AuWqlyXkKpyV9ID2XCicqOEhB8hCwBsKsPBbQm7e8VK6Wt1y88M8zrVwaYpeca4d7oo
eo4tRFXkYN3wxob8ejwcPuTU50EnoA+oohbT2q6ZSTTkqHSZ5QXsNNHfVrUoOYq6Ac7hg63Iw7l5
DQPa9toUDE+8/uB+BA1Tnhs4MO7/yTOv47S3I+3KIDGZyK7h0NnX5p+rC0pWXB/zFG2p9a6rcvYZ
3V0j8X2cx05Sq0pSQHHADOlbC/pZY2U2EGBcCpgU249Plfp/mzqXWedrNFYusD0nsrDn3GXRKpD8
PYTUoYFCRwKh2haYsxtus3tPrLSlEBCBpNWu5/tLBE1sdtLxpBWHc8v/EzBxnem+FK4UE1ERhfeG
ESADFZFPpqClP6ncQjLD2U7xKGONmbRzUXX4cl9UjG3ZBmTJRTvOpc2AA5BQhbXyUk16jtSLiC4h
hvmMOG03WaYpymeUMSg+MaSjIYQdObuusIJiqNWjYu83bnrUldLK4/0ES0G1rKZPl6lWELouRfri
oEEOR8zZxKCdS9k5wHRy/FrVHYLUQ+MIxjeFmd+AT1drkkXIV6ZEeXcCP0f9HWJLv7r9EeJYpTBz
Ea4FX9WH2F49Z2Bj4+/y2dLc7wOWYM8XpGz9oxS47FMeVdD19ZK+uw+xhPCQBWrMhjjRyz5Lt+SK
z7Zgw5dqyA28vuQKj7Erma1ojohtG9eB29fOpjs3ngaFAkybxResmYKXtW13Zi0mXVq41zknxjYh
wtUvT0h3HaCVyRA3piqKs7+ooWyp3yKTMVn65sGU7oyXmtEVgZPenyxTc4QLLWyzLXUyuyiUXCcc
P8sl75J+Kat6TOo1xqsJYbApZOzjPbyGnUT1gGQGsTYgP4gcJKwaRdft/6mgKvS2HeSirtujNKDd
zQEPSiFPzWf6/SVkwfpkeea0aHhg3YUIO4onjTRIhnH1w9EAIPBVf3d9Jk0PKkDndjgWvRjk/g9j
Ca42NHDmtriAg/IK+2AW8/MotlecEvoy46/VbaHcACQ7Ui96/WFLSjsL/lrqq00mV7q0vOyEBadk
7SIEgylDtnGeTalhnBEJQba+V9tGdi2Gh8UGXMiP+OT+AJYVQs319a055nVVoPLstaGdhDTh3/ry
vJYNMbDSaE+oFLwRDjpi2N6hhbRCcUagiLNmERHBEJCf/WaRipFRBaT3uJGAQum5HUEfYgFh2Y3n
qXgJP6ug222WqqTV8XfPvrlqaxf1VzVc3KpFuXjQTjHBov5oN9o5o1err9QVfYcounlaUyIV7Eyg
UD8wUPPYqryMc7m9cMIJwAHvhk9Z5UM9T2zLYg+0B1xB0LKYmHj/c55wlz3ICBt73utL2yQgqbnp
uA7ndfqto2kYYxEXYIYs5S5UNXaBJ1h8vZeaO9vytyrfUoeygi5eHpGc1JKxlEifyDqO4phHSDv4
jESPW4h2xSQNUtL2DZOIDlGPXOAtymorEMNhJa5WCTP+qbjW4uE7oDI14iQ8krGKcZSyABOjwJmM
YfOfYFPHaobWw+HsRkBDeK60bT1axMETvH2CUrW0xQSIZpuzNYuFMb7vWs9zgmQWwRfAZkZC1dnY
OQI+vCd903YIhyk95O7j66SZPdrna2Rwx07PmmKayi1K2jN+zCIXyEAOVUhaA656vZBL9t7jTTeD
uUMlWu7UoZsn8QIIPaxd73Bq4fkI+24T3HLlnyFUwEiNhWPEJW6EdBA3mXy9CQgSsTiRXcJyt7tL
w+saOZ0EX7p5XjZglVB+WksFVScoat5WfoqA8XsOFF63eeCdXPUcWi0BEZ8MkTOe/hIJ0B3Hs5ap
g5xBXrGDqio0hKHxonWZxeqJTwHPiNz1EabfOfe1u6rPBjeE7FPW5ncot/ck+P1d2qh/xFLaOjad
LVXYS+8uPQp9M4TRtahrqRMJBMCz0NPDI0x3PVNW4YFY5/SDuUOQQ/0EYakxtvIII4kmJjLzQS1J
RKBSI9YQwLv+8kP2Oo/inQa9Z2SwMp365Uh1ALJd0tOFg8MX1Q9DBKV64TdRJ7EKzohtGwjCKII7
fZDggcBbixF0818VmVbCLKz1nFXlEra5d0w3YJttr06XuBH+Tak7JmGBfQxCvRLId/8eK/Yw29Gu
dz/NgaS7rLDeBGQ1aWDcW9UCWFBiyZwzhw84zGEB9mtu9EtqTEJIjUBCWZ7oY2C6sb/yE5Xqu6oS
YhfzKBqgJthKQqNAXvkHrJav8QP4lzHGq6cTfh/0L0DbebmVdk1R18mUjRScH2H8YcLVVDeB50V8
Hgjf6tM0vV0mFSiL905ZZVYJu+F9ywbqMlEtwKNcA1lVujYsifJCnf0PtWF9feA0XTOpDjuUJh97
ppWT/gaHZx3qgnyqlhom3m+DgOEu7vYuvo1kV4BoycUjQLw7gHuCvCFKKCw3VhPPrHBEQ88UkTjT
nnngrAzDAaX33ebW+UQJyopbav3zW7DIBYueEzPgd0o/cso5aIiQBThzhsfQtBbleki2e5hsnxTP
SV4GLrB0uqKHQE7JuigEIFNGQ3+tTM4IMIzrLd7988Cyrv6M9YHlDLromIMSKnDGbkE67urePInS
XZOW72lIqOliIMHDUTvglqaS5FLKjtzAkE+wR+tHGLi3g7pY0nGTjYpk61xf8mAeEbpXCexE2dIK
d0FhfbIpixMmEQHU34E4a6S5O1gMKnEcCj7L7LFmLo4rkfNe5PR56Tdz9peGMXvczqYw5n3Zdkm6
p7BMOZMiPoqBUxz2xZ4FFxZp2QJWbkPYOuYH6s+HlilK3F96iAE8mX5vLG/jhmoVAvjhP9T8trHO
H1M2nWGljFPrUf2ZKoH7g86ZR6NapfPmej9DADZXk/a/AhQuGDeseRGmMSHLBwNHIXrwtIA4XeNb
15UJKTU4JuErn3vHYC3hjXssVcp0lI4k8f6tqxiCehoOGMVLe+ZrYKpQ0T0eHvN3VGZ3LvLH9+T9
LRWpyNHAwfp24yfZp1Yfp8qx4KsgqoCJ2IMkTJBjLR5XZIeArAJ9R69pi0c8M0iLhDymYMI36ucg
kJ2ft6MeUaM673ht7H4Ydrb6eQJG9ni6ilKnAEBf+1+Z4Jf+QfgSQ69nkgMscew9B+MYYb2MO2S7
4+3+OCBaPx09CzC8q0H9BYwDB/T7GyiCBSerYf/d13dL9J+vTjBRvx+re4NN+IdNfAYWV81qO7fd
DjxLyqrVdcTG3f0akUl5Jk7a8On3qNBAPj0V4TvxqUxR6GBsBOby9vvFOFu2y9KPhKfbHpVQSAeb
tA+GIfjttDDs5fBO7enD8EpS5QSxbasZkKEbsWB0a/viiwyqcTxX+LCPqjJvBd0wZ+NT9qMH9Ug1
OaAZUwsUkrWz/t6UJHGkLvkS+N3NOs7xf6IoqqkgOK5C3n4+N8bOuza1wL/VYfupB7v5/LYipp8O
oCdU1GykWEcSFQfB/AFxVTOxprG2Pk9akcL39FIkUyB4GZbEyHTNpYRO1GEg2I0JydT1naHWWU3D
sDEHaoVmD7ykSryNXaS/7/zVonLyKsZKWLCbSKlspAiG3P2JGXnGQmWv0ixKi2OxG84QYh6griH5
XDNRwL8yTTLHjHynrM+q0PsxLixXAbeJQdQS3UJQN5tGVvGRJ0cnY2LAHLXvWumSe1ZMxyULNpGy
PIAH42b/4+yXFMXba79zsXMWWXUhhhsKzK5vKau/+a4rZeRxsbtLW/8wIWikfZteQgKA1LnThSra
LqsQT3adabB6UOeqd7rXl0W8rTuP2AmuxEtSMNQ5IU2bYMLn2ReRaB+eeFeP2vmrDfQGdpMHbWu4
vPkEkW6gf1jSXqVJQ1OTCYzNIih3+3IevMhljHn7H2Jv+AGEMUQ8WiDTRmtQ4e6/WwhCa7zKRyqt
ZvWnwA32iQ/MhQ6MJ0v631rcgR5YU5ZcushN5/lhEVY4q9PZaVE7wBd7nK3QMMnFzJiXwQAzB8cn
IefLK0VhYW1I/KuTgDYSGo70jMa+fbJ9Tcv488m5avQcAN+0fcVV7Hrfd8z0k9yK7m2aZF4vSzQa
MMX3+rt5HB3qFgp/ol2YP820z2WV4yUlgGwWZMb3qZeaPHgS1hZ0qxG0syt8BTa2swpfRNpyJjY1
Q3VTMrR2wbfKJa2PcGFlazIrTnggIrmhkhyniewGXL3N2IU3Sli4lq5VeTjOTBDThRiwdr8Xewvm
x5lNO0e8lnjSxleF12iXKZP8Q6B+O23EC7oUQEBgShFl6q+gWKGVM5BQ4bzUF71vtNZyFx2hn/IX
MDBLsD4RtfxBwqxLQXJm0fy7TBPTMVoRRsxrPQ94is3iQ7YxkqdYwuge2pT10csIqdlJmRBeBPxW
7brlxbHUyl7RPW28EHkpMgfeWpbaTYEACu+jkRBAAYqVW+I2w4Mc40KvDD5FFxKm8nZFgr3gQwx9
2M5OGR91ZdEI18EKxvE4YAGuRvXnYTECnkUxz2dnrMM0JNy/zstlUqiHAaqfEKyYwO/hKxMmNou9
/oTKHZWu92W+nkvZydQpx+3k3k1dAuK5059aD6hws+uiMoxYZTH7ATIrlJSNXzKCmFlN18nr9nNa
Sjy5fElJpM71zXNNkD85MOy+UOCqFQkJK5DJK+MWochqACfRyj4/zNzHJe8dJgDWHFrsfO2ncesZ
AhFBGmldXE1o6iOIptYliuYpUyqrudjnQAwExpFwJ6yQ7nss6A4TD0+qyakRP1OReSHUI9GCi99K
T8PaetHTxug25OYWUu1XNoUUorw72FIuIpD13jcGVaLzn+qTHInbIpxmEyqlOUwF8ZUbohrCs5KT
//YrneOJZSh9WiiSltFrF2iLeiCSNV1DLI6uqzXklNqHrKjWGXMYKf7JlxZdctDvYNodM2sNVQiN
V2fVi8kxozCWMadnH9FXenN5YYoenHNZonCqArKTQaKLxKDW09b2jcERe4i1kP3umMif8gOnvIE9
UtNU4IksPdVCsAPLC9avefJYtgd4LRoYptT9mont3Dt5qybsfgoJvpwqJVC428wMfO8wdwzkHbja
ksBY9eNvRZyW4TSQ/rzeNvzd8zRsZKNG23DMckEYo5XKjQqZGQnNvx9SG/HBPn1sRgcXS2w2/2x6
FNbRBhd9PGhsMyY1fGkPOP5q+SXdEyaLIwhedT/Lpo4kWo/XOOBLmCIyL6Fhwc7c64GDiE8JmZ3h
ywf3inR9+hEHNf63CiHUDI06x1ecbrDSXzpGcsebNCjcGMyG7uPI6pE+nI2smo6O94meK6lXRVKe
VknDIGATvEfs6WkQsBxJoEmPxuSdzAiw6h/nzyjAcbyQcMKKo4u9wR5eyI/YeytFMg1gsBuMudgJ
BYRPydaAREFUrjTWkxLXJR81EqjeQbrMN9ING09VD+sVI41VzFPpu4d0xNtCroXn5i1tCONmMdWC
LyeoCvkVukeM5W1pA6Mc0mrEuXBp8P36P5uMUPdy/6OrMoYPO9/k3c6SjSVp6JSoT9iLZiHXAbqz
GOO/YqN8+hdLa38Cbu/AC8CE4c0mYmrRvRHEu196sVSJ/p1qOVIOEdghABi14QqfVPYgVgcoS3yV
ZmY4uCbVannTFj7XOeXEdiOjPSI1NgFa61MHHq5jpbu5Mq1J6h/tvdgD1T7/JgxhhojV0Q1wXk0S
kC5rtc8iaPiCdlqPY7wy6WANC7jgLdinY6vBxUHlJwA+OpX+w0zXT3we4d1niOTJx6Zu0MXSMt2Z
rAQWETyz74adUQGBHpPLLryH9uGRbOk7C8opjAkFeJdVtfdPZYLyi+7S6JMhBUBTO+2UoiW9COe/
HQ+uTG497BTlyKAPQg50cYtqdvm3wtLIX/JbJtvpnipZFNxzsti39eYS24c5oYv4wukNgJ0WLMMN
fDtR3gIy6O2FWWhPpRAo3BSwATM2/XErDwoT3AQ57N6AQOmtAL6v1LSpV4R5gyIlwHRuros9Lvi0
diyBXNM1fGWlyUn6bxEmTNNfEfhPAUT/8BN18t+6PL31vTmF2XGfQ5C5R5SdZ+1PmHsj4K1WDT5w
Ccf/elq2nE4ishZp11B3HzVFEFTMBY6szJ6hsFrOFEDhUMiG2Pxcg2yop2C4tk/D3iEWjM7S85DR
vEqA6J/sAaZCKyVEi/ePxCAVjo8RanEpFntBYX/cwF6bOZSgnBqJ+tekK2tf2LoAfCWzYEggzBOZ
7L3bSe1Br9Gp6NpweVdT10Asfxrp7EGSCMX0sSBWY7o+ySxg3YyhfjuVfQxjuuY1tGJVwgwfc4lS
WAN2qnhUSsg7p+NZlhGPl0Kfw9x3WGYZ19bDS+j9NBdxlgzLccBdFej6grUoYnlEseanWQan1Zs7
5w78pA1TGcp/nxq/CU5iXkAiSpGu92850dqeu7LzeXSL5jCtYsBHpjgq8U7zEzfkGoe6jXjrl/Mt
TxJJ1OzmCIX4mStiBq2Oe9dy0XtBNcntEQpCO6RD8Yt4NfldnwuBmXa59lrvufioK6bhCk1VG9kC
Q2NBF7s/+mng1Jl1eztq/qKdFR8V8WU/i/N+Q1zSygvhhSEvgGw6bO1QdsMJ7paoNKpzA+tY437E
DPml6fKb3CGm3p2jrKnwAUZ9//G25PoVNLX7UALdpFcQJ/JXQGtlZaxDLBvr10XB2upOYlPqK3ui
lEbuTiWMKdPj/B7/DkxkyBRWQFJ+aJrnHJ6p3sOlGtC4CvxLNJjmZwxbVUL3npy+qgxqAB2hhbUT
XHWgNprVSRfHb0DWqKkitKrqvnTLjfKzHC3GtDj/fHz/tKygzwzGO4Xlz1D2iry6n+EZ/T77sLT/
CNdJzG/ecC7TsoKa3q5PyXKIsZrUlh5nemNqcHOQoovM54JXrJz5q4dcpBoDuN3SZ3Z7h5feLKnP
1pnGSysl6r79q0cKzz7XkD8CtSG75TeX7duYLKxT92xUy1shlIVRd+tVtXLx72vNtqUHozCGY1Dl
59EtMGQhtQDmwX6d3R27X4PH86VK6t8U+FFwpAazEMVqtLtHEJfEeNnkRWQEoQX+AcB5QDoDjzk8
mcTkWd/BCNkrcqENI5FiCZFdOQgUmEBkxQRs10jyBzFxeLYOC4GV7FBNY3o+HlKrDj2iKeQfw1Hd
MgfV5lMncTJMSOLeVjPNcML308RGVzm4a2F5DonCDFf1YCipdFekI7EOTR11/HFkCfXAedAnUHnL
ZeYs0iF9Xd4QL7pwOfyLyomnYJXHeYQMyZbl+/ZXeCdc02w6HD85KxexsejZ0iMxsNgISleQi+If
BI7Ny+xyOmnrZDfUvwZhcAJbBKOTpcAB0anJJQk9njtg5a5JuaZ0OY264XhL4ttIM0ndeJw3EeRj
nqvEYKdPPcuZtuFytbA0vJNg7oqLuSoR/2TLyHAkpkhlnPSd+eA+flw/SpWbLDerVQNQM5CCqUq2
iLslq8v79Aa837jzOBg3y1WVsFeKtRSjQ9sn7dE+2BVHo4hn33AjCdEHO2wWJamZR667vECQlxk+
xXGqLp/ZONbex7t/5sN3h+ufSMsN1lpqSZiGEjLEYE0BI+yKfPapiBxEiehnk3OCBbTohT7VGtNx
xpShD/S6JIUZBr4xJoUyc3og4u4lOhuZXBlD8LcjQMxM1FttZ79jG7NzTsiWRrIwWTMtR1COn3Ec
DHeENy+ZBi5J6JkO+iy2vciZijly4J6kW2W5FsWzPbvWVIVwe87zlyhuhKxuQMu9HQs0mzguzBlN
TBEz87ByBWtB8m1K6fMYSt0MQpSdReqTY6rramvyFjuULf/LcxkBy4gaE8cfsFugzWESMDHd67aF
q8JQcuRqAsCzKqbZbYpcwrT5vzvMcDvSbVA/U/oPLBCRSpBoWIV7erXMzHNdQ66nxPQKPTkEld3j
nOpp3n7ZbRfQNHBmbEswBeW7hSxnrWO5wmXs3LdeavS7daw/c3llVI64MQbK1H24wzDSwP0ldO8J
NNSIyxscBrUVpzGy0i5DXSToUk9HGJcO61x0kUfmphY5JDQJH5zZqCKmGh/00GFRu+++seZL2ivU
B+Vv0T7ZmxAr8vGEU6BnLLO/p3TZGUPPLoLi9xrE+geyCEhusBiZ1HA5/LXH94/yQ71m+9E3NG6C
d6koJEgk1zq71FSjAfK3h1Sa+mfyCnPaOVAx2eEFoe1hqjYM2OVhGqaRmKWDx5D87os8dWQ8sbXO
l0pjcLYzy9oGaCGMvF8wxd66jpNNym1f5gpqo5kqwxGoevpWSj/qsQ/zrgxFl0pHl2B3aNoa/FKY
YKf588w/NOkvsya8evWjNp9nxNhVDw7D7s2FIfvKYIZbRU8CTbWGYxsT8/6rtTwnjEvjy/DsfyCH
eDimcX7hysckjMlByIZFbJRVVVA+vKx00fB6hkip/U3PHnXxc4LQD0F90/ivPbi0zx9I+IeEhajE
y0l9cBE7oUuRG/a0vVSOlgQ+jNCkkTU234st5n3Zucetzzn9VrDZPg5Sk7d6T4lMGt14NNLoSb4r
45U5CpGstEJ28Em3RumAuldT/9b/SthXM2rlkTkzSdkE4IYYfxPU4ehRgr2sOcnh1mxVWthlOnny
p5nd1TicOFkXWDQK5U7/pIGUIek5pifYwEIqXvCpUXsqtwciyvB+XRS/rM/T/W92cPlb0Ji/mQ5D
kEpIQZLjz3KOrDWuZXst6TLS6xJY/rX95fe2l4GaI/eR1776GoC/bMbZtC6yQDe+4vNEaTV8tojS
FuJO3VsXaXpK5NIOda5jAM8RjbO4oE9BqrwxtbJmPPSjz9SuPUvEOJsj9UFzy0Nj0WXfpmj3e9qh
FTi0ZWlGItZJif4Qf3a4u/6+fPqJ0F3I1edLW79gaJzFRz9SU6kOG0UA2nLn1AcnTjwZI4ns4tDK
p1Hwa1GvG44+wCa5NTtNSPMtiWIuYAbfaLeuVbAIdefqwDaCg0kB8ozZbQIABy6WV8k7c9/kaeF0
0bK1TRMPrrmtcOSpPSfNiKR+5YX5vQXYUx6lc6w8ZwVlKbPKiiGKE3l27xYdpvQ446yaPjMQHhaC
tTmUwUtGt2FEY8Sb/doCJLo4e7A6CjfwsvBc/QwQ6weF0EFTjIJ5hEVI8C1PUG2ut87m+oh9qJv2
RYuDWAEfc0yt6TH9bqxWVMeSYZtu9yPxC7PJK1+Kks80O/qD1FPcUn9Y9K0xP9efI4OIkueeRcWz
vseQgFBWNT5AZZBnSkJX8KuY6FEfYqXfAlsFbc/nqRfdZZfiBAlFOXgoGAKrLusIzm0Gwav1a8OH
e0UEsmZNwmrCc3vQ0hOHyAS7peylLMeOiB1SEkisS7ZoyJlOeZCO2h52TCqjKUr+6C/fihjOjTFR
yr/VWg1fqQ7wXRVKaLvoHp4KY914dpdrl8bZbX2yj802RgPxN8HupJLqe3570GRzyrWr5aaMa0mS
5SPtC2HXM8JZ+8aPiFXyLApe4l6NWo5AW0za2sM3w522rmUIXgTVOanQAkNy01jbP0lfbHRdbnYL
hBwcR/MbxqDE2EpPHyL+18NOInuuUae9je4oupgid/zQszElThXz6KLdODEeRkSYi0ygfwsxBDxl
aLCt8c+8cywuP+KhxhPBvrgYROWecWJc7SIGTbRTBKmu5IUf91qy76B421yuzvaBbuymb9feJpkv
dQPMCK+O8nTUPgKM80Zz7+uhAx5hYZkuQ9ymvi6C2xW4iSUswdAxQUn+eBV5/D0PVwgLT9Boykdo
aZIPYiCzROlNmvNa8aOduVC4DeAmp7l76YAu6uX3AQZU889WcLcCuvhceKDXD1pgmM2lnmacoXch
D70tSX9oMoVjpzkD6r8u/bJqEj3lwCOmGis14yqD3vzXFwvdNmcWweYRbabhlgVxy4TDhE+VRSVr
shwmsUm5hFq7C8XwLa7VhnGakl1xkiDmZxP65YjKv8To5ZpV4NZ0jEk5WCkbE7FA60jU7DlYaILD
tgaaRmwuqaTP2wTn/WyMAAeo+9Yz52utQfMIk3RIs7mw7JLCwbWuHDkbfHK/AhVH2p8cWAqSthNO
3VbBlcP3+pFyjAwp6QMLdXHUK8F0IgwskdDA/MBy2DrhFZghSk4GXybgv7iOBwrzuG8Z+xysotfd
7anS9S/giaJH2MrTLEIID6dMD+Nv12A/EU3j9RcxseZFc1UgvIf5s79qK3k2MHns2TNPEalkxSiS
ExfkmWiiH2l0clwe2qSvt+J6r6G1/WBxmrA9+HAU2AVmLPXuZXbl2B+D0q9vuS9WEON+9tIbYWaK
dDdw2hX8HcB9b2j2puDXdFpvRVP+eRNFZe2Q7xT8AkD5C5BLBaaVTcSHsoXmkZN+8/6NnvBU3FMS
70rP3WSD0CXFGAw7Y1jKZdy7MeVDWDmecGScrQVF1+pj5fndY45DHPo4zu2QdDIovr+5zkkzV3Ec
jEjpcT9NO/snKSeoWi07qgEQYYDgUcZ1rGJ5U/1EHwr1kTVhwvr6bTrS5XeTTO8vvyWfsAKf1+yx
rHWordXtYuEKBcBopmdOiqkw53kvP1m9k/PVsDAGjORvM4P9I5Wf8mdXNAnC+V75y+rgcPfmL/8u
IEv+4zntov4VrgEqT12rYFwF5N07xj+krKDdkgMhNR1P92j84DwRNInbd9kHsCMlhnkM1BHDgdSn
0UsUOLzkprbtikaQ7jaa9DhvhCM2HMcO4ZvPt36gMOEo7DdaSWZv6jHsDEd236RaGxpiDM2SvtNM
s9YB/FTLleuVSCKmnLRuREKiOBCGmvyb21MbFakkqo8JW1Yw9LKjiVPcHwpk5Ab5B5+FPhfJO/wF
BPkZLDjmuOa1y0oH79KFpFw/vBNY1qVPUtMytan7UJlScLxutWFvssApiFN42BIa5Sw5Gm9oBGw/
/YOruYeNHI7/pc7iFGVwMOtrC8E8ohoN4SNAUU+FlHOBQE7g4k7R/xYzhfWmksYq0rKBzy+/A6g2
GG9eRDb5i4Z38/GfUMy9unfzOCchUCre4B+cInRn+TiasCRqRD9VKyDN4SzC93Kl63ckCN/S6OL8
dMXEXseVU+Daq3BCkHCMu2MSjoH2N05OPzwrR9O0c0PrT1r0PG3LkpnLN128rGR1f5/ElV/Q0Kun
e6k88frbH+zl/Njewnz30buO8P9+sf2xQCB1esv64n0GXFuXdlblVOoBdBzQR+cv7a8ZT8fmSztY
Om035kw2jjWh6xIFe/wxaha0LhMSq91xlpKamRqmu1pwmfJhOw5eXbGwX/9vVK8+rMStcXpPW7Se
KtaV92zsrn8qr3CZ1op/Q/OohIWkR6wltk4sjSci7kQRwMuda3CaUnovhTA6RooR+4VT/P3SHfKE
OrsxJdEVlbVBDIBYK8sUbF6wQJzBOi1uxKgXvJvIiEtRnjDnd4CIasok1IiG+Xkw5aUJlg9IEhQr
4CcC3qDn6v/wJNTsBrGqwTzRSgMd9q0RWmwCTDSDUqQvbBpzYqF70G9Uwech8Tjx1JjV+d47f1jP
tUp9uicJO3d3SA37wZTslOzmesgyW9bU9OV17RPHMf7LnVlzXFGNaj4tVG6u97LKPfevhqyNl7yR
hWcike5LQF4JNOWk87+JlQmo4sahy/kn/CimZY1+0twc3Fv8tAdw1QCWTeHCLKKRxbPcumbDGecC
Abq0mGkzslueJ1gG4M6y+9kxaGAiZvj57407tYfwtPt163RELKYJjZiFn6fEvkNTjJ4CYnf2u7wO
IHZDEXIRJKd0b1CJV/wuOCqVCVGTUzJ9Pop9h5QaKYBfr/4AyFmkfQdkCTC/ZK3s4LW7LJ3AZ0XT
OVqiMws7e0J9ON6aUauS1enDCvEuWg3K7Ude41MkOQpJ8lS3uBJUEVOqj3vD/QiU625kv8QS1c0H
mjC690Uq3qGUFwKd1BD9Uqr3Yx4RV1Wih/RFS8AchSWfnPpzo5tVo8SrWLwXN+6SVWqQXcDAjB9c
CYh7qsNumf9stgiCHPEYUFdmRa2UCA1SYuuhs7NQieomvFd60gpGwVZ7WXEdSEa/ugYcqGzbs2l4
oIEKcgarC99ZlUx98WC8CjexNkF4k8GoHZbnwbkrZs/XMamDfCbvnPrMF6cMJ1zr1gPDzKRHXVf1
JWZQdcm3RsRMBhZWgiOA52ypCcTyuk3+4xMj/qGJb7CrIqZ4gfPmtx+lHWp9BtljFucblYubj2EO
axBWJXcILrAldvTCwnZF0NdnLTMm9/T6N5X+U55pzF1Fh/2Ag/STwMfhuq/9ExsbI5CdfRMlb5fO
0I2DEQif2AG9zF4qAKSpsLZYBzgEongb48M/dTo7djc9/X/rMaQZpfs2Vkdv92rwdUdpaxaVIeEs
UPxe2Wn+3lApv6e0IVPXm48EQXEpIbonG2tnV5nktI/qQlfRAWiAamX7pIBNB97Uyb2ktY++I5Ok
fLXvFtzIaKq7u/cBmzmUnYNWIVOsWNMQBAsDW79xeIM+H1BbbwZPEorSfhe8w5CfCQKsYvv9p9mt
Kerb/rZueGyeE9ABdRDZtgY+L5BkcAxqt1os9cmz3j3OOxo27UovhnwoBu/rKH8wVL5jNX+EJNrd
a+HVVclsHqqki6ZtisAwIjWHxbiJW+xMZGZVtI9B26hMrIodZRarLARmkrEj81W/USmR9N+PotJA
3DZ+ddaOcBzid7qQdAUy4PrHXBt+ZrcyeFJqnt/r0WmLxU0IMPiIP0LV/b92CTCc0xD9hjQYKlNH
Xyq4w20muotIzHmoL6Lv03dEIFOF4M8kdBp/lROYY2DDZnE73OovExvz/oC3XLtnWpLwciipiFg/
m5sdGpXwEc8f3qaBhC7XxPak5dNJbymryj5i9XOYmxH1+mxwM2b8hRszJt2TK5j+7o0F8X9OnzIe
Ry6fIfGRtU9+gYPdhpz2QeiYqQYoSkwOR7AQZVOVfRZien/ibMavhrrB7aEskZVXA1ZxVLU/TNwA
dlR1vlfdpkA3KrSQOfYD1EuteXj1JA4k3nzrrtw5/7IOeJbo3n2buMLz5sLBe3521BnTgUUlyId1
7UxBZ1Ahlksb6qZCRLzydg/mSipAiD8kjeuG4ivb0Whp6oBQrSDDTuFZcRNhGgBUBpkaBNj6DiUh
p3Pra38XekIzddrVt9dQkAORDWdyc9ejE4+gnNsMUCU/3IWpBo66XZGDSqk0oIr797K0WENdFUUD
0MFG4X8+HJf+rFPn+nuw1Qs76tuq5b6QFh/BxYMKrJOFJVO97Z9P9ctPxqvc0jRDfNMDvsYTxRSy
hjVP96fmzleBH9Mi5kjJs31GZeTnYNNbPpgG6RRXP7jjnwU9kpRfdVQaiS0s1Ym8EAhSGtKS5XSp
DeDzIaIMFypAXR2jrnFZd0mkRS3KhYsuKwQhdNgyM1t1rw1FIAtLJHn/R0pv/jkh7ZCy/aXQKUIR
ksnlWCangw0nl1ewkS3VTi0ag1zqFWIIDeYziSbXPe9nQDg1eiHza8MzKZTlRb0kzRx1+qxhWyeQ
AiptBn9ktA38t5kQnlgj+iKxsKAXuUllmgWB1lihffia3D1DJYfixU7HE3rUDkheRNI73rpGEH0T
uknC+3H6T9joTOC1EN0R9dm1J3Wv/meoFIL9/sTLIlPyBU6id9fIK1l3gmP5WZtOjb9/rIwgVx0M
M5GBsc5wqxwS6pESUIHj06/u2huYALLozgAsPo5PrX+MWwcjnV+y28VzQ3nH/Hb0eDwYCR/s3dAU
HrcZEghURTdBrlrC4GXA81XbjU5Pa4CL1pXlji8u0eHuctD1Ndf7vyJxgBiMoSE9bKGbaBt0FLyG
nVGid38TjJAHx3fQEWGe6WKX34T3o59XC6IB/DQ/foKCHpt2iFl82IGsleZE7nmjYLnj+gNmVZYX
cQZg7kZHrK4Buhcl6Tjvv+lDPkEUzqO/DgPrreoEublcjJABfVIjud77ZPH0QEXoTLtxZ4MdniQs
gpzGv39KErggIosBMOsz06eBxC68oAWisXYk7z2tstkUItEz2URY1dEAnciAhMJVBDewKiHUShkq
+Gfuh4jeYEtxdINemzdvaqvKwK0kjejysQxezRAQWcCb3Z0rQci+ieXNFjlYoMO9xQxUa2sJFh55
S+8vKGZ7fDt1ggPEtLEEq7XjThtfknuXuhr6nFIQ2tzYXb+2SpttXJIh7wKx5BCtBVXley8bTRK0
+4lJmb/4Wlg6PAwT5DTBqx2CYDaEliCk0RBzgIUyGoDZ2d1IjzrQKnN3GxJn/gpqG/sB2nUhzeMM
7AZgtba0/4cNYGcoAEoDmmg7hbNQM48twO5gd6eFO9aj66PYo2CQ3fTKWrch+OIzt7nlr8BLyDmp
B3BDKPEy3mP5lfi34dp1S9QcGB/Cu8jYY1PZYPFDgc17MeLA+c31xSAXl9pvTpr11XG54NkkVwUV
ibVFO0tcmJVNDnfOpz5zipouz7pRpGXxnzxfEJqgoQ9BebN15T3lYI46NrxNKNA24h8c/Ruwwa4Q
VRJKkl13AzZBx9a1G3PNt+ovWPv5IQ/9bmRF2yRY2rQbp/ilEqCGEBDjLNxL0EW0jpQBxWGSSKLZ
lCOFAoi/yQidGvtpNv3rVPPheqDkAcxt+Rnt9q50gV9SUVyiOzPzGQskqKM0VydW2EVrCZ08XgRy
gv6r9976PPT3v5iOZA4CAU1TEF4rZKwE+lap4+XiUyo69oP6k7T8lkTOiUo5d3G87Q6leYZH0m78
3VTtZD0QSd+yXcvf/NSERkKIMYJA5uxqkAFXRZZd9t8DzOWdSsLoTLrFcG5syI05cMyyN7BFprlx
4nfmLYba/Px5RaKKkauPTklpW4Mr8BN/JPIDFfnOIiYRu5sr6bl9nPc8cnLshH2NUlJdoRFfG/Ht
WMm9nK5Z2uBvmOamjRghK8hdLo6GakrOsBjplbiUhbNRLR2B/JmU+T2vuiSxpSzxS4Eg7ssTO9VS
4xeycjrgGUP+c7crosqfkgVkm5DryE0KCxdkRdc+KRQMwrvtZ7khys6QCM5/l6Y6JGjdRFG/eT1E
c4V/POQSec0b0Y3B0xFI15oQvJxQZTnxyXtLOKdnXhOFqFiqDcnrq7MTKjosEQBH/bpoQ3dxqtG8
T07GJP5LqXdJpRY50cWf+wMXD2XbQ4/19b4wPJDDTVlo+33AUq4RFRzYTuT9XgnUGdS4ChMeOd1k
7hxZJ64OwmI2MDDF4rf9k97boXGemxkWuopkznHNEmQaeWCMW1Vk5Yvp/H4qu2Ot4gmYW5IqVcq+
ovaKfDmivTBbKpk0Hx/VRi61TIKPQWFjvDbm1clc/a0KRtjSgwLRAtGjjW7kApbUGSX66AY9Yw1j
59lnZyUmlTsQRUVgKdjJNqZV6PgczO6pRYQJqyNNsm+aSZZJq+KnpMHJL8UcSjcPvO8Dmiir9R8Q
GPG19M7JFIl+WWGZzP1kAcgJIDRyWASkd+HiYhfIN7JlO867zhpQe1gXapvp4QZd7TjfYD5Y9bf2
oe8YFsrBhJNTfpcHQaKriHQkUzddrXmTtYFqxZxeNkoRjPRbLlPo9Sg3B3y5/x0F858NDYpYKB5k
Vi5eFpFuruWKmvnYNwbq9o92df1AKeCfbVnARTDS5ZjqtfYfsJIjoaeBUj0yI886ZO29IrP855Bz
kJgac3MO07NAObU+BcQXf4uL7FPxZy0YPvkghXohU1Yhs0PbbKadUFXOXhnu/7XL+joKt5RCFfWj
uwmweNoaFZcEQcL48dBeqJ+LUNoYzdA+ea4jCiheIg6WYCwIk1J7eDTFBFY1oXdU1+7jCK1tNq14
/t36U1kzyITvZdX1I9cGMxxitm3PTyoMfVRtG4hpCgZJ80ciEFevi6RbOd0Fzuen9lSXYW8yGgd5
fmz/QL0VS/TKatf07fgWyBKr2U3aLPtwK5xtFhb8bfYQwXd+uqiZ0vFSOy0JsTUcdflEcQYHVFaJ
mM2/2ChST/3rn4wg6dVscTgnhbkK2d45MA1BG08CW1wHZtYwYBYPWVV5eiicOyL+UXnS6OG6REE9
DRfbchRwwifhX748ZDZgVl75OSbsyYAiNNX0PHaB4VGDidOoZAe9n7BoKugcf91PDq3TJaxmHAYi
JV0mBwigAz/1+n3zh+eipncIswmzjxGWj5H6UsWfPFJ+pyZGPKMqA6IUKxfh0SrjvZGTjdXecM8Z
emxRe9M2d0KRpGkGdp5yfPgGsHdEIufSj6tskS6CqMcZyetjfetKOgJeUVh2eTrSSg3rDakCcLnp
1AX54OEbeCAdC7o0IbeSGsIV1yHdnB/hmZbGmqsOK1lKfZsvIyY7jOtz+iLtvRdG0cIVCK9fuVHT
cQfBJfAKpwDFAH+hbQIPELCtzuC2s5JjOlj5+9SMtanEfJfw+AfdaOaXnzwubNw6VGIabevodJbp
BL/zrN22h7aXM+ifA5MDJ5jdUykYp2K4HXH6OF6/nkMZm1gA7WF7Ihg+gEbo/2bjEmP6PkhhC4bt
W1BrhKrl7udGIuU9nXePh5tXWnJcFpeYG2lOD5kjwnNUg1ZI1kl3gHXOWZo2RHkaWPvJHnuw63dG
GBKN8caOXnoNgemle1IAdftdImowN2j0iharhK8Ol2Qrm6MlQtVj1PELgPE3k8WrNnQKG6BBkDgk
KywYWFI3wr/nI9zxOcGbzgqbwc2ICtcyooFbch0S6t5n950Z4WxsXT1BqCdiTGJNZSNG72v0dZ5/
KyB584VQmLQJ84ZZZsV3YJH8yEAeAfU95Va0wkFf8EZ0AoOg15LP4hASJFDpqKkJnZUUbE9uZ6CT
SYYhbi8lzqTiKxoifxsq0rF8HEYNMeaa2bn9gag+GktK2xfRbO+41usc9pV4HjMYNE8ABLlYGT//
pXMcSRy7m4pFuUj85mEi7jHC3Lc6Xlvv5lWs2DDDo318jDBaZwyLmaK53GQkZIG4EIjLeYK7uk84
DzVXu5hi5VDRXiS+Ks2KST7VSyRiw6K8Lxi9GtlT/Ft/7SdKd9hiuR1o8Wbt9ADQqgBZToNO1hSe
zDTje4WesG1ywOonu8SUWZlE1W3gqYBtZurktsflfdos1L28dvCJjyE6Hk1X4DCjB92nP3Gbbfe8
lHlDCNkELTFZdO4KS5FDBdTBRrRddPTVxS5BO//zAZzF0ZiZtQ0/63pB86ND/ng7X94ugNrdpoxo
COJWL7xezBO/vdd1Mg3YAgVzCqcjDeSMY0jvftkUZuBSOU9LB8k0qu4We7egR933ib+IzMcRj4sC
80SDdxOlEEaA/IZu5ninaYht9AGVdw9tXZJsU9WjaVp20cV1hOG267a/CESrrdjYnttzxwuoX3aC
JY4hRv6H1/MijDNJDNyVJ/pfNl8AXLnty1tLUHqhNCAUBjelvCGRvPgn9QB/7vpo0NHK1CW4n2nO
UZAzbLFeTuly1XrLKqeGuPNDT6XRyny1w+T7ySM/0W5ZG5bTeUr6r/AI5FwHpns0yCD/4HwdPGLL
SNOnZN94S4sEYj1+c2iZ6asOQYcB7SpDpU/qKTRUFiekpQdS313tU/s7/MYWp+2Rls/feRG3xXZc
ZznT05IhDOGWehvm2xGZwgmg2QyVFO8v1eoUaUXw2XmYTsiiZ45nTH354+l4LrmqkMbh0EMEBoie
e4hv49NkX6OKazgpAkETSA/doZBAWxm9qrjFoic0NKMx9o1Qg8ItlLD7fJDJOuO8J8QZePdoFkZA
8qHqS7fvyY+Z015nsxRW9+Yg3K0tpAFmMlRe4GQKsfsHRQqLNDlxJEaGcE3fsYIoaBI2Mk2BWGYc
111Dt0F11kuiG3e0Q6cl6ASrL2utrOoxktdrTOEapTrDO9FBtzgbhZiF2JEZNDHhtt4rqVyv+em/
q3cUEDOwrPbd4MBTfnADZdnebPChgYVt6NmBqDwlfse0YmlZQF2Dk+zemg+RMJ6zvd47YuOYmPtd
UCusjM0nD/gSDSNTCKjYYhZb4AVljpxm2a2Gt671VRsCyYqN4/b9TTamBcRC/DILAxc2XsYS8LIr
7mYGfghFEy3OIkMHiWqmIW+KBhF28xOl1pOrm2CH50ZyszmV83thSnTchES8t6LLNYT1ZX+jKPtV
dmRxix0HUAe7+gm1H5pWskzHs4q6a/u9SNpiwVMuyjjl6qxzSn29NI2JD0a6503/m8PxnHrHnZq2
CLFEQCICWzaV3SQD+F8dfvVPwIsnPeRgzjjQaUddNZQO5GDbwhmy3+dg/M+kI4bshbRgIPdQHNuO
78yMMxoBrPDVnD1jPQLB/pM1An/l2WJhRrD7D9VlHLxK1b8E7Wy/G1Kk5XL8L/7FfpcQOTjhKYB/
QK6G5pQ2x4NRWoN8x/3NWMl5LSJHoopvu0CW+zSIei8YXHSGzvl1bAGvbhCgCpAQM2BnF/nPFMQ3
hYvpZv0D0bqN7YIPEo8g3MR9gXp4Qb0fVheE1pyIeIw3zlMI8ofqOBbECNbpGwLjCYwn6MbEhrqF
c6Fw73cOw+cFm6E62r2jv7TqlTkjGnRJ4sw9DfxGr3gNDbyuZvPjgj4TKosUXRuTT2n8kSR6vcSI
T904hMsmEkscYkeg2uhYxdAgpo96wcv6+o5ynENTPvH6PvVs1qRnYAj/TvZt9JvblWUqnU5lbS6c
tmwdiCuNHPojAwhhQYYO2EhN9pvgruILpsRseNDaVVpEbeeGdv6J6RERPh9WLe0cEjTirCR8ca/U
98jAhhuFwIWnVtK2g4xh10r5EnZKbz8xsE8tW+9NCBzzC61NqqJqDXEI/CQILgc38p7qDxvlyEQf
4WI5D2SyoT6591++ipQobWoBUX9zqc62lz5pzyEKKh1/yT1pPyf+LVe2RWPYq/ZUvhPOjnjt1i75
i07SXRYgM9rfW7zJ6+4vFLoBNOFy5scPMmjz6W1E8C6QT/dPLldEwC2m75SkgsdVIeyICL2zCq2T
HnBGTdb44e0nCxgqr0xu8eb7FNKHH7sQ7Cbm5ITVoaUz67zbaQT/Rz26xjb0JwsHxGPewBw/Gkil
YIrMaypS6c/RlyVAFHpyz1aMs4HFvBn+2yedhKPtApfrjIuzrxlhS8HvdCpDoVpWGzsskTagJQDs
jJWNT5ooN9apABAK5Cxmc8vnxwe2SfiiraYq8FixvFwTby4PkntG6Bx8/T1TEjJgy3p+GYLXHxt7
siEW4dGStcwZK+9ZGW+vxS7j8tc+StoShekZgRymiurD1utlsduQKSUvmajYsCzaarPB3C47m93E
3JthLyLEEWP25o56Qf3R9/w8V2GJkpcevuXDSl3VsyQ2Pq+h/2pJzN5kQ2FVRWHSisuJud2QdxWi
S4+EWtU0ldQ6pg1xasyeNFJQRs6f2bFNiQcU6XxwjOkMS+ny4AagMj0MQqTxwxbvmKQpZdxwYLXW
GfOykGrTX7cIerlL++BEe9UiIDm/6dxbooZ2J6rt6ueekRyvD3X6UZrEy0oLAcFk3yBcsf6Imbmp
5Xhq9dK6Qml3h5AcPM7+FA2SN6aJpSZImYCe10P5Q5+cSPOyShJKy55gDRPMs8q6dARIPwO+kC5y
E7VrB/Chc6bh29Am/pwcsDQ+PQPwtjiuOtRXoQT4PB1L/IqrylV+Bto3f4mR8msTcXidz8pdAm0/
V6xzjYFOgoxy//0LwHVf/QrfLSJooWFkeJPtNX5a1XqQ24E+TMWXnS5xGAxPX16KsVVSAGHyYJcX
eMMLFfCk19vJ5E6vn2o+UiPZZ+qJv7IHHBunqn7lmNWxzICftgxhIbFEZ6SdGfBLKhPlESIaHpAe
weyEFVbqNl3FB9gV6Z5I2NxxdMYynY+wdR+8W5UnDDcHpJngha0JeRTj4nI99r7e6eTZAMsm+DrP
aouxVF3h+IHfRMZ2LoznmR6RNVEdcFqLmek0SWajYec0rLnMBcVNXh8Mu14kiM2PhBnw/mQ/E5vH
B50rFpxCqJUhD37Uyzhy7JpNNPkjjccGvltwxFCrzg+LHh1ZTNqktUEP9LRYgCbQRGb/4Rwydp6h
kczOytDRBYiVoi994Ge3QeSYC1XddWa+OEAYep/wmKjHmvgtKe/Ll6Fto6JciC4nxbay9SjDslwr
KzFppAM+vcwdNUDMJbryXHyLlyKyWMSlkWQMUVzgUdi1iXzTLcFeMUGNtVW0ud/DHCtK+9wr88lB
TPApzVPtftJPxoRWLT4R7S4fsdPa2PIY6A3BMKumqAunWKg0w72fYjjueoo8K/QeYYg6LoLsy34A
dn02AzXf0ku0VbN80y797WBuR51HRTobv7dVDj6x/hUaAFgs6nbJW63z/aRpMHqiV1ahIlGVjaBv
SqI8kM6PTHXCTiDZdfGfepB+SQU8YpntQR8jlcvDQKNQwzSKAf9Ptm2HPcyQ9k1Pth351GA9TTTI
Fs7NlDyK4Hg+kW96IF9qvTVA+4isBV850aQrDE9F4QY0UIfdAR7hO92cAG2LDRIQNiBkCtpNO26m
zOgcZPgKxownYo2oOAUK9vKChUWhWv1n2Aabg4NqjZ4XB1MdM3kQT5MXoJBEHwFy6PdtKrG/rlOF
HKlpXO+QbePIpfKuvOXEPDslH+uyS50olVvzc5uxpddNT5M4Q2aKjZtnHW10QYk9SBWJDiLv5NzL
A1LKYcvN8cJWU24hWUPTqzhke7QG3DCv1xuWtnwpuz+VD03fJ+CRU1luMNJPXcQgHUGS6AwYpepe
ojocitUpHzrF9YRcempY9wgP9JH8ys1cUmtNC+bE01PVYGsv7JElHkfSJG7Ai+6Fw3HwM+Afl7LP
pHXOmYIdgxi2hziv3wvL8OEcoomU/71qAna3YHZOAoosJQcCqJ7YukergEvf6g0pgTLybxdeLI1i
wiHUiRyHOqeSulM2NWGw42nBQh9LfDyT1cRH6270hSOPEEWoflpYGcxhIRbCYiMkTA3yW+zxp3Oh
n98z6WqdF5jjNsLZWs9InvqDsFzkX5OU+bPiqiiXDJOITin8OMqbBozWtkTnDhLJBJcr+BsDrZCi
zZ6hlFNnZXzCkxiGf1jNcfO3pgdgipSqnvVPtsVnsktqu3/N8n2m4tsVKCAe5HOZ6hX0bkZNyrf4
LCkqWgYST3BbdYz12mH8+jzb8OhuZ+yBqIh8mjTX01zujMKBf/3UJ3e5VK/6t19sN5PGa5Rlhl7H
lw/Zjjru3rCAcZImueNQpqjjeIlmq/Z7dMWf1L4b33uvXiN+5DlOYBGdc6KGASFp6g4OcGJfDaqm
P1+ILqDQ94KpTd11Z9hQGxAQUWaeyNhHTKRqb89Ri7aNTBvST9S6xyRU1kSFTVDHzRbUtvsG1mzL
g7LEHlH3oPXTNddCzTLcjVk62x5tdHcTuh0yCbdScR52qRkuq2Eiix6xxsJpUkk26eVw+WGmyWlR
BxYCa0X8o4G/zum/bboBq/08p5ICZ7JBJa0nfmhVrIv0X816pTrgyhZD9pMczrL0znWwxyvzUCMD
RupKQ6KqM7/yM/Jy9Roqd07rdSNHuN3udyeP7VC0XEDc+F0eoxaHs6KhhsE4qc38FEmDgXpGtyBt
xmXbGJkGd8WG00O/mZkbDMvr71aNTjnWywPQxkz9LxWd2EXpHObf75Tp35NDioQDLMLhtLWIwNup
biEOlektWWBEPS7qgEQIGFP04tNXjCDsBfA2NjdRF7IQREKC8T75zTONX8bNPUe5XBEVqo4nTGpa
I/zgkLtLnQE3VyCyCax9axV+mOkQeZEYJ9U+ecQltYGENNlRoLzqwo9Pfam2SFphSPgK88rtUSeX
q1wCMquqNkd65lrY5lQqFxYUmW+4nsuHLKMfjW52zsU0EsPxf15Ib5nGPOMsoCfrUFWLFt16Ul5i
IrWbNdWMQLGZVl6zCxoWoIDBZ9/oJ9Y/p5FgOHY/k6PRmGHckHkbnJwodUiS4WrgvsoiTtjR8E7M
J2TTocbiv85e8sN9GCilyhD3T7STxQarOtYa2BAZ3g6m4jZEXE0QUdoTIXIw3RcmkL3YNdYpmMcE
s8GJIlqsH/1eTU/o+J4bt3vuJk+zDghf4jOkwSn0V9YC0UL8TMKbFMJw4L93hq4jFKYMbRjfMEQy
IfTHE1/vfG8vtzf0sBUrzriRMt7NSk5CD26PSWGwdpxSUF5wqKt+DLz0uRXrdyGrFKnsiMvelhWX
kSzPe5Q+8hZ3PhqWUk8dbQ/XqdiZsvq9e9/wcu4ZRL5zt1kwx3emO5VMO3oYXGH+IIlE+LCtnm3v
jb3KJan08JfRlfHYwOYTIYrY1a2UBi7zwbxmctG6t08fyh/NLmsDUMEs7+AyF2DAfMSTom322jbP
c5EruTvtj023pi/EThPHDHfkUpWGNfMuVmYUdrACpEcka/EA0gCx6quFl/eukmtpau8jlxIeMbSI
ybSUjSeDw5j0EEvrusKlviHNiYXlMRLUaSRCVjGDo7JdWGl6GxuybtJc4dDfS+GuPgIGnOVhaixu
5Ddwzpa0L7qP5gO9/iE738pz9z4iBLYQrbh6GewO0gqsh49D765lL4zCqYY+8DmJXSBN98LfDjKB
2x/vAovLDtIUvcQgMeH9z0AsmTLlwRNdaW9S/r25NqsKrTtTzCjbwXbFPSw2NcKmHARK8mWAJqZu
HNGkQC+4s+9Jtf73N2zxKKVraw+vg/41IQaPdZYLffHide1vsuQKl+X4Dpp0tL0hKYUNRJ3Fh62e
IzlVM37m+ZoQ76ubWnMblWFKkgNkRc3aBbIgHJ5WAzLXmc5/p6y59rxQ3e4slF+mJQFGdPzw1K6v
yh/JPuvzM8yMXy9soyV/bSfl4mfN33U4o5Wni90SLsM5HxoNBr/oyaHFWCsi/KNs/ot+KTOupjJ8
FdzYc8lBosMA9/OE9UhSxCR/jA9rs5PEwYeyPfZrDdFW/ItCfuifspHD8WtzdTisEXAr6bC+Ad19
/HDRmqcPE8amd/j5sG3IUgeSxeCt4a3nRv9MxxGTFWHiFDp9cF3qPYZM04jyb0L+xo1g3TigziVf
vxoZKpIKWoJBTEcEKpRNu7c6lfaL8pUgwovWX4BYVdzsELsd1ZosOKpu8JYQVpBH8kA/5DQPDDlN
x5rWFo1TdWgQEHmz5z+gcSmb5hfOoot8SIdv0bAo/l7pabvofsPrtw6PbvliSF5UdytKIh29D7J/
8Q+OFurRwuKH9/X+bc/XGVhGWPSRHKwqPGuVpcz7pFeT8GqJIXJktNvZvKRQwplz9F/OXacKYfPf
1wkTjxry8gEDkrgkodxglxTUF8FJLz/d0n58yHOhCY2SGTQznd5wGkKoVpsSFvCWjKXEH9hfRYt0
uctoYu9PjNJtqe2w6DhtxOiLxCjyiifYjTySGv7kzDf/kDsguvs1net6P5gaDzoTaDdhCljxtJR9
nnbG3MvtA6xsEBBLc/HKvdRG8Hd+NZ6IGjn1bd3DckcKFAHTi64lun+gnGUc14JqFNazYAyxOB2+
bWQHvV79yptpNwy/zMLYktIQ54RW9TL1mEI6pEXmEOfdr5aaAY9ZoUrANfNhDsoclbfwpQoBurDh
F6dox0ua/OfcasmrZW58ynHqNoIGy/5d/IJmJAhZF+bIaOTqRVWjZFZsXS7ey3mEvaYdoci00MY8
osgpclDWv+tqu6Yp6AUUsBcg0tzwoWU95g08kDUAyF2ZYWj6HJDFZRY2QOJD6A5u8SWPey+G/SPL
9xSPP8VzI6pk2uagEUO6S3NZED3sau+kdOZrKghFYXRnd5xFLg6KXzz9qOw7hLD5mhVl5nF2Vi77
e7d1jEn10on+sFkZve7M5ULLe6P9BL9rg/vNuKAC1X0ylVyzdHyGRj7ocbhIXcik8nna3aYaz8E3
xa/xbdFopBWn7/lRNpQ3zZFMBzI8kz6QJEAB5MnLN2rFXgBLY9l9YEF+VgvlM/hVJnxyCguxBrPD
4wV1QDQFyZleYb/tjFrWWrWc0VreruUH96SXD9vIELvUYsuqr0YJMA/aToWB7Arcy4+SdA0sTSQO
oOT252/0BcotRCUmKaqqqeVx9boEV5Vu6NdEPTwpfMju558oN0id1bADQWcp2h0k61mO+FgfcLRP
PlrcdiYOtcaqy0U2bgTmqVU5LF0bCEIHy2YvEt07MWKQgwXUeVGLm+5DTHfswzMRH3Dj1z0tJnMz
ZofHb0LkFxe+TuEgDpxx3LxqpKlM/XtiG/y/sAs/kgOzIHHV2UsoXaYYngpQi8KJ9BYc9RSx98Kn
pJoiHiIzD/u6B6aTKliEaM0m8B+qy4eK5Z8fh+TdHPc1uqttWDnLZ7EZ1qfclIzcoRzo7tUIZ22C
r67wvUrFDJgyRdY1yE+pHcX70s5LANjr30seHzzhRtuBwtk993FbFauTxTUBucbps90EYX1ydGdC
J0CpAtD7gs46+VEsvOgBrXnMxmnXuJd7nr7oE9Z1ZQH+vMScxbTHxyCLT/bR7bqbqVVa7qcmvD1Z
C027r04P7wTQ57yZb1sjxeD5reWjcgJvjBW8AU3c3Y5fg8tfxZpdtwuU3yhVUVjKUCzVyzy89xG1
KpmBU+FcaXsZTomWQvUBdEwfi+MEZlKMcp9AyUq8br8ajmm36MhOoU6yPEeAETM3bq/lnYUjMtus
jZaxMnCP2KjjYh9aQG1q9uLHS1rLlwYRvhVv3uo3DmsOE6AfIPSCL+xoafE8ivCZsTL3WqqFjM3J
eP+YeUqWcjR/8vVrwJc1FLsy1OCoCiaYjl3zkIvRtTCCTitE78FJ9jzMq2yPsNAOSzVGBUZN3ByH
rDymQJSVfql/Wmihox10eymx042v32kQ4qtOAHLcvQ4Bzq/+KlMU9tQ8LgZ6F+Q89GHr0f1Yo/x1
Y73TNe5XU67AJANqxTG9BcBCgN5io49W8iABcYodRXM6UoyBr4sPq6Pc49D9m0+XDXL/WDQpQG0f
iZh2+tFl2EyK999WvBuEYTEJVwxEcAbI8sVeZPxlP1kq3kSl+H+DWOKSEh97/PBa32TCznABOuLZ
tgR+pVtxC6VV1NyGjWkr5apFSVPlBVJVyqzlmGvSw0D3gDebTGze0ZzShLSabDuKEDOMIwZ6kDeD
LX36E7aqmganHl7PQib/8Z3QYeegGm9ZqAt+5VU6uskY6j2sO6N+QZdKoPl9q2zIsTGAirEvt3z9
sE9jLK3z1ENFbnPx9qzMxjMoFzYhWFc+9PLK2P19H7R7PJhFy0X97tg07wA3kH0B5V93jwwuGfh4
0SHHPPnKOmCY3OePy0fzUSxfUXKRxEmLjgvJK2PQ/nDzhqz52brVaZ2lvW6qswI2z2lUI4StvTls
Qxo6O4dDjuSeiJydsWDAuja7pIkm2wtwEUORfVe+msRe4u2FjZrcd3NjktSHtltBrfLSGkD/HSqu
uWZZ5eB8J4ZolFhgo/QzRgjoRk7x/4ehyAfTcXzWxz2cdx+pnz2vYkt8HVUgiwR5eh93zhhtBfx3
GMIuIHEjXKlGA/lZTTHyDZqUZAk9McblHu05BY1Yfm6omiwnISlVmZyz1D2SimAeDJ6bvr810azt
K4CE0VaP3iwJKlWY9WA8siCdIOYZXD1B0bPK/gxk3RpOr1ZGT39AzZuaGsG3o4PvaK6FtCoOjObq
li+I7C/6fWjQcxpe7CTRXQfeqcKwzZd7yjxAZ1Tm2gRTGGrNMDiaRoR2eJDi9YQaxImtZC3PSF8L
uQEbD8k1XUCERjpgIKaaJf+xzV7PQep4/Z8jf9AXnEHL7Wtcpms6f6fndv9tq7Cy8pUJGOol7tJD
tsiU0Fv+mmiVQB50e0I+Tx51bntXxRqkucwIf5Ad55IcUZ/pnksbfFjH8JXkdqu5Ksbr4/vzx1et
BvEI/ClGC1Ze+/ntPGbT79YGKFr3e9cqEDBddlbWmsaPQp5M+BPkwiDXQylgpyBT1OwUY6LPo0FR
xzxQE79+zZsP2uorsf93QC+8kV3Al3a209E/A0WCylRtasGiDRAbQZGKyt1xZjm8Hmjyr1VUbWv1
FlXWeAL70eNTbjNUldiFIMUJ3CUO5C0w90Aq1Ca+Fu++yrlEJhaTv0SCX7dpaWHHLjDXgNDB/h7t
Hcrwr8UmaN/n98ol/xmIbYy6x0OluI0yxoWwpcE5fzO8ohun29LPox579L2THtZIRnWeULHWawyi
iUCuvWUHnUMXmpZo4fRqw8cB3tHyAOdxDBL/hayT1+RipBb8+Y6ix0AbgqblQdomD38cAngDKB4X
DDBTM6sPn+vMlqWptT8Zpb/yUaySVn4TShpTJpqLZ27b9X7wtYthc1YJaCvZ9ImsoH+CnSYB5R5a
dbzAtRG74IL3vnA3T5FNTf9zGuh6RQsWBvPSFoiw/Any6TXRqqyBKH/Qfb+GR/CCwopYw/2NAQe/
3tYC7NBiguTVNPEutFGKeCCsaDZ8pwCRbBpsBq2ZMQp54j4rpZpbnV/EcA91WG9noxGxciLRD1ly
e2Lq+KKgl3CxOpa/PQUb7zqx75DFa5IuERBZmVPwY31oyH/ZwaP1SfF4cYYEjAugeeswvGM02lA0
WlxpoLmogpZo3/Z7Bs874bEZvh2f5kEs1nBwC0kebQ+CAvluwrvf5s+E8ukWijojqYBkr9gSEqCr
J+UWpNqzFcG561bgDzCNVCQaF/EGxWPbG4/L+U4dJGYEvfomQw6kPqBP3tXQWvN9E2cWWLIjhNMG
nF8vCU3NI2PieSGi3Kyu6uk7asGuEL9AsyTU+XrRj5CnVZuQRYzqdjo9Ea4n4s+nalibzl9YdAD3
Xo+U6dEo+1feNHP+Pt/8ARlke8t0GG1HTUJJNwzuvRpUH4Nk0ZcKYfhgjbsXXv8a+Tus2zXDGAOB
IgFXINyeIbtl0W1oGdkTI3x1P6P9ChNwwGZ77aB/v2gfF2ROXL8ThxKsemLPjdMU4s0HjIr8E/A6
bSAbdAvKEJN0KWf2wFAPEFS8SVb2DzeaGVT3f3/5unqM2nGXQsqVuH9z4T6EOziJYZ/vDH6vDNaA
tC0TwIp/7sLGjRlWDcEXEfrfKbqCPbWeyJnjvWpiUo8QAJAaaz+e+eVvYrP3B7E5gZFKvf5OngTX
Ep2d54D/2fGFz8zI7LYJd00hElbVrSaWyb6eAcNWJHitw+lMvzFKV+suB1STXkhvxNYww3AX6SUn
Z5ZapxrK8KFq6bwMekUk2WjNsat2QXTzRQX9oRzJ7IB7XdPXzW7mUlJjiTc98h2WGQcoixhYervr
xFwe7TGKEgiL7VnLTWdrNDZh5jUaQF+pIyx9OR6PYXsvTsMqwtN97yAZM9dbu/nduz1eOgVRl9Sy
mZ1CHnIKjFy2opsNY+zLhqeP/Tuv5V87zG8gjrkTNmOkz4dhi0g7pI89b6tMKgnznhiWlXz4yguF
QSpncaSYwiD3DZiH4/4rWNFIp3MuGn5L7hUxJWkGJvA8Sod5K9Dyum3UTzeo8hzvYCarV3vIOXRX
3jyk5RQiPTqGlRX+hRlpg23auVdORHHjejFjLpVVtBzfaxhk0RDZNtvIvmyQ1w5vTP30Ob1dRoLM
CikKH9hSAe2tFSb2FEEv7dpsQKB81f/bt16SIwQzwcxD6uRaIeYPHxLmEF21aMNvBhm6/z3sWCXB
tVHgoXPeA6+iOrNul7rGwK3CDwjUv7laF+Zx6fW3z9af3MXs/i/1j7idJoXjpHfmAg6U1ZRx9Vzj
nmaODhgqSe3LBwlJR9YvUJNvYKIYqWqQ31oDKYPJ9i6hdCsa9c7TndvyA/yODDRD2GsBVKr7INLU
vnhTXYPIpK5CBXAeZ9q0RXaiv2PYTaXWwNq/AgICX9fYgGdK5AO9/81W3b8CiHSLSLSHDzHpzlKd
EMTkjDHUZ6M8Fl7KEk8KpGriyLSGM/HXi/+hEg6dSyM1kr7oJpixP6ASoWiUEwCn9mn3J5PTfG2W
WTurakmjDQ4hLBGzvEOfRnIXfa6VgI4iuOHByWlCbMPsEt+E016raq0A9ozZkdD/oZtuai6iYAaF
zNSftJPp5iLcIlQV/YCGlvomR/wKnij8MuDUloqV1OJaXyCtM8eFDfM4X1Dt3RwS0pMzMWErowVA
nd+hf38mYLvCzWRflBVeGTV6E2LtBBPQtDFIZRcPyx5DhGIAVBOborD8vCCuUe6G5n/bf5ylmAbL
q3VxTqgMRdnN+peSogfJfNDHtrV+wXZbYxvFldJtbzp7KUJCTznV/awv6ks22MIFrY5If2wXviTt
4LhPS4x3BsyibjrrX1dCaGQky1XQS+61eM8mFa/FTPyOimvo8GPC7NZDIRtEMd9VTnDjsvAXBl9p
91o8HaUAQl6t24Zj1W6q9vrh1VJIW/miCIHoGcqSoWwSBit7KhyYvQbhgKFJ76e0wKf75R6M7nTC
ByvfbEqZEk0klZOV2aKvg7ZXCK9pxnx8AbmXNx//+26DlBy/d0SSqkswYZcy888xxbzfkFccjQno
cp+9klgIK40bNvb3bG4G2WlyTkMcX6hpeHUVmdcQUlzofvAuL3o46pNE2aZsr/aSGTCRNjea61Ja
GBgna2W9geezySxaQVxIwyQ8KFJP3FwoDyh0DoxsrEqTDj5Sdx8lp/u7FYarBvHuZOeToEacbULu
DvFlk4esAg71UVn92zPCbxpBtcLiA2b99lKqMqiMg0mBxNy4sTflFPE1Dlr6zBuUJS/Ytw+KKGPP
jjeq1L4B8XzSHCFDsodIyObHWEPmQ2mUrTuK+baHBWn89U8sQoBjOsTLoYZDnuPm9LpfypDvFm9G
Bo8GDBIxG0YZVY997v4+T/CWsUr9eHGISSuh3A7JTElZUHB5EoN7637uoUCe7IwRM7xALeBiMM/i
UZuaLuAU9lK8bA5jBCstny6iWTtRpcNTV2mPgI4gMDts3TFH8yq7wYYF0EuM+XIZVj8Ac9rn2tbO
ZsOqFsBe4Lbv9na78j+BgwSLBc+TnYAJcH6r7m2JeM4NsYL+6kJvNAusC6amALcSl7Wc0RdekJ2j
XjucKx07HgxBvJEdYV+BBzB1lWUC0TZ606jSqgO2iulxRRtVhxwENoKbC1ogn/iDeMobJp35nhL0
sqCzhGTPh68rcun26FS0dKHr4S1cP2IRxfSh1hKLzUvCHVFUie9rKeyR3TBZ9dJJ9M9wJ72Qn+sy
DRV1rn1//GSKgvaGZa2WsCTwJltYO+HVUWLHGE+kruKWFpS4LZIZFIsLSaGj8lubTRWqQzwAcvbz
F3iyF4fs8qHLK0SCzPd/NT7CZYfqKTSUo2O2zuhQNfH8qc+n0xvNOWGvNV1vSQfm4z6Lcfgx1IHT
4WUktOmV7OhclpsxUmYfiRo2zQWCV1AHW/PPO4Pqv+CsqgUlmg5aUzuqfnGO49Ldi/3y19RdC0lv
9rdp1kxXId80fd9c1tqGCNZ1q3C1353M+ckS2PH574qK2gbi7+tBytDhEzApG+c1Bp/AfKKhEBSZ
CEEnOcpb9yJHG9Rfj7pjtn6FmuvY3FG9vLk0U0lNol5GWRdh8C1yvVCY8YLdRweK6yD8feESZqT4
UnDnOJy+mmGRPZxDfED0m21IrSVPaAxAOxyLfVTMX5L2tHfYlEJw2q5NnAkaxZ/VZZMFPwubRnQy
7BYon1Dk4Oue5hwGdwas04RZoRU2wifa91v/0YofwOeThn0KmUucQ36+OLJqKQBO460PWUGJb00A
eUR1+nnODU51l6JfAMtrp6uCtloQBA9TlYTfPQFFP0bklC4KVa0ic/tJDSc/V65zeaFOQk3FdA2k
fIBg39e9N43ORafQjJA8riSq1Wz0Jwu/8IV8vi51qmbpQwnusWV7efnFFr7Tba2HFPx7z6rnBDwT
KscDfMFxPiaMUrtZvUkLADodKzuSkKjrnMhvW7vVslHHCYgqDmo9iSFiQlfuLQELdvA50liSIfcR
MQgiZoCt2YJKlJOGWR+57XbEZ4+ZHhBQzy2dYBlOUBKCdpfgjjlPpWZo0tAN+EM/+zvg5j1na2dB
BlWWhnMCiRUaBooJZWRxt5OV1aHX41hzQb0v62hnwP6NjEJkuGPO0LAXkRQ4mmNMVNZVM8HYfXbf
0XTRwNFqJ3xRT1rGEthhsN+uOH7jT4/rzyZcepfI8YPr2XTzByAyqZDyEWYzq0/2dEoUNo1h6LAS
ubJGJShNeZ0utWQSos1bjhOg7BHux228NP8Kqd8zs2FwzPopMoApbGgIYoh5FOsvKoSONBievzy3
36YSFdecddQTnHWQjQaMAHSrW2hG6RHYgIDEU9jA/MyOZ1mwmEKBuimy5YUpRfNLHds95tNK+u//
ZqMyzJLuwA4efiLWuK6fx/2EscOe+4YNi0kWHeHQjDF8BKLBo0vYHyXlWJA+4TBSgE/LPzbEWncd
FrUNU528QpoMVh/t04KuS0oG99D6IHtOk1ZE9fvymTH4ZnR7tSqHo4lwqBx0EymVf299HVssHqHR
56seFXwRcRpRNB0o0v8xDT25q5xkVcLT5oFRWMzE8qLnA5BKxmcI1C/pxkoR4reQtXcYn6I/Joka
/DAagNVy6r6bSPmsSAHtmwiVS3T0Pm0LA5ClY32yj8wiaKdz8us9TIbrkFy1H7AwzXcm/khL7Jio
VDlpszybgsOTPSjL1QBKOVpTazA3qF4/z082Ux6nkx2ADLSfRqJNjbzAd0Pgi6iEa6p/j2a3jHVO
50oSxQ063aFpRXlkz3KggBaSrkKGHXG2OsVzdWxQ0UApHYP9agQTsUd6uL+NundgxPJ06WrgEMU5
0vlVT5icJM13yb7zncf+CcYTuuE1jHp6O9j0JmuGq4XNXKB2fHSxmsJ4Fg/Qm8jxOYhfIUXgi2Xc
l1krF9qFogS5Zb/mhZC09CN0f2T/iECkBOw0qHg0z5QEMZXek4vkjbIRyOxo1BzFlzCh+Wn61kDi
pTIAyWj7DlzeelHIMYnkwRFu8xTvDQXScbfjqCDNLp569FjiiIaHtjERSY4vxSxNW/Phsl//3eRf
YfZxV5CSyGYaq++Lchw9Mp92XLILkqttC88yEKk3J85oA+M8qSiHIIa53r+zc87EtqfIDKmpAoxW
FfNyOob0TTBKZnWCPwhAQeZQKf7cXr/OO1lUpc2CKsbacQZM28i48DNCM7yiONH16PlL4HIUzN+n
NqNW9EDhlGR94zAcXnqHaCvltKSFpp6SdjlqNuFQZMJgNFspGSdtvpqali4BO1qUA+QVJX8rBcoq
uMeFNTvuEOzVv8oAqBMk2O7DPyHAUgkOpJrZyuckuSCNKNgb+J4Mi/tpfU8xbn8Lw/8xPgKaifLI
Va+Ux5/bsK79dvHlrK9NK07vNTj3w8wZBXK0JOO6vS2bmKWHy6QwcgVIi42ezTWYAzjVIy998bcH
4jIdwNBrTyNZSZT1+3dM1QuPoTkbzIweLKBSBFS+yNHyoYbqNg1tY5nu58wvVcNtDLmZ/sTcu5VV
4kUudItNT3/NqJtJRs6vDWcJBxZZRADgK1fCRSav0fU6NIMnIrh3tQSgoxJWG01qmrJ/0ByY91Yk
B+NYmgw07DREQEdtddzXTUhU5gBbZwUQo6MLOGWT7I64R67U7pNkzJTRnteqXiScldHRd4zUxbCe
H5u2ubqlOaii3GwU65VX8frE9WE8AUn4Wk45IQhwHf5qiSh0hPrKhMp6u8R8ch3zZ6zH1kIdxLor
B2r2hY6SMIV42Lv+LDTAntSM0TIdp9awed6KTGAGw2YckIQhYztWTpwbiBo8Tz/w7jOSHepoXTRq
ojwlFpLCUgrC3uGW9dvb5fW9xpbVfiaVIrp/rikRLaE+Lin1Nk1DNVuYeeX8Rz5gx1l+5IZU9sgW
Bjebsk3FYcUpDhFLTO3qjvLap+rAj0E7ZqkKO2LRp0dMxLKEp2vg1zYOImEKnqGodFrxaLTZWy2I
MvCGWk/TnDVORX8+9hKntECMzt9FfRSEC5ccBEQSmHKnjNeC3KZbYBklCbDVu7kufW5Ke9XtQ2EO
Yyh1Ksp/tR+YVzCcbcGTqHLWolvayG0T1UrglwVPYh+PrT75BERPD5sLE8rG3OyoW+9k75KiruwW
gcMg5GftyvC1hCY6QPsRxMU+nhOIDMaMXIIBoGAEIYI5t8REZWjQVkya/35zy3T9L17a4ZaPHO+4
BeNmf0nNXBexcVZ9KgUFeTJYO82N8RZu/gBA9psh9Q2nSW/Ma5M6F7daFt61WqkLAucaU9/G9NAi
JjOhs0lefuJoHXwM+AgrrL+CeeW556BdYfuVTwJd1czHeGf6NGKYJ2rs7LFjj+fnF72JJRkSCITK
VsSGyluxdNolQG4pLQJYlMI2EWKHH35rU5O4MIzD/z7jkeEvEGm3KSK1DlQc1NJIcVBfY+Z3Gq6s
9kVp5aQz5XAJ5irK8+tvvF0TG+q+jy2oJH0ZgVpJzRzCVJ0/+QI/Q7fgbiRbZCQcl5FQYEsKUbmq
ky26ClqkwvpgdEDRwr7yeCUYDHFqj+KoeOVGgqlm6D97LWXR0DU29mk+M7yLDaBddc6oithbCzZb
mzR1xHsyt6pcixndco6lJ2QA605tj+z6EncOizudlzR19dJ8MdTE9cxefgS2lxEsw+tOe0Tqa1R5
UvIWFZn5bCvCarMIHeoTF4RyibJ380UKrQDsq8IhdnKQUayWKwG89/HPBcciL9CdJv9MvXIQGx/c
eudtNBASQMZ0E4v7u7jnSib4pA9vomWZ+SbR+mOUtWcvS3qTSMrv+2Y7MG9vsy4vPdEg/lPyahMd
0ymHyfLStCaKXh39mhkeev6GHP6r48ddP0e8k+aiozf/6S+3rdJjk/nspjW76yq3guV4un7xydik
oxp9cWfRa9D1DMRBTB2kVmTVMymEbJEdUymRobRXpqZscM1XCcFk3hhiDjoXyGNpJRbj98zZ6LF0
ZCgPlReFHTaNDFuWVOdmhFivJbmqIfivCrJVnwwBAng3jXrK1QBE4kIxvsvzo1p99SIES9iKTH9a
mCCxwmsI9Wt9aGMxbt/D9rZnKYV4wURaDSCZhBSZLkCjjmOdHeSW5Yx8Ldf7M1gWsZoD1foSceac
diPVsEATdU2ZoZJDupNqtJEyuLbMMPkVkh57jc4R84IFp8YrvYkDbZpBQl0U3zC8NgYW/Lb60ZFR
UlhQgCFRkTUfypMSmPyY/zCNM8ksQht7sg+fF7SMsP+4UdNVbJRfkeLV+dz0xrIzkRWRaXMlqdco
AhIiCdZeozWkcOBcp+j0rNZ09/0U9xfoSD5/6ZcJH38ExWhMsP26+Z2zSD56kXSW7mZUX0E7SRrh
aPU0EimP1ZmuvwWPNilqim2tnSojQaRhwOxS6fVnALXReMt7m92DhTBamrC7sb8M4kqeiHIqlRsD
b79GH5IXzS3sWpTIb8UzjkNQWBgldDzJ7qREztcTAp5pQL8sf1wV6WTgLjdvLrG0Fpwk3rmK/Qd3
FJws8h8CmNEKJDLcg+43djadr+tsq03zhKp0ZjV6wSNVAWrlmMbumPqK6Kj/DTBNAAcpM7MH+JUC
6Eb3cpV+DLRdiLlizfbXLcEYuA1RuufhurTEyWqEGVqxskdwkChBN3j2PHSNUHc/q5htg2zXl+hi
p0E+cA4OkdM3cQcBvVgooRYLbM0BRTm6+bBIEx62b616L83VS0aXD2eakL0W4AQTy8+Qx7COySpB
2pCx9Y9zYqqh0cIPkUDvACj7Lha8tjTjGbaOXxq5c0JSPOAQnrBN4IxypP3/ap09+bZQrGvnYnhD
YjCYMF9thlf60daVlhnueMk5CQJudHC/nG+apSyKZiRhgxDy3vfD9gLCins0pM4WtjjzB3K60NnX
m55+aKgB6m/1K2oTcr3ZA7CB+ARaySFIdlkIISLFqK7DYHn2Yev5hi9rYttDLEgvBOKc4xxKb4wu
dME5bwWvMxb7oS2GXmNiZg3Uq2CkN9x+N1HlxqnmrTJOzTE6o4t4gdLkJpigDh0wdZteXqxAWQL/
nP9LzSxAMnnNNhtuPo7sWmWYYIO3BW4xeDJbaySZjRXVomXoscHUDcR5nIvjfZvmKmbUJGAHn561
RG21HrfwWcdyytP3KgvMS+Fmi1MeyTPO+Q0en/Smnggn0aMUH//lt94/7G7+fIfJEg/io++pYZzm
exqU4mB1WsH4aEGZnyMgd6rcLL7M2IFcvnE2cCENP6neI7mx6Qb+w41MhSYocEkZ5dTMKtpUUsi+
EqU9S67tYMHoMCrg2sFs0Eq4olT7Sy3G9m/dh1sIjxDpm8c9F561wr54g0jPcbU7vRNqVvuYex+N
hW/+zpi3yXgQDLZtD6uGg4auQsvZnMtcGqGIhyGGLdjkY9c7NwdZLuVRgWTzth/Kdurd5ehR6p/b
YRUS72pfRab2vDTqjYupCJ8eeDiJsdIowOHvpFr5XJjcKvSapuKVBijqnUyA/XP3MSNZ9qhtywT2
Qm9TlqjfGy40AKvfUTLsHATDwf9eqI3otDcU/fDWyGjs7gQSYxOMQp0eeklPlnCGJolfN8/eufme
KBV7V5Lu8En6+JgJxaGoJ4VrpXYL9O5YUlmsFIoasL/rrQ5VUosOHo/+NNFbHtSK2dBsqUXEvq95
jIEc7cpIsAPWZ8irUv3jdII1tuaWB7pN2IlnPYTp1V89tGSdM6c4k/8XSvHe1hq6EoxQSO4npvn5
4du4jzfGutLjr+hyDm2N8PSW3UaKFSChJc84dAlZzCkYHH6E9OGloVRtu/ZzxSX9kRy+QP9sJ3Td
3KdPaeoLnTr6wMS+5RKZbFf0hn1stAPDBHIR4WKP/R3nIgcwFWlSGARTwKZKlgDfu2M+iz4zvo73
NsMe9gWRQPDBDbuxO/jlkDhVcuHVXf6OyaEnRF18nSPO9OKMtzhY84syEolYL3LGrSMaZHOtM5q3
jmUHv0F9PdHdB7weyDQIJ1F/+KniQ43hQDh9rebrQW5KZsq8LYme8IJYLhAET+HEFQ14dE+b9VwO
obN8OEIHC7XurTUSNQ8j0EX/LMWvL6efEflI2OVyjrpwmuz2Nm9Wl+a3c98qws2aVhj35S3+fws4
LW2ZEdwsEdduci/rB1FTL43cGRZ7vQCmrzYsESVYLfVERx2eFWBGPfB2TP0fReamN0X57WDBdFB3
GUqDW4Az90LejApHt10ki/HORrsJKUtC2YyYOUK7IrNSU7aJBvpW6VF1juOjW1FQhIzZVCNVLT/A
8rLCgXkItVS6Pw1RQFzdOy7U++Mab9ZuAi/5Kf2UvvcYI+Fl6mE5cnq6wHWKSz4Q1KMEKodj6eFM
sD/WN3sAU6wpVgzG5XY7nPbch6mbsj7LK3goOJz5Aq7xCLu2a1t4AqsWM8ze/OlgM75zc4WF4rNy
EXJrAg6Dx1yW7qO7+xil8/1KDXrQUcvU6vAXhgYO00aNF6t8k+MY4i+LvUbajii6s9dcx91UrLQt
CCYt8gc2DvJTGcb0ier7EESd1X0eur1BSP+FX2OALqfObi/rweQOqHROBUQWFH6hfIFUgvF8bXqI
ndn6qzi02Y4L1ID8Op0LTqJrC5hwv1ev+Q8YhvrJgb+/erU5c/q7A8dC2wXkt0ees5j7cG6nopvE
NsH6ma960U0etc4CVQ8bnRKVVcyZfLMw4UP3z2IHwXdkFMd+Hx05UNLw/uB3Wuh91iKOBNfFwt6q
9S0AYVFZwEAQ/LIbiC7KJ8/2FbomfsvkWdOgWFR/MQLNXBtbeIBhd7U+dyzjEB8Yd18CCYO0grSf
I/fkMGQOkiCYmEANytwqiahC3bs/PIvJ+m4ADmPv5pLl9/8dBchQEeWvvYr+eXLOp4RgvBHqhi89
5I5tJ91Ht/fPqrviw5ENJlBybmXfvQx/+AIETSLyJ0zF58jkwsbcKwd7plfNzBcwsYx8sxb/HMEf
fDUY1M/NA/l3tMbIvpqskInknfLTwNjuAZA97po9gkVsjjvodeyO2dtME04oqG2JfNjWvzXPfFNV
gm0TpsV8tbQor09U3Y480VkSjtCuYoS2zrB1xRszDtFoEXBL4l7/cSgjNlGDTrHycFgyeFtwiHOO
GDlbGeP7oJ3tSSLgIDz3QGlE4HOKYe63khXZ2vLugZFLpTun37qlz6xWq025PZq6fTCfR+Ztk4KS
Ghl9qQhvsXvug+N2o+GhKz4ILlf2+qxZN3zQgG23TyY9FLPN/tuq/k2wULGOtttr/5VLiW8KaagX
uowlD+4DJk1hL5ViS2cXd7XCD8VlVmvfvu2KTUPspI0SgZVTtFWrH1It4klnsTGoe5d7qNdR4hlh
KmuEZy5S/MdZviTDX3/hsI9Ypu/sgoN4vSby8QsFqzfxyHc+6TezVavIcaYMjFIFKijA1kgRHgdq
1VX6gQ6D4gDi56SqP6WZkGvYOFhu69qmKNnlYBIb618O5Cp6IsPMEn6xu17aEnz6Zs0Nlx6kHOym
/Tpc2tZgSdZUUewiLkU1xot6kYhBPBbRMuIrVwcmXjPYRm3v9vZXWdyKfbG7jQVHpb6kZKn4EIT+
UAI/uchB4TmjOrecY2RVeomU1hUDVNoY2naIt2L2bfdapGdVuk7lNvptoLLfu27EkAXj9P3NWnPi
NZZuSe5gSBreZfYizQ/Z40mrvi1Q5uI04/KVLW/zlQ91SghaqkRaWimkMxxshUXhF+TFG+DGQrA0
O/QFwBfPJ/wlS8+lbsDTlnF6Y9twv4nPwCcw7xExFHW8z7aTq/OfmQj/Z6NHXpahD6Jo8LFYYLVN
59B3v8FH7XoxCNyaxpZeXlo+amZlTkSBivlBR3oD666hm4VsHzg09Mgw2gOhjSXXf/k6xg0fsWQu
4hekbpf1tJ1fkhGIatAwmVmYRMw8opQzrCIKHaVvbYU922OiapZXKq7uriSlMRVFBPUO8X3/X7Am
dODK9DGTY3LSwFpjbgKvD4y1pulATxlkczJUPXC99glcjpuxu7oGE/2NhvjhLH/46OaBB7vOIOBz
Cv/8PpKbTfaxQisnI6FNV8xxDw4oS0nPIDCKCZm8FOIdONMPYez5+tVxnmMP4/lSwxvp3OiljoOn
jEOTlHGF1y4xa+h/p4KjAX5bzCq0XXAluELAL1xeRXItIoy4fNE+RDEq0e5liKWFQ3vC6lelGrzZ
bP4FTE8UoE91EwCZ5PjwtQqejQdgbfnbY3qFjcL6Ond2Tg+98zqdIKFut9WRLEgClWZ2VxaiNYh2
WAssYJAZUJwbF3N8qjFGAxqrpwXUmzjw9ub0NjknP0S6kWTxWDAPHt894hRnBAtbEMPMEPRHWch9
Nj++f7XjGlfsxWH3uOKkcpGY8s7741a6VaezwEW7Z8v6lv5ZnbZKzFM4UOutSIREmPRsXOtb5Euz
rLcYQBBlfXNdnu0pOshdpnZP2WltHuOSOKR6KIop9d/it1WdF2FIeeiNUTdIxNR1CPgO1ed1cmSx
WCFamDcRKorCTJigI0wZtOSO6lx4gbO3hp8NmKG1iog27e3uaw0Lu65dyvRpeyfpPOJHZ6Y7vaBl
yRPidZMNr4sJ7pVmIwaeKyeBp4psmFo4Ssv8Wm6pbu7DjnBn5G3phKrdUHcupY49i9jnAWfMVIsq
EtPObMfnkqHSB5AWEgQJsmXI4yf1KuJxSwYtFEuybI5fcmiMgFbyq+6iCOsX4wSx8lh2oBOuICG0
tHVo1+5BBlBw6FZ7z8VxzARsZ4jR8r/G0T5seGx5PiSgAInwbc93MJfn0siS5pR95ljKAe59slCq
OePM4CvCY738yJePxHb5BKA4LqPUYlWfRC/gWNxwEAUziSqwqcHHS9DMXRWTGF6+xiKamt0yANgB
amywC2iJ52wdI3uZqCe+qu7awYPavFZP3kOMGVpzWapj24B/BXtiGhOI4yKa/K0SOkb2Xhjbtf6w
u+Mtcs2vxBXaA1/HQKh2bE7AX+Y5TyrijQr5g1SD5W8Swrr1nr8/SMt08waN3MBTqeuJgQ1ulMD/
G35KJJoq6CmeUvDwGYfPXs8FwI+84BeDwMRW6rdvK/C8infrNFQlpoWoZFthj5aFx7aKEFV8i4tT
CY1gvcvYUKP6DJqduzeArq/sQ/cnPp8BdD+M96JhZBboY1QRvI4Z6OR5bCEMUNF/jVJCZaEtRm+n
YNhJqxiXUv9rK9Pr75/PksF6Andqt+pyJw+BKUt0Hok+svw9AywB8rCo78oxwgORnUah7dYuEOGj
sY+qOmMJESaPyrKplG85BNNmGgoenAbZkROO4QwbdKoUQbDBAZUphf83qZ9iDk73rTV6ZbEwvNJm
I61nmhR+mxopwi/8gWXlecyRbY3/U+OTg38jvpE2VnUNOMY+WAvqCZOxThFGaIolZMvHJ9LRLBki
PNu11sRY9/VUT2dXKUjgVOhzAv2g490Il6oaFZVthuqCpfplv4CjXGSmsG2wT17ulmkc7m/rcmrg
A+zo7tCZC0UUz3tDDv6DgFfInl6BrFdValiNBd4fAnG6Rx3gPvyBOqnknrFBWDkTAh8TwHHGOFgG
R5k7mCpHRkzb//N0zZ6TfDSRmy1HOl3kULtdxceci5hsZndsPtN48f25XwG9dhPObYPHZVwPwiw1
t2kTqTiIHJ1J4fkNJ/AwpPcQzVCtD8IP6OFqw1sLmLqejpBdFu1PE4ScgG0xX+Oacfq7rwoX5L08
Yu0Af2LZ8nzvEt3s3TVNA1o2vcYElabZaqKQMK6hHI1n/gvX4B8OrkxjxeZQsjlU2yzY6JlYf6gE
lkLfICLTgjBtArkPH3NtB9pyRR2RqYS9kNnmxM9OscqEBJ0q7mQU6WhhqwQ9vmQ7l2XUkmUTgEwj
vl8c+HCNWbMOjmjKyN5gp79xTC/qvLwXgVIxfItDYSQkc18Zm8lS3vsZm40cx8/Gb94ZdSoZmylV
TkWoi22HiEr5KwmiCklZwADFWrPs0zDYm+7udpz2CjUE0np+tcLF04jMgf0COu78WXXHY5CGmAU0
dtbU9RheA9sGeGSnLUOxXRCS45/6VJS04Es/ztUwTbyCmUXygFyMyRsme8oIjseY0gXbxTAHZZu3
XvRt7C0ZcHE2VXbcTTW4SYgY+nsI3HqrhKew0NQfai1kRG1sRBhLCRBQ0gR+dOary4UQMcs5ymt7
I9qqY6spbv0aRqf1gF17x/oYiwn41hysoZtVryxv0JzzM1y4tyARmwLLptrJ4srVSfSyr2s6jm8g
pgmq7BxE87YTib28Jnd1k1TjSX+YGXlVb+SLSaB6ux3PwPS9gJCc0yGnFeEPmFKwhc+20DdmOCaU
levPkgbcsagoUYxesIFf0FCQbviESBvBJewxuXKYLhkqUC9ZZjEE86KHfU7G/vyt82Um7pRXKn8k
XsiLRYbCOWtsMoWdx9rKvjNfaBsFMG3+l3uaGwuYTxC3spHxFdkdbqPYVTSGMMD2RHIiu+OnKzC0
sdcBbPOOeq7y/rv2YgvBjBucZN8Rgj17aw6gRdHX5EQWFfKazWy8xUushBZKFW0ENKOiTz8XgDN0
xPxmORsnH0bJMk6YLjcZYJ3jaMehsODl5bajNg57SpTUKg4Byl0pQq5K8CPbLO20JOoBWX6VJCWk
44GgXhHcMX7BZqbCosVmLw2JdDNEPBTSxlQilEGfyJMww7qYBldPbNxSiR3NYazTonvRmDARoMN2
6Te/7dO/mfFSX7Bhn6cRAFDEeq0bgN0u7FdyHle2CYJoZg6D1iaUg/TQA3+pKDfvul2r0BdeLhnZ
li0o8DpHLgpOC/gk3RQfzsxbOfBuZXUbXNIzvtSctXLsOzANdGD5nMTSC9m5EWIR9MZFKGQNQ+70
jARccnL5Q/Vz42ZFCE33uHrUJ9/uQwDhSlE2fPioPFyQ09gyY5ffIbmg+xkf4OtwJCl4IbW+TbOn
MwRpkRmW0nBiAYzE4ejMHViogzKck0iRMcO3TgjUQYz2tibOljsQPXIwLXEAko1Og2zchealtY1e
/JtsDj8nptB3Rc/IW9QfYQkFnbVhKx4/qtMcL+DTh/TqHHYwzec6uhDIsWu40JjYy+AgaXVYhTab
aE2C2CluaRp5fj8y2sop8RgTTk/H5+quffrmzm5u5FtgyrRd9Ph31ohec4PuI7uDhuE2qluaooxT
JUCMBEwJTiKobRZCJbFu31XlP9XC0OGIIcIS6qvWCzE20zfj8T8kjL9byYboU1NzK8n0FAER8iVp
qr1iHJv74OR5McglB7j29FQoGt6wDFiZU+j6AA2IFr4UkGKd5VUBCfbDhuNwgDO5VCv9qU+nS6Kk
teoaasdRfMa8e7e3V1GtLVgyB76SYN60/9cf4MDl+2ZRkjwLkdTET9HM2d6iL9499Veix50MTGMH
liEKjRHC3bkDQy1EMIYLV1Ex2Kk807xl2edb755EKpynbG0vLG3QMu4Tjfv/ruoEU2ounRhENNPa
+uGob4l7az5AVa2W3aBm3m/1MGqQTCiKJ7/OOc/KqdjGfFCF9Yj6Zq32RrOOoQpzxwlTFgAMJts1
goXKKnFKW1d6ftUnOKaTA5LQAvabPW0NOgEn/R3YN6G1rkxNDq5YrhSZc505ioa5/bNy+7SInm2j
92pamhUbkKzNonmklB7zRn0SEIL/Rl2JpfT9NoeSWfLODO4Cx07GGf947kCBQPfoNmyNDZVAiZ8l
euQ4wAjQLBXG1WP8JeeiDn/xg0CLVf2aftY4ttXuO2Waz20qQXNigZUrZOBqfaqNs72FxrExQAHB
iizjc4FymC+e/1SEO0kr1g8IztpPOyFBF70/Dco4dCzTCMVcgNqliHUDSz7OJibEy94h+MBTRGLa
8geOtVjYC783nxBIOPpQXzRj9QyYlyaR3hhITzeowNKofsDDlv5EzNb8tfkojjhqeKk78Fugxgrr
4zGAQtQdQq366ZXUszY6wwac2ccZDR9Qe63Xg65tMH3bzpVo6JDlwnHkyA75VhwlUVl6eH1e8p/7
O2QROct+99itogrDwMgzW8XaJzI7g2/Yp2l+n9z0+4JrgsTMy7flTdqdpRWlsokTX2rl2WKz8LRs
6wtEZ32syXFT/hxEXOZIAe+6pylXRKDot3Rgdk3HfJCNt0WaGsPcg2v7IEBJUbbVE+ZuAzJNe1fC
Fggd+bUZAPwadI1vxeu8ueeg6MFldC1Q8r20j3iQHMsrwU6rhXi8ObF0QCd1jy9WpQhOgspjIYiY
PA/nUPz0mBnBdnQmbvxCw9E0VapFwOlY6CHitrSd0kpvgrJ041bPTTOvyh8Uy98Gt0a33GmBkXkH
2yc58dq51eKZ1QihzxUMzlX4jOaLqNvA5zC3Y3LnreVXXu/R/oCHpej6wzlTiWiTbip1C06qvsQ6
fakllPSO8B/D6iGjYBM0iaThf01CMgniN/JBQz7dQBBzujMr7Yt79q+wmiMiviCczoadDacKFEzm
kfInXQG7j2GXQs/9kLl+XyZkbaJC5P3l5balIlXQdvBwDaAdg1DAjeaqM7+0KGUqmq6oQQJsITso
OPC9gVxbNW7g95NZTq1E7juVQ2NF4bCQgk+BQZVqU/9OIq26yAdzSqagHMcfgbO1U2uNGsovg7EJ
olrgoATQgU85IvAFzciQAG+qzO9IOztitfNikViSa9EqrZEXY1rqcIvkA/xQ0yem9GG/U8ST5t78
yT7Fyaab0BlVl3eNA2BFl6r0Vow4KfXA2ImoO8Oh4yVrvH4a0La83WvG2owtNRTqLAMPJs2VusZH
O759EgN9yUyjmKMJCr2zdwMPvsXraZtU766T7e6Fke5e0oi0iMtHPnaxVSk/YRX+8kKq0816aGRa
WZCRM/cDiR8r2RoBn3Aam/Ddz9GAb+/Y/4cjnuT4E07iBZL4ROduvaA15dNMv0z4zmpEHHbE84Hz
H3tlqpY7zkoIGdQc7O+TxlVES1NNUIlFYlc6Gd5xhx4Ec/mekbEkuAjQ7rBUIIGNprDqk34KdPzc
tS29s+/Wakdwtk6E9cToxTV5D08r7uGDDZu6imtLdHIMb3EBi8SPYYx8yc8Gm0lYXMKToTwoDIcL
QhxiD5Y7/Ofb/GJ4AzvaugH+HBoXLJ1VT82DqSiLUp7gCu8WVG7oFQ07SAgTE1zNIMrUAOeq2z/z
xKHS71rgFZnjjBoL0b0LjkrS78RV3Tm9mD257nDQdVkn2MtEmOp3rXYhlRhonz4zFkcZzh3ZBCel
419CAEiJP+Nn1bgfW/ZsBtj5jjl9Li1ItYhehUjg7yTfFrXAc7/bPke2S5suhnteQr/m7WjcTvpT
f/4Qy9itRToHK86vyGxcThSL2xEKL4IwcvS18h2VuvdD13r92UwDY9yOzTTD/2oe/2wr3CUvY0nb
ABNhsT/N/Iriij8fS3xA3pQj/SMBT+KHJfX4QhK9AnPex9HN+bHz0xoNjAOcDdrn+SgJCGLXUWMv
Eia703/FLbk8VpzZdgmwlrxAVHUJY2Pr7xfQcrg2Y1OlKtIB38LHHZWx50uMCv8ED4qRsmQO9PbI
aPs27tv/HyeukwocfwOp/ZlpCpz40iNEBepNu7Im5QEb9JRwEx9Fc2S1h6kKKWd8P59yJpUB483T
pZ3omb799//gfsgdtoVEHRSjnFDLiNwOTfJwFLylUBn1S8dKMuDz/+QRKHFDGT0ENUX587n4TcVb
uSWEu8qsvk83ZiGFJx0oCEeMhdK9Hp21/53J91E7IRc8WOBSGiJpV+/s7n1vOtz6sqA54GP5ZWfu
cAVAXrc0YmNnbOikTW70wozxaMIsYQxgd12pc2rRJERuOy60kbv2ptIrhWM3xYF5xyAM6Rxhn8T/
4edwD4JIQMb7rGXmlf8mw/RBsVZQTR85uK1rCoW7YtVkDgUiNsCL5wcjoF4DpN5fm+NajYz0Cloa
M1jhffHiTPy0x35Ilh587/gJqsMzpavuwNkDs/BKFD8l2JwOkTwhteGFSWxVEXfGSc1YHXnbOyaA
dPqMyvfkI+Y9sJTGthnCxIdnispcKnOPUetEQI9GdmiInl1pyfgSLKcV56ODKVFn+OCgcJkbTKZ3
2OUNaFQQWUlGXZwTmAOjBpZ/qLnqSH5zs08vktSe6xlzH5nWkAPmvEFXkBbpbxslTH5vr6RFzToN
d8HkdBMoWrx4VfCjs63CnmXpo6LPA/hA8ytI1oz+nelfCSY8lJ8Dj1tCplCS+wsDW9uQjMuU2kqz
mLxieJRBnkBNNkSB8GyMESgPUM/z1MASrHe4QAU59YyUYKu12ipKvAKx2IG9tO41sYMMsisldZES
hUyZrIPEMojeo17tx2jd90vrLwR8GlTJU4qW01T0DcMopM+grC8DOheb9TXOkoaj2Smo6+n86z6L
OGvf+uxG7BSpEIqja59azwAFmBVsbpZZ8MqX/97zZ/PuCn/wH5Y4mverFvTIDW+nU0qH1S/waNXL
2AAezjLaTkTqfwFQ/ludR8+NUWbXaJnK0bGDqC5/halL/jhI8c4/Uq77AQiM4yK1PRSOAqE0fyPD
V4g+ag43iEH8wCheEmkNGSeBlXJfW/6DlnKZdm+p+xAjQmo+E2u0P+LhogGchLKiMOibdpwJzknW
DsD11L448fLwd4FMq/Gh/WXKHueBIrVBQpkGkq2SLQkO/0n/1ZaHlHMnKu8hf2GKYWqBMrGtja95
nGcuWrg90vbAJkctqB7336uYghPcVX71KyjQOVCdXarCOfL77LusLI0q/6xBKM94YWEXg71d/Iza
WLxtzjOjGAnD2FviG3rkf0LP5O7qk5IAvcX5qqBolEUmp4m2KBOGn/C86joX1aEMQ09Z8uQCrLZL
f18ReoDMVi71AeGouCqUvpCfNueZWp7hrBXpPRTaAmodB6gSKuCAiqcPgqiInZHxBHyxMiuxbnnu
tCKgkYb3X+IzIrg5mayvZxWjIgu9HhvEd98VRJIfl7o2Js1TvCeyaUus81TvUYsfk9CsTuV0iFFD
uVX3a89JWG5AwryXQ1EbPNwK0LVdo1A0OXi1x6gtZPIVseh1uJsbuLvRug1zGNwfvRWxvj+10pxB
n23LusWNRpOjnaZwEKByxa9lh6HjPe0BvYW3AtLgAoio0yQPkyAKGVIojk3n0AmfznkLj63T8WCb
UkNa2i9+5+ovLlVCXgeVTy9yM1XgjBGmuNAEqawuAtdeWz6+ThgUC+63AOG7TeCx8Y8fBRrvho2K
scRSVOKc2tScFrUNHULKMmR1D+8Bt0BgcrBVBalPka+9L9nBLUknmx+HR+PtoxAtLq1s5a33xx2m
sHL6QpiCA00XmP4k1hYmCHq6Pd34CMBYRf6gHDnzNxFyBjvbs42PRbM8mXKOFLCN6s0tGJtWyWpF
Ibe/kcNYrZu61mGp+eR8uOld3pEmWuqidMgVtycZvOTdFLFb9B2gKHnGhWcEiA40y6bawStii2N/
hoCZ9y4/zoq3mkLzNIWxsOaj2S/9wlg86W/s7DzY3R3KlCtjgwu1zd6Phk3EZFSCt1zJ1oZnnaXO
2JxLJ/MdMqYR5SxqCkg5AFZwFRB2hb2doiIHZ6y3UGqAFCCv7mOewBEFfL5iNfyDM79Re0KWWIW/
Rcw7ERMxG/R3ZppMpHXbsdEpI1yA1Llw4c0LPPzhHnhrEpHT44bhvrkqM7l1HOvyB0rg6RnF37Yq
AxFDuSInmX9O7BnPY769AsJpizDudLACFeZb0nuwS0aMsgxwOkQbxZDPz1QL+3463ZSglGpyBfN5
XnfX1V4tLnEyDpiFq0UImCz8f46wu3yDcLZvAI5U0pEixNDk9myiSO5mnXjE1M+mLnD5eyi4yY+a
oj+Ihe/7eNrK0Cyy7IytZtvTzZ4T1cJXiUpympIdjLof1WPogjj5HF/89AUucE2F92RhxD/YI5Nu
FIiACPpf+MMsL0CoFkF8VAP9nxBjnR5tDI+e2ibnVNYE/MYCEJ8Wv4yPu2/BYTD18C8yA7nliOSR
uPbESr6eAeIJBTWl8XVnw+xfo26b3jmpF7ogxfL3o0+I95HDYuZBvjpKVkuwdlHnMLJswTqtwidc
QQ8KlZdaPYTcV3myHJOxA+jWUHtau9ZRK5EPUBagg6ZY3etZQdliVl4i0U1rSsIxnp2RTeU7wRza
YEfj/lkjqhbK5xIokmQTmbX/agFbPxmdwG2yA3TcI8cBFnJtEBOGaglFnNDRLhOfMUv+s/JE/65L
GaFyUCvzZB9+QQYiBS8CNY5fcp/haHum91E4QFoxbHkBvan0bm/qNwvwd81S8cRG9E2BPw49ME8X
YyUIAgi7CQQ4WtowGmomfNKwbMnXVTsTumDagoN86UtvBXcxuRFV/x+ZROj5L02vxmz/wsMNQ+I5
Bnb3pzBKJ8HYKBlaqLGCF0glt34wDjt3io/15Z5wPfrCYyO5S8OK3GQCzh9n6ce1UVlFugxv0gHi
WU51L/WFEPWSOeoBggaWeNPmwkS6xYXag3Qur7XF/NpI9/gO0eDZRT0DGkUhOqPZNvrmaNoEeqgK
3S29YWewOhVaAQiBEl76asqTrAKGpIoGAK+9oLm1vLFeGBaa5hjbZGkJ/IYkHgM2H0+Zi5SSm2e7
kEITPkKSD+hnyPxfEPCeC09Di8cavWGNIBVO/LcW4LOr8+t/VdY9hI2MyQa9cPuPPc9hnoXft0ra
PiK+LBSCCUAg0TcSwncrscAEGv/fJKTMbkYrz7d7o85Yk2uumCDmjMiZ4sToypnf5b+c+rhMZg/C
hDETS/QLwk9fUVDF8POuKs+zW6F1+RhxsTDCOTLhsN0oeXoPsY1m2y+HJI6y2RCYBs5yyr6TXYDF
YMyE9Y4sq/JNn7CcuJ5XCrwFE8OABVYfANEEvsul633i1oZf4EDbOHUuoHM80DJgutpBft1senAF
ymHDWLiefzrZxg1Dum5euM4QYaGz2egiSs1fMsS7Q0+RvliVxQO892LMGXmlJNtOyPHljqx0UldB
nUAul4GOYD/hNNmCXUBvwbvypE6k0TJoTWMfEKPqcu03ftxKY/uf2CBCiBhcwVKsQtspFl+J5pRe
PceqcQTxFFpDOdcTM8oG42Py2tRpehZmHKXjmshqqxljdOrtIvWxprGwXYbRy//JLL6y/6INNeOQ
qxYv7gU6YFRGa2Qm8VJ1qLqHGoHrrVL84eUo8qOasXee4OPRBkysPI7fimxygql8fNXLYtlqQyYY
6L7LCEsCn4xGp9Z7tq4zqKLQzVPDhuUmbNm1xVc6TEJFZsGNZT3lY59elC2aIrff2OzH9wm2Y0Qu
eXPambY2Hk07FRfyV8c1vwCNDrlb2bEFptyXVWGidz9jw1qjoDktJoqGf3cv8MvJfITOTgCkf85n
Z/b9tqk9WY/tMsm1tl7hUXOMztwKK39IGQbvagMoE7gfEv0Frk+0x+NqOAMFgbWaxSkmRYhiLVkZ
Q9638WLtzG2klH6UWtd7Xi25jMpq0QtRbVf870MogHHNDxAHiWWhfjutqh0jhMydgNPNdAAysgo2
HPuobIaKfKlNMYnXc6kZETAcn8gvCf7Ih2YqOj/OtJEr4wiS1tmc/I65nxw4KIknz//JvTz5HZ6b
i7/w5sHvGKUCZpnqgeMh8o//B56NqxbEoIHPX1inf6K4uRXJTLBJPwlt9WHZgT0K1FMglfIzrFEZ
7Pgss9qIdJPGxR3KWxDveJCJ+U/YsC6MaxM6YZGt8VxuPGJropdyweKFFCn+V23ihmRJD6A9zwFY
poFKoTvXJCxySuvQgPm9zd2Z8yQgViUre/t/TC6jBbOglHDz0TdAlZRdj3DRMmnBxSyPrQqtumLG
sltnYQF/1a4+oW+AwqqeRZgq228bdiAR8VfnpXLm+a6jogGbEIFYdUa+agxVsFXoox3eOw1rsGg8
MsgCIGTfqSacgo4V8diT3G0OuNJKezEFqklLAEQ/IaLhg1lFCZuHIFeWpqGwKeK6HuwlVCZ/O1Ju
bGJhOHq8K9Z8baKAoOr8I9jTPicsd27aEYpZ5bv6p3pIZ+fCeU2nW9U5vA768dljJtcmaHK4X1Fo
mcEL6RArjTYdnSToL0yRVFFKM+EmiGuuIPw7TkOhSyZJbdAjEUIJeT1hH7OC4PWv8hJpXREQdYjc
6o5+fJdUy6jjrOtlbkVWRp435Xd9O633HM4daLjS7Ek9+xetrV38bCqCPt10VxA12K390bfkvRtA
BbeBYUVOn+ESDz8rckNlqV0XqCyZJYpFAD1p9OGF0cpXdk0UzCAVIWAEjefBXNX43fraWCsYFOEp
yRoK6HLS6nzPZaE7S3efcxRO/JQuAGcdhlpomjJsNAvOQFhCdMzMWbLzPxbuIbVG2ZHjaXj2fKPz
9JsPd9m3y7V39fhwp5B0s9OS5BweFl9K5eFN9Sbxd6TD6WyQsHENTUxNb70ym53QYkmt5o8LHVwD
OHsQS2ekCi7jGqeZcPvwA28g4ZozlYCvfsHvXMAVhl+QIVK+Ig+RAmZCDEc+vyQl+M7doq8HHZ2F
GlDGIuYnFqu9N/CRAs0m7MLPI04DFlxjl2jFFhuZu9uS913fsCjBmyzyu6ITOFq4WMGOGmYqTKG0
89NdFgYZf2u/rRLKfovDzm0su7M2iIF0s5mCMnujNq42CjWmPcOmZKF1HwX8Qpga6VQR4+vWx9R1
TX+WEGB/7BPFZQSWF1i/QlFXkhxtEFM3xm3ms4K1XgF3V8V1jwEcjMSDBhPiYiV/nCbqzjKzuyxn
Bf06CjVtZExQ0CpUzPuEB03OHirAv2iJFoKBelDBy+foPVrkyN1gWecNo3mic4gGrh09WxJ6PwFv
Uz1kQ+Cp8eRpqpRHBJAUz/pHu8vTC1vLk3JuPLEGJCwSfUKi3u8YxwJm1DwTPUZ3Q6o/3saO7i71
z6c31H7VvTBOvBFO0c+Nm1SDp/YMxtdQqs5wTBr/zwuyANEFmEV8Nx0Jh5svoxW0ulVb5Y6uOGKS
5RkvCwRVhxyqHxFX0OgWEAX/H5Zm2Is0tANr8tJZk0GMkhmWX90ZRX2fXsPyd0eesPHiWiMNGDUX
CfCrjSYyeKfLrkv4hq8GMXp0j6jX20pv9BAdBA/F3MVpVdJQSCIvBieRtJDIQO7r4Os7ZyujdAMs
KrENMkYvo8FQVgJTj+UQESAQGBCoFzDV8+0bSYKbOY7Hw/s3SdbYClDrDcC5ZGdyQRuC+zNmgoY/
9bR1gJNi5O5UOhLfqPuZ5R/MBPRpYxjDwtfO1/zBJ23196MD3Ch6j5sXLtnDpSTsQsky/k6atr05
Cwh3mkqLnV5HE67J9KcVUlKpeG19Tj/SLIMoMrX2gs75hprxCOMGpMn/WXEEgqirVsI7Az27V+ta
eMt+QuZednctes2tzZ5VHhPA9QY8DG0irIQE80N5rlCn4OOpoMgvJpkX2q4oqLM4n7Vpi6QNMUtU
04qgREoJkw5qiH9EdNPcwI7/p504H1U48AZ+tfwpi8NiNSc+XNrWA5ZpIIXqDO5GNUeh8M1uM+rl
w8M+kgPIZk+NrI3cDkIkSxNAOO9e5nXKRL0p+QW7Fb11TbD1R4sqosTyWhN/EIwnQQ40T8DHwgvy
D9UCeNISLe//g5m8qYrsQbl8hOh6aDlCU95TZOTGxPk/DZT+3XTjNEqOQgcmZmPVU5Z7INE7xuYB
nl5T8W+inCzG6eMw8KhCagPbE4ps/q9/Zw8QMzd7fZx4QF/S5vLKzga1q7NvsEFM2ipjBr8KdI08
ODHTsniOL4kriM6o61n+UMnBhcaazJGtYEO3bLCkS5xOsEBakLPMGoUok0l0d9sghejtu8FiziH7
65CPcl2QNx4xw2UblX+qdUWUQqXfd3Gh9THNidruSVWGEz+4FnUKz7gyrFvYgjAK7fK40dx5Deqo
UgabiO/Y+bXyhVZWw4c5fjvqNAlPfFjkZXE75egpfHdib+Htc0+7K6AYD2+S86qYqjhYnBSuVCvd
Y6i2JchNlXKtpQ3bBdaED+kZh5SG9RYE7VgtlLSaefif8RcNIeLKDEXR9MpwGnT4tSqHYD6x9mMS
iqsz9k44jfhKvbnXmlmzgvlTwg/PisFw1HOKGaG4p7ijZ8TesDZPh0MAcXeSP5lTQMz/txPMm1SE
fuE1gIx8fmu1+R/nvRHeg+siEuE0KmYuB6dQcrpA1Y0xj65oI9oF9zvE7DQHHktZV9Ene7lCa/Zk
17RxoS3yxCbwhULjhbXDWrCvv0moXXCuzqNYdjL4RB98MQYcwkbIK33ZPnrQiMrGqwV9L7rk4eO0
nBwoE7CTqVXDUI6ZbFP1v3flBHdGWQ3jsvq4po3bnn4w+jZumdYRT/fgFe1Xk6fMbJ4OUOG834U1
7xJKGiOnkqzXTChG4ztP8v91AtWlcHT30cbEzPhh0brPbB8KpATFAHcziDo6EOVmZyYp0iHJby/4
xDNiTYtRor3y2p4DFeWqKnuSx9IAwXU/iHAotcjlS5vRAX/U1eGRKw0sqxj1bV9xduGFTlDee9Hs
EZP55PePyeSliyoWWI5LaXg9pyQnkg2SwtO3ktF0WP8HOhE3gtnU6c7Q/WdDYUaXTfTxxo7G/WOn
aBDqasaNSpxGACVaaiiN6LMJw8+GN9bSKXDTOQhGKuAoMBB5bI83biWUKS9qXGmwYYg0b1uwi7+V
zOgQ/fYy/6UfYSdvATeNebJC1e2T8gcWTRwntSenpcwFdbwEWF4mjgGBn3OterPkncGe+MgoBW3p
+FdMoxjKP+9O/80aLpyTK6WIWT0dbO/eJo/j12oGgL7GpCyV3qJhsHsqaoM+Y/OtAEQkZv58Wkmd
Q8YBVx8F0t7lprtOubr9zy70f2EzL4HjHS06NbTZJ7w5kMKicD61yJXeBmv1pmu4wByBB84uHCTE
lAMt6anFKPW5B6hBMOqDrX6cziRt+qkJsIB6VlCNkGYnn/KcFovjGpto+BUriL9HVbLeOCL/hGCC
Y7WM85q4iQV0LGL87kl7loO+6UFLQp7d5YMLbhpKeuuvgTeAxG5OtFVOLT8uOggkjqE8k+P75osH
83lGgnzA1eHvMW93T7a+WyBlOLht14VNy3hKXklFbgjsl2L3um/vqqvFQUGYkG7Cvy53G3XR3IQV
KaCY/ymBCSTmFWozIURTVaRYaIEeECTDdqD3yJaAMPNGB8GbKlg1cPbnyFNwjg525ypPuOkMDNiA
Ur6d712wL9HSs43MPBJvB5j3McTfWRfv6WS6rYwfYLCm9nSL67e6CEdsK/ruRga+hJ91UffnzhRT
9890pwoi0Ztl7T2npvjpMp63JQeIZYvFiSetjGg1WN651g+OBjaRC1Wg+87s5v+q4EobZTKjt29W
Kd2tzpavjTzr8tjAmeqRSrG6PBausFarfrTjvoClWvik6sx+Z53eoT2T1Fvpn5qc7RA4WBYYc9te
EkxwGt9eXdMIOwzy8sa66f1ns3SloIDTjZkT+XDLUr7VPMXFZV9ja8c3CMosJQYPBxS6q2dk/NV/
5RHKwDoli0ew9DrR/bzDWe3fvY6r3G6GQmhpexvla/LMQULfBOUB8AgSASg+BhXrOesAsB4GD5Uq
xbRt1aSmDNieN+vN4XgQEIVFj9Od4WIfhGYg2lYsnahfye0HY3jXP3V4zvPBfhSiiB5CLGFxvnn3
YP9+VJ1tk7Eh4Oui16Iz7oNbS6Ev24r9L1WFC1/HeGP3IyD08Wrm6xixZrzGpZYdWux1DWI+Nhtm
unu/ai+1tVtS5SplP3lnRN5fuKi7sD1VcFC+HGfE6VP/M7LzYDuEH3f2XeS6tU/PGORbgcojyNZ2
0a8J2DrNXQeNFXT2y11jWQyhfPedjaOXCxALJvxPVHi9Sp+bvZGbosgqsAN2uoASLKijsUZyko3X
Ng0g0tyZFoIiWsDp3oLbOkx8D4hMxVVAznU+6IjHMnfsufUVqppILDRBEET90bF0b+MJRAYPVsQK
AdgUQXPZ7AqDv5/9kF6UDVsbvFu874HmtM8Gv8mcErrYcx1Au0xXiq0sLwLbqaREv6cmQ8R7LGOc
w7TPCZg6BOL0/bnHkVZELrTE1wKVWij9FT8WtIIq0H18FLs1od8VyVVM2VzPKPUrXtqFNJbeVkug
MOh6HpmMfLXPHS2VUmMZgl02q/oZzcUmuNvQIdZZ4JeFb5HTQOvkMR1PYVbAi3tHuKvIMY7mUR9k
j0lc2GOTQc86iPeh0U5A8fVOYbuJfjMq8drACiq1G1Xz+RVqi9mHs1tYLV58lkXHOIW3yn3dtzrk
FFUCGWQBvXsAVOiOj8mjtxlE+vGRpIJxsn6bsADFjVJ2J4z7GKDtRz7MMrAq0PUstHxWYRIHduXn
B/2Nu9zHgirLKwIVgGpRCremB9Mvrvw+iP8uvPXulQTkULzBBBNZBs0RbUSOeUfVjppx+i7QcmJ8
nYEhwdkYcRPoLwKtlpKxsYn62/e02IHp3Q0uXh73MJ7gL56mqEe/21Q6WM58m4c9UJmryeKuRwBv
XznWTtPHyRu+sfOU1G33+05LgnxPkGkoLljBr4cbmHlhNJLT2j7vUHqOjTvdAlI2sZ6UwOcc8IkL
fbZdxfACxi9O7kDuUtz/WBh3u/CxT0Hz/DoZ6Shd2PH4G77yXrHTWZukq4ZeKI0lFPKPFpJgONht
0sCU9C2bAVH8FOmC84igq0Olv77F0pnJfJCr+9gYyx4ZXXfXBS9OlkpoSXXjAadJTOpvCI6zUi3N
B0RkVNOkIVuqiorTZNMQwEfgQjCKNoKeKWBk4UXX1ZyC9tH0ZrNzmYXQ0QtFRmWVdb5NAsuoxOJd
wjCneSXhjZAxDMcDZ51cid0/32TZ3LYri3S2LLV+okNA+ufZCfuB7vrwDS88iFPduerICWjpIYZ9
GZi8Lu45P0UDcNUa/oFZKdpWFlH5MfNMtxUJu9qSpJJXHh1X1q/EmMgRzsmQUnDmldvY/lG5AdRj
uHSsHnr+UuCFAmQf03XVeAVe0QZkgrsGgTHTwKlh2kRHVEI5IQSgZXFIttGie6FwQhZSMWCQTudK
xGRa8l9u2kuG5kl8sg0PF5MyipxctpWVpu2t+BdDP4DWxTTcv65NATSLLnzX6AEPJcGfVEWBx1do
L3AR3Aj6cgFL1+cuiIr7CNJBa52GkHzmo2HRznApIipUpltfG4OnduDs+RWG4HIWKrUc65upA5N0
cMZGsjRR5QX9z81PR456PTGdVILByIxmlQg4n6bRuZcd6BtN/Illt23ZKOzVljO0GdQwXDGz9J9k
kezzQVM0vxlbz3hTpMIX/YaEN8zQ1bTS1Nw48Bq9HYGoT9V0l5280NTro9KlZT+z1nlaeUlOA3e2
2J3QYgM/upD8AjUPL6k7gSWbIYoVL9nHFueDsyWvMYWpUkZ9febHuh5QfT3JqGl7ra8/jGzwi2CU
ALIal8UPQGuNUHV5YV3oyyJ8Sf4+6zeKCtcR/nh7wpA4/ARZ1eNvuj78qIuUBotXp8gtxW7LchoX
6lHidbbea1S5oO+wtPV9ru6y6MSkYkoCKekbgbxiXAGg2ZVWs/wSO0FB6H1gU8tq6cOrXLCfX54t
QtMkmJhS1NXXfRNZb+zLh+TM3IYqXyv24NJAVwN8Qeewt4BoZL+lv+qJht/JvdV4tmrrnY/Uqv4C
lstvHFg8eAG9oxFmeNME2b7MwTi6fubZYJVRLMpYef67KkcTkzdSaHBsnYpQRIRs6+4Kx+T4MSMD
OYJH6D5O4591WZ1/ZmHRQcmmgGUXWPBhIB/HOZq3/imVYLUP3p1UlZVr9OIZIryqLV1vrptbJo9M
KBTeH6xxRRWniyHICMxStpx7H39Nyzu/hxoUWTBQe6lJZfqQ/tUyFn+ZdoYNnqDNOhL7KJ7cMQGY
Ln7oTNEfpmoLiRvRCy+zKhCN+mj9+cooy/2GUGwfx7NV5DLrx20np6H+G1RZOesD774+EpgWFrTi
biOXnLWo30gIkofbO1WxKiuf+XLKkcN8LTg6xD5HmAfTok+GwXdX/1+AoeNVgSxIM7JFviNUFygi
ExR5bKuD4StMR/qZnK/OZS3xkZzLDCHAT9Z6v42vU7efsG6wLQSg+jkgpxKpGiQ3/P2342Ouk6XZ
VwZX0HY5FplipOBNcxO+8He03MxVoIRAqzqkNGmgQtMk1j63BdNsgD0ih+ZHTxZytMWKdyM4Uod/
t54zuJNPxmMlB1mxR/xNlQthheeBh3osldM0Aazut5Y5deRKz0b6PPHdFwVRe8dq24Vvi1TRyA46
N2D60yKgj6NSPAwjkcz/AGx71wDDxzxH+8I55ljpR0iWhDQncZZYOYvigd2oWhKWxKm2GJAHgBuh
tgAoXAqn4+MB+VML16XWYspcMxlHCmnpkGQyDUl+0AL4fuy0q5r5sYXoLKoe421CCRtZLlqUYQex
75MueNqlmqVWKb0XxCngLR4bYe9AklpEBeo52ANpHnLEgTAzeqCU1ZMghrS0z/wnsEVOD9s3jtL4
erFIH99zinaqp1b1z4kHF9CzEBQrytyw7MCGGmrZ0hr0hRywlv7Ti6PwnWDaC4ZwijHcZUDzxK+1
sltBKrM8L+VDlJL5oog2nPUSI4z9mgvONxZSlsVazM7yuwbIqG95Wh9JmRizJaaFhuS6gOPz+SCK
tO9ECNtHzkCutfVqKJioF77guS7SUD5GZVZ0dTe3b2IpVFqbsSvGNaghnd56CojPwVkpo56q/BdO
0fuS9J7yi45XaRuxBsflMw1W3fbwUqA84lmcyFPFT6Ly/+Kv0qoCGdPu2qbJYFkMYBXEFIY9gibe
IvXX+MZvwzLFZlk5gu8viE371/RN9qXdfzjfPicVrfndf0Vev9DB6pQ1kRMwZlNph4Fj+gmYKcjG
axE4LigV+CXH/OK7KuE5d2CvJoJwzRxhR3f7xUgs6yezcvEeFYQiXq60Qm1qf1fyW1HjsUBuJxKa
ZHvFg2iVOvQnVxuMSyDDWnG4cb02+og9TfC9155rKBSe1pwDwPF9+hTJ2QL+JjpZBaAEosI/szT2
pJfATIwLgUpqdtACLb4/NYf/OfBB/jjpoOKLAnNzk8zpXSfolBzk6zeMIJR8DdGuQRMcGkXT8xGa
ZK3Hod9bI7i2SCowTi+mEmFS66VqFc31HiJfE6qW9IRFNS/YdQWwc3oUV9mu5ZQ50GHfHgruMBbx
4lU65vcz0mOyQmSIauBP6x8m6U7pN7IPXv9+C6I4vcg7NLZjXMoCnArgAt8TmuuKc/0UeWns0ZzU
ybg2FF5j20FVcPNQrrCFQdRfUupoQoYIKskS9+5TiVr4+Erm6FcujrXAsD62ol3RNcCFvx8j5DWP
cEqz7m31HtHSXAgm5DHjmQW927g9bWQ1FFqcuilA4bgVpuR9CYSv+Ccumu+RLoQcjglf0ekg1yT2
OU07Q2EoCgQ3VBybb3UR9HliTGX8uVH79DLDTSO9co4LJbTml5TWwhuNwTza5l63QeFJ0v12mVD1
7zj9mJyCdfk6F/ghIRNWuU7qTvGqH8fgszFN0KrekNUpTrfusLRiSaZywjQjvoJRi11/ImpGR9E2
Ofo6XfnkDAVrAjP4KqJSKNGI2YNBijOZ7BkiFDWjzQpNY2SsxO4kza5yY7XLuuu4UOvwr4U8VDnC
oYzdh65hsJWvK8RZpY3FbPRihxAVBp/uuVQDp2VM25uXpWlsOs8wjCXDZi20ZS9EiKw1x738xEKc
XSP3ygSBRzmkXKKlzjcNxwik/NMt5WLEdUtvfO1DuhOoPZIxTGl3hTuM5NDyti9oZOE1cXQWSPVV
+16YF7b7h0Tc1xPNycZT5rzM8O8Za2HA/+A40dCZ0j2FVMArNxA00q2qV+3akr2ZwCA3ORQ1ZyZn
kL808Si4Ls/2MqeSB45ceWdLjNvbd0nHa8h7xGrb8tfLUq/vLiYbONpllF11geeH+I/aU4rWBO3C
4zAKIBXcHOQLbY2me59MJh3o9dKBDa1RjxdFqvCvnX6Dh9BGpIxXn5OaAQby+TYYF3zjLBBVeUYp
rDLk8uQJANhELjZ2o5bVQj/ycM/4mFDb0ddVEGTSrWOwqt5UCwvE3UOvjRbPfIUItRCrQcSLFldu
XOE8aeT2Prt8QUGt3qJbfdUD+XOhXhv0gHRt/kYedKr2c5Gh/eb3J9lsU8nra79fA2VhwcDfiQHB
KITXARrWKRUG6051u+g+lC5pTN1DR7UiQCVFyT82H1eE5D8xYEFjeCF5ZnhrK7EMF7tSAdBTyKpb
C1BGFkbwrjcPXku7GqwL2IKBh+fkYWt4MJK/pk/WJ4qdCFSs7JfnWVX97FigMOhbA9Kgp7nNYJ99
Y1a05ch3np4uCst5q7cUm4w79PZsS+uo/OP22RdvEc+tT7Y5n59gjXPSCkdgaQhkYnb/of188m4S
fKD3AEYb9eALj3CJfD2IzKSDIXjUqf+N0ZorJSWPyjbqobajXs/r0+vwW9bsyYi8q5Q46DODX3lc
FpSRcI0oxdaxHG2xGOuwQySfvCuY1PEAq379wjdIAziL9xKl+G68IEvuxON24ufxFmQqoGsJZK1Y
gZ+ducr2TEaG3cg26wTYfU+BvR/E7B542bdPREZtwcNnw07Z54hW9vqktkXC0HPq4aj2630hGir6
0khl4mXkeatkMk3n1QB5kac9/NBsLLpZ1tL14F40Ya3EDlNvOe86YtSm+7iPK1AqOCH7UR7v8Xmu
qNDAwOf/IOyjRCY8kjMBJdXAmofieLIfc5iHVduHTyK+lsnb8yTyJ7XJ0QGtXQJHgBVG5Wq3JXF5
BQMfjiUebkpJpbne1yDsuQM2h520oAbUWDcQrOx8gNK7NMjXiLDKTRNohIpE2BxNuyW44Dfvo3MP
VPfNsPM7PaYFxW3ipBMBHfx5yIYDQFdrrtURP3k4E2ti2iimhD2Ibhy/B5i7sZAmQV4T8ZUQxiJ1
bF+6kGVLqVwitU4f2OLYKdqmVUNj9gENzcYpahQAePsCZidfBowv3l4acCrxlnaNv8eKugS2YGsc
gbA5xnhxxYCcldL7hiLrnVOxVus6gzIZ9T50kRKHtfZAgXE1zOx2e0QJpcfpPlA1VL/DGYuGCyoX
NsoDdewWa9wt5DRD5jTCwgC5xAFd6KObXnrEouDqVPj4jeTfzMC/Dug0yfuffW6mIrBfKOTHwj9Z
tJzyWwCYUiz8xB/YYz2s9FS1VCsZNFMjQfDJbtKcnOcNFGCMdn578OTcBAIhgMyTnFPtqwqzODDx
f5xFms+Bst656yX/qmRxNatkK9yXkuOAOvDkYtH1KVh5dZNcLvgOD3L7S+bWHf4Dn20mWRLbjaRH
VRGt4l4a5lWyQo4khz5ohLT9RG1v4SBXGmN23BJQFLdg7Fi2R86xX29cO9BSHj6BqfvTiMxtoYRy
wFmRRQgh73mS/6sBOdbvmUnIbRkHpGm3wJgsnVXcpkmA9tzFEW6QLJJGjKB2ZzJanRA//LkLy5V9
WrkG+98TLkbfrtl5Uq9ChTxK1ac4tRLJYoZ+GFAPjUvLCKHp/n7V64oWgIW0yHVlGyIooFPvM3jb
q1RPcf1aStgexanmtOLYLYucWtWn9dsbF+ZxcBF4hBUYaklbpt04Uz2VM7hWJDG5Tgyu+eWw+Yq9
UiJ2GjIsaJPfvaYfVbQfcZ2A6R8lY7MeShWxxWUEFMIRP4aH5BhBvBe9AgPC5H0tqPNBKDlj+9gK
SrVrJXaUDwo5R7HDFez6xyFJ2cgVkzq3vNVrkg5gKmb2Ex/lG8RWfjz6amqjdOZj2fLhl8xoL5oh
wfjeazalvGaV3Lpmfq63B6XNaYgBrFgbWvWEnWOwdeghMqBeLT7Kxhm9rbSM+jUjrQwbsIVzDvrq
NQzuMTjTpT9jO2Z6lRPdCXxSvpwl6LNOcVUa19lgNM1ns9VbvYF4hP01s8KPwwQJ4VU1CZdy5Hwk
C2O6K0+kxP3yTf74d7+4VNR3j1SofcBh19yOMpuii8t30Jyjp9FUfAdgKbkthSapTX/s410PHob1
maZCW9f6WxGZRRkyzMcN1hSS5dkpD4H6JnlDNE/fNSXAbU5xUy8RBfT5UqLnysGfbS9G7cUdd98j
rg5NvAFTuyqHE/kRAufkgOf3KM8TTvSqt1vw2GHuSUiYRAoo42DKgrrTPJK9oQ7CrYiiGqDrgEh7
iEXn2GWkXu+zSLZhNS61ysfju45PzSb8pmdlajtmZt+17vdfLzBa9p2aY0xtQtPuQa6JnTnfzPgW
uS4ht5LPgBhJbi8n85RrwyKHbngWX76shwQAUEbBKXiokPGNFCuIAfelW2+B/EPN9R50/zox2RPk
OEbpYn+1gET0XAIuYlRR9PCQWQalZ3r7KFUfyPonIAW1N6QxlUgWGWYb4lUMCkeLukzOmQam/67X
QVTH99yXAlnvOmFkwQ1W5ITumuvN/6RLFu3TwrLMf6dfJnD94q5nMQekb9uF9NQwbeVS9fezWehB
YN9GG17W6F1NBKw2D3QmDkhLmr5yMagHs7DblRrhPMxikczoovg45ObKmJPxmCsSSwlLt0MbqtPJ
m95b1eD2ePTsPPBAgkN7Q5GXOb5UqK0EDTMezwcOF3053ZyK3aLv7FP0wFc+0sLulqrHAmULOfOJ
cZxLuER0uSDT28xXS5DNRVRi58yjjWw1inFEWMGhvdD96fWIJSXF27ExBi0OgASte5Q4zhAXWAD3
mefNUyGwj55Ms64q/c+sZR8DMjwHRg0PWZww0qzBel5Q0QlOoZqcZ6sJDJ8uCQwnIiMZmA6GeiJX
YmQmL28mvUVEhmPn+fis4khlNtIvjNYkwJ1lGG20dRaUENC4lX2XdxI1sV0I0sqM+XCpjbOUa0nl
7CcNXXkjZLH6WND1TuTqiwI+53w6LDL2P20Gky2YF6Od0If+vEJYe+NPg0lmQc3U2DRjh3wbmiEQ
6wySmRnfnYeg2X13ohKS9zt+3zaDN+Lsafo/np/b/39wtxPv1BRsEexoDQJTA/F8Xjp0BGv4UilI
gFo+rUZ6D8eaK/W469o3to1y4njeO0aB1IFJFZydaf97xWwLbDEA8te7aim9CpHs0a8ae8/N5Boz
C4rJievwOqAoMZqUe9JSBFeX39b6ZyjWBcAi1A/2Y3J8e0cRRdjSUs8F1UOCYF3pLp0LXAslicMT
YzCZenWOoybI0q7KzO7FbCsFLYDZWTpJIMHzq5q7/LAkJ9Z70nZq41uMRz041XzzAwAxwMtF3nDJ
1exflTt0hwb59s75NRM2WxF/FkRvj3Mlg434JYXzpoRTdThqlqlvEK8bYhylwHYj5KukTA69VyrJ
nLRVzql5G0BciF66ik5bBT2XsOH7OrFBiXcrad7misN+qZdJ5EXkZQzPt+sq8ZpNCzdSDBZ6Jdih
l9ik7az/Q1hx6EWHDF7WcSmJd5JfRkUTUsfnNFPJ8tOq2D3AH5PutSq4d+zK4TCEjWfj0daPzF7Y
XYAgeFc0m6XaSwkS3btA0fycAh8vlsvck5pOCENAVjC9VQ0dGsQFC4+cLJ2mBHZ6GlnHiBrFTdqp
RPMGHt4VEyO5m/QwUOvCxbTgeklvWdp0O2r2Vv63F2S9x1qAe1QQ1RCgc+s9As13/bGgZHu9bygM
AVzwS4G8eeRt9gGYDNzSWHH3cjex241Dp2DBOKiPguB+79c6eMEU96YxSh+DL1uiE6ZNBkpS40B5
T/U0bY/zURbkCsJx4dBrnJ9Gxhe46ZZDrigSRtN/k/Yx9WbvFfP4P/MKmTXP97dBNGoajKTEBr1s
JIgcseqZQvWSQXVeEFUWK3NuWasBW8ohb7h9ti+/ThAPQmQxzR9OD66GvJKnOegB6sSHwgaMNvD9
TUKV0sXONCFwfP48AUmqsrfNoDQCWgTOvWI5o5PFsYyG8DSeXAEjn1W9iFJ87wTr9lDjTFiwcqQP
dVXY53cpit8gbUlWfwdWaOwYUM9VLhfgGjrsbBQjquCg1utwjclZERs4fp0/6UqISRxmhe+g3UZk
lVrhUapWyytZCoEbEgkJIn0k+qY7Fe3mp69+ZrUCBhqvUII/hAiR5buYuX86Nbkgz2xNbhxTt708
gxFspEd9O2y9d7wmSOKZid35OzK9D2XKuJJjWRYD02LdXiPvYh34nVmeWChmHFBi6s82UyCQM5XC
7+ginIVqe5umTyTOnT/wZsQtAMkh69ElJEWDKu5qds8lt4nbj5RJpkkOZ50J2BqT+SYbamQlwEdY
KniOzpHjQUHOxuu8co9T8QW8lanIIgv5SegaMKroRZKQYQggL9rjaQMPii9vzhL/i9baSzMsRZBx
tbx+XEaSeWoOucdfGIk0LrWEJlu0sKKLIqBonS7bgP9EFJxMo4UMJ9RVndlrgTXJ4jHWRw1JUiFw
ckfN0PIqN/NSQpdGyAlBtR2NZYJN+MYjtyBoHv90MP9t6OuW0MvOwOfyAwdOVvZp/13NBVPY5JWh
Ol/5vNfIZI7xcWQddL1UcTretj1D4KkdX49fsHhtkR9J9O9JwZR9QfHyrI/bqYxWbtxtk5McAGeg
MbQ+YBL40Dr2aDmgMTdX2Kn9K0+u28cj2xHYjSkGX6qj/t3lg3S2PCDlR5WwrWr6FCWN3JuuThaZ
Etnu2P9h0tJgLciTtJjRkls+HRe42uhe+YOf6/3p/pbM2r9ZQukuaymXXQn+hJf7rflDfiQRpfqL
FbL++iuggryTiM8CNIbkX8eUOsTlXwZOfF4POCIDWZy5GRQ3+VXtCy0mdhzNhvJlMrWG4sieFA1m
X7xJhEw8zmTB2KoTnnL1nUKVSMAGhshftQgrNgN6Xif9V4QrSUARUqOXGZe7RUil7bJExmdUlL0D
yvRXIcIxF9vGiobJoPcKjV5jbdzZ3rYu/B3qPvOwFURxel2CAIru2UcXux61A5mLoHFu6qfDUZ99
UJpITcAiCd/oiiNnWpPe59r2vWy6dBLGvaJLv5XEz1rBcBlHfdXrNc1XSd9i7GHVmmQ5idDzZ5Jw
xajBbOi2RKT0U3MoPXyExVtPQpAQs7QuYNU+RlSMdA2D6LUA2/klk5aS6txhrAEHCKFIRnSvFqbH
AbNLxQQFqhE44oEudemwKzZPw04aGN5+wDGQ4vJ62MrMWO7K1kBa9jEVMTXOxKRO1gYgw0OzGLfH
mp2cweJ+7RSySz2XacfcaVZQVuOHnh5no03qcidUmHNgAzq+TgNgbkZPimHVMb3sGKKflx1eqSFO
qXmSe9ipF9NN//SoNgpWcVk30rum3/w40hEwO2oaktWta5vjMse2AIbNIhq8nhZMFIpQIkIeIlRF
vf53xJbbZA6fMUtwe9786j2XnFS9tzsT6oAo4r5VTaz3OdiHgdKXWk8vn/5gDNxRvZcPV851kCvP
0z6049W8hIZFePpWVlO0r9G7F/dK5cYz5Rr3Lr8WGjUfCEQroX83BbgxpGx+AnW3rW0nnMzVaoqk
mMoYoZSFoKmAnI1YVZ3u5WMsdZvA3g1V3qOzdsOdz9gSAgVWI/BLNBXXtnOqOVaMqkUXQmtv+bt7
kZ4rvQuedrle2tp2uGcE8TolwOhL4f96in6awqGx6A0T+mbGQViEMm4WHwtdYEaF2u0LpJ5sU9F6
OCtGSSIA7gYlSiEqSDTlcDFX+dsFx2FU1votvijN0LGtTI0Ez6XLStH7qjXpxpsWtluUPssaoJR5
8RkaFTQrPdKLanz4AJgtobAlvrRGreglw/d1P34qmic5KG+85tIZVOd9xK+keMN6Jw6zgBcIrgDM
CcFHEW/XT/rqyuxorWYJCggFlkeZe+y9BzDerrLMNws+wTFF/dinUEhcR84yDlKJnCypTqiFb1X9
oo93U6rr2Fsklk3WNJZRS07hx90Orvnaj7i/cMmzi6sxNPQTPiofFElAAAeOP0SO26P3hyR6aPc0
z8snA7MEgSqoadye+2A4NgAWm5nFz22ygKzUaFUCU+iw/pRk4BOZidcLu7XVeynGmg9MLT+jBo6O
GTaG3eQzJO+gBS5ypd937qDrO6ulY6s1rzRjgLLxPcqfhvjz/UZGp0ktVqoiyH9mhfpeX/1+Jm2V
/Vn03ZtZsH5kLx2+TMkEg0+WNkjAX7i8cPCCeOs227empTeOEU6M0lV8Dsm/eZ6Yg8RTRRPL4GsS
11CmHoDtAHzYFdHS6weIFAXe+51tLwkHFCTXRs1fRrloNm/DYv88QFgrOaucShoezjX3os56o1pF
EOotK1jFSyKQ/y9QhQ/Z6+raZP/QIzRe16hkAslf/i4UFPXzyMU0pVbYg2g1uKiGHPFaHLJIt06S
Ex2QGdn8VBjY/lKntlPM8yKDP+quvpJElxMTqn8yyrgow5ILpq68tCMPUBl8CW1FiVryFDmJpqR0
YfKhVJSNUppxkHFR4QTHTGnCiJcb2g86BeophGLHXxeKH5QML3slult0vmEkZa6qi7eX562K4hwe
7iX+euIGoJlWx0FjuJww1NenURPwIeWlTfR5xVCSp3jcT5mU6O8CbnLaWnSHh2BBdXyBwQ+cICWF
HomhLW1DjFKXc0eJorh4cHdO6a/W4TVQA1sA8SBwxDGL2LQnCc1PUnnau7B300J3ch+4xnTWVFbP
BXLT55eNA/5gc03ZZ8mvvXkOxT90fAxfhg2v2qg/ayBYC3s7gF2akJBbHZ4Hrkcc9TBeBPCiegqd
30aEsvx1sjqhUcWTqD2aPOaTswZOWXDhEZ0SiBAj7CY5vDQt8WITS1XYNJHsBGmFwq5DQ+e6QOB9
wG7F0YwKydFEFGDEvVP0+4wUPZuKBZz+lzWeU7fMLKrhsR9BtOd7bIdVEIKdela2WDTo7gfmQi8b
UgtOEVeuoEl5euGsFazXzz0wB7yL93uRZUJlH/UZAKJt/I7sSkjrIhnoRNnzSdrJv/M2YCeObA1l
EJViyl0i6cnr11thzf3PHukKjXGNW80r0CCOrHRjp04ARJqC7RczCxrJhBhen9TPOVX5iDqc5DBH
Sc7LmpZ/Qu0ZoTIVOsC8xVrGbZ9/ymfM+QssaEZGilwYVZ0F9ME85zSlpYtU/gm6ztS368d4Lc4v
TosimuDkI44Dwxd1xJakxhXfFuELPg+VsKbgCJDEyer586U6wNiCg7EgYQWOYvIPqfbmsQwH0+Pq
1ZpBP+eQf/k6NH9bV2I3mUymC34al7Lv1Zt+9pZyVgRmFhBnMSXW90dZ50S/rhmMwJ7OCz4zRsdp
Ccehnkd0tDAZzdz64wc7oP0LQV4g8WdkErsZCveILpHPRfhWYMk1anq1lcTNxnRrJG07bVhaTy9/
ODydbzv/ypHX9hrGNleE2Ky40/hZJlu5h0V6mej9oexjG3nIuDy188vNodR+fnLMqOgo6lklFbtT
WaGh/MvixK0HpZp12sn6kmVftVsHcEX91y1kteIxzl1AIdbapjpgGV5Y2s/0UGT24EsipfK7zL/n
jxk3SJC37kppOn1AEjex9yQWWVAYNI+OwPsewowqSYQpaCuru2EO+ajG8lHHYu4/D+LQwf7kdgU9
UWztMsN57cO97lWzQOm/nKDPU/0dsxQCU8oAbHRTjx45XvjzCP3swD1L2dfrWEdf93YgresliEM/
7OQuQ/0FDW1OKfhWHpPaOjLCRU2qG69b0d3x4867dwMVZSxAEl9klulMYCRbJCh4oRWyb+91hRDp
Fb7y9rlG30tpRaHgVGSaiStATxXPPFnmRisvHD0jpXHXSVcB5MzLWFQqydK0JleuN2T9vaJnc4ER
WBnUCD9rq+pTVoZoHWDNjCFPPtItT8QDzCGrTIi1Fcip7ATSdr3yBeHWpi6bIbtZ/esU7WAV93PH
5c1T/1sfTsBcqNv1ZMs+dJxAq2bSMuFCxN4F4DaNl5AZTit5JLch/de4OuFK6+Ne39RYX7C4tBRI
V8P1ExWdhpbZb6/o9d7BvmkMBW/HSqo0QJey2bUYYICEz2hquPILJpP1GiY8hE7Ycfvtbp137JK5
q27MQ2hS55wNHECQbJSV1cDtX7VAKl0xKIQ90RJMkhuvp0rwVnNCXvRT8CjuZYnRvrBE85E15Umo
NHL4hM8bWdDKMLPKGPRY7zmsfYS6C/QOq4n6/F/AgL+bNi283Dih0E6m9zP5YAEmKhLjABxJdWLZ
R3cH5ebXPxTXrTJu+RZ6DdIwIx/S+n55JG0mRlQzJRFbeB07ftO7wBkTWynIIWsat469d2sgcHpY
p86JNtHCqKb1jzn3TL1V+iD5t/+Fx1nGrCAAZftGjWCkxA240xLMpT1JGjumc4zZwhKgRfzJ7Wmx
1ySH67iQazoBXuf2ylQf3FMBy8LGiiJgUO0Jz/OZ3kastMBpxBUIU8Z92A8FMdhc9XyB28Qsq7Co
oLB0T4YTpmTENGw0p8+PbCmS/kNI7/K9Z6o/qmXLu4Pyl3eRsVG/VWwLoI4wnpZe+h37H4KpIVqW
8cHB+AdVVkhx4YIhez1Qnk/hG8xXKb7zZ3lgLt9KBm0PpIVJuI1ZCfV73bW+1FfnBcN3dcknzHP7
DcUMf/+1JvoLCTV6WDscwT7L7o8uaFSNIfIy/7SMLHcyZNL9xwXcOhgLCfEnTPvT2mUDD04MAqn2
zfwTi62XRbqb4z3Fpc07ti44iEx5Gj5+KkJbwKR1TAntqEWRJVAZnTuAavEw8khZSjbv6PCdk7O5
SrIKDXGWNlSbuTu4JKkBXjaRYvDumxZeE1B4pNQQrGXK0J0FBPWulX6NqYlQetRAmvnu0uUnBpod
lZbuO2Vxo55CshIvbCe6yrMWAm8jYl9Tupo0jODf8/JKLfmi175bBLOF8dcvAYRpp94lGG2P9Cbp
k1ReCJVl2YojNVI/sR81sxEKoswpS4kSkRvybQeCPUMGgJnkLErlK6hBhhnLdn38NFfcMKu2NVBE
f4Kaombbd5KXMz82ugrbO08QDAjpp9QX58qgGc7C+UHHJQUKv+pb7fgYXvvkW5ys70fRCvG7utiD
rJgDG4nehvwgUg1wMnni+062MpikBp+8YLo6k8ge0k1cGqf/OdkTLs8B4ny7MPjR0u4f+wYdcAWq
pEWUG/vKgLFxODyhYJ3y9eEoBhMuQKlMhC7flNU5ORHfQKfRgKEhQcNX5roUtpLptm/2rNYjC7pC
DMoaiORtrRjZaSMWuYAcv1R1mscLmGuUbAn8Fq7x/9jAycJWxVoNN/13VnuNz11x+hJN9lktwLsy
cUhXs5Lqi49aHu+z6Yhnj06AVTF3BTJut9CNuhjtlU66NbQ6X/w99GPI8uZp3Xs+f99/TNw7eB7R
//yAC69s4h6VGU1b2anMZpSYCJSPY/lViSYZkPaytkkxsehEnWs4RhF/u4RLK8CG8S2vKlKB4DZX
G5a2kvf5vvFYHUuAxPLJadOFC+Pv5rqTROpGdFLSDxeq6QCFHhHujUf/yWEnYKLabxgzwKOKbn0s
F0ohEOdBrDSY/f7s1f0I9Ieu7vVkGRl+9SHgTDs7ER8tyGXWATzxWo/acTR66OiZhr5g+Dr2a/XU
VGJbthqszk+CLiufPt4lyq6Zf2jXAqgv3Adw1p9BK3IpjPcT7STKOdtoeiFeagDBmVXmUMzm749o
Re9T73ZrJi0sJQ/+tQOaOSYipsQlbtThHFjQKc3HAUb07gwFmP0TtOffzLBTxbCYY16eE3AzdQ9B
2BFh8eLkJF3U7EGBYKjEFAliFptAY6WJUo+UE0jAfjMi4/FuezBCuAIrwpcYFfhEG5wbcvYFkdyw
dfhz4eKV6ZegjIQ+gimxzd9VTqPnjFAcIf3hg7i2NG4xGK46nIU+yiV0xgB5Ix+1OY0wspN4KGga
N99NCVqF59WLaHj5qXglJbIqjKaWsgPTH8ideikq2TFuQZ42YGu71rWjDLfTorOHV78xpZWcIxer
1+sWU1J6mVFZKzxr5bhG8x+peT09ucEsfPZz5D5Z7xCwNp3f87AL7+r7hlXDIqnzv+0XheHDj9o1
Nn1IMn9eNVed+wlEMzi4Lt2InBeL2EwTzValsozpOGUNnVgwrQqOsxrVDXX1jhzV6OKkuGhHZgNE
tTjv2lpDUxxl4+n005QOfZarWS0hJT/Hk+3BKNmSGIYoMUOzUskELlb2Lrp+gowhYE0H8S9W99UM
lnEBPkUWpiO/nt+W+JkrnZhzHxxzyFaVPz8dPwr1qgJwV7kIcdAESyl2nb80g4tIXHL8N/euJM1Q
Vo7J1NqHkN7SVpnyfkVxl2FNk1iWeIka791xbw9E+lbeFCBvdlvTK+ANuuE9k7A7G/ZdEqXU4E0G
kOKwA5LvYb++VoIVjWgHgqAXXvC51OCDPSsEOEoI5YKmGqbYLi96m301eHWsT16/O2CenDRd5WAF
cID8OMkOr6Jz0BE8C/CN9EK/qzyNlTC7jqPf1OhyU9vokwVgkyseZiMneiUu1kR0cHNJhjPzTtQS
iZfpo/+OW/ftVpaUcqweTd0pnxtOCXonLbsEjxjjjHxqdeyjkEqz60Yl8LJlEmYfERJv6dwa/MYb
7QjGsPhuMrd+XKbn2FTUeQFxJ2DKxUusV5FRgZbk4uo65/2ZCUlgSxqLdqbFufp2vS2kZ0YghZww
OM9UL0z4cNgJztLs/MybYLOxOfrw8bwRPrtLYhjUVb8oitXYyLp1pg68GytXlJd909RXEVW+gRgF
kkqNT8Efn7NZU9hgFiRbwD2NpEedXbWbb0OwgMJvRp2X37SLyi7IO6+bWox2dwql3AQMjulLRyhE
VtCE3jZ54sMWLSVX9yyzt2dByxhUrfbAvb+xpMlvo4H9ijaa/5YBLfRSgr3nji9i1q38E/byOJlA
zWjcXzM96LwoqEEbmMrFwey4ZUQvIjgOfvVD0uGSee3CEFZ89KARzc8vRP7fJymOVsG0XIxB45nt
0giMVgbYZSpaaIz+8pP/OMVUR6Aaj0XP8GmN0nga/JqheTz7Mu8MVuzfUZbkcHFMPth+/tcxhUiH
nsZvV0xZUDQr0DsBGl8Db6yknk8lLMbk+yE3T1bDKajd8UCvdHJ7DmOF6JkER72lEerle4nrRehF
/HFKfpLN153R+lwtlzmyQX+T1TDvG8cg9dB4eR4ieXt/FILcSq8CD3kXr2QGNx9N1nFclQpsT4Ne
nC5l50ZByquTIumORXMOe9sGn/mvusn9/eK+iN/+xbScdtAM6BwhIAeK4xfl7PmiDYAEzyROxKnt
IB9AqVVRNOQVzACzCcb07mYe95AiMqFem6N8PvWC8ywdLruwWl1EobUz6diI5aUiubvWvBrQq7ES
Om7YIoYhyMPtNMAE+Nu4Mqb6HT8V/lXsXC5DVlNbdi1jMkVK9VlC0R2N9qrD01F/LIAltAq6T0C9
MWFHpQHO6H77J5tJFOj/+0TfkfHX4fjjgaNUU2aFWiWQqyLnlQnGELvsX0LL96ZwMzMG+CnzJA7C
Yt8pn5hzmMXYrbsBqvq/gTUxMew7MvsudXyZsGTDkDxCBhJt+rUQIlTA3uOmhTfriBoVtToI45h9
b1aCLR5l02Cn/hej/tcMk8zEdDt5/k81pF8GbtK67e5NFF3UNyv8M88EHmQ4oh3pz4b/UesXbwvB
aA5PC+FyGETDeHiMawWRFbxXrV3o4k/j3UtXay1JgY9u7aDIq8P089wmLZ5Y97+h3WsEILZl+quh
El6Qb1JkBth1gLR3//riNwpGM8XjSDg0n0L6JLD+QUIJqAtLjgKlhsoDmF9vhh+t36aOYWtib7ct
AI5bS7scpi4iqB7TLxUR34uQRWw3sgkrLUszmOcSNi93mzqMkuTxeeWuLNeLhRWLXQeHAPmMaTfx
tBbKVHA6nldt4Gvx5a3xVorjk8sJTFfNKaoPzgLn17hBi/8gZxkDYcAiFkki+T9zU5G4P8l3siCG
w87F4Orw6a9hXRcxCNNGK64yi6vtrh0frHJHH0lYpVsBO7qfNXGHlwXhcAfGBSC2MA8xxXdMYS9B
VkmlOAj/20k7s3xHDYFrbR4q1PdIHNpNwJh1gZKx7beLgk0wkDffrduqZzN1QujM1Jt8gAxhjROo
cU7uG3cO7MMKHUP5+LGWBEB01On1UJHRAu991tLA8SQ+RYrI9ISb/dkT9P5YfByiVAakX9whZLrE
fwsYnaxl18M8xyuFWAo+b6X19woCSwFSazOeO9g4MMGYMPP5DNjhxpv9GCBWWjAHPuqFa9O8VsiG
nt3hJF5hueS/Cv8GkWER0WrCDTO/l1CfkdaYVXxA8hH9rvEyi5xowSPRgPYOqJP9bsT6f89k2Kn6
UiYna99G0BoUAF9rqwECY55wjWVTlVYH3+fL2eDDeaEQh7LW9vWgjpbR+eDBtGosndGxTNcxaPqe
UBTiN0ZGwbYnc7WVurF1obc76LHRCRFuTum3LlsGH1ht2iQKjXsz7DUjUK0YPq5bBEPSBhKhwBoO
yI2gYpEi4ZBBvcD9zNREyhNcbIsB7WXtUR9IRyO/TnAZPx+y5sVSTg/qfrisYYyxtgIIxThaCvOs
qsenaBR1MvOvuDCoMaIGAHGkmwCxp/t6YO8LadA2LvHFiNRGw+Bxk+rkQfqpaWz2PKXDzrmICPGr
1lGWUwZS0IE4u64xWso7HObG+uTopQkD2uYRrqBqpYvw8CDblMnaU1nHYpd4dIlKIrGE1+Y2+Gb/
+E/reai+3D16t/4vihJ92j7MfsrC1mNtSCq8deg5gK3H4PZ0M+d+QR7hFaQKrEZr5MEYMCQC3dOw
RRne5lfp5hH4pHFyB+osWxdi1gMEvIxqJj4pyZ66NOy1BKnlVehZyMY2mqm569GlNWY5p0HeqpEH
7p2LN3RJlyBp1F0zRYcKhwD2axt1feff9S/8a614JNugCyU4et0Tehei69Obyy3uFenlqEbd47DH
xi2o8aEdPt2cmFYHPzAxbhXTxixVPv29R/AcgfgXpFydtm9+PUdqLLDH5P/ph4IF+aRzHnGk+7dZ
Ayx86InMkBX9wlVGTxtMBDHn9o/5lp0fk09ddl3Qo6pM1igJiOJLSuS3dSYF2SWBAqO1soYrIfhq
RzfFSgU9RcYczNWL7O8MEbIbzOmx9FNPoL9dNdVszUJew4yDFieYTlWgD2QREVcamjchGOeEwUYS
kP8dA7wjuGluyGvt2vPcmgG0gO2xYpd9dM10+IsqFA5cvNJHJNa/DT9kALBARJ82ji59ufQemcxs
Yykxg1kVusyYZzVgD6Pr2a4GBGXXcVPtzejWVIOPOBQl+nUc5mLpGl57QuUcz5qe0UkuQYMnlX2l
pwZWTGH4/ulSMW1YV+557GDp4gC4PEsA1RHZlZFgkKzHUG/IFI0b06BNLTlG27U03O9zLr7h5pBA
v4RNzUzyeL7FGOL5+7HQq2OAnZUrXRM6FLjfIzuIEs7vzqhyDaYLr08I8GylDVc4d6LTU8sHZTrO
HXrEBPcW2XjJpRzEmfziDkobqOEBca69pKaZfv9O/OB33lZiCG9hE+5sWjx9LGkAsrAtVUoZvdbi
CHOpxqqk++YwhkJoI2miJJwmE7AJbOqZjrs3D+VYtPyDyS5zICROi4itlnzGgunySTrJ68FDI9Um
9RYCdDYTTDm5PyJod2Ha10THct+F70WUEHSets7OWYnpbmvUWXNTCPm9uFnCDJmjUGhWTVn+TA/J
Pcnu1dY0KV5aGgmEEQK3AeNbhHVGjaSVX6nhigG2HtuIeXSmdp/kC3MwsgBeBS6hIYBaegNFr0yT
naI/JSU9RfaRNLn5KZphaowlJsnaSZw7YkOKonq3hKQ55DVsjjh4/YVLimZpVDAM5Nc+RvAmKsOR
7R9vbRxy2TZZQPN9QescMXKG06PKOn83T1yuLBk4CdCPxAyBcD5khB0jLUWE/kJXTBi0vEn4r+i2
PHNBtDnKXkrTdKiuwMupiTNTc4WZmWTjQaLOkA41hl5j1IQlwxw/OTM7okKucTsSt+88cbc2IgUN
AmRoxZWP/llceaWGKWgsz4bXQE7AK8rk8CPVUiTWr7krkHrViOZJ6VLgFXztWBVZof7gm1U4umqy
Amr+h421K4bcmu8Fgr475C7/jUN5OfOa3e8UIgjWsVaoc+yILXnk/7BEg2w3xag8KTLgvYj23j06
/BZZjCiBrJPZph7A1ZAZhBJ07YYEz1zFu2Je34aov4NFjkoUkNHsumjcdY3s9EeBw5hAtN4Zn0Uk
QOUrPpBlzR+Aw1t2dwbyRjvvDF4JGDmJbnrJhjjtOeqXRvZf9IESysNzC7VF6g9XHtrt7XpcgRBQ
qk6nlIaYpsfkJo5PsO+C6XFjzdKEXsc5gZZ+K94KBpkkW+UgRV1h4ashJ357dwUlDto2BiR2cmf0
Qkn/ci2PVdHPKCgnWOrmLoCL6kvWxfKghgSlCNFaTzS2XpP5FFM0GtufMPjuY+LLAPXiQW8CKCb7
ISqeDf0sJKeMCMxAaXVBA+ss1yrVlnXepIni83ZFJD2JgrFFCKdpuR0Yaup3qE1Z7eiDriKQFaBN
Ik6wCQcp9BIuTf7gRXvR5s9VFUFop72bkY9l6gg7e8/VWT7m5CKjnRZZzuwcdNb0ER6n6PbqGH1E
CqsVZbs94VdVQI4NFnaOvQhls3YzKmzY6LeABG53oXwCsK+NT+7Xb70jSpPCzihLUpak6enjOqm9
2hf2BQF1I4/gimZB/PbWaKjxlwQI8/lvde/ZcYdZiVCXlCkWyVwOqqAj9tc/kXWk5O3xiamTBKhh
q/brfHGHD1SDVrN+mB5VAIfmyHa4PnCdFbFP48C6NHVYIHYMFjq8QZVZ9EsKvZNVWvOEVDob3ycR
cqQxaPMkhXaKw32fd6LQYTF1CQok9BSbCFB4NBGtQDZjwBJIodgpJI1DEJFEaG9StWnpSNxkIX4k
UrCGAFgrpV9DCfmC6B/jp3hDVF376RNEevZA7kRG5hCVYKwB53pjXCgFELMPaOGVDYyTh+Ii5IbA
WjJGLz1eCZwNK9DAKHHC8kHhIYzmtR8MAy0+mlc/SlvFyJHGXvqHE8qlBjkQlr57eM+LsHu+yepc
L4Da0ub9P9mcnbLYINBrWCDuV3c30knvVGnkAbGgR4kYCP00BO2Z5txxNlOe1EBqqyFZqUhVRjo4
VM7yhjLr5L7Ny8iT304w9eQm1416ze4kDKNKZbPvPcfWlf6bWSX6xX3+rfCI8X+dSKKtZ71YP7EC
7hCBE5j8LANfhCQVb1SVaDQrWVR868BtlDUS5paaudYmzfotIPeR7zH3o1gx2CLpEXWwhlMTvNxh
mvG5pVFXRMA5w//WI7PHPbIAjf40cjFdBXy08RACSdlHH/qd/LMi1H/wwNEG+cMkF4bJAbicB2+R
PBrb6y7sDKHJjAw2hkOSMD+sUTxPk9dzV+NGVGg+d/PW9vkQK9aLisBPT2Sb0qe+9XgyqoG85HMa
kj1fCIom/ZqEH6wcrNVb84Klx7/J6CoKEc16dOCoeG/DS5MlVioqlywre5j8BbZztz+X1doWcQiN
HRGIAKDWmYfqvMmuxUcONci02NQ2UkIoChMIGkUrDWC9KrIp5984C7iksGXXxcYakSM6cHkUm5nO
byBx7eYGLkBuxr4I64UfE+e2m7TXy4WQVecKE8vlaKqanD43lGC09JsgHaDbUfBvtqw04MmkcLzk
nSJzFI4wEdvAl5vASpH47LttZT0Y348Z8iCu1syhOf0XQj1FJ1aXzHxRgPTesILITr9j6gmVoP/f
t8cs/8Qjc0iQSkNMtBzT6fZ0I0QYf1qfg0kaqsgg+hnPN8I0CINjK2G9rKCpgjW0GFcW9K7bbIcQ
IWZk1ZozENP27UFnapwKKABubMbL+EuLY5glvRYhxM1gauEsNZrBBDleL0FZbgN/0BXdzcS3SqM9
WufJ38lCg6PFl5IhH6uDhEGA3mw7n/djxoIX093BzOD88ObCxaIgl7txx8h1ya0YLted3yjrr6aG
05jfdwlWZRvwrWa/ncQ0nYT+u6MLMfd0N8Y1WnFOY30qy2Qwcp+bFNOev0zT3LyGSCP4e6MG+5O6
6qAUuLgldGVaauDYLwU4Aop1GlxfNCHJI90LaFY8da3QQasW4zu1G6QTdZBpFMeaOf4pxMu/wQnx
bzcAcBScezvE+cUjZS5MSnD035GO4qp7dLPDfp93HwaP6xog1hl62lFk6ZOIx8i9UznsAMvM2UMt
ahTgvd3Yq3BQXDhKs0L2cgzfzktEFv5FCPCsLU1M0+IOVprI/WfiGnCYjTDuaT9WuSN4h4hE2QD/
Yc58c5z/6yrIRmCphCwPQ/YgOqWfxxvTrYqx36G2jU9JU481+05x6g14qvTtrV9WQKF+hoYY1/TH
KMKobZImV4k906GzwL53OTX/7wzxFgfrXRHrGyJVtpafCozam6JhWalYHJeIWmeUgIL6mHMUM36B
R9jLvw2HavFcm8OHt+Vh4qDFHkLcKK3m9CTEU5X0HuExzSRvjp+pUEnE1MKMS07tUEyBPLmnd7Qa
fYn7Qt0nVXYYswr6N0Fhx0aVz1CZUs/4EI1TRBsi5NMDm1Aay+wS9aOCULw+hiSyOxXjdNfOjoJ5
MYDCT/44j6qOduqofz5tI4J5i2K0kgVCVyV0YLEeXHJexlA7z7BxVLv2dUYCsBBu/i6uNfau4o7N
frivZZyEo5O6tM8HeZiQsuBSp5dHfJwyQ5zXg8NZyyyhTecrx1ZPWoE8WtzivuzfP4oHYmc9u7wM
o2Ac3iJFeDLiV4hDO/hcv9XKVHNI+MFZLHlFZdGOX0/n6GfxVHP11CmjjbOPNpWSGCrrebRl+SkQ
IPijC++IZWACMdTcDdF+BiuVcow3Yuf2Tb616CMSCXdFWit+dveMHvASD9maVYtb9KiLWOYV9Cd1
26FSrPdV83FrUYQ1EMo+oMgsGzk4owUSI9Hz4d7MgQEzJolbZoxIDsER42VbjbhVhUhNXVF9RKnH
oaUfsnGMqHzA6L8hpY9pBZ1NILtpr7nsP8g8JLdRFWUuo7pNIcjkD9rJYyQbtKR827xPOrqp2cAD
lY8zuJeXg8Ggmgq/zZUqNAR3KNt/NRirpkvGB2KVeTFPl/Ybbq8Uzy0b2wFaR68PG8LLCMjrLxY4
2s7yF+fM+RBwvuc7yrQxpxomf4wvH4zRDf4j9rHmMURZ4orU/qfD1sEP3iNoLnHzrX5LLMJhIdDU
JMrzm47svwHJrNlBpPieWEDjelQV5us2plaXMfDgQytfBP5ydrxSJ8SyCgf0yJIT74fCTvGw6SbM
xY2uy1/JGeykHKubHNETgQJgvj0+xQt+fQXEmteDCts/QRCvoDwzaHDFKYLnjGqnzZLgW5D90Vp6
mvLTmncVbvJC+GSpJTVqN9p+b+/WQ9SSyr/NTsTfvJENlhxfUK47kHXXi2wgVXee6uhqZt5qo05C
jc6z1VvmjkrlGCch9TF4N1Y1jox17uZKwljtvH7bnvloK/BWu8kypr1JIKpVKRuS2A7i7AX/eTzs
qZ7cJOPsAPcGinZi2mNha+SP8nSU+mOCuTK7YasBIkK499XDFWlw2FWJAj5h9E4KVfOeBsHEkDTo
4IvB/8/39CvGClzU2Hmozf7/LJtp570nQOU9RcNkPqtEFJYgZiIEdBonZ3YPMQTittGchF6H21tB
F5V3RCJKkBEiGiHBheRkIvvQHw/5Fpyc7iHulI6Y78H6+cSRi8DIl6TWhyvCElO2CXQthTmG6NNj
QnojvgI4E69DC56xoyAFgBLUFadzTq4SmvxjfIXAkFEBfHbMoXw7mxh7L1YE8Qj3kXOF3SfIT2kP
ljhpOfZ3ygnobnU59g4iB7jcDlbY5TDmQEoV5KlUBjpzonEW5h7NeWW1HCX8aYFd9shfR+X7G4Hx
O6/nlkRIjvJy6AfT48Aml3g5Cdffd83U9sQ1vnq2D8MOvDeDhTk8ie9k4WjtULfoHpedItRov96X
TxBQ3scc37InnwvC9bnmaFE9uCggw6dkE9rnHiYkWyso0wfRG0sdPx2oo2YG33CN4kJ5eLU7n6vb
ZdxXo97Z3K7r6aCm1jrISj3bjLtIer/qe2iKJQlZTx73+9c5T06eahY2vr7Ukk/kL2O+uZNBRIy9
aljYSsrV17G+YMWNIm/uQgu8Wy2hFoakn+KzDU1XJiJhElP4oIlv1jW2Mfm5Qy9whu/yyqw6KVJd
lj+0eB/koFe8aDQe1AR0T6kSXAM/HouSM4CMvlaACww3FOVptPIroSZMeVKApac98Bx79xBHw6hR
HLmlpZ2uGVezyWZMEIS/0N70QJ/Pm8m8aBBjTgHU8djAwHMy7gBxep7Y8bAtrx28mU9fVu0OPoIu
1FhKxGKv5flM0tn0WOB0tZObE0k6gxOKxTAaC1B0QwUrg/vWbTuJZuT23IwPOt8KDoP4b3iDC2W9
brWbxirggd8ihuid06Hqr0ZUN/XUA2p+W0kvTdAryo7CxVu7cS2daatODWv7DYbp4+gXDh5P4Ug9
6CXs3xMQbj6l5B2Jir14V1VukGe8U6ZAJ+tmhEn2ZII5bSAy5EQLx4EzJ339ThH9DUPSK9ijyj/a
Xt+8zCVKuDqDAeihH9XoNH+Skfz6MLLZhybIcstXbotVHxexTO3cqcpzPse3OJQZEzeg6Dvn701i
QhLvYHVaaiBTl3my+iUo4uGYVMEl4li0kHmvrpbNBBxwjY1lDE8nBfprMxmECBY4aGd0hn9LX3NW
tnmfjAQqxHQtRI1aSjShRpgHCa27IeV54uvEEA0QFWIQu802gRrjfto1wKPywv+u4N9P8a6lEqjH
SWAPp/gdkx1HAJ1CRpy8kZdGzVkSS6PpawCIulds/+boyI2RyPrRTnzzURM/St4Tx8GaTnn+/45S
1sTiVZi+CQ4keNhoTpv5+cDSwbsD+bb3dOb+9m8tyDLaN9ybLrObAPCXlO5t2wgKaGkGfklsF21C
cCo2B3P4RcVvvVur/AQ4aXwVCdpjuckqH6vAgpIcdTVCxrO9O91jONpIih4ZUOm2suqDIvjtM6MM
N0Xn/Z4GMZTJadCYgVfJyJ+iUVBUDmfd4t66yxXYp6V7Pt3pd3E8EnQ9a3Qy53DR4kIC6qBdZTfB
XvNBzmd4diNGtjz4uZda7vlhs2McEaGHI+NYwi4ZPllmR932dQtEaeHTpO98QmFcKJ4Lh8ANv2PB
CGyfj8yU+VDCSu5kBbofGqjUpCv7AJYw6y9CrHPr+OlqPiGeFExYV8gJv3C6h6jTyBbPRzIz+CPW
8NsGmfqKIvzdaIl9smO+Ik5mQmI6B0t2zEwWiSktNLve+VhDtf27wcmH/uJEA3fW1vxzuLonDzqd
t2bbeeGsOu0S4FUdA9K173toHOmldgFf/YFBIdyfm4B3fr9UGWeqJju/lIHOeGeIOFEqiS6JpQZQ
GgUVPpNdp7xqcauKO+EUZe/i1mfafbdzCvoJ4/4CaMnljZ5OQtUlu8eQMBAU7rlF+QMXXAVDut5u
YvUfAaqkPDJ0BYZWK/49AhrNLpOVMQIgYYuiJVyK3LxhlvF2w8qQJ1+pLm51FXpL9GPTHsuwmggc
IFuiIoawV0ifneTsZ9z75vpnHwmBmVvuernObbTOoYWDpz8GiTUTH2f/VAvIi+3gZQ64pFqfPcJj
i0q+5NfWcbpO3vjhpGhHX7VUOKhIoFcOO7xawHhJZgN0L6waejgzKyCOV3E39ixR9zLYRa5r0NyT
451W1gcVwXQ3vwGdOvI1DIvAycb3GGmBiGr98Alynnmo0q1IkxCtQIPis4HXf8QsvwDxorsEELCk
GKVfXMXp5vKINrqVoVAjTopZCLZrmexgFfumeOTzsWZA82v2CLNLA1yHj6Q+9mFJfwF/tOu/JZpb
AXiD3U5JzJI4WjebTphMOuavaiuCThza00Mi2L/15lBb2vwpxARBET3ehcrXG1nznvH4Wg3iwGC+
ZdIwWy1RRIv5TrrK4XWzZ6JVaF5RcaJPDxitsJL2TKWlVrqafgDz3puSmHUcHlwryJBi+xaXXDa8
IISTcyFWXkfySZ6aJxAglIGzIWYwageEROFnP4Qj34Z9TbL+9yrlqBOx0LdbTgbwRqcWPueialeC
fjU29FWd/TcWKlO3EobUvHkNs2p+qmD91E8r5N4gimr1iNbwov07L3zURWbwG8ogsSndNxa8QlSI
etRe6vtKkzA5kLeZqkpeVQ1J6Cff9I0q8A90g32Zo0uyn+6/S/CwhoUi92zXE3nRYFN4z8NAU7A4
2y2n2rRAG/NDzCJCu5TMw6bsuMZ6HWhWThEqNWGdXltP61UygpX1K+zid0jqy9D1sAX/3qUFWBbA
b2DKbxOmsKv/bxG1/xa0n964ZtNW0Rw6Cs3DfNBTQBCfDSo91X5n8SHvPRzi4Y0wEka4fAkmueZn
sQ3eByPzYdRfTdGeaJWjhsYrsFUNN3bfGmMtEgrIAS3+IE9zuVnnN8phfbWIO7mOXMLx2ykHIu+5
CXulU3RunwqOIxQhHd40KEgPa/MHAEsTHV2MITish+Oyk6g0GC3fngcDN7CaCt9qxgPbLSvjaGHi
4/umd8sr/Rwq7iOpYKfNu/XSGbrj0LDDlEVZf2ZXxyBNmmztNxJ6F5jznmukZsYj4XPwwMpITU3r
nLC/J2ZTKAlMfu6lqMcU80yGUmC5LWOaoMuAyQ5PRRthw0gzFi39oVRw6CfVtHFw1l9FwZHd5Zuj
/+/zLplnZpL3tcm6d/EjXhpcvA1vKPva+bmHGEqI63NvYiObPda+KRYiyrHOqNMJtZVIb/21+kT+
oRvhFNEQSJoKcUBhAOvHIL4jIg0GfeoYlrX5wDfZKkkbXHnrfBvQ7unvt1ETS1ZAjiNdysLRiGUZ
ZxHs4EExbYesIcXOSUrooWZijqrE6RIzUM++Ps/mDXZYkGGVKg0JqjuPnSueylc0jxZ1tQcl3pPb
x/CsvG1irnjuIzJsXNz9NDkqYtrZTgZ+73vXIXYEsR+dvSSOkgUm9QeoZ3VyX77/ura9dneRRYD9
WdrQ9Fww2NBkN2W+7Impf3oVO1raMFanou0p3fExdX3yjrnnStv2yH5Sw6VikW29SO15ROyPcMkr
RZb8B3QQ5pXtKL+6WnAf9cVRxHrtYtBG6YRaXBZ0WyW/ANPjD0LuddAgsVvZnrASIWZJwpWMLLe5
FWjd5mf6ClkN/fPA95vTmfUqVl+LJl35Nn1GBG54TaRWVtUHqPQwzZ8JsNAJj71AUSDurtN8RIwt
gf7esOoNiBw3JpTUEwdGSPnTeidifGTKsBBkgUnyVU9uIV6GjlSW9usXEou6v/91kiFpiVyHshC7
eIE3vSU+K3wSKorxw3vwItGX1j71Arxzl4h1YbtJ3P+Wo80wkHotYqvoj2T0aFm9WIqhxHcl6PeF
gR/SUk6B4xlYhBFb/aKtayWdzXsz0hSoYuODQwJhk8zgzcmgzK84AfD9I47cCsOQ+HxmHFXbGAT0
zEFCugV2jZgWQfb5QhIfCkwpV+UAD0Yact/kOT+OyEuaFiWCBBzKGzD9M9evuZ1qLyTJdYAEyByo
DE6ql8m/x46Zn9xTnAoA4elsp0QvtVsOGX/JeyxaH2ZdhjXHGchGKx6WnM4xfU8oEU/HJcXN+Zm0
mO5b3cXc8YvzAF0Udzp0sBpxjTPIekEeqoCHrqKBou4MApBUoVDXhJ1778VKqXUHsZWuOWwl1yku
339C1B32qvLQ+NWNiv8z7oB6cF8d/rZunyrwnKU2TQ9k0qIiqjEhB/Rj6BiCNUQ0JLcTPqpgBD6r
jaPTsJ/trWLS8JGvjUDiT69pdeeg2qq8ZOMZlU52pZJrehc+d4if0r9YRi5D9zZbXEViJuSbwHD8
9Nc97Npw2bax1xIWFP+ZiRhF3BY03WR7L2y2zFN6JXdqvJ6Lubs+03guCCMKOYvd4t4QRumNAIwP
4ZHfLpJTHsA4vK1nFw9gUSEbAq1T7sfCjUdqatPXYdGRC8zF3JkNEg2e/ScKpyl22+PPkUrLFUu5
XstkBS8Ykc47va+gJFv6VtG7jFaJFPe8PMB1yKRzH3BLFlTjmviS00PVvqNSShrmrLDQDC8/+9Lo
+Kqrn4JvgPq9WoVhz3B8+W8OgTb2tIPhex1/C0Ui0dRbZdx0779V7EktB3UHIPuGEaooeixaRECZ
eKtXkOzTlpVzN7Ss0XhRXkDKu7wMxWgr3PjtlG07SvJzumIV+ofDmR4UvEtlrjK5IFNLeZK7D9bT
orLbtWUjNVIaC+fjRKWPl8OdjQcNfUVYtkFHtgKxLuktv3o4L+cDtvHvQ/Q85zeLlVl9CfijXxIZ
wuE1HnxLzu6PcQADOwQTDUoDQ36JHxrKQ2PuIy5o0588rQFJj3aQFxYrSN6BH96pNf7RbmWV05mJ
yADVSg0HR1sIcUkGMc9U9v34Ja1+VGSWeYQq3AolldftzEIq9X/m/4fUGZhfmuF5gzFwrY2plGxv
k89ni1+4iXTlxG7Mehr6HNPuYyv6g7WKFAuFJJwmOIsJUCEQVj2RX4QcSpKf7pzxuhSsBQIZzYCb
U/sF92TEQ3AsLEdg/zG3EZfvqyMYGFzJaslxUlCDmSlGErySEw91Ol4SpOVvvOW6Q7jbEVnHXfPK
gIpKgsHZSxK3VLuHoL4v5Mk5efrCiShvhEtalvjq6+iGtaOkCPE+UEOLgMUunp4Cyc0j8Pu54WmW
7i1Hhitc3SMg3XH4cdldFfmtnCeGdXC7izfrrowzxdkoJYNdxIXbu7bikXzSKcsRmPihD/gVJ1D9
dvCjloRl0ZVmCXgkpLEY+TR+lObD6i7QpdzVfHiARpUkrxSHtPzA/FbBkLOmYPoynwWiweWsCegZ
h9JNEaSj/5AXJkHKATNtOH2oO0t9v2kLkO32vfSzUHTVxGx6oqAqRUeb54jniw2ugIPMYR/1mQfu
a+84TgA8rMOzm3gUlNVs0OcIqBEdjOJCO66YRhyCPMrAwPM2LHtpgblFBQhIRHhC4yMtX8ENHNUH
6/S8tQQRNIW53KWx7G+NLZ1YxmOHEmM2btGDfbPN4hSy3cE4wWWJx+rmUwjo+8jJ0zccb08LhR9d
cBjHB0lcZOk+e/TbHKQhgqb6tUpVSOvQZEfarVNTqfhAzxNxyQqLKW46rpRN4Oe2Bip/6dW55RlU
vCGYbWRS6LJnv9sYef/qOdeauZmGbJInnflthE3m3b2HPO4GNezAxpzTkIstJCWgLkzzkUm7HMUC
un2y2TNkYbkD0F9ugnS0DCddvDGwebGVPQsYkrA12wONPw8O8pAk/jagZg6OORC/r4kCq7PrTMvj
xE/IQjdb1SLmsXKQuhPbK9j3K64xfRVq59GFD5We/InrCNQQBrQ9oWy9d4kaBWZ+LUKPonE5wPGM
NCwPC9Qwg0h6mmKXGEjqSKLZte+ns4cHBB8MG9WV2/s5jQFJDgpPTYENnVEQtngNYQljfZkqopWX
rI1XL3hKNKOh+qeVDlik87eKVh1ntkiKDsuEnuTcAkd0fIS1yrdnsGIqRD2a/Z37IMCmTag2NChh
mVAnXZzoIFqv6+8b5rKthm5xuceLwQWURFYtANhE0BXsDeS3vX4b+JPZWAN1M+O4ONJEHpq/qrbQ
axyw2YRHYqgSrB+4RnKSi7u4os0m+x8+ZHheAXGjLGXTFz8GXof6zdC9CdfaUDgPqNu60hTCfai6
mXz0VO6kpm3+z1fw6x67x5RTGIg5M1gxL1AEAvVaggBdhRmhOJi/bbi51RrA2CJG4zQ6H0e2ZGd2
xauSzLdVrdLH83VqnYnCY4er4kaBmRj5XFRYRByOuOKoq7yGV1K+9YfqOotC8FnGFUs6uEHnvXGO
2BRTgfyv9BgJK8EP663Wpi1cyAOBsihJm7MFlS63RTgvuNNA6089VZfIHlzvFc7aJeLHDboW4Jta
Z8lGXHnNoE6wA1IslLCQ5lBh/Tlo4d9Oljfz4ER/K6rbuSm4Tibtmf3RmqSTL+aIkmcc2kLB10cK
FugBE9fTunrwA5p5LtCQ4p2iY6kphXcbBwHT3LdByl4w7VDOhJW9k/OyX7VNrNuAX5dSAlAEfG7K
6rSBypiztNZDUP9WCEmErDkR38v8fYMhsGtVoqvLtu0DxmpFrZIxKo9ibesWe60OP5Mj/0fA72iQ
BmWP8hc1MxuS9VdpqMlhmrb6D0FMCm2PFuHRHWaZXPb8naYCJXd8FKRRLSyQ4ZBgxOqw1OjwwQTS
GTplTYXvi07zwjFa9D3xho0r5V9CAHbW+8ldF+//XKfKxfC8ykqBsw9j1UdISodutNKcZdCV3EWD
91kwZTavUq/PYosAfEiBTgrGUAbWescRtN3KIMXjOaL5YSS4Ocofc+ykg2OLQ+RYmZZFZXsxeHQc
Pe62V268LTV4MrL5JbEeBuovomCXBHF+zzun+VO7SOpnBEDHTVn1el8/Irw9NlddjK6TAGzGhQ4Z
hbULZ97b1O95EBX9ZbNFprLdjQzVdaARZzTH7anEsmq5TV+ODb2AAACXzhlAI+aKxlDWnEaMb9Je
2lCBf8bcQ5xci5mR1tvz7tZ6Q/OqGrzIp+SGdVR1XbR6RbmtrEB6KdKPMYGxfJJMiLLv18tRkDa2
X/1/3T9HX3F3qONPTaJLedNV6fqDY6wG1sfPNwqPHOs/ghHywa3MVZJGBp+Wk4ZUuJuIAiIoAKgq
pvnsQB6/P6WLadBRUUBBJ4m5w/Ek9c4YBz7HTKy2HQ+laS/nZVLXTFS/DmRXWkynVdmX7sggDB/A
xv5q1KMYzbAR/WmRXe+dzQXu+zKzD+mlGdVHpGfP7yZ9gdZrPL8JxV2ooNDbCQYccsdEDEXmWJ6J
abZrkzkFmlGejL26j0LRSUBrtoFjoEYvbbvj1O0za4yGYNC+KIrJBzr81CZ3HumnxKu+596GjGXc
+jQu8DqnV3xWWfeBshZzdeRRl2iz/bXkcJT1QQuQ1fA4xMvUJkODf6HRmb9m68AZ6BjLAOzSCev0
oZnUeb1MG9/WFRurCHiY71WOAi/MY+Ok5EVn0okcGe14UNOaO/4k3TTaZYnIyaEZdkf0Bb58HBwT
CSSdevsDIF7TJ1DVE1D2Vyj0GtK60/uj/wlkYwCEDE9iF6nmvQFD0vRjfz1vDSAFGYU9+d33yWVU
OXmkLX5wkOpnszivcKBXCpTh9a7nzpSPpm6GqhURY+hpMMmLTOZKCu9sV7+M1PISmsHFQh+mimjL
5DLItlR8QQpZD13ovmSJgXUsiCZ7YmnG9A1ldU/zCPNw1kpq5mpH07btzhklngT4vIg1hCc48u+Q
2p/alp48XD+DWBuJodwtvudyhb9tOP6qfgemks5zUn+UJ2yZDQbATesatIPd1QJWv/NUeQ7zk/pJ
bAt159qnFXGGiD+tzTkxGaQCaKPx4e0AyPo5FDGPIMQZCnIP8l8jPe0306SVLu5J9oVaaaGDebsH
gAZlCZSmMOWtYijMPAlNLGqX1JWxNEdyWKRPEGQFlPnIaWrvREsPacQhVAxj3OnWunBcoLWeocS1
Kt39Od9jdde+8FqVMuqkgP9Wg3b2xXgd92L9cWByFR5mZiU0LdEVcexN0rHdPAZolzrvGK6tis7L
Wtlv3DNyVk2gn34Rw2/xIbncoGwAdYr2nEXcEzP+hmCqO1mGE4BKOcHa5NJpknVOyKVN6XtaRqZh
jJ4zUEz9Lh/LDrotbXXGeM8RWtL1+GmPBKSfy1gtkx/Bqd8VJtr1v+AHdrp8KHhLjvJvXvP8Dm9M
guSHEMDA+KnIa5xrWQSvLAHbV40RXgPeN+GS6mMdJiuNmcUGuUrWUJSlBSih/qayUJiI7n4SbpLC
tZ9JEIfB2bYTR7ajDNHpz6TNoUpwxvc0eBs6PsoucWjCQ7Fo8cMJ2IKhHCNjl/Q3MAIadQYAVrb6
KQReTn9+FCaCrU6MKBAaVBoUo2sh3PDVXBw0wi93fxwFLorMT8dOow+rAuH12hE9UyZ45eEG+oXj
OurDkdmqO40aY3o3SJyXEQhIKRKtHJa3eoykgyTneEzVdmxoAkdzniFFBhkp8xVOqCblvcIpSgLf
ptqeA4125S+cjF0KHLjRnc2cutgWaHEarfYeEpC7UeyzS7Fee2v9NhLzhjXqwVAsz7WQ9CEiEj7W
H3SQlmWcaIYY4jhGeYRqC07LPKqj6KN9BODroSnj5WRLyr/swJk4twbYmVugDqNCntewAhbMc0l4
yDT6joc7XhRAadDEh+B/8sNjMVFdBuudJQLhto/OOenoiJE5DZwTyClxxRZehaR99ufPMb3fb044
7wHUeP4gCBcD2v19/BTTUtZCeFUGFhJRZ6OvSghRNXWROYbFcfD04G6j8ALZVaQB3VAueEFPuZgR
qFBUqP4nM2a6Gt267c73CrlpNxXPR7wfOr6dDvZ/5v3+pXR/CJ4Ndxy3qctYje0PNYRHhYKjjbLA
vHvHthoPeUvnUODQyZ2RkLrOiA1LumZy7tj7omvWWW80fpcH8lLEdEI2aTQqXeDvMXA9ys1axQwt
BRbtWxc6gD2Mv8ESDC7qW8RlGL4ApbyJO4gHWhjaPyKXht9LllY5vaAyij638uq78VpoLbncxxi8
r+OmsogF0hktlcfs88x+mQaefUaeWphADuYCw9MnxoKVwH1/xR8A5MGV0Kmm7AbUk3Oo+zKnbiWE
XPZoEf+xujsEpwsmCA8/hiKdgBZmU7JbxR2eHN7elzfJUbrqGZb+XOsUKO4/0U0vGg2AMADB5Lvu
TELf2kWlGls55nAq4+S5oOq95AHnHEuQP7QjFNcm70v3vZM2KfOY/SexISrOOYrc3UMgRaacTuJU
3YpumR35bt6EuluRwhzimelkea0n/+OQ7wNk5lUMWRkZZnTW+i7YachSMQ7hYv3vWQBPYr8dDo9B
vPpfW9G7cJAWyCVVZxmOauSlP1AG07xiX3cMDbVGqr6SnsknSZeZjHSXX19bZcPeJAOdQEudovJB
dCbcV5fZPlOSGcmpBAu4O135Jk7w1XeylDS+Q2s5NAWE8D5H3Io/bnU4v0ABGmYKF42etaoTizV8
E+65xc+w5k4651twEjpTViiZBxQDisXdVO+jqKv6XxXdO+WvJ0FFph+PEZOveiXpx+cN8I6z3ebm
MgOVul4xkeC3In2iOOvnAiagD5cap7tpgETpuJsTEVRlW8MVGVKFja3q0eYTjWM1QpeOFro7QnRJ
W2X8NKhyU4qaNTRF1WlKG9gRer5yIX1BvTAfAwmkVSyMhEBjlerA9hQr1TaYcl0VjO5j74FYZJif
qhvOH8qu1n8ni0NnacSleJl7+z20X+XQmuhWpIkQ7eIeYX3IQ+OzzMQVFJMJTyuAQTWbkH+EmDj6
VlOUB7sn+5sV54rf5SXp43otiF8I3xF1ZI3fVVz9Afpmn8jti8y3B2cDM1KKVGQkcnNV1TNj6Dh9
pHSIK4w1LDQiUkZNbGGW7BurGBc6lJswuS07iv44Kt0P2GaJZJNmPp+GvpcGb2MLOkXi17xqH9jL
p5FM5HuBlCvsYzZx0e2A2P8CG7EluoIDs6pfrX3PktP+fZ/8Bpc573C7MSOfZqxLehM2dN1W4UwI
OZD6lEgqex5Nz8FhEE1Al9chHUkFPvIb+p0tOdTV/ka0m8yG+Gcwb+TTUchdwiFWlJ2s3gEtOqbf
Q88LrJtygQajxxxoiijMj8P0NaP9vLE7RGHK9bCLfICWLupNhvp0rwW0vi8d87Q9rblnPdl8U5Kd
1ciUsHGvLQ8nbgUlpIpIEXJxFO/NlBFkjvWG9td4WE/iIbg9RE2rPeg7KfDQmHI5PQdzq3nU8p4G
SOtVClcTaCre9BwfnPQ9GxYU9QcR39K7l+3UJljT8oqhdaRXB6hkP5ZQnp+ajc08QuwnvxtcSPYx
+GirvSDifngXZGvaXSr+b9IQVHSAIjZzxcDA8JbH2DN036eOlXw0CbitQbbo0gMjbKoWMWqSluN1
UU0Id6j3guVoz3HKM4ubgAVsGZIK7Rmhoi+ch2a668PZx/V8tbZT6l1+4AGhfrCqcvIGtlhelz/1
/ASEUVlQY3MzU1QknD2fhtwCb9I2Bok2Jm6W5dP2tvkYn90iGPcW8pOZCED6ov0HpS47bueBo/mh
+agZo9RX5yjvZZZ0AZFMPSSHoCdhQ2MDHUX55J4oNhocCcfS7mG8H/gVPcipm5Hm+J564EakVmu1
XrqrJCk6n5V6n6C4Xj+xzg3pVi6LUO/20HjPVtci1N+uNoxacdwLgicBfLgR1LnLYYz2A/QSfLm8
W+WvuQVnjR3eRRlqMHwLViUf9wFmhTX22nUyXiIOZEs68/L9L6wv8Ug2uM33ryi81YScn+4RTFcT
qNEwTndbtLHnKjzP2YlqLZT5rCD7wSHi1SPITCAiJ7oCkpJTdxzNtSB6qGQFxhx1OFL1qnGhzB6z
LsdyTOUMLD5jZoVC4z/uqd1K/9L+Dc7PxnIXaeywtxJp6zrkPnnLX9hNB8d0YxuiUMnpIYwiXIqW
rXGGPsv1mUsL07m7OqXQEDM6M4dHkDoR7a/8Rc++FA6VOw/EZq8Z5TcYc721hHEXnrnfKIhyP6pG
uoDJSYSAxyHG6RVrtPpxb8TATlJn+XV7+wY7VqsqSeCQWtAzGPw2uZs9+QQGln67IiJbmO8CEPU6
D1CcHT14QlXYUTjOPDLoHKLx9XHjotsFeii2MH4eUuoRJhfwewk/LPi//QaSA3zBPZMs00Tgyp1h
VyCR4owKpTBBo6e+UoZ6ofb/PX8IyOp50ubMxywbruWMkjIjaUUYKoZIwcFZxU60iVgQWDYQlvIm
VhY4upLWgwPMqU7+xzpiQlXepmZgUxfDs6+F8pjHh3WmRFsW9Y7UyV1IONPx0UtP3ouNVULq81aq
G1m8yKmDgUXkUDC1vslXy0Vrp9T0R1LzE/R5OujBaZ9+p/CPKp/a2oHlL4IutvbqbTUBF3r/Hcil
33wHAIPL+LkOereSRam+1Ez+Oqg3cAk9D2P1FrE5ln4YH7v8IJW2lPIuUEdlgCE+eq2xxypWx31G
P7MvXumzCTwvKIazLfX5uREm0uwORb/euc/h11iiQO4oDiLDwzfv405mveMpRYY9CoCqUMOjZEIR
Cq++Yvt2lQkiVLWCESvloJi6p/IiEqxRiZj6tao2XAYkNlC+zkF3CnxekRg9nKd1PvXPOPwdAd0v
uB9KqX3DnsVYRDVXt3mdyCL9ePBcJvTut9fxUuyxTdFQ8I5kcdTKjnhQvY0ow+gWNFf0aacV6eYb
jJ5MxAO19pXtl4y5UTSE8rRq/l/mPUdbfph4JlkiP24Q/q3XSGFSWxpjvcjvT3UXZfFPx6twURRj
Xv0/2GDMBWTcDfEG1+JTtPEsGbF81QiKDExdCP2nS1yvhYNH9ejZ5v90uykvrMQ/eUevrclwoUWZ
3vSw+HfzHnDuUR0IMYg6OjY7n791VHXbHVJ3nu+7VXJIRYUX1GhkuZH/Z3Gs4tdzAzW0kWXv8EbA
ho5Kf3OQ4eY7mTNW0M2CSzz8heyaZtpIf8NyFFzBaVknyIGFHPKPYxV9jeWTXc3/t/qln9CRtY4E
rTRpNJNaJ9OhGGdbMPsaTQZePI35aNFAxGMvQ3uujrvyquh2ht9uyrrTdq38y2a51Eggzc6Irb5+
ENAfWth5BUxf15NZoKa4NyPA0KoN5a+XAnB0kGy8+FDJJ97ACZbZbe63JirmUS5gyC60nrOx0N0o
Y5d0/XNif/UrsDvj49moTLK2WSX8aXNNdgjV+n/Y0XO9pv8sNV9ajBFUtNdvZJjhHzz9GohLyEg6
+RYZ/JNcmXeGIZU6qDARVgn9tposbFgkX15afDu7f2o92rzbZN4Zhp4Kf4z23FzV6pP0TvBybvH0
+q6n/FRY4BotAjwNNVYhqWCXgjPD+mmY+8Wf1ezxwBo6mSxm6tgpMgtkEznRxW60PX9OtDXRkJHA
tMVcYjVpt0QFTG3ibOX+Gpmkx4RoD5ZWdLzWUq+c5z74ffn1yJ5n8XgcaObewj7N4+gBEvnSHNLJ
5o1XEQIInJ7Z/exblcB8Zf26omHsF494d1eshhNp3hTjSrlxxWZZ6dkFE/rYCNmfJYgScfpF5NWG
UFx49yxaX2BnRXrDrl9F82MJeCIZDf/Khf4ZyWMl1pOYPvyE+dGOol3qeXOWCRx89u6fe6PnfFAV
wooSK81ZMrTp3elQmuDYyLQK9KFePxTd3PgRu/Gs1Z/8um0owLXphDaPJ+IPRtVT1akC5DM2+96E
BDjzmFDx0vTBRtBlhRYyC5LY9Jw4XBi7V3Xf/JFsM3RxTdWyfYLD7RsLDonhmv5glez7igE2+CJA
5ZptIGhGicCi5J9hfpq7JvhHzRJ44gx2RqOwuFF/FdemM9I4WnVS+g2FIfjyoWH9jd0ExkZES+st
YTcuhnsk8Q/hd4DmrsL2Gq9x3RDgwCuRYFRiWJvi6C17AGqJzbq4zCoj3dX3/1js0VMZvgruc0g8
19VN2XFpuY5sth6dWrA3ZcgU9WLerCFDwDmwcrkZYx0QUDnpHwOvhfFJ4Dizo/H4SY6q25QXF47k
ryqFazhBX6qvAqas3SMmxvKiKzQlLetZAFhail0Ex5S0gQG+mxFharj/QpYqs6EzqMmPt4cwVqzR
ShcQ/YnQYA9txLJeqvrK2mID+wFOpi4FP5Lg44QWfO70XdzZ1g+YhODMh9bXMpjCJd5dHDb9zu/u
5vQO3qXjNdjFCVRfj9nColzGfD0nUJwjZZS+ndYlB4QlF0veWYcNtjaFOB62cZaJBmjohyvBDtdk
3X3CyiU+q/u62bbhoykvWwLAW9GwefyDJWfA8WR4VF12zZEPi0LGoQlTTxWuTlCuZilIgqU1ieXa
TUNDsZ6Ibil5vTqP6VyXDts1QpQQeYLQ7HbvrxwI6Fl0+i0uMlhz27e6R8DzQUzd3JYamy74lXKt
HylLKAQwfPiNA+A/OgCUDu2zNLmq/U0qyxDyPcSpm+fIXnF7e4DY5gQHCINpVlBwPp8PYoJcfUff
yuZPZWfFsi8G/FJiR0jrbGaAxwvGJdbViC1llgFjOiQDYns05Jv46YF6AM/QTk087V5giLO73E37
xxOiLOChnbFKvNqbWaxvQFIUZ2DlVCd3HiTM53U3OQi1JHR1Q3cJxaDM89OUjGTR/wyujQyaV9Up
2D6JqAgzJS3zK4onTpHuIWRKkNVGRSg5CVukprPUrgAjSA5WY5FpQCYTS6GIJ6e9yhelWaRbkWW2
PuOsN9BVYkeWAnbUtGdIgNn8wGD5V2WQQmi6p2FkApJMvAbszxdbsp7/Tl/EotkXTYp4OchGzG63
1zU9Cq7ulroi9FU+4+xA2Vg72JOEa5bp2JAImbYzrVuEwrGd4/o6hCaJ+ynmYkN7gmeGVc6TyfL0
qU0CdsqDPoKJ0mA2la+Za2/mfvu2h1BEi/5CuZr52SLNzllH/as/TD4/BQqE0WuWvWmTdWZ1lOSN
xnKxpbFkCZcCdfAx3an8ts7vzYvsCkqPdz7VXQIp6Z+nQJhjMotAzmK8sAXQ+i0L8GfFw+12Rfv6
F5O7oGEIQAb5kEAkC46eB9oAyGQl1tuJ+REwzMhNXrCQXuiw78xhi/w/xjTxTR9JA43mNWwJZIKZ
M5ZXwZFU7J3DO6VJclXbSiRRNIO0PrSZnlvYCX6OGpxaCVwnSEl4hRF3centDO/ZAVijVkT3UlSK
iEMhI9LGuISiEqPUKK3nD4WDbzDUGXwGvh63HRboXC1b37ppqnPtHUlfYU+YY6UqSEOkcBTkN+Gr
rrs5GRjai7GvR2QvfElMiuXft11T/wsueM9CpmEFkJdDK4bRXtqtgvtbfza84qbiqhvdcEJjPSNd
l1pMq7zBi0guZXZ/P/m14cObJJMD30Kfd9Pv1lPPv1O0E50s15GGUxdZl+0maf3bqC17+UZPgfRE
pjHPZwJxg/EuQksKdDZyLOoSYt50D0XGzSZTiGYuWerBhBb1JsepZssHR2B042lcklkREoXZQnA4
mNzBtLgB25ciV9kOUFQsnwqgCl7C7FWnLyEecD6Y0UHxaQzh1obnjDkDJFAEdnuVMfsXlwqOVw3x
blbH2r7iTDKhKGwgr+HG4XhfovuILhHgPCOIoA5ByGciSfR637N94Npm0KsBCEz4QqAPBlKjzUnQ
VQb3iT3TEqFKb0tXE/DEq1KnvUhbCNRCZrOWUfJ+pGnwyxmkw3GeXM4GaHreNfDhqCdWDdvjbk+L
Ha1X251el1u5BY/QPFIm4+AyZgMbkpQHUrwPNeH0LEKxb6dx012LfQz/4kM0835OSpn1AjRXOfSY
xcb8P2aQvZaYdT9uCD83oaaVUGC0YcJvoGE+RmlYdAJneKxM6QR6dWrpgdhXj+qDCjgnHYAeHi3Y
2nIYQSsFWZJET/iImNyRRJyRiVutbDYrXnZqocxg7MHDkcIr5rHkyPZ+FV8NXSPO+NPsPALIU9qr
DCdoT99w1Z7xTRNPGjO7wHH2H0vx36wGDxwVSWVPdRvxJYFV8WFHeDyMosZuNmL4Njmkndhj75+H
7eyR8FRHyzQIVuZxREHsEWbAJq0h68oUma5Q9fIW/0ikvhuNXHn85QxhIXrzrhQNFLEmaUSCQ8Om
ZlPp3iwGu0C6Jff4WMS0LfNUgxO0z88Mu8UoI7bspKXDVw+925xfSeR8m/NNtWN39952iSDuAJ1q
uoRQBMIQFWrPJe6l8b8JFGkSL5BZlqkp9aOYEsz4D92ZHV6CuQYA0JC0VmvARHu//ndN55onmS4p
1CInTE19Mr44ZyqRfGBRHN+3g09pgnGT1U8FDGvZ9e12KzZle26wzgaj0gULIHLkkBymn/EzFEkK
U6SfdXOEX+tV0gLYKqwkKkRtMsGYvxwi8EOT+jCWuWPnPPwJHw9tduDu2RSfDCwyiWfZiXn51mvz
AWSCtvQSZHSsS410VPqmpEtGz+PuCsEiphed+yGuGMqmR6tqtn8rWHyvHTBoqLQOxlEYwSEgL/19
CD2eTIVni9H1ypkGa5AlNat0YuTENk77ptlADrP3aD8YUzNR9p3cGEyyr4zkA4yueRpavaT+5YvO
KMN4O1fqyW9yyfxQ/ZpIZ//ZzU4anFbxJNKF2qmPtChQhNpvKLZhT8yXK2WPNoF2Zo/rjzX8dNux
GKThsta/d2aVlo/1T0wV4RQ+pxSmpeQN61iuDRDhIW+8Ft8PV3QXXGsb+8xmKl97CDJF+5SnFzot
gejx8qfKhZlojpFNNAVpKwwJvh91ma34C7co+tYfukUKwuqB5V3fhEXpXdN8livthLk/Ctd/a7n7
2x5wpYwSppVLCcLwL0fx04x3JdbsY7kvORliNaOHDfImiAIhBAnzXQtDyrYG2Vp+qXHZbPEcyDsG
R2XR/eaItkXeNlPS6EmkUTmh1ouuKj97mt4f4yvIhwtwGLzF2nAiBANcZHa5JSiZR2GiSllAWgB5
OFJ9Mo/mk6ikF8iEisb/s4HpwGQXStboLibGVvA9gu8oE/eqYgHL+Gm/QPLNlQS/IVeaBbhXuO8T
7Nh5gNkyxZPa+ShusIWelY8zxpCvrG6LciUQHd9nfIu1cP23zyl0ZxdwTB7o5Kc6nXnUp//LsHPh
99xMtBpeqoQI2mzwM3JMLMqYKbKCpGJop7fIumocZJnYd3CgrQKPQmULDTh0zu1MNsE9FiAV+y16
U6DsIxXWtaNTW1vRF8oIl2J4HaTFcO99y+5QsuO0zcOHY1CLEHnhF01zgDbBCHbk3aUq/YvUjOwy
VsRSrKhtRNss/WnYw+tp9HJSea9HkHDBpcOKk0kKclYPm5LG5dufRqX/2XNDMPqMFYyLwMBHAf2z
Apnz8NWdD8rB/M5/q2cuHsME6hsjQlXg8t3XfpXKR/8IfDQUvkbtTq0xfrK8yHVZfEzDMkQAaBWY
w6WxJIb1kPHkiI+qrkrLiYNlOvu0obLLxPwprRR4+S+y76hL3Iri6QFqyRCJvJYtHanMeh4OCWpm
DUwpICEkn2U+T06GfItuSNOi0uv9XQZVLIFkvy0sH/KnCcedYl6qkjET43LYxq7Wxt5ysm1mE3Kp
RRF/1ihI0U6xCIUdrfwJH9UZZwqIx8In6KhyNSmibSemdXOF2W1P9cJh1jvzJVc01AZXrXZAmiLo
O/+Ko4+MCONR0YqVCokKdxNiHpsZy24OCyoSIpeMeA+7vn0yN+ikIUXkJneJx1GjNJ/ovJ2DMCpc
PSC1X7SM5Zr1oMzv3ruH1t9A8V9MA3CzYyTgbqRI8/5IiPVdqYZZmJjwdw+hGt1H88FJBnhULj2L
T9OxWDXHvmXHOSIkWWoOLhbwj7GhSEy9tbDY0kKO7S0wrSOSTTUr2WKmL0KA0VAHSeDvHGtzTrwK
1g1PdfYTJJim8wsKwmHCTS9jwm9QsSC5++1Kk9s/5OEuUz/Y319PXdGO+6ACcuKNx+VIrjZ4W9+g
iuFuIhyIyXzYmbnR9phqRSsSFlALGqZqrbpYK8Wt79Um9B1kX2HZ720sR9IjTzRFWT0+XTi6IOkF
46tOC2yIJcs/OHiAl/zP7f/ugcF2KqxyOaADhJEBPNWW9Gvr85m1zFBP7MdE+NSZwIdN4wedU3pv
3EssEMoPc+WjHKmFOCt20HKSI0KDni8ctNzsQkTtUOXwCGVxIxYPY2VWq0SfKI/TxFM66Ws+PsiD
iqMnFyh+hSlzfMMXhTrB2sezaVC3LtXfhszSa0AyKcwuOzWwL7TpXGUszjiEy5irDcUM3uVxokdV
06skgFNJLEeF45cCExIZOWPFkUgccKlXsYUXPhNSPuye+JM1714cwWKRje4DrwYFRdx04yW9GeVf
El9Wt8KQ+gLlBeXDH691llptRkxNrFV4XZ8KUUkXZ8EMbbCq1KFeehY9nKsOAy5n6v6w3JawejD9
SvDrQW6eVOHZayH6MuVaQVkiEcExg0W+633g5Da6XJU2ICuX2TEl9t9bKjWyluC4ooaSDMQSVya8
ulzRDCTtAIaae28zAiSWbQmrGF2puHKwp+177xFHmQe5i9nwTK29K1O9RT29F0gkQnn6ZEfvJlLB
36w1Jh5lgZnOZtBn5+mmcNwPGRWOelUGQ6x6QlxksUp8CSKQOwOAf6iKp00flvH+AW2Oygub53Ra
WlW0ZnvEt5rkgmuD/7vu0OUk2FOhjqS4nGLKDkQnr7dYUMpgfy1PLt+fp1n8DSULZD3VsUMnx+J4
D4GbcSG/0G0/lq1hHDdaZkIPBF/ArXAPwcvx3mMyJtaVbotBs9qnnF93wcw3j0SZ8ZZB30Bvp7Rp
YhMdlM5B6vxsBwWuWyxgX26hbjt8Gtcg72UUuKI7zcGpX4rmSJsbR+Wu9L5C4ueOCNmnAoqBdyMo
s+xgEuekg9IsKcJzRrDT3Z7n2dbRYbZqrPCCqilM/kmLSynQeTCxaOFclt7aXZJafGVDgjTQD0SC
2ZpyUAC4Vutm9C6op73vi9IczkwbJOQASAGWFFa5eA8yCBzBaUnrkY6RshkfysWQJ6pkKcDQnv37
7Lfiw6I3DcnTKE8KrpNZGlvKeloHwZWASz2HiGnshGfNZhotkGDQIxR2DvauLwVSnJpS+TYpnOt2
+36jbqNk3NoBvXH50QtZQI6IdzTsZdWJLa5exPc2noJjmxD07v5CXpH+QD0WcSocjRLBuN1c5LoL
r1ZLsbNXrPGyJS5AvAmWeQRz8UDqwbuird3cy/QjF07+EbRUsGQ1I5Do+jU5TrzXvHmvxX82jHD8
GH+b5SC1/h0HHCTLvDVCKcUXo+YEdzUXzTfHbgneSp5xYpBR4kHbYx83NhlHmWbByFIzhuzASwOZ
5wQFWa5WbpFkN0zmqQTEvL028AISwr5QGv76RV8274SRc78CwkRGqiI3iTqBCF9jAdaQJg8Ohmv0
ZLzRSso/kvDQTh4ugFjLgn+kZr00tWlq/TO3TTYY641ezf89zlo3yNFO0MnOEDFC/0zphBCMxSx2
ICtGdWst5vs/ahDUEyzDE/zWt6dYAv5lBuf7DdwhLhHC14PiI0GJxEDc+5ziwD7Zfyg/lufD2AdJ
3jaf1JvmUJC3+0zm03RvTrn8jh7I2MOmRXGMIbAJw2CeblGTBE3PTLxQFq/xWNF/GquKMk8KytDy
H63RqFZdjgNbAA7iRcivnYh4GRzxOoDDFTKmw0Ao79Erv2ovZRho1bsZpzzGxfuqA8KT1rMWmO+i
fayR4/7Lr4vSPGR3OJ2RH8xBsoH5/xpCida3cuaCzmJhubKqGr1+cl3ECC9AdvMictQi6jB2/jGu
jaakndGBwHufSRWDn0Ge3kI36sJnQxXckf4pWjDTDI92Yjc1IJUeI0aQksbjdpc57RGgJMgIkXZ0
oRsCfZ4GxP7/qeycIG5PNrhJZpq2QX+Yd/x5Xj8kd5iB4RySvLgFKo442UqGkqzvtH6yWU/zUB+W
tnZnBedolNOvSIy5T7fa2yxYCDNlZVLX1K8X7WdFKi3A7kItVnklxRegw8p5+6lTTpGmI84ZnZTr
3e5aRlMHKZBhDffLhd/lwV8b5Jc1pyCY33KzOh+8oUv35DKqXnaeYfNYUfG7gGMwEeLeiSxcW+zd
+IzyaBDSoSNjNUUtQqbxQFLMFh/ReFcZXXeC+kTWpcWIMOeoF/MhWeKQWSyYWvIeS9MWn9ZWk+uI
H9xe1h9nZGnxtFFGFU/yAJlJtG1qc6PJGB5ySvDSu64vXVLdgp0Erg42lgJYeS89C4rtjQovKP1P
c0UraamPp5rX6qM1+dqzKdHLDIgxd8W6niIdzbqHlBb0HDt71F6ePv7FW2+itREz95sQNO7d/aRz
TzSY837XJG5unutEgKSm01/IERYNGI5F7lWxy+9PU3wcdvfYcgVOJq2JnRtxBgX39g6yodw6g/Yj
xDQcdUyyyf/gEuPJ6boT74JmO5r/l/So26PKy2kLiBmwo2cPymVDkcw5zgHUIncCZXq1ByqpdqIF
kPC4Mrk4+/MeWsedBPFPsBeeaAgbEgDqpD9mjRbXfKFuMD3+334AVtUJuyk2YpzrG9X3erd7dokb
gT6cIvfSGq1ALN/vbucgBszM4kXDGi3gEA6ipQPGSI4xxsJAHdRbHFpTdcaT4/Tzv/9jfkEXz5w3
9rcdMiGYvFAJaD59RFTsvLCbTUeDX3HhsNJ4qtvf8Xbc95MWHQDkSbvVOd3M4eaWTVaytndjXhXR
dzuzcGam0prx0sz9UmQ58D/Mg5tStl8l5euckVsek1N555qMnKzFdsf0dCHfZ6j5RHdOWS5InaCg
GRfoOB1dA9hnW4FgBMUKynpiZxjz5+u6EpXxsCWGL8fazY1PAROXm6y/ra1j0vQPAmfhp9G6Fxp0
S4d8d+Hto/J/OwRC/874NLdcXLwwNcu511KchLrQaMprG57tkHCAK4KuKr0+xaQy6OJyK3vi0XS0
PmpRHEJadXq31PDAu2S3UFIyk6neWI8DCgMEAs9z4zNHJ6+j2dStpP35HOZ2aEgbp+1Vn+BL17yd
Lh9ts1jPlKbNhrIWLgd8UtbpIdN//ne+H4wABiWy5Ra488tnwXlXKHKogu+iH3BvbAbmoLexbsVz
PwrTE83jR1e50PvMixiHZ4FnSrOaY/sXxwto3BdSSiKHC9vAH7W9O53D+/r0WtfuikbF+/dT1noj
Pzc9NIsaUc0PiV5bvBwe887yaBj03EJL/DwBWmq44lLUnKV8b+/piJkqPXrmDU68X/lrAuI8ZcXU
pH0L76smhsYdsXM8DLvIXq4OMsIbB36Vd9FMHeT4GprfegUgPIiJwnNB8EIh4mrr144GtNW2mecK
Kqw3Qy37vR0uyy+knUBiV12jdIB19G2gkJqf+K7Ow35L7LaCwiuxpqNPpcJqLmkaCvB5JcHQVSeI
pDPQ4rka+iQs1+uWDGPCWKrOoM7DEp0ti64Locd1T9jnAryamaLlZgsGow/iZz375Tm7MLvR+xpQ
tRiz10iS9h0I3jW1SaBbbg8J2CtE9pQXvBApVh4+qB3j+iXAcKOYiQplF6OCAGuAfN271Ags4tOZ
bNwF4sQyf9ZSzQENgXDQcd389H/bkUdCgUbQQ5+8BFYFWcFFwIHfocpUIShAGHbGoXI+1W2tGikv
cRMnQ55uZSiMbqfws0xA/UEeMy16Sf6bwTbQOAdhgC4ux5FJvku4CkhUcPMoWBZTGLXTlj3kBNK9
zC8vVs7zCW2TvXiobd9czSa6UuGSUChFkRWsC5f7OLLKp0uuV2wZsWlKBnziZcO3cAfa0a4RH0gx
dZwGgDePL0Njm01TA3qRLDSS0uFrxE9R8JWKeOMkK63TH+4aEiGO8AvnFlhnHHMTkjbeXhjoDocl
xpkY459V2ZH4SH6SCL4SXHduo5T6KSJg7Q6W/kPo1McoI+cqiw2EvTmds01NB2qx0utuk/P0v6uY
rgz58eX4LsADHN3/l3DwFEvOE01QlwvKEd7vwFJDvpIYsqJjqiSWBXMTEJZI9tVRpnR1Lv7fcYg3
BPwmcD0L7A3T+YGXdpKMeNk/F3GJ3daEhQ4kcZNv+vUws/rUoid+lugDWGy26TtbAvewEU1xVMXd
vs69TU//KDs+DipI8EnoDdqWuHQClZqPCxKot6Gy853CIgYLIOYUwAGpEyIsd3FK0MqngXaFbFnj
w47KD/D7KysO4I2vRXwXoBCBUFHgf9uupzOzMXa8tUI8fhSzTe1YY5hUuJq6Fs4RU3XDlS0n1CLm
pqn4Wb1MJ0BeaOb7F1KBqn7euoNuSRnYy+wXO38W+m3EjhwH4C05oKRgsIR3BbQq1KGI0ac+BXeY
vWZI8ucMbSkGIT9YkQxdUjKOnNXFQ1M4alxRuHPbXyEOjO6WT1mH/8zwbdcyVeBJY3FlQrU2w9gf
3VXNTcrV2meKeul3vN3VaSuDQpeTM/jj836k+8WRcSQkJj0EL/GeB/wlXAbKlBrKCVhMqSiwG98L
mPI9eSgwIv6AN/ANTyYi4p+lF+tupAk2brFAIaB2iHDQpdZGCt/xdxDUX4n3qt0SFKuKeqrbs5E9
C4RAgLmQ/Fo6WmVZORrho0NClqNc+gPouz3Cus0hwxOg9ggBDJgZwq/5iw2PRueP+3OjHqG3NlNc
7h5iBdUrHGQRBc7/SAcnAuonAwdvRsgMtemDBmvsublmwPvutLHJgA8GsYqU4B93xRoyjWQclFvh
YM2153/vwEXXNHqj4efhKvkq8vHNbYOUr91k0ngXxTMsgWRk59u+vkdLItRv2wI0XYrWpLze7i1z
46AYXBFheVhFjHxdWYXVTuT3NB/vFJvnEhhboAR1vTmBjoTeu+Sdrd+N5BEtdBuM+3RBTfpqX5hk
X343u9Qe9c2U3ws2t+Z1siVgiYlPG5+u1+W0NP3YxLkJYLxAlklf/DHOIKgqGJnPKH8xHUn3y30G
Tsjyea810X1REDnXpq/65XKSIf8UvsMBTFUBerK3ZneLZPDUJwmjk9z1qMhBOCXJMO+qhPE0QtrM
D9zPKi0vUgQGrD7HvjwDKbv5hEsyQBJSf3GLxirKVo4eZbaP3kUuabaK9/UyfHsvRVBn6VI2sQi7
YoOG2pOegCopt6flhWc9EVrIyZ015yva3SrwafrvsBaPcDZExc2KAju2tB0/5YU9WSJTN1Uh4en3
LRJoRZTEoQSFSomqKBJZaQ1dLwiTWXnyiKEiRhG9lcHwZzlC6sA/riG6WOvjPS5tQt3ajkfCYUhG
6TuB0fbImu7vcceKkqqQk/icQhSmagdstwZeZEhDItK7HRuUPWyzHPn4U8GaoZdgZUuQhnc+pzGk
jRa8Wbj7KET5ZTBxjyodBzBThLzAlv+KM8FsuhHAGKX3XO3sfdLYPEc9hZ3phxdVNCUMewk/7ME2
uak33K8f1nsGmFP2IRKu79PZNP/foqznrWrh9qUejjGiOh0NL7NJWtOof3cu+7njbBwLE+uk0965
sVVGP5i0a9k7VmSExwnM0ba3kSUOzkmuvP7TL/NNPhKiF+lkKU/ysI+VoNvVYZxC5qLQQT02KHVD
1x6JdIbc+rqv829XIqEHzuS9Uk1k0f3IwdNVMvmok/jNIgPgQq73A5n1yvDuYYPiHyWg16pBG9jK
gPXbCrOwerVXa8lepnysCkiSP/2T2af+RgwcCEcg7qqnYhfzH+ShIgySgT1Fha3Mqyq2UD3gyde9
ys40ZF2bTVdsqxeuBqwdvIif0MGnJZD2TTIOs9FI97miY+AuKFs2B84YkkZqRpTHYsh57JOCKsBa
P7um9vcw4mFZqLcIRxrHLZAPtMckNUnE3h8jA++V0R4QWkaCrk5QXtpjLhCB7qWbUOBxDrmYqYRj
HIPI82OlFibKUxHW4Zqqd+EKiEr41kGQSu92b7xJKDtUkGB2NN6sDz2FpnAX4qqJV8mSilgJ7fqG
BWFSnvqZPJKSOGVaSKkjeAJ5NEIIJXtt8qiapTK9DsiZc0psJLMIweVQ3B4gLULlILLhys7VGe6u
RsAKfeAdmS9NQBlANx8hcNV52iAPF4hcPALGxQ/1zbJBBQDcaMVnqpW2CwxBC5DkQ9RJQHZerQiD
ayyIuLMKwxXq+UJcpHCCfdTZ4CieJVTaKCP4MkDOK8yIi+XYJ1RvAM6Bl0g0I2+Ysz128qpRFcie
lhP70V+itswn/miJtXuSMquAHjL9O8LZxTNtajsoiPxYzd282Q19jskGshfWBNWK3bXBvJoQkcu3
mNooQ9KxYc6y8axQFKgal8f98oDudKVkyrrZSbygZnuYOHgv0hez3cGfVjjin/YiRaz0ACw7LpqW
UEU41XLVQiUTLDYk5BCx8LEciDSvBSPDHl29gWmkUsfXhu4JWTHCCF/TpzfFuXTUcN2jLhGGV3TM
f5YbSVzsqNtEopErKTzP0ZBge+tEHdhTai+jaLYsUezs5ku2pV4eaznglli/LAR6LT8rmGANVgw4
UZbgMTewiZyKWJJfMwEkaCdrV0LhRQ9vmmHPryKu8NLPd45a3FS3X3duFrmQcrwTVVgAzkmHcsRt
8O9hURKkzuZnYWnxpwdfQdfUzFPwa73MJ+bUYwq5lNzr+xXlUKWn6QxJ/xQ01yJzV9aHq/rmiSmG
Zc29lq+MibfFCC688ephORT/WBRUIKrbNgpvuBTg8yarKo5U+Ar/BJZCY8xBoVwES+LEc3s+ulRN
+lN+Ptlmg3QqI3D+hF79zAlx4a9cAsxaXkszXk5TA+FOKzbjxnrPDRJBfxCrEFQXii+F+Ddm3uva
zy2FvCYeH76hlZm7eU3ayv6s+N8TXE7CbIxh5lM+EOe3+UBFETIMyqOW7xZ/IvxJCBIsgouYgJym
cP3CIksf9LLOl0YCMoE6VXqs01Ss1Te3LZWkBY30/e5zXaCe3TUDWbM9Y9RbNp1QLp0t7XrraZbb
T9nkwGKAwPIrCZNt28j4bEyn/AFzHqhk0tNht6twu6AL65xI/ntWqw1SxdG3ke96cpzlkFQNcSOm
PTPOg0xnuB2GKu7YQioZ7bg8762xxEE1oFhuq98hJdSenv5N9/RFX2Yo7X8e/fvxn2IB3R0CDKsi
inRyWzo+8jhkENfmjL3M6jsKyszG4Rd8VKUBX1Qo7HjjOKPw6tdYLiWMi/5z2lPH//Kg7+T5Le/d
urTunwJ2k29nL1xC6Q7dAs3C/lGfvc587H5uIbx1VEnMmVKQqvcLgmYH9Lga/KhbpqJShbfbtaFt
uVhSlnGI8JjCaTR6A7hmlthRaZkoFNxmyudZijmI3ZhD9sGDvhFxdqEUyLX0lrC2v0wRq4WnLwZj
4VOQuqIniF4MYv2j2z8nn2N/usH3+XnOEslyNVG+3N6hVQ8esksmeMnDfvn3Egob/tPrNNoMGPqp
3VsHN7lTHjHR65yRlLaIyXaG+ec2Fe1utupXzopT1onByZV08r9iBrFb838Ef0fpxGNMDmHQc460
fs0lH9TYTJoq6ibk9qEoZW/zwgs6OILJXtP6PgmTmZ8zPvDlMUbjn8TxmhxJ+vGb5UTtfcpMu3C8
uKyaMyZEzUz3+QQM7OwZz6j17J/UDZL0+IRAXufWHzbrj+3DSlaNhb6O2DGzBozIJHtLmjg5s637
9dz+/dfOgA01i5I6Ci/Bf/7XX0a6mgD8iuYkfCJS89WRT8on0peqA8HKiriGQg4AW/EEJKLiaS1T
aEpI7Ja4SFl+N2ydHn2ZTAQ7Ts3Fhb8kJj4PIUUPsD5wF6g8Idgt+ZanjCwR8RxkZGRtuSWVbYRt
7LtXexsfeLpetSljgXED2QrUbp8OgvjGvcZizTC7v/JnfudQM5CtHRJV6BmfiHAzGXewXk2Jg6Fb
I03nTgRD1VaYkTdQqAjbElxs7XxCHetiRz3ir5wl2vVimwTJz8zeoh91q79xvdzEB/vLe1koTtha
AjOx4nXcaIKWofQUjoPSwkv5a+HcWoefypeMxWLlS+Q8DvXFH5HzA4/Gw4YJk4bgipcKIhWiR1Nx
udwfCmM+3Fpln1vBGtdGdCxyh7NaTDFYJL9RoY4s4BJZJ3ki3a6donRzq+3SeedOrbTdbh1M8Qpd
BNI/tU/4CcNdYvvLvHGoC1hK4O4hjM/iQUuq1VSGLdY+/AMRVehVIQt5cJ5iIVwt0UfeHh9opLLc
4asdJB2rmUdp29d5cUaPMLnZHXMfSxXPFPX03319xbBJuaScACzLhENXYhX51/Tr1ltOXp+LviTw
70Nn9UXCwfde6DuLfXuuneB1if4yw5sJ0lKu+EogbG0cTmc6Jb8uzmPbFNcsMnh6BR6C3bpRgOBt
tApEJxy6+HQXRLNC2ZLsr8wmtFp0saLunY9v83I0IQ7zEwhv7M0e18te8v4Mok1i5uVB6w4DARX1
N2z2aoeuQ+CV3t84WzLsJw8EBHuOS6S2S4cQds7XQVU8hdM4aSrcdUcvbrTStOKRvOfvCCTQqVWB
ilcVEuJPSuEgaLt5o2krGfFXRMQ70sWnhOFbLxoXAzNCEn8okMcx9R8U6keixoXqH9rUDK4ZqKf0
MKVUxPZmHd4bloJNnTPU0V7NRiQHxMqX2S6IitIGk3d7JyZl4lxHc6juYfcwghcIUks6kSRKSozs
cgCsnpL1gQvng27N7TT65qLDf+yVRxqrfBiqbLEjPPv3LFhrEc/p6k7i2WiqbDwFeOOSgchPzLe/
oT9pOfVtCMKBdrvMcJ3sYDk9b+sFsalms8CAwpsMPjRYi62wsfBVrD89vdRCHZfNy0XG+lElIyrg
Kd+TSMvfanzxtItaOrOTqfIV66sEex0hTUVw6jLUoSZbN4DYg6IsT+WRvGiIoInlw7E6JVJp/u+w
OMI0pGcR9PZQ3qxxGRWA4slQV8Kcb39V294krrYeDlN/D9gZ3soaNzNWmJxqo83KSjDCb9kEk+Jx
YQROVcLWpyArXfZjL9QK8rQjJfV8nzYJTXO4ly30Ag5W+PPHcmDI7oJCcu7GFzAsGMTcu7gmpIaB
0NA99jaI9SwaPz8jQE+NDRP9uEPWLet4MkJ3D2WzMMLpYdGBEcNwuYfburNyfMK1GEeIgNU9nCOl
qaYqPKItqUDXdDs9bXNVGAJ1vaBps+xYSAjC6PfxaHBKXwab17UN5sYwBj8h+nEbdH2Q/tKziIds
MlQq5KlamBG7y5m7VIoYnioIIFcl7wEkh575M0UZfDcmqhOkcll13juflD3nBYuLXopZteNP2dSu
zONHjTHD5CYlr+nO2+Srd9tyx9f1AUk3WB6qnTbsVpq7hsvEH8xUpUb8zg7bbh5hHGGnAjXWzr6U
c3zSOyx7xXrxqL0HPTIM4YlfSbB/K3a2wjw9kIQ7pyCerbSPJOLdi3P5DnY43+yKUGEuDDkne8qh
LWsP/bqJdkgNQvHfdZ/rL4XAIYby7ivpEtjEXNygynSlgZna8xhTq3jBBOyv5NvqxZGitLsN2hdZ
CXthXH4GuYlGgq7R00wvX3REod/rpjkswn2cwz7soGdtisCOjPnwAY7jGUhlm7kfUdR41cMI1gn4
0noVGkHGIXxFbQ7KlI14/NTsz6N8zdy9jYwN0zBUKAkGCP2X9YPDNi7u8s+f+G1FHKIxutWJeGj8
eiJvW0IiFrtviPfZbmgCwZGjnZ60ZyFteIA6jLATytrdtfSqJpjmrKP89WtdYBgOMfeQ0ylf1P0C
0iwxdBWZloFN1KL9eFLrFfI/z78nJ+BxTtK4RMmkGJ2KEaONsMrjO+lf/Jg+FxM1HAXeNo8Z6lpi
zEzt3JCMO7CJyusK4WEpyzdibkNAUsUXV8+r1Ff6q8tyuoS6CGNhuRMoY4BCTedcwRYhjszu7DyV
R/TpDPHwtdgMNDo4778NuvU4yE9TBI/10xzxPtWF+Pns3JpWpS1p6XS7asdubvFxuDnMusNtucnU
oRJehNBAoMFOw3g9sXqQaYapouE0VdrnpDOH1VG5UxFWtemApdV4Gve/FWRXWEGOya+JZGir57Dw
lHDPdhddxyBvordD9gtAjkLtbhS19IRTjdupxJB9zrrcVTuRJFy5pd0X2Dx14McAYLcNm39+i4iT
gOLqi/I67ff5M8exQosr8J1ehuc0so34C4/khWUK6nLreZ0ZbEp4yVVJzfaYvH02wkof3OoVcB5e
jKVkiyShq8QFr5iodTb8UucOQHJPwvwRey2UCT4RyZ3viitGq4wZo+u6x+7kaFosbhc1yN/RSAEi
S/0t8fTnpr57XzdgbcKI1Cjs8CA9YM9Z+otT1c9OaCQMXW/sE2pheazmg1XkcUgSitWUTIKInI6Q
7dLjFAw77zGDPHZ858u/S2V9RJRre9GptMaVdtAkh2nm90WY0HLIaGBQbZP1vGpBCImZMDjuAKLj
Gy+mlQeFJoYTcBNOmCcwSnVCAM8J/0lGTRZcjHHzkSpSnBqbnjzfZZmb/WtwHy2UxytUstMQWkxH
TFeEYawxqcBl3nGJIVSuhyQKGcyh8xqurVYymyDEZCQ9bTG3S+89KkbGGEb7rmmd+7WdkKpnEspM
n7AyyWDI8kfUj8QXYcd/8BFB7mXSrz7JNhbpVdjW66ee9wJevfoDUsj2EwikWPXZ2jGAplUbHBXE
Ew1uP5AFaEsfthptktHIlo/pFhrf7b0+xBXMYvDiVVtYzfbJN5MPotvQlbV3V2NNvMb2DMTdCuS5
2SEpRI5JcGsnnXNH+DbbPrOR0UHvCwtxxH8LXr2Fsppur4PX80+Oh1+PexTfr4xPwchgBMeGbnGX
7nDzq8wLUJhJgCFUAzSPGK6VcAoPIPUkDCl1HKEk4VpfussmJjrNZAPbm7XB1OCP5NNAMEAz3na7
Xf+ZzMLygx4lKyrY3MBe31TdC0pYa74L2ovNTKzpC0Id00zxhiUSNNCCItM0Kek/lyjydJm/PLek
yJFAJMw7CeKJICHb5kqFeFatAy0Mjh+3lU9NBaYosGd5LXURFVQJAsBca9M0tzGDCy84OPrOslde
OP0pnKw72Hmc4FEXmvgNPjhGIHWcuJMsIGmUZykaPme1NPY3IGApu77ErDjb1qqUCqNb6V+A+ZIR
OnCUSpUJKNFdQ2uCE/YUfPVUTEEu0I1JMSLkjbb5Sb40YJcsfyoDitrLRa0wG/ef+o4vlujNz7k6
RKSdMKawUaaSs/BjcRkW16mqpZlz8f0bgqAJopyArHuQ34YQ5QqnOCpPoYi/E2BqJE5kBGcwSwCj
wRlcWRIrpaV78cjg0E6oMNMuaM/PnrPg8UVf0RBfJGeI7ltHa0AWUnC2wkr9eYl8ECWxfvBsmOFH
q99lLn67K4+RDvUu1pmMLoW97F6vbRuMM3SuPqUTH9WGLZiqbMPSpaAq4nimv32/D36IZWxpDx7v
03cRCMAzE3VLLvQhYh/U56tYBzk61jjvCQjFsPoTCyb9Hp7C72ZQif6d2iZZhrHTBioRv1LV8kGE
5ybC70yPQSu1hFub6H3FzkPYpS5WwVqRaETRIDxH898i27ntGns99+mQdMJ42QaxJ4dvNJaf/M3u
aWmZVqW5aSo8ShcEfOV4ei7K1gXyb4dLa5M88Zy73fIb5knK1AnLczCBNWo+pEbKeDA2fSKWAeYn
Nh/llmzbIoitv5dDppGksjq5S0Ic+RUnwWOxTbxk602OM4ZAInB+9HjrcqGsDhaFZd8jpgVSq5lL
6caAKnwXpqjD+RymljkaFjj1wCCyi+jmagSn4FQqy9tQjnpzRSX6yOZQ0mGYoa/O9d3ez5Q/Nf1l
YmnLnyTUkeDEnI0olDcv5etCQTpkiSvV7SZGXnyVuQhjoqnlIBSr2UTgzwMKWVHVMOktcQehbGQS
3ffwRCmH5Lh6nJSGfPK1g3Vh25lfl4RAZ3zyChfI4yptKagRKPGMtdH5O6e2LvLsq4be1XAPEYpm
sdrZn9F2t0tIUsQ79iE38T9q1M1mkDOdv7ngljWY8c7tyHI2nJRPIKu42UMjRLYpkvhvD5kXYcxW
fb5FsMtV4bcE+mz2EXuK7CGHgmbcXFFO//oaOlo/iby9nxFfGPgkrYnGwaAH/ZOU7tInBdp2dkAS
yLbIkHQuEZrw5jvrmiYWvqN2rD3/nEQ3lqxLiFrcXkepijTB4kPGAPATrPvxjwEpbhbSgO/jXDiZ
5bKt1c7KrtWZ9KWnse5WXNo5o9P0pS0HWjC2h03Jha23uTNxt+l6ZR7HQUk0dugA36BOxFtQbD/h
ZI7cj8/S9EZMOxoKuY2CfvAqnPM6+VFdHYPUnRLAKgGXEuH5CiSHOUducQh9i36xzIx5ydeOvQeY
HbrCbK0IYYEkFOiEnInFP+yA8ch32C7nQTzYwtZQbmjTp0F63R/rAtHaefWfh21ceYHWgZywVy98
cLhZbhLdYAqp+1oUy032KZnzH1R4UwIi6RvCRdtKEybg4xRpVPrCh0crQmKX78mrrZCgQt7ujmxJ
6VWAyjA2ngghl1Q+iaMDhcrmaLKcWpz+rTiOUrOVH1Z6Xm8ZnK3s7vkCOdfnBWh+J+vySfVQzEus
dR9weX6bEbpxzQkiOjFvnRA/oQES+CqafrUYP1S2t1Fc6l+RHOUAzvA5lesYuTDNcKH5vU+EeyKZ
W85JCXWle2JKjP+tODdxDZ6r5nvRm3oi7nSACip/2pClDfRX0v0LjDWox63h6vBDxrjKv7xDTUMe
X10NHyIgXJ9iB0PifXUcepk88jpwmMXBd/4+i+YQBHC6Uqvlb17qs0mUZfwFH0iQf82SzWc8oT0R
1yx1vJwrpeVBYfalavZ48lVDqTRhfOxoxJbPrWA2DlSwAyQH/01Ln+CQWsSyqeVHVHw6i/KYlQaR
5xQz1ZX9RJ0q9uEoiS26SQtrHdqkqgGwA4ObJyqbIU7xgNRw4DVXJwCbh0miaa7orfTzZlHZ9Cu+
+H+dLnusmSp4QPj0T91FKwlxCqV0vGp4P8lXt2+j7pahOXZbhfSDNTxpZZ7b44UaeJLv9iZPhxm9
NavUGJ0zECqUQo1XnWMvd5AtwbhuE2a7nZKoRvm0/cveaUps042aEOWh9jw5RgTy2Aw2sO1iNYuC
yUleh5GM3TIPO4+VAabEAANeqcSKIaszOX/mqodO7ZRkogVTdINPCiW8gSFIlgv0/H+AxWcVfxV8
AQeN5DkbeeJHbOYgn/pGQ992ggCaEIY6+ki7ppL9v7O2m2+TLsyTY9zSzD/K25wG4rGUVZIBFsiV
IlBSQhwUglp3Apti6wMyIkWnKRLnI/2VDp/MDteKESqwYRWMQ4CWxZqZfeLk27Tls4vU9SKf0x6A
8zfhlr0NGtjQhiKWRYr9wV0VtfPZhfAcDTjoZRrGxxLug/oUT7Npsw1Bznv2K62duBJHjlBF2GZh
CBD0FY1leIhA/DskE9sC2ra12b6R5wPhCyfLRTTzyFTFaGXvm695K3N5ZLB/LzDOafg7mOtJMOGo
aGqDquzvQcbyEgYAVbyWMO5TpcToT4E5zZSgv8MW91P/vJScH/QOmammKIVhk+PX02CDHG1QdljH
hYW4qwWLyvUQRo8gn9i+Q/FvtCt8rqdeFzKqFJ4705EnGnMwy+xd/NsfiNMP1dVKXxT5bQ0efgJG
+Paou5opbxsE3nKLdXkvY6sfpLOBY1OBrmWQHXcSDUufG/86q+36h7rNOL7yFdfye/fPcS1XmF7n
CjbLGOYQ5L5l+v+49COj1gnj4PD0IDtk9VNipWU3BzQ0fUyGnRA3RPTqOep5D2Tow0qyF2LJg2uQ
/Vd2R55FLYiRrEhKoUzZK/9mxusZr2b+C83spmWUOqAdOWiHA+mZH6ycWC11xhLNhSPvlgKGSb0J
r4dIeYErUg01ziYf6DWCDXyrtfZfAxAjUkYu8s3kU5/kUwho6ZKub7b43Wn/LdETIF2MH50w/pbR
eD9hYMFgA09Ncl/BAApvOvBlSNtXL//AaxPW/x9obhKpqTtsEKQsgg3kHWmn/w1ZlCSEI0MvGGIr
IavIG7a0+hzsbrNb9ugYq6IlbIVoIYFbfXa8eVm6yW9mRgrFyZXVwgCOrbJ7pm3GaBBAD/ckfUiP
ZmcUbsN29vJct1Yj6f3p5pPpMiOUGIgP/0VFN2OThuULth/qJHAeykp6vWqtuYERcpi4Oi5n3VP1
z1jQYMTM6nQlDANwmdDNS1CwD64BudVQH3VU6cNmgu9cFltz6p2rFkve86d/ieAq7DolfACy4Nh7
I7U8w+ls4GXowF9bgffDVFLkyhicVYkRh9pK5E9BvpCkZzBNSj5EBioo0tzW7kRekaMMc3A1VQig
Wkdr8VVseA+GRRsb9xGJfOEPmZBmTK9ttpPHMrZ0TisHsArJe2xYPySmITLhiNy77o0wGGFsKCJJ
b1eDnrwlSB6MQfcOzd8eo38P4Kn65PE6UojhROZQMj2sWG6BH85d6dRwqz5QypMhWNVKCj0+Acfs
3uiQxxM2aUsYwngZb3EGjpmI3bWP8efKwvEF7O9kkfNOfr23D4NjSfJe36hxDD160pLWUcUtgS+H
XWHKBvXWQ0vZVnen4NiUkWph2v2ZopBObqpqb5LdZKfWQSPsRjHOeT+9X8HFWTq3tOx/bVhECPv7
rKZgYVBe4UuSioq9wmn8xaYRAFShBtB6QXE8fHO5JMshLPX8DrBgPaQ/ko53UEGL23uIpKfEeVMo
byFe7M+nlNAXXIvYwpxQrZsJjwLrWZtO1R3yGfaS7K2Sp8jAFPRC2u/FY0aPNLNViQT90cletGtK
fR1fmQMBktkEApn5+oG32OUMmhtPjSTPsfKSgy/jHo+x3RXWL4fyOI3uaoEIpM1BfPcP4dwJwK2T
uGtcl0rEnFDKg2fhv6z1WV3nWKgBerxvVneBFtwJEbI7szpAn9F+02aIA1hfgK5T2opnUGYcggYX
WwEDKQ7S2xibpxMjjkwXRd18x+igcXb3modVOoWXWormGeV50ZaQ0qnk8cGYBw4wQSQ/QoxgvXrx
HnJ7qbJWHQDqMglOI8Z7qZbQTH77500G3ej+cKTk4EjWzcI4SIM3IYWdzecwOE8DG2Nx4mWlMwZJ
zHU+FSCiL8mkWHgE5wAUmovc4YcjbPm1RQ+ZsnG4Z2HG3RioTNag48xy3f5dhN7bttuCy8OO5+4W
J8CsfpRwpu7dwj7UYpcH3jmFRZgua72xnKJce23arABWnoxj8W9zqwLzFgcij7iOjBj4cW0O1xAu
aITqIhkuuTPAodch4ed+eBZJk7S2ZREFwYriURaropT6sKWaG6fT/kpjKdkJnylukJRxQ1N1ZwB4
PehWtoWAkhLpaT7OKgB4iKL0kTaTYBceoQcvYQOva9nuTj/lby7pd5AwgQ8Ku1BbbqXZge8/b0TU
JbSlNiRwsNRHXbf4O8fwd94XrOK4LoKX3bnn+EyJc/R2wcSKK20CTFaSp1A7JImpzb5dzKq413AY
EgQVTYsZLOpVJjKbd2bA/7SqWb7QutLXTqdJGagHKgdXgmX6tpPQQRwSDDI5AjPr7Vb4Hahx7x5G
EF3yLmcSUFC7Iloxr3T2UjCYacHLb3enrEbkI7oSJPG5U1uJMsZKmAyWPwY6APcC25SlzkgqTIRM
SwhR87dKgySJtOvo+gqSEUh5daKGgVP4GPGFVxbh2WIPP2Qzg7HARdvHfTs1ZL0uJEGRyoP2MzL7
xYFCK0ffFK//6mI/GJ2em00ntyyoQYAvEavH7Z/R77bvOz7e0hakVkwJTJ4cenEv4ZUl/5hkQR+l
wuNaWcpZQzp0P/ZWF7IN8sVU6g5YwAWfZye3FQxHUNh5qu0nUGm9M91Y9WwbCbvr4KfLn1N4JybX
F34FfRNaEPIr2ffuROOT690FiPQmpl56DEWRsRjWWs9fBQgN92sjb9adJ0nNEY3lZlKkWQF5ShKB
zTnEDMb527o04amfjeKz9Gs42GOnV5StcuXLaMxgQ2rI2jh9A9T77iYpAUZxXcWPcH4tM0EfF85d
2UO2weu9i08mEYN3WTFCvDbdKCkCBXjvy5SY1l2A+bndo7g3FwgayGXruFoEjcW7y23jMOf2jRKQ
nje6SNT6ccyA2TZ3XHcvzZpzhE5Lo67Lyd0C+uSKtmpzgt5qKR7YnoIZ/NrquT4OXvWyyNAJwwgM
rNUeGkw61McBbLzqJ6p+9fOMKwgJLjsPhOV1yl3M3ymLqNamY1BOwARob1bITpy6bMlxci7sXpME
QJ+iZPdjW7f8JHYoEAPGcEHH1grm0+YkTsRhP4QKE2o97Mov/MTiOpH1xUljKcGekVrBtsFd/fxB
bo83aJtKbetcrq4sL+8rFf0rcFt3jrIiNfrM0xE2MLltisapVMaW5+roZev2Q3iAebZijl9nyjb+
a4u1+SSRBLk5fC97OhtWS1lpAWoj2rKzGfOKk0hqtabWHStQ3riyqRznDPlxTr/IMtGkUWSHHpbH
4orwGKuEvUd4cP9Fp8x0dLnogDGqztZdBEsXqFWUF1cKzb0B58Vtu5ltuYlXiK0P+2pO1LxBHdAw
wwEjNpbWsy2oA7Zt0IoMrW0NhR/f3IThf//TM+90kbTk5syU8GiBsnbqhsbsl0hRGoIU5thD/VEy
jARwzrEA3jwKyDsFVapR+V5sPVkmD2FLBGu0fPBIGr2NNyTYkV7AhwVcHE0J0njOlD6VjvkaS2Tp
Yg+ofpfWPtJpqFm2Flt9GtLJtsk17LTkicu0cQ9wptoWdQDHYAkh5KA2Wh0SfV5IFKhdMn4RcO37
GqQELpZfOM/MU/roAqBZ+Bqsz9Y8O2pTICifJ+20kgPIvOAcMtk+SXdZAEpanFLYZHwSu+fBfk2N
/ccWWIwIIeww8OH+Y9vHrJ0wokGyaKmF1gDnU5x0NKJHIrTeJtHCOENy3o17vmgQFTvIt6qr1eI2
kiiAjITBcSZAhQV/AEnzkZUcPg08KlhSKHnySplv04dD2omBJNmk9UGajUC4I4hvjGm2Ac2lI91+
UsRy3YRtpzj9XhuFKFKCrsm0HzufgbZ/ZYIydSH2yvNsjMDZi6JQvGhpIBLgz3hfRAleIURQeZnQ
Lw3Pw11h6VrobNMM0IYiD2H9Z6oT5WYzXGWE8czU9DF3HyI/BnsTzD7iBYM1oM2P4Zj0YOirVWG6
ionZINf6Rg59MxXlXODFFIG9OkSJbIjOl2cdpv+O21EtSJIKuDrw2rLw6r2CVwlIQ2qtBdEtURE6
wFEAyUEkR926rWYKX7sQI7NFvtTLL5QTu8KnVMyJiGaRzoQEEnAg9pjG9RVJTBcFrkcsp09NUGGH
GEF9hJPeQevIZss1nhQcDmCLGDRm0XM4JW2EzxXUS56N9ObIXwVNKijLQSPAcchF6vOtg6svd55T
YR6uqww69kQLeryR+axRU5iATtNYJRTV6W0d/NLdx5VuuQ46dI9E+f56IC+/lBQmaE+hU4lotnb5
li2YaRaiW8i96Mz2lL3QWsLruL8sUbAX4dt8dj+lid292OEVwRp0+j88G3KmgTFxTJiRyoXJGtyG
LfBrv+m1y1AVI1T+iqn+bFqKzVXz7Txjxwkq2gMRtNTRCAtEC1EDXSImmEPXFb5WpKKpHwf0B9py
gD5kptOCJgZJctYgTq1Cd1xVfS75TmdW4n1Z28q9LNbxvsfFGdB+dSzbyoNz5GOsDeQbOqIRdZ8o
WvZGeQRQHu04/DcQmASj4WwMKLEwBAOBmpGJwZHD6hfh/GZt0/MZMzY8zuX2pAGo25lw0Jr094hc
Ywt/S+6kIZcodf+rzI72Ne5j/ee6k8tTsORTTpZcSb5PfVRYJ+TcYKcLHxSWv8DuDnKSOm2GW/HL
m62uq3syBLZdEErlVBzvcq7yl+jN/gxQB34x0R7sy7qDQDkESI7b9kGByYLGhOuUzeJmb5Kg5+DP
QMSSSiyYHgZrXhQXS0b9ZSkTfW5u3uS4bWMYKzTfS+Ef2GsCFytToPnQR1NDn+k+rUIs6NEYw0d9
fmSmk3Ttsfp9787f8OFd4izYnkgkrgWWR0uJigfrjYt6HZAWStx9p4+QeYxNxYGPsgo5ufzK7fMG
z+J54EYUXtoEjLtan0Gey1yubZ6CFUy+ZwTZJdQCnunowuP0yphcJmG5UrLO5JsN63jKweb4lSAY
gpS+4Se1Bbdup2B6/Jb7+D+Q4+uo60fl+byVpYs+TP5qKCZvptTemvZEREN6ZRoaj2Lh3deSDhsb
mr5/4PBLEwx1EpHWcWJESDW5gdfNQZYIs7xaIyn+di04N/QK98ElnwoC/GnNGfMfHUH2pYDg+Mxf
J9rYgGAblUiUTk2i9zGAsGpdVhRCE++otObz2EaOy4ACAm8y4ax/3JXFA6xmYDP76qepICnE3gU2
H6WT2Mkg2l8m1ir5Ek2OoWy6sjD4gwx0B34XdcwIYJhURRC0d1TrMOSYpQmnQoSh//NP17jPcsdA
Xqziy/2hBAbwJdXnvUvOQLtJdOMb4qTM+ebHmwhkU2CWUJ1a7pCtcVICaHM6C1aTForLMUcGGqa3
IfBp5mbbxyDhSbKOaB7PCVewdFgQEqPUz3CwWwytKZHn6xVPYzGuO+igtlx/x9r9vClcyqAKIsAi
9IdP2jvBpoFFXDpWsiVvNygcv9A3zPyiwWW9umWI+fI1jThOcQexCbdgKLf3oJxTTmgCsDbu7XCC
r+43TlPpQDjE5pWUKZGTl20ec+7piILFvBC5ZlaxibqgqqH3OXR0kZLxANNejTxDcoAxVHNz4z7E
8KorahSj3loJAA0CM13njggAL+FhLKz3u+PMXMdMtuKmCUSoGTw7Aodtsc0s0QGWrqGi56m7DYWT
QJFuYiaNQ7fvCz+MeeW0KkOmrjUq+CRCtnPKmt5OJ6DUYojobwzYVEnZ/fy0Lu+lAFJncHt55kbx
luwdcQF2dXUYoQXlrFeRkwdsXa+rD9W3Xc1FF7yYdIDv5rvWTj8Yu1nxsk8PsIbnBzOR7TgpsqkG
bxkbGqhpAjcDdOyqXo+aiaFq1x5ZRZICKyspQLB03gqhXzFwvs+vQKBmNxG6JupHj08iahp6GD+4
Ft+X6w9cUcVJ0vXGKsBy/B+PVVKcqZ5RZtuLl7m0bvvnbBcVocZN/q0UvC+Fv5Sa3NcoP3HrE/Nb
qPd5nBWfFzFzR4wdTfQXDXAYIYi+Ji5yHXgqsFhXzG5AlDJvYvLztzZhLybuhqikVUSWVma/kObC
V4CfPH4C/fCtPaYCIEJ+rN+DI58AdVq4ujedizfW+R4QR+XyJ0OYl+6g59hxXBTp0MN+9RxG516G
7lJM2nLfnwScUrwrWwRQAsQa6v/22zYPAJu4g0n9hLKhKCiqYS6F4LKbaPuU6zTj0+yan4lzxRo9
1pqh876c79LfG0ZOY5AbE5l2IK6k6SpKFbpG+BQuoHz+KhfKODhNhHH5RL2GB2OSREn7gmoowdQv
a8NvoS3nRd01HZLB0UfxYDdG7fAfi5+bCeS8v9nEh95ZLAEYs7zpYPVvpN7A/4wnBrrYTY5YR/oS
KNdoywVuusBDkmf2poU0TRAozobtvwHV4V83ePKTLEBG0RfVafWK4JIM5zrwCC9cDrtodSrWyyPu
UZLwtnjgK/ieZ0MJ3fcwOZ73y7WEHU57LigcR9Ey51Brxk9mNM5u1rEf8orpHT+9WViY8irEZA6N
pYk7fm6/DV0DHRqCG9sQuEYqnkKHKVVynieROVYz8jPeU+ghWC/g0NRVbpCgViZctWbrxieXWvan
YiPfotTr6+P4YHa4VcXx8Om1QjH8LqGCGNLeZRYx/QBdK0R1F87nQvVHDBVbwTx5+KGnDaPQvqh/
BRj+cYMtBPCYpc2/6ovdsjuqTqbjf9wmn+Ya2dsQmK79ii/7Nr6w1Nfm789Wdqe7FgscyEg1pCIw
JWlgp6tNxtOI0/xkuuOjN+P7hIdb7hC9mFt2yKXGGwfTaoFu3/mAV2Wv6JqA0Q5Xr5jJuqwptxJN
bt0k0DodYq1UOa6rU/9lWADHGPNpPKgmoOcE4/gfoSdWAsjZAZ6zUgiT8iT50lJOX1z6h7UovBLa
RqBkN04fGRWaikorPJat0pwFcJgI0nuywDL/Hj/6Z9POnAtELobQ9MVeP6XvHE/K4H1GqmeTK4Mu
2CU2BbFk7lWSWi7vtd/C+lk+b1lAceUQoE0MHkd+mA6bn+WsmhoKnHtM0vV5R7B/suvr+iGWYH/y
1pwyGPhlTXRtlAqt3vM3ZpTsyYGM+QSq2Ba1WogT9+ldV/u2VPwPad4Y8eN4xh19xWLsrzrY/M20
xwswnH13Cil86/b03ezsoT2zR3XiugQ6B9dk/j7gmpEjvkvTpC5R7g+K9LA055aSLQs27QG1c2Hr
wPyL6PNlzEiRHvVcKYkLB12I1pstoxaWQqVicUxjf2szxV+P5C+MNAZ+l9jOFMD3lyYjy4RD7CXq
ZWVNrW3fTUtQHEDtFS3vX8fgLvnI+ej8CoMpwo6V10x+DgVskL16mEm/AfkVramDkNpd/P7ZgqAI
041xizYbZ03h1waKXf0poqI61r5EPEZlkzF08ObMJPrc3MBCqCAPdrV+1m/jCDPCPPd0FiM+p73t
kELqRoT875AsV6T6GaQXSip+VOAsxtVLHj1kHYsJYOQOgC1+dOuV306T8eFSKd7OfIN4C/hjTI0q
Y8ppJpkfp8t3QOamWHolwkRgLVTgFTEGkCzxtz14Ys8/u03Y7TW2k6ysk8dhmR7SzXoxeqTAM3CW
LllIZP7FlWQnSMrHO2WPWcJS1JxnqZyEmqlfgp4adCQnc8H473KBWbGZ1LdaKGGmEyMnsEvyfpwz
4NOCvJahPXSd5T+Mcf5ffB2oQd3zm60xWSZrcGt/0rOLU3NB+9MzLMnjclCpQWen+GwWF+ktADr+
EnnGhK8QQoWTk0mRVQd2kmyF4H915EDX5bwm+fNcNJQhij3bY7cZBx05bipVUcwHfewl0U/KQx2T
YkJXJJt/HTGaibtjNEqET66KXmBhzHKCR22c6IcmFHBwqGng4lmkO0azDDQmdPjHNWoVk80s+bsa
6OHRxy4Upfb8Ic/2KybocqvOkPIuvBUUWOm/nPoYS3IYrgRlMSnvleXqcCk2twLlzGYTGf3xthtL
3vC+LxnE/S5mHHh9PWy5lbi2Q5FJzirdV4bf2UpRI7+PM6yEGpH9CG42TyBhWET0nRCRHsQ9NrwM
yTPFcom6i6WO2IJvqQYUR0kp6jTSC3d7DZ/ur6T4LV7PYivdFXE6/A08xRdjoI99rWA72OWd/vSz
7ApAJZNiR93T9OZ0nst73tPrCuNfUvrNc4lLqm48KNSZhMiW4d+Okkcj46tAmuFFSkRklCMwkzyw
lD1xUVfmXvVqTecSQ8ul9xBDdAogWasyuKVbzoUmkydL4V1V/mnuYR/dWTppje1KOaoeFHY6rya2
duR8uGFyq95SYOGjQJOIf/j8GsZ8PcILiv1j2CPfGy0v9I4ogtII8W42bNnq4JQW/dyzd9FYhXRP
6uGK+osPA8jfB5gHEy+NhnwcZwZx/Mt7diFMymWsuobUq5K7ecCwHN2ljTj3Lh+GSMOrfb0tUrcu
LkBl+KX5ffJEkgTL/YvDqdM9ldlR3bqmbipXOTSzog4VvPZVTZDLJWzV9qjr17BnXQr5Cl8UL61c
mvS0tj/VaTDSzcw6T0XIxNVwoRZ0dZnj/BHqWwNJFxg79zvOUZntrtd0NJPkemBzzTCSwZvY/yn9
84ZIFIIJTS16v6O9DnMTHdVg65kxKnBWoDgQZC/BPoJ04dl9syL4ycFGXSXyJkSlTNtcgInk+50f
g4rlTVGbrrp6+9Lm84vipYnhpaV6h0wQOdzuCHZB0tsU8SdWcKO8fTfRlQ+NzeUFg8L4WfUz2LkW
yLvLve85Dp9hFkptKfnsAJtkAFVLYPkBzhUbtYSDr5IXMuGIE0ZJ8zWzxN+ZBD7Qc8Th41js2iqU
+lYZ/Fza4axYsGA9cfG7sX5fbU8MjeJl9AQkAqYhUNw2eHEn05qARbQr4bRuCy9nQzeCvYIxO+/z
qQ2YNytaeYTVuUKEOr/v5IsubwCuyLJ5M97co/FkkTQEQoPI65jFwfoH1rY4ptOmbPRSu918ro9f
TN7nDa8CqbGkjvoyoYSb8FLr9JYUZT7zK91OKNqJfhGXTtypVcbU7zWp9Jy13JgTxrAAfoynYOnO
Na2/6pyZFtT3aEgARZ7v6Wr6BqEvRruLrLRCFiLbWIb200Zk2SMe14Dr1pJ/Sn+CjJPTLWV5XDyW
Jg45I5MS+HyAu974wjAMFcc4SKGD5WuYvRrSe/ffnUSVrhWr8gdNHpxTx0aiZb9E96MNua4FNEY/
/tXEFfk2UdMSPvuC3oIRTF0cAzn0OM6AzoCRED7B7V7jJJ2s/WBTvKkHxTP5l8nW29Nl1Ri1Wudm
LiLOVxaLn7wXXSYD0KVHALKAysO4bVkHQrdQzkEoLgSdXcEk8AMczyick2b6HY0uJo9mJ0MWgW4z
oGcChjVkNe8FY/2jfj6IlQXSUV03H7vpswHdyTggp43KKs/o+8yB7IRlqReOU+/qMZtFVFIYau56
NBRUALa1QSRlgzNcnSQwtF4ZjGyxJyERLNVPDPP/UpDjJBcOJ+alpGurnFFSA1ZPleDi/L6d5gZU
izIYiUZ1lZbABE0o6yNG0GHbRWopnCDP7wVyZ7HZjlljYQEbVyTBEICR5m2AoczjMu5KXtR708Zw
vMLFl7aja+dl09ytEBjWtiv/YQOvtZuGKaHyruauAfQOCIAZMAdMlkYJRLHY8sJlHCRZnukSVLZx
amGuXlTLIsuJ0OeED0/vW8uxZHw0Cgd1pl6SF4BA/qIwPEhd5OLQdvauuJmZiV1zKT6Fqvrre+Uh
Hjf4Rg8iqpXckV1qgaIKD6Ss9hYiLATLJQIJChqbDPelaIrJw3KyMtAKsxNPUpfWtAxCeRbc7742
vtN1spjEAjTPUIJdOEOi1+y0SNYPMOIIZwGg1HBTJXBgbQHLSDTBKMLT9eJ8d7678ewjMmKG81ZP
IAAFOvpKvaLkqWNUujllQP/5GKIIBGcPncIt9LS748Yw5oZiZXnfd0CkmHO5U80Cs1k+9WDj2l0R
NQfyJgaxliPEBfc7U2udMN9eGqvZ6hrE1LTAIIpDexgUzRplQ2/rY4lONn+oLdL154lBvN9pYLUZ
utooAgMiZJ7YFzFqOD3IKA/+Ro3xfAhyUOtGjPNfLW9wdU35pXC8B3GWBJZs4ZsqkzW2U9MN4mQ8
hrgE+zcLlaqDXmZFGhfvuD7/ed3+JqT2NrCCjevAZ7Z+3SHCWGl4liA/bMcfBN5KInhom/JTtmOt
Anocd0eJ/sX5wGyWzDItn7ehwy00LbgFO+xg3e/Y9D8Gb8SCp1rOGQxyf4P6437rC1ydFOBnkgc3
qDVmFyt60SfA+aVM2puQDwKldpnUxH6Z/Xp9Hvcl2OE7ai/h2I4vUcU68M6ODMOJRL1hmQk7JIeZ
vzYpEhdDKYp14rWDoA8SQ4CChECtwB0NBtoab/cu+C//uE1UlU8W7qc++UG8P7JGZfo+/GVgMNFg
ElFc6nXYSyWrJKYvSltLcD2kal09xGogXUo21dB7DGdXGp06cYBJKTXH4AnUHBiRRDV7uWK5AJxP
FHeVlL+rdGDMypSuFow88ev16KSa00r7/7Ks+tfQTWvRkjsLWgUFbTvm3jIdSOR8he5SErK94yQv
AUkEolVdEJimHVLO+Yr2oFaLD8G7FGGK2hWHRxMsyupMc01SX/sLNi4ZPQvE8GeR18Eu65cxZuPb
eAr3Ylmiq6aqa3784bEjgWEq9s2RQLwy+M8xtBdhCxHSOuVV+h1fLOhae8TKHQycKdwY2jhkP56R
zQTRflWB2cDqBum59h3JwuR/3a0oUgO+9OJlBG+UBJMAD3KbRN8kXKbI0ypJf1wxag3mK+dsDOdT
70S0zCxzJxTs9uEY6cR4EDC7BUKdk7hqzuhRSwcZK7fVNvBIx3Er+eKgjoZOMr/bfhentQ9kKP9S
ClsJLq314SlMNPrDPM+Gd8fqTR+N/jnJdl0DW5ifG+7/so1ehhI/VeU/1zuD4DxuPZSNWln8x8Yh
dkl+BMxc8JTD9CutaS/tFTGlZnsOlPn58j4LFaQ7+5kwkn8GVzZnflsgFXv/+d4vDCC02hX+iFAE
lfw3zcU0Ah9UbwW+FLchr1Hi3BGwL21P8ztPZuGrw/UfqQ68XZ2SRwQfuawya+35hUKMpIWFO/KM
TrqtWCje9msiTuPS6zT3DGQI8/3DiccPs2RTCoFf4Iq48fQujNgCxM1P5v+zn5lfkXSNZWIym6QD
ctbQMbKHJ92N3yI1GycrMwQSFSpn0/djLWrMECh933cXpKsNTlpXFKFz8bm8fBXPXjqLL2aE3ARo
75Lxu2RqwsYVoFVYsCP4GVt0lVE2RKbkRybYNo6tMrZ7J7pKLVSb3bO1H4Lfr6p9CD5Dj7uSIOvr
WUU6wVA/iSmrxnQjwVg4qJPQL529EI2dJDXP0GnpwUIYTCUs7i/UrmmNchZFRk0PoxM+4qiJWX1M
9NXNUFKpJC7s9o0CnS3g9RLN2nX32aNSbOpgxNKjVcLh7Yo0M3IBj1uwv3di0ywstxt30asO12xP
Uj9XQjL8ZTcKyVI87b2ktmETS7Op5Kmb2lmcxfB3D1BJWpNj52CrMgQlDX0EEKEWW9Xhny/O6B6q
8pIBkmoxA248GqdpZ7kxulTyoYHRrugwc+omP1md6GBjkA99KeHr+xUadbJxL9wyGpscOP1PTv0s
UALK7yPqwAEUIPwjiqIYkhotPOP24UvQn+L7EbVnCmemDQhScmZxHL+hIOF9zaJi3PQFYwlHRcbf
aVqqA74MA0+HSrOOz8Nt22vT4fOxWU8GNouZjWR+xNGO9/ET6g6/DYQFtctCn2S37P32ct1ljx7E
STosyNxpTnwLXZBYDQ3lql9Gcz7iAVXkxpX3XmTmsEWJpFsexEX0VAZtXIgVrJNZT4h9SSFeaopN
LF1WGvjKr2K53smzpKvvdHGCXSxa/YNZFRLlgCZSlJBLNtz1xhUzwD7qz20fh2/SEgSQ2Mbbq2I+
4aIOQZoSmnKb8uZlYBZqhP2CUVD+o2WulXSgDBi2DlWXn9oIY761M9aQ2SSRPyGXESJbSmkU+Pwx
JT0J7YrduDnJB0IBOcTRABJgeOIfBg/Lnm4/2ysTAnzMERhzZFAdyYf5tKxyiB581EFCXj0XGJfC
tSBysegLsWq464MBBtt3Mjmpi0r0iQiyF6TXOaDuR+4oVhWNhscDqMcDB5+C82Hql8KaGhEZztmo
8t4o5aSgq1jBnEbHYIsg/y9n02DwCqz519b3Gq5wLmKYZIvIjSMTEEc43GAFIQ+pj+GGDCOGp+qh
kWYqqQETtOiNvDkqoCGijaHJ9udUVxKV9jHFuZWMrQ6VadD+6sUDlEytJZ4K/yyXuVnERG2CfHY0
oqEftZYjoUvvvXsEmo3sb4pmExp65fO+pEGfR0NkQ65cKw+QD0LK2cEJUvlAzpUwjbC1c7nm8tUa
urVvA5ulBtS1962gHyC2kVztXH1/hyx5g7/FW43n7FcjgqOOomm48Wy1IPDFAQdlr5M8ELcbr83G
xlvxO+F5XIuwd1qQstJllCMzfcWxfWfvCsoWJXO/by+gJlJ40ggWU+tYOww6BlPqsLL4wuoT+F6j
8ziGK5Mf3TGocHyUthl16k72qHix01BGsh6uXzkxV7guibKTX56dfLWD3XhEpsmw94S9G+dYETp1
MVkC7RLACphgRhxIOoYxm5Xy4ocD9i1ej/YOjLoX8RqYq1G9cGTU6eFB/zzaphrfdfIgKsdkRiR7
pphMrKc4faDEZQ/K9XeTKUAHia6s6f8Wd7y17Ez/r+bCx32Bjy/niQfyJy4YSfhFsBLBegl+iBHw
7//6eLGJ6xNeUoYiLOOWhE7BwXylhqtxl7tVbfqnLnERoK+daxUYXwZwyTuk6pKF1UsXP6vt15Yf
z7guEQbtb1ta3JpkhSOjshevnYh+f6fTUMe8h69uTgRivDjDYVvX9oBNAAe/fDtGpkw+Tejld1+L
9UT/oIyCUypmZ4/0y3A7CF17CBRGb5IMW+dS5ubs1bTSixvcQADduZDgUNTbkgXcxNbsNwh8smnO
9ux2aU17BXdGcE0vRaPIMSdf5lnHiCqxfW2HfZX1IBIglh/p1mEFfnhaCEDJUhU66wvPXLknVt+m
QFxMySpMNFrK5L0CFTQo63xd5x54Z8Dp35KXp+3L2lwvMZaiOMGSRMmgt+50DvIE5S1Ka65B0j7o
WDkOAnOD5hJf7ueOL+l2uYxXBPSlW1Muz2RqFT4kw3Uk6hxCw8dRwRZNO1VN9Bv9MI5kLSBJgdWX
18x/nrBhPqAPSfAMllXAwOg/xqbJ2tqQV9q6XRB/FXoBXWg3KFFp/dl/F58IXvWPYyeF+j3b5EAH
/LBu5rQ5kZzsTiTW5V2nh08fzJ9G5BZxiG5DdLcGEruEvUuewJ5MN8by48q9NqhubZujhvFfCkYr
3SDXXXKP69IQfsQ4jERxkl8qPZ/6dPfpeZ71gavh/SIvEogIA7iq3FbJdvE7I8rAnKbowI08PQGL
9UUFOWrkMQI4jWB67kdoGqaIvufkAV223fwMPQQSzoqohSD+nM3TzhCCghOgOHKiQXHHw6XV/lTl
wzgQT+FmXEtHdm9hBC5yL7yKVlcKA+29j83TqFkU6DNe7tTl1suCgxf6MelSMRkubNEoVhH5cE6H
tvhNwk/XlAHHEFizhbZqZEOTbkxMPGZtLTdLxIK+Y1jm5cL0tGclaLhuFRo8Rg+CJoJxFMcG9ZCc
xWJ3Pbal/N5Ryr5rWzpZ1wz+p65jloH+tB1v9vHDPGiMNKa0rWSDjNBf239cPmiy4wdxLpF9LmP+
qQjbNQlhuu1P0xV/La/GuvbMi7/gz1VyrAN/WdzeDo1dxpDwpDAQs2fw0agCrG3Qi9s0BM6JYfY4
3FwEDK2VHP6ZyjCXlXKojIn3bLMmkWm4i3+P6M2cX+L8MCkADRDTARhU8zb3WzYI30HTIerEHpie
3yhhfHBEozN8KyIfCc5qUC2JeDdNT284506FUaIJx9DyxAicBf28AQLfB5zgsKg287916aXPTq/W
LjwBTAIvEsjqd9wpGo8g/XvEmj10Wdgfl1b2QUHDJc8NDpwggmytWp0rOXb73RidAyinW+pL0AdF
LfY41PdX2cQl2QMsfuDODxfSkFyZN8a2iEVfWGUotK6aaWbLbTeke5QBTR0ZV3S+RO2ngJCcshfl
R4iPqVc8n7rH8hdhAm2mdj5jrDAHUs6uGhp6vEsc8UYr9nEgs7wVW8xm45JMHLiGx7ENyReXJwHG
AndOX1lKlzxvZGJByG9b6NPr0DHASXk7MCP6l/6qcZT0GJtlgV/5eZ8tqvAnW79DGc0iLM7k3XoE
p1zWpJ6hkztC6X2OFh6xeC64UkZvUBUdG+8pRTczKsMKE7pGKbjj87SgbqF4H/TLhhREMLtxDAiB
LfhayDqwMPzYOG1zegxG5fhD9ugDnppu7o/LQtq3QnCaJuhgRpFrOkH0NaMR3W+q4GgYuq70+iLl
Ad73PXYrmDVRvsltWg5oEiZ+aqIKAd1jIibREZIf0WyQGJDCwbNxACN2DboYFByNVCmXtF8zEv3q
Ot+DdYviyCTHVkJc9dnp4zvBxtHBnQhdTaN1uMr57QDmKz1DW2AaW9dHCNTHpHW5NMoVGML4FLhA
NEevHjO04DlWpUAmX3pGNKyttCDXjLtffzmQ4LOHf7n9NlpEBV1d14MGmH1vHzArz+7s99XJG2Lm
sXQtVYWxlAMbLXIGWvlTykub2yiaFV9bfTjNOIXp/2EhLog3LTml4E4xWDn7FL+cT1ViwIkcKLqP
RmgNOq5sG7HJYWb2Riq0MMLOF5rwTJhzjVdXsCD3mOjxOtCTux3Q/WrWAw/LXHvcI3aGhNRZ8ELq
12vOnV8XySIutgHBBJt0rTlIPtkOAEoHMaOhi7bY0e5+/dmLUN3iZy/z+3VL61VQmSq/k1/edHpf
qxCBTvk/tKYOVXrQ0u4XoncmATxcYOyXQjJ3spx/3TZL0OaCMkHFkADVd8Q4nSMLq+0mo6laynPl
FsGmgi/OMXcTpW6+ivKVIanVNuQV69kfVJFvMFexSaCb0JzNqxpgeMQMRI+FikC/WGPP1KFe34ua
qDBxrfZo+mirgoG7NMCLgjNI4Evj7JzVtC2qsx9kgbBv5GpIJRG3NrdpwzaIY49G0ucTJhSzcd6Q
2j0KRiZHfa90f8yUulPVphjvh1QyenKO8w/4TX2xTA8wdLjks+3xgowl7ksA8Lj5c3GZ5LEnVb8e
rKCLqOtln8diEATT19ZwA+FkqK/lPghct2Q4v5ThsUSRK4/XoE2tFR57EAmDG6DTxkRrH7TCTJ8v
KzEDJlABK0+AjD62UMU5NBD+JfunAcNKLPtrDOWwhNW42DhEv+VILWs6NCLCEdE2ZE5Qe3poIJ6F
ddt2D3h0BKK2vgzMLoApOeXJ54zrowJ9iqfFEB18XFTaq8pi3BWCwvwrVoC8sNyiSeGkYCEcQItf
ydkCrCoQfDou9CM+6xQhiTwybTuUfn7NbFPossB7LrLlhhmKuhmMvg1fGToFi2onYnaIaTVqIIDD
KccaXwGW8EpQ2DW9vrGoy68i0TojDf1XZaLPAjAikgMeFpjhPxHP4EYrehz5schLUphKGxpFJfFL
VwXyhFoLqaucFcLRR1evnBGe4pBWHXlm9UyFeS+RMTGof6zbjpOtmaZNbM/H3L5YurCzKVu4+1WH
2sOwcez7SJzNgPfUWpvXq/FwOgbEt6XaCOigwpgY3QPtjrPEb0NX137QzcsrrAyE+3ISU48G654b
ji5iP8Ec4jHG9/5jz7KuBweqEG6rTHXKweQEaXa83AKPFiNDSvWJ3smy54ctql5mHcGIZ0dlYPOC
WFtlRUCC6xM/xeQi6tK0uZmBuF9szklUcBtr74zL0/n5ZDFtmBUzRCyuidaze/fpE333K7XhCfKe
ueDF1vmBlzCB7Ad0gq4G3yT4+sJUYKOVOq7FE28WHFjFIeBBYReDsrMaRx5C9w6np7hiZ9lfI0L1
QEDEMDap1PuBGeif2A7pt3GgkrNUQf8KAQz1l8eQiEGRueSKPl2oApo62w+P3w2i1iJD2vX2nK+2
2qKjhR95bdP749LWZKEtzXaKC6zaUWzqTGOwLPD8OkSAjKZ2tdi2vKBOfklWfeGLIQEzEFlfCafd
7/jCYN8JOidbQRAy8xlUSLKbgY8v3TJBLGnNeWMF8zEuoj2jUElKX0TmH2ufsxqt0rq2wiWZqB5l
UUJT9akhTbfQJvOagRLEo27wQFYFPCA5L/kSBbIS+aMnJ16mCKR+NrBJYDGxyvf9YCNz+YVkBtL3
VbMtPdA+IgaPlHQYSPsDzlNI1ZPNYsLJ30kfVA+jiZd7/rxCDhWeBB3QrhByqVs9efm5gGgY0oVI
h8Q8jtGOBqZQDuEqlc36uUVp/wjcQ8KmP6IGD4PnpomeaK3zB3VqsY0NAUWfibA5zlY7aIi/xKjW
vNike987UPdPYxDDGUAgfYxf9MACo2COClQEq562W+0WYHQWyVVhcYGvFFN8z6MRaTs+55qEtmts
CcATOk8JnXMoMrame1aWyHx4y5jfPEnA64GQcQJwsM1rP2mx/CwtFz/v+ja2dOJk2350bDyzWagL
Q9tmAytEXd6fDnFPG8BrL2/t4J+MuO5oE+CmD0cnUfjoRwLCdFrlsvr7T+HU1E/aRswDVhI/qWYG
B2avsdTsoqjjunaamhkpKNlJsku8TRtfNezVrm0L4QEBgoS06i+BNAa3yQnUWWnYc4p34RqZgV+d
VvaZJRYAC2RxYt8SeHqczKYEI9I3aeYn6FOMOSss3c7S0MGua4wR/wwFnSl0batQTpMs9pTofdww
jg8YezECB4wfVBpz8ga48Wxn5hApeBq9bMXl8HE5MSw5kvZErCsuoQf1rS9igCAP4RE6KvtgR0M7
T8TKfBDWY6gHHye+0NVFlZW/2Z9HpF2RgwjgRtedLSw2hx68QlHBtgOrmMLdXR4BBsqcWbigxJ5K
84JKWEM2vPoXnRabMWZFBxWvZ9OT6y8cAYKYwlZ/vio+Pj7SJa5ktmaujKwYLWHEl4smd2DPpKRN
ehr8BLu0ahAvJsX9ULSh5R9QgI+S/XRWvojSQEmk1kYcwBZ906ZnO6zNEhgOM+0WElod7/+trlM+
EG8wdQojyRO9NS4fwIhN2BhAeq/cZHlGK9strs+7Zrzy+G753uiVfs4ucs8mTJcRQBbisG4l8J1P
xebhUgehIZPfEiLeA3lnMB7RsDxw+ijtZW7Qsx6OG+ZA0rOwCmzJ+12EZFjOtt+g9mNIGYnOa1sX
Gc/WBmfCH1qTh6rc87C670nYbu+Dcka9Q6uuq5oAI+rAoBaT7N2+Zo7YsdoB8Rfob5IFoz4vAolJ
ndvYsp/T7AftnbIF5zEae7sB6FixLklX2d4CSsAe1p86cbk1ewF2QsVGLHoDwl1r5QAgPXD5u9LX
jz9d/fTvKCu7wcdETZAhEYCDS04pepa3zmgV1iObLsbTALPi6DcO6po95F0yZ6AIXO0IuJXPJ2WC
b0eEcvoOW/t/6IGg5k1kz4k0QLLsntCucua1G12doaLQ9U+QWH6T/tMIF92hL6IGjESgiRj2fa/J
MXPy/sEd+/LHXdjB+G4hlWNg/h9afMfjbEdPmZqL7MDTUE1czUc7a4YNky4VHRJomLipwUcreNht
Wxj4CHw3vLfiXWlRM43ab9PP9tTuJRXa/NWiso2uuGWQgy0kMXb1m59tyP+iX07xRd8ZIyidksu9
M/K+3BuD82aDJFGFDx7jd1YfIwji8Zwsbspw7Q4R9Ehu3KTGVnBQcfFDd8AVl42YazwWk4OOBkIX
ufTVWhV75hwB572OYD4mDtF6ZisKaI2G0gGcL/QIfwZu7lZs0pLYChTPLObzVsTs0t0ZppBTmYYK
WXaqcyHaB3mB07ghyWs0EcdW0Wystuv/ypaYx4xvtgsdd8yXHFBzFUGzaGIHIKTV/08zuZauZ4hM
1UGvrSJxmwuKZ0lwB/c+t5Wt3EzjkJf2yV3p6zaQqxJnynhcDyUCkWZNnPPD6zw9O/iPc6yGNpaY
xR301U4VkbSmk9oPoGOAFe4vLEbRalw7cIRdlROQgvnzuDJZoJ0Mme+Ibq4HZ4+bRkhk6jm2ISvB
+7mhxIfPeu3HCUhpA44eChrZydz7PXoxPQEPvW2wXPgyfAVcNlaJTrSt7CuLjRGkmlVH6RiPzLXd
h5hNjc4Q5Q7PXMmcROQoQ2Mc9yH1UQAIVmhQFVa9orz+i7qrujmqaPKiJltss8A8VBLvy56OUUyW
XDUFZ9qq1QZdULPI9eM4vgMKQTrrM+9IkugRM1XeVBu+RB/L95mVqlSXJtP+cS2mbVhAcg7OiBV/
vO2EVRjxL7y+DmkZul/6Yy5MA9YNBuUTr+y+FtiUxBKdYcSXYjeQ6damK/shMAauP0Xw66bXgB/3
VeP5AQneUrNXqaIrMxNzGni3YC5L8eNA3nzxiFmwz87NHqWSMDPgA0qC5GSSAEJYTFVLzzTVQUH7
1QRkIYT1NQGpFziy26RM9h7MdB+Ap1ZzhpvDeZIX06NaARhkzQc9uAzFZOldSWn4RTCCi7aqLa1+
LxAFHaA2HVH8U+akQA/jXZg9crNfjtnRmO6xUahSynvLGJohB69/c9ebbnP3wy1NjVt0yXUuLsYh
8BX+C0UJpBJZSw9JKu/HQYLNBHNLOPcrlN+DlKZO4p4DOzRM9BTj2Yyssb4EuLZ0CO+NbYdB2FWb
ES3WZCPXoCLUOGAmuZ4ScBi4O4ZeXj7DE1zd1AKm1VAxkaaLgIidFjx8mM5O43MzY3AsxzeT8EY6
fIrY5sTy0rToERHO5/re4c7IA55V98AWUoHo+gg9j5mhbTudcgW3y5hTtuLE4Z6oCnkwdGOSAcnn
K/X53z1OM61P+TBGUZKOxdsVvD5c8jA0TYyzvK1HM99VSVt2qU28FZFFk20WzuN3q0yqFvdMr06N
MVLIBmoYuLsPREoV3bN5H9YC54hPW+75DmCy6mdFoRYOmVpe5a/okfu3verzpADFya7y8ujcSIzT
u8l83qi8Kmge7Kp+AONhYZbLurh13uOz/nTAIDQJfqYWVX0ZqTvREA+7TD0gCGSBeuDXS17Z+Dvd
r9aqYy2rGuiT8jw1OHR62SwarVOqWecY7/jUcf9iyupiS1L7XpGzj/xPJhYLG92GdaeKud/eZ/hD
GmBKERCkaOeFss+RlHfGYR6mp9XlnTLmLEzPUG36dViELnY49f2gyrXIumRbHMiS959OcVjjAP35
TO8k3w0tkTaQnnGj05KEiXTFw0PgDSQFwBop3ULT4JIfMHFl6sGwabGk4AS7Ogg64r7LLQdpvPSl
daOK6lrkL8Eyvf8vK2vRN6d7jAWNWbvbnPhuPucZI5qcGJ7iMgKkU0G2k3iBVrjPicKe4cCPHZUs
+Xw9hyUq+kUw8F/QhIyQJs6hmfgZIcHK6R4i5xZ2vpRGSHjn5YklzzBfpjVNUzxTDocpjJlLdW0W
me3ORpZU0++lTW/mG1b515W6RpFf9fdfH6hsgCx5GtAUXWiPhHZDD8Hw6MDPaIx8rXhy2hGGXsqz
Ez+RHDjL6vPMApXfv9qaL+6UVMdSnEPAqcQPpLD68boEm914FB8bCvJHjCvQjK2vdljACoOVvSZn
F+LhjycVLlXP4w6yEOUQAGerlHN8GHU0bWe4v+dWZntn5IfnHz3/R7TA3SFVlL/4/rKB1rZyC947
lB0JajTolUo4QAklzOu7rqw5/JM65sOVxh/UAMbSJ4nEpQsVIDlAsGaaMkhgPmIvVTmteEdZvPCb
7S7MIaxRlPebpuxutLNn8B3O8l2llC+VEr0RKR5q4aKpGqtXvmCVFfOyvE5bBL8BI+00pj5wGweE
GOqkVtzP+99ZK06/qKSk9P8/AdBnR2KUZ9UgIDMm83r9mi//+sATEuchN2Ve1Sr+OBE4jN+DicvD
9GDsGdht+9ghOo1Z7fkrE2kHdWKPrUiHebvAiEl/TwBOK+h7wrTclf86N+nEC1ALgV4u0YYqLqis
GcEVG6PvOpo6V5HmV+Ymyhh9/fddyax1ZDsKQfCD6kGZXRO4YalqxAAgkozyHN/aI2XY1fHqLGlX
qOth7nn0ne5+mPzh0i+7vgxdq4aIHyLyIgqCsUVmZDnbAHk/WIjmBrAb2OT0EgT7pI1gF/39TUgz
3pfAXAuc5jNX/y6w4Ts+ys8Y8vQjLKjRHgKO2bxxXjF2nIbjZYurmXdkcz/x76Bqtw+BUnrO4e1j
7xrJWdQZGI5v47QZU+dxjlrxYI2WgfCM38d2tLrgyqBwljaB5h/ROFYxVXLfVFHvVPBBOepJziB+
J2/VmP4QVaaL2jFP023BQ6xcM+QmAs4oLnn7octhB5KeLEdo/TGEY0JTUAYXW6ehWYBNfPb8l+Iv
xt7sC9RLUwij62cPZtmIdqly1WP07Xk/AjGpwtiJXY3YhjDkpvprbK6HxfgqrYtEmxAuHgEdmg1a
hqOd5IxqyQ/VMEICK/Khg4xL4EJ1ER3JD8CZPCw4GqrKHs0CvVvLHs2+ID0f41W+ZY48uvNo1WJ8
/nowW3O0RIbutqPyu/LsBJMK75STk2aCikERaPghrG+4e963C8rbkHB9JYCht/n+3EsM4CWJsIaC
kXSxRqs3CX2WpGG6P1765EuXJ1qXRT+oQvAeqilUyqW0y6Q7eCnCO/saHyonj1DdEzWiF/nGUwOX
jlYN6HqrW9HQKNNJVS+fVIgf00qj9EtN8yRd1b4bbhwU0vUNGU2x69eupoX/kBymMIfprDWr8SI1
ghwd9niBV4TMKTsuN1onqIUgVgeuwAeOfdNNno9OK77b/NYFnZOMwr5K7CklF5fPfyoXdRIQyXBp
olX2fclE08JK2R/94olIhhT1mda5R/EtAi7M+zfy83zbrEBIddCp3CynW/oWZxV2QdoAaSVBwyL4
vi6Y1GwEA6CrzVKASi0SMVE7MAC10wyWc0suLtadPTi2vEq4eVRvuLVURPt1ykVWo2QI6+Lbq47k
md+bgDKwQagQaOsj25GVV91W4MOMe2Y6pgT/l4sgD90IU/sxlPWW+9tQALZGoKwaSqFQ25I92ozd
qDFuX7oJ37pBAvw5DotpHt3LyDy3Xs5EGE3aotLjihGRERQJLDAQhblT26IeNtwMBvvA1SJdquaV
jVnz0HIoxuZSkp2iqz+rnzhr82vUSUWlHZqiT9JftJRPbm2y/8Ay0wexkx8g1JxWQVLI9tQGfG4o
Q3y9ke2DydvbEHnMAbbYrtITamIfblciutkCUetNqXYjYBp4h8rEZ16WhppHR9eJXquDpU9QoDz2
x4Efk0jUla+cFkWlAo8Y5wAqYCNeoO59s10u0u8ZRQdDf/eOIvyRYXZDDiIqpHI4kcjaPd5DKTgc
uMRMOty8DXZRAxqDpoKTwEYBSazRFr9HXta8orTiw0KrmZz8ONBEM5DqRD3jqDkftxcpu9zJSqwv
5ZNbDwdTB1/JahKP8Zh8/G6VWNmZSOfeyGBj6bTppyLdY7enfMjy+89+0pEiaJHQTh9JXFCZIlZR
ZbvJz0oHrtMCaZYhJyhHTi0ErX85bJdzy/UO2WnziG6ztH3gwkmJPTWxG6l3qdp6vW5qfMpycnN9
ZvugWfTR7lsdJRa6rry1j5DyS/kvp4mojQ1x8y5tWKthOKO3i8D9np93xABD29g6Yj2w0Ps1C6XD
THTBdLuyQU/4kBmtP/BUTlSuLklU4y0zI0iHU1sDhXmNcWbgdQzqC3SkbgBw81FWT4h+2gorsRu/
7ub09A6F3f60+PYDlIFNuonJzcO/tgjieR5KLQXkQ5Z3sbf5uwgPQQ7VBAd9NwXTXNc90bzciMSp
cM1SONPozbtqaBWi3JmuLvKVK9OV8+pl8gBLoXXJJlVMKZ+Hoxjpd0Sjh+ZhoQhn6Ah4mEWYhn90
R4XiGQedZiT3UO0sx/QTBqMqd2alj97kwUb2YbsfGKjA10BOogT1nNOn+z670gBfYPf9kG5zYDDD
WLZiFic717vG+Eghmfl8H14WnLCMuv5Oss6tzjomyRZ9akz9TcOFyE8pF/PhLfxk3rqn9ff+KrO/
jcmKsrZ563Ce/OoQONQnM19KrYtVATTuiEOBQrHWNv1TSJH0Im6JoC/N06mvw+TsKsgXPZ81DpGV
bzWVPXXxKcSGccIAptvmVClkPyAh3AEWZvXnMDQ0HEDWUBfPwqbrR0E6aTFdbqz3/MvaIsGeKr+l
aXmrqBxJmmN/rl0Oh1bVNemyLjMB6WNhnJJQXQyRa+/9qvZmTXV1nYYyCZ4YY8W5/sk4wfCtd4Cp
XQhrkWJxebo2G1D/ZLii07En29eOwyvpk5NLNFe2J8ITIESYDspaQdUw9rIs9/9EcMjr1KhO0v7j
68RMnfYpPQca4PMd50pad9XfplBBjGekJCwYzjii58K6Awa3lBcpX+czd5WYp1gpCNp06Ew1TBbp
2wZccvVrpoyCCIMDuTYx9dCsq8GOmqyJz7Fhp+YJho5wEVsL2fDjFoMv82Wp6WqfuFm4p2tg3BJ4
gq6lhTcb9vgvLnDqg9vFaMJhoniko38gG9USCyrL9JyU5XPoio1juA9GlEyAJG9Jtf2qzIesDART
MvL9f+y5GjDUaLXiXrMgwp0T9KwaYZ6gREKCV+0CNEfOiY6ySwpNLyu9T94cdFREtncHGNwwQhRl
I935ZztsOnJEwxgc9GUh7gRE6GHkvZexMinCSWTGUMPkNR47Fz/HqvsbcZjvqHQxhKncpdYjWEXc
TQbR8INBh7HS5svaewTVZrz3ibkxABD5Z+i9Ku6cjO9J4Nc6s6ewnoFrYcJLXdG5bY2CRBJrFqkY
r28FOXNM6vUrG6nhMaTIRyT5Z5XiWLBTfnZzBkgDkubeMTjfPy2z8tRpQProrYS8C7qkpnGCJuvc
p3DuppJAJ3rzQ7ypnVMzx+3sHe++gRKntE5abPDmnUKRHsbuxFohqUO+NP+v6IX8W1nnfTPaEhKm
bgHpDeOEa2v/jKnwky1APqQPuDaApe4LsCue8r46nHu8GlfrhqsCvKJq5ug1cUfehL//wTgd3Esz
g4dptUnJZi/X/Nvv+qOIfq9n1E0srcgE9JgV/8evSKmJEJ712HHltvcd44JOLxeumKYomThjnzKx
Y99Vf9TF+Ff7SXUXffAYoOAaRVt2y64UY8lSI9pXaDEgrB5YSrEeOJf7pcNuUpIXTcdXqCuVFNqB
m7SWaN7sMHfIusio38kxrYuCVYFuhl9/NNjicL1viTeoihIg/JUGoEv1XEbI4VMaUYfGWdtUsfpY
AIewu31rzdXIgQ3k2dL2dmgz63uYVEoT/rZ97+Svkj3UGO39ttKjOhYi8RDa2Bsw01PNrqI3l+26
81ve4wU/hw3rcy4LcB2UJoEr9F340i1H1RvZmlFSlW06RRqlpUISPzb4Esm65B8JKwOOQqa7ibRc
2piMf/lOHocHILJRUCqfztKMbUGNsoKyqDEoBqXTpS2TQM4CZDNsYOW952KPvPEbKnvDHiV20LsD
bw2EQ/SljBSl78zlGjE6eOvBfJZ6H6YwqpWVOj8lLMK/kpQUUZYrBZaA8Xr2f9ppmywxsKYV093Z
l/6TWG+EPrkCWVGnMazZxdLxGazg0h5xudC8rp8hjrRYjgQT+EOf3uCD2ruXxOt9MafjdLHg6l5m
DZVsZWKlrbejf77BWKzZC/hg87dZHkj2em+Tm6meH82/vjZnkjgO6+pr/B1dloA+nAxGzDp2t4sW
iE4EXErq8zzrRw4P3xoXSdJY+Xev5HXrm2sHW5eUgBvJzjJCM2JjMIAexHilKKxtZDRGsk8ovjT9
OotlWFgckhJLDFwv5nvj1Wfds56axJQLRmRSS7+FpLeZ0/CuH/Hy0dDIKCOUsodK6kDhCIjdXhQD
ZA0WbvL9g7JuYbGCnIteIRhmeJ/gUM9eNDuC3JJJmJ6USF53KZLhu8jtq09FHRI4IWxc45iNLdNs
ydfFWwh1pnNRkPiIfF+wdCZmDrlig20fdlYxsiC37lS4cMCjBQj14UFd4kflOM3Ji/bOwUY0VoAs
3pSUZRkCS+wD4DYgArb23qVy83+9+FKIyHimYu4NNXwFce0Bt96cv1VZofrdouStA670tyOvujRk
vKODJGxWZRP7pK0dYCneUTsNLqb4/qDvf2xRLMJVPr0InQ1ucavn5vsCRbKQT5tEetP8rorSTo/R
snAHgQCRAz+vGfD6JfNexZ1dxbGckGhfP/Vp+6SC/bbjril4+sr7ywe1+oHUCTaLiLivYc2Hn/aM
9AmLCiMPoLRP1m0aQOQd64UpCJzJkfQBs/I/NB/FjSyzwsK1DY3/B7l6cemyCcmQIAKHc+qp3Vs8
4+5UUXoEg4DcgG4giw5Qj69HMZmPIRVJhwXDcL2VYP3p0xpTjAx3dJafp05azGeEKDsv+029zc+V
npGZZVSe1ObLjnUTf5RJI83umGzNgh2Qt4QKGyNceHdYkz5U6bDHS+hSdflBRqbMKEx/KiG6JOqO
LKGvS0PvMUTOTzTUoj+McDVn1xZjb2CJ8kAbVocybFVezUeXYSbgcZ4T+Ax/lX9FimvrMHrmMYTy
wO0VB/AnKORp1lFTTPf7mwSsJWqseokIrtIHJ9kpBAz9wod9b6K5AZ9AssUQclbNUv+I1sfsx7+Y
Jqc33WnkIAxnoST1NJrW2yC6K6lmV2LNCcKlNjTaAPpqmo1rd7cP+Ho3KiN1BTnVoiOJEJy6MZj5
5lKKSKmQVVLDEqBe42oYxsuWzsngo+9qq5YJ81LgGLkI1HClNWfB9ThVrCicrEQ+RTnoT7rFHOwF
Bqqc0sYePCTa4cdnZqff9tcOp8NTcUhIOGAjc/JuyACZWclrvpkYzniRDw/JJIbZm1r9Es34Hs0m
p1WG9lUeSM0OPBCjr8ANwAxEYQjzU4dMHf+ovOmWL4l5HnHbgsNyzxoIhHM0QchhqzK3mbDsdV4N
XbOCXGuvSE6BYem1gt1gGbMw2y2VXdooXWf2/UgIhicH0c773/0iH/Ss3m1DT446ACFRUcO4w7uq
d8QvczoQYe6v3ZL0gD99Vl+3NsIx7TCj80mv4WiqQ2L8xKOWFn7eP/c1os8oIjjocEzXIO1yQcfr
dSGHb3Jsy1QZs/zf/dQFPmM7tZCKq4dpb8XvegUtoIpMsTicNoS5ettYV1iOZdbcYZqQc+11FMwt
Fm5VkZQgaDoo59rKX+KeYeCUOang2dlXvoSpus2DVLs+dmO8MJLRB7tCjJm7Y9QcU5CBRiF0PTUY
mmwN6m9g1LKHnFCG6BQdlaHSFMAz6Q3L6NfcbEDU11SHwkgVNlagzTRmga8gmfQeG/l3u1vzQQIu
364bKF6VOEoiGrn7pQzjN91nZOTRK6Wdu/RmnERUrQnRFoq1cNwrtq6a9bCyAEodOBoC94my9HtB
SLyduB1q0jH+BKzZyQfOHWq3MnUnk05phyR0DaVMREa8co5JJmCCyTx2yjEVO/wBIE4DKDH67lqG
I1CyU5RhYaOpowFydqW8hy5BOcQHoi4dRl1wFYxjZRs8MQ6fSQpfeRUgzJakRgGZt6f7ASR2SwTi
1GOxP2EX8xf2ULDtNA+6461EYc7mT2Pdmb4lJrDbgxy+P0pHkUxd8zg4L/8WzdCh2v3JiB9LZ7X6
R1egGAt+wib2fFlqsYtbwEC7ZPaXYy8GTh4rrUpiuacdezA2VxSR4ozRfw+4DyHqV9pacULjBaej
RyCbmWllebP6U4jhYZio4JcxK+sccJSY5VOisruMhSEd5WEQRUQdIW+X9a9Xtc2QWFjYoyAS4cwU
9xXG1gW9e0P2HapJ4jElCBJ6zKX5qhrbRGHKp8DzdUAO+kXfE8llgp32idp6RT+thzNklCKevIjM
Ki6OHSnZuBKeckaSTAdkRm4ekEE6kiFjjRQDv7hWle8zDsE/7SiQPtW4Yqn2Ox/8bhgMwtc5GXWe
n6bh+UlwhaGTsUsMXNwYmdEKScc+/Fu+qIElIfb0kJZ7iGlfVhi7L1h66HBLWVuoflkqyfU/KSPR
1AGmH5v87VvbTkPOqJlsW+/CSsOuKbYzf9nVPBtMWiLbKl+/zvS4yuixK4jKgEbBvPNo5QCr+B5H
EI9minRGEgJ04kZYMDml0BWQ+BmFzbrR/oqWCBL8IxV5KBPpr9FCnaxZiqzBq7zdGzW091P+Obk7
BiGJPorKz8lakIY1ug40Y55y2w2TzxuO+azRl6HN7JpRR1bj+UvJpbxvYioF11XABMAj7T+bUmEU
ngJhRxKTpjL1qoyt8gOLyTFkhXFwVJ3D7VR1F45LJVRcvdJcHV5QqG4cD1HbOoX3uneOXxQTsxFF
TAuO967flYTSN2n5s2RWn6FO1FiSdSnbPEC0YcJDeFg9FOouNevn3cGh94zx88B/Je6pMeBSS1UY
escw+BisHQr5LMyBozYAbkfh+3MsANkLy2U2txaad4qsCUIuh/ZKzEr1uliNZ29kdmOUfg50I6y9
Dn7nn/hcqEplXTmNYjBrVoyVq0R8RqhsGEcMC265laqETAF37bW3tE370QTwqGpLI68aizqUiS48
eZpYtjC9CF/YW4D1ZsreoyyZzNw20rQGvhAUNe18EBe+SQmiwnM4WwBTkZBYAENV8krp4VNxAilF
JLC0GYqN0E/1WmxddbVjkPvTEOKlsKVKtIMrsYnckev6g1aUyscqeECKpDI+d06U9A9S//AQQ2DN
0Wz28EB9fr+ApWoX3fRwgqirglxLsUamo+zSIJriiTyMH/CZ/fDP9t7+Ll9m38thOZneHbaNaZoq
0RMmTX0N1L7KlVXHCEr/Uc0rfF0ZxQW2ducT6YnSjv4WmbdMkte03vza8IUD7zZaQjCBO+Vzl6oG
D+IF1tab66/8K9wQaFMAOQN64hxduc0vBBynPrREjQbbLyfGD979NgLhRVOAxBeffB9y7qDVnpYS
mhqph2USVStbR734Ptk1YS4OkM59DMiC7sLJeSYK8jWdwJpSerYLpNnGmAb8uD85VSRjelwQHlgz
Fy30EaihcAXNiQaDSdJrFAFevfDFnhUGtVXWPrF9QOykngwsmDQ4R0AhMmkPc0dn56W7+EQ/5ROt
xLbcLyk6EMKq1EnhkPeaZIxBweQWLT9MbUmZjYG8FdotA2zyHoKVTyJXih4eyg9j7TPtCUyS8lwx
2qWL2BBeF3kGgd+cl6lG6VFodJ5atRlAAcUVCa6nQ9jI496ycMuVRRNzAcXpNiGG/A5DEYXlqvmA
9C7XzVN8vq0vndCC9CGqn9S4qvtKpO0T6kIdS/o9rd86yWednoB3VhxNUPRPwk1F0rOVFPFlA+CZ
9bJxr78rq+icPI1uwLmS+WZp8ID769ifmM5pOeVMYg0ZuWK/49mDSdOl8ho+znU3elbELwY9dN7b
p+qrgr4qWeHL/pnEUUjixmxrAZqTtV+2+wVWUv8CyQD82v9fxDFQ7fZTBFkmjWbTeg1pn1bGW1sH
rbTd/r9snLopckrjJCb++ihvvV0XMqZgv82twZMf667Vnr18td9z6ww9uQeV0IuicyXY2kaSQE/x
bWETpOWtoaRaOsiEo8G2tqXkK7LMItxV+6vQRgvpAZp18EljQ5ptcilTnYM3S/aE16ckTxcQ1rM0
ZhjK0eOQpD58ic4wVLnzkUK9kRbwMu0a0Nb4KgnnumQ/qj9CSJ00jawSr7a6DrvHtipx08L0gyxg
Uhyv+bUfBRaLcbE8Z5LqBcecSIFNer32Wg44JICn6U1ioUQVvMqdTKgsXTMZwd/44gjJLNV3919p
L8EJ5oGJu94NpCN+LnnUclFSDa1xi0tyJ/raUaSi85ECQ4npLmvFrf1Z+hlXpe7isVnteHh+Ta/n
PV1tgBYWAzYQm5JY4v4FM6nBODKxtbJMWdGPcWymdkVUvIJ6PxRTyNvmkRyQJQZmkHvw194GRFcv
UnGOcrcG3GK52cAlAzyxrWDCxuW/VuYbqI/FyEnR8J1akuOknWxqsup19YnP1QMn52Hj540upBHg
WZmyY6Q7Wp9fhgqaqlbgcWJ/aSwsw4Mpl3sVSw2RMBqYkNgtdPXOO+OZr19PYyRNtAJBSU0U2DVu
Qv8pggLnpuL+pxKW6q4S1KFoC+5ZMV7H7k7CHca8IkYqbI1IwpeFIOYkd4nhDywh4Qan4MfidKZw
9JLx9JMtlSKOHGtNHF69olEeziI1NZUzkxXwxosJu7N23K2W42xQJupevNiiXRSALPsCeNMAJnDx
dHW21xbC30ND5nWOb2wIIV2D5SWaQxXeMRR2tu4XTew3BGxkn6Nd+ojPPn4PpyyIem7YdXiCA1mV
mNBOY3W4iT46RBSVUwDpaf3XJXSp2TlUEIWDWWyQBkmJ7WfD4vvvv+PXUtOKbp/rxhXGCQuO3R0J
zZBhHqki2TXgq9CQxZbW/ygndGWVnsuFKHqpe5Zel0VyuIHuGcPli6x1Q4py2y4GpGtzbRh1Rj8B
2BRUHK/GqEAPOlQ59H0JfkusP0wZ63Upc6KJs3QYgbyBst5OF2caWBslRNGuHhgIwtkAboXQ9IOG
UBvA1xQLP9xcJUt8AYOz70y3LTeNqBwACfjEHrUNGQoiC82Keh9GwoXnS1bMn8PW8UxawHdkPbtv
ULnU1QCRYo8P9iyUqdW/18wTCDMFK1+piG+8uNBSIPTZ3KUeDNCyUfYEonu3iiVYn73W8ckSbWi/
H/nojtmAnDr4s5e30kKwiuWp4Ei+AcEady2QfAfdc6GNcI5yTAvg7agyZ/B/NZyOZeVYTISYDiis
upu3p+pRkOjbtpQ6bNWvx3xc20IOFGPxy8rspqinwCYR1eXOOVlbNt9GsCapkLeDdTAv2Tw+xI3H
Iy2cO+vFljMESX/kJiptT42YtdnuZUheqt8KKvG8WxzmdofNcpjX0Cy+Kxf+Xdd0lZuqLjht4JA3
pUxliC9CQtUeIhKNa3uHjYcT7kOUiIzghBLaeyATU8IvrOHuIrhXKg3g5MYnZd/U3ntPWCVoUJJw
Aq3JHgF3zlvFxpN+y5sdwNFCul+UcH1AcPJtsSvEJ+zevx4QH8J3jbMaPVQexzpEZ/GClR4FOaGj
oQ+kha6Y9yzPFA8MWzdx4TzdzqK5d8L4VgRTfmmjZe3q443a9XtqginHmSoVrIKqq9Flh0yQsyX2
XYQs1a7h4ef1cMBEzNw+dR/XgjeNyyjrZ3+EW2Y03nYiQvG7GQlJ2Z7t4nR2OE+B1XF6q1XWu+tD
zhDawZsoRmwA4PAK/COnR63SobuzWH0EUcW6FQpuv9/WG+VkXAWBw13hRl31M4IaV5N2nKFiWW0d
ML6VFjzt8I0PYbawA6X4zew7cwZjPjNHp5dol26IoR5KrOM7uYTvGuaHJn0rOnfCxkB3jpyX8f5N
uMAU5I3fTSC+6+mOubLPSUwVnOU5KeD2reEUeqNVurtsEfm6Rs7KGLCKxasjWalM+KLcmXtYUpYM
i3CW62RfVtIrRR6ET0z6IHqoIUieUMcfoNlV6oIrKqecu7UC9wYkpGxm5LpzVQhBo7gCbRa7y5aQ
IkHbpT4LXKPUaYiV4+5ZtMWraZvlhEsEVOPeWTHWEm6rSZlRjDZDqgifixx3art8o+bzIzJAudMa
Gv5HwYNuOLW0icfFpvZrVoBJFH+71rpqo8LtIebS6hqgF8RdPYREspi9La7pugxavPEih+lLYq2m
13DabUjAXRESzZMfq4HJ9f2/4C0SNNTDpL/D4jRzbFuzQIrGem44D0gwnHPBSFm0IGrIRWv29kfj
sNNWSw9oJsz8YsRYl5M4rbACGKqRp/RrPOwL6pt324y6WeZKptDR0ADOlYcYsjOotE7dSB73i/8v
p7eNR2O3l0LsSoomc+Yke1HUsS88lazTubO87mYQVPMouhNHSSBZBLfgvXX2R0+JnNl7f3kGFWTx
otqr7vgmj5XhhzhYw8dz8KYhaB1TqMFNZZ0sB2rAAF19fb7bAZNLMqmRRswJvnOvprTEG7ENC935
5ubjpbPtBN8jyAVJMaW0wpfsjDNzLC3N1NmCSw2JUEJJttqlgaZbzgeDj9cChUo2NaCTIwjygvBs
2VpzkQz03+lySKcj14GG7q/n0UBabNbITt6A+TV0vnd684tQtJPc4wPx4+3togMxwuUmCcE6CY6J
p/2CT6DboLJvqxVqVkXnztHDmAiJD4EbZQTnYg3HZ1gIwDlzjCscC1z1QRUe1VRtLOc/+l9qdnyJ
gTRCwV4g3/ROGcfiGB82cIzmowiARdM1oq5DKqGiwWDC7LxLUMRdcQLwPytSI0HnAhgkwTg+OA+n
3ih1DbiJ4hSxvqHliosSoNoAAZbHeSWbmF78HIKO5idztItA5VKcBOwqJqoFqgok2Z99Mc2Zu6Kg
JuglLKnSLKTCn1vyqgPnOb40qv5B74Y3nUF34On3FB/ifd0PLV0NoTtNSixUY8I5da4mZyh2h48N
SF42GXYP8MM6aEt3Wj/NgHthSsN2/IoRcGI1+GBdtkMICjeRuGb8TbGtJdbK7W/Q/YszLCFpkJRh
V8qvzPrpaMLZMlo46kIm6CJpeFJu2GU+llE9k2oqzOGSQ8cZH41p4KJczX+XppHdMAi80qnMWBuS
acLPvXWf6dF6+6GG1lREhxvl8XamHrrbpMzjN32RQyrLLR1TxMEgyQoLJtsE/wMRIr7xIFt0QHox
/lgJsfdmOHi+G1GV8MYRtl4wz0EPdekB9bmRJmXxI7/g4sw7o2anrnSwHc/Hat8+uBRmPCvxB9ja
rfOhHv/nkbPlqFjw6STrjXcPg9TxiQw8+xUoKeH2wF/xJWNbYfGHk6GROg3a8H1+9APbvjQoGwVx
N7wFQD8HdAdVJdiSBfHo+i5snMEO6d1Vq6fApr0b7WCEufvkU4xSDFGXahwRc2PaynESKhrAZJMJ
4CB+I7cKtBastMIO3IlPbgdFCeeAPP89NeRujsD1cbuskhNmtWRT+OS+QWYbawcoG6Eo8frOkjoA
SvoyZKecDriDIc/9vlfpnOZBqIoZGPTU7ah1y6eAJO5XCLxoHURq9ingNocYMdVSLJHINoy8A869
O3QrvyzS6peagubV1KWfFlJZMMlyO8qjgeHWHa7LnVaRFzsjVS6IsiCZM5ieZyGBeyaFiKRi/xR2
AgQY/+6owBTxr0MG6rUyCSTX837n7A8zuAt0AVE4HoNhs72dhgzHHfVD2ROxXECEWNDVaVbpeVpO
+qrqJ3+eD91R6tCS8WyawhkyKvMLWVB5bJiWmB2WfI4NxbEffL37gCh6rc9Nj/0RZklypATUa3rR
zeg73DYPYInp0muYTXI8pc96MJc5laO90duYI+lqMIwagDjmtHm+f79VR+T5eQUf8u8I7VGp/r+l
4/xhCtJkzrUTuRpMakQU5bSP0Z0vm0hYGqEHee+h0DQtdNtEsEfNdR2gF60Qo/WmrZjBGij0kmh6
eM4EPAXU5yuevUrj6x4hauoq7j5+3Lb0rh3F4AB2o2aw1rOmEGCmVmIW+5C1Rmq20kCebBKjakgP
KLjjUZjopfawZo8f0DUBfjOXT87ciL/zKExiVoRDbve5vscToXInEHK/088AcxnrcS0YTkyzxrLH
Ho+5CKbDbEzndFyBKQgl8AQtux99lgpyVzHhjuG2c0FMyNn4iZObPpJxyJWDv4tRY3DmT+TlzrVL
HnkFO/Bw3M7yZ9ze1Lc3HQUUo7Vg5TL3UYrRXEUPUVsig8zUC/EY4ssHTY1Lj8af/+hXKzRacgsQ
afZZ/Zmeo+vMHqeV1fBmvsJ0EGL08VrN7E2WYauyxSI4DQzZhZduk1RME4/wntm1+0ePlzWeF4ms
0+HbcqEFpfFZJrzUwEd5USNvQEPel+tebM/HZhtuZr8wNCPYt9yaCdkIzIVVulVapNxiezYczQij
lz4DsOr8Qoy/pXKE41syAhZ4z6ns2wJ5YHhMrCmwOiGNwY0kizSWEWTWGkQJ77ld2yUcUV77XWSz
erL45NiT2kpW1lrYt8YejQBgwNt2C85OvJ1n74epK72T70+df1MQV0eHnti8XaKYzOpsOdDZnjI5
yPRiS4D+oWW4UlZx/fl+Na9CJjMaLZjy4Q1PkMZXCW9jieQdrO4vRmqknzBFmUp+iSnrNmKYIuPb
e0xXgwyOOR0Z9AlMlqlzOFSFF5FvkYHRe0FyQWxs+Bc8Y/QYhgIrtniAx/y1ORAdcvjXTtIvMQEm
p0GABDdQL5/H01u41sai0L3vWxJ/kYAmCbF5nmqR6skMAgdZf62JKcJVTXv+X1CK2h6fQ6Q5ltPU
zGTLwEb+/7oqX2xCm56itVO2utogVI+4sEsYMbiQ4LyT8O0gGQPFNEvaOxiP4MeFW/iPAUl0nPBd
pORGw9bNDaJGTHQE4CYoIwwKL+qTDouFmxhxAZ7Ph01l/cLcge4IcJbqysNFRbOvrj15KRz8sbB/
8ayUABbAYhvrB6R9KZFPVfY8jb8Qou6hSqCztHwZXorJlOpUbx0egUv+J0pMdIhoBhERCe7bYu7B
F87n37yClttxwgR7db0oKWiPurMNu04Mj1L1xgB0gz6HVV7DIR64j7XJlIrOaeo1Y6kfANlE50a9
Bh8Nj+odyfojkF5HbUnqw94OzDi6p76rpvDtPwsikymVWp5WwSnQNkn+beJWPjrIlF0/W52qSuQB
35R5R54MeK2Za2Y+gguMd8lmYg2OoqYP4amennW4GLb1pM7IByquuIgSwz4/0VkMHJewYvRIegwI
8OxSRqjExdryBdUKykdxjzTCoTOoFhuFsw+XyYC5HGTtQK07NYvqbQnR+pnpgZUyVSg4kAMjaNDh
fNGofYUDsybf9iVMhXdPu4pUUZRFyccFeJuTvFR0SknpPkPaz3+5SFmHVVrDvz+kZ1Fe1HsMBgN+
csNJhtKP5xyULCFwIgF7yehchOft39Si3fQchi0STGUAUhj7YroTN+hqX0ZrB01zN3E5NZGMXVAf
E4XPedn7udpDGdMOGTcqUq6zloySXeOirKQf53BYUOqORTmg07nOd/F5HpY4hrkJGvvH2vWyZ53L
IUvPwArrHXC2BTUHTpN9HCVTes6ksRrxo/7FlUvnAoUbPEqeflmRNA2EIM2htSRWEC4gKVh6T/1Z
G3SuULhHaoj8vXPlVdBvEs76z69pPAZSimnRVhuCzOAEwdR4/hyNmbpWHa/JxEV9jX2dOQM+S5/p
Iwhkhq5gtTAnviL8qeyZZmHbymLBlOjOqPwOWfgeXVS6/wXGkYjWFdjIvNp/6uSaX2BAgHG2eBqS
GAXHiwDxDh4A5YvDo04NW0S06KbvmstEBXlK8bac3FZIQ5Sst0m3PyJDT7Fl7mAhyDbU58ZoGjC6
dmoRM23L6RGaNV6rGMvBXGtmuetsleJO9tvjHim4wybjjpFIMzLKJQE8WAf7wTLKuee0mKxQUyQz
OY1KVxneW2CnSkEtNGauMIXyCgOn0EVQyVVZQPRBrioIWTc5vtnN3tkcwALDtH1dU9Tp3t9CAxk1
H+ItXIepEbsf2omkSPL1XsyMoOTNvf4qqre9I3KeJQlG/ksHtUqMtPFxMlnQfu816+xXYPx4qAMi
nmYunxt1vzyihm68DaoECZLE10kmp/IwU5gXJPby+SQl6xueMDm3NDqC+54w2oa3ScXGfiIPVD2+
Ypo1pheBVvMZ5k1Mw9MvnyKSNlHp0q6iAwGZ2rEV1W5MD+JrM44QejrxyRdR6aNrE3rbyhe847ks
uN+sU1xjHI+fh2Qd/Ihd+++nPYbUiuysyqvvYKTZL+ophgrSQNswmv80Ylm6+6gcNyGjkEL8CGk9
YGLCr/mbFcdkrX8jF6Rym+8vzRDcxIMYY6GGIVRIXXoge2SF/Au2bX4mfrug/IwsMVL0bH9vS2Ru
dvQZnPfSxxYiEzPMS8q8PlCCYPFxkQ2M0AkwWVZYBKwPAqCZajEmarDR9zjWg/i92r55R+jxaNaH
FVHwXo5TKTrm4Kvfzk0rLB//a026CrJutz2sygNYQdeOhgjgMD7H+Yu/sNt/Xb9smp/e/LgJLS/V
N4lK5FuEMRq94La7zWBh6GNdW462LyIHFzSEkPA6NeJqZYd+a5gmi6GOhimdSxTD4MgCusg+NuDc
kOPHZL/776W7Xe2Ne+Phbf3yFCs0WxGPHEEg2MfGWgxsarUQaAcM2ZzXg+KzqaecoE8bRe/lW4c+
81bwIwgqKSKQ4vK7jWE4hnENdkDJuCbeY2aJttGIyaeFfaDorKLCQKBHN1ynOR/zMtNnfiPBRaF9
N61FRwacVV4sYN3b1wS5HH+HNO91bAWemNIRWJm9At+7suSdkiTRqTu2eYlIEKmPvEwdcCPkt5Am
+8Tir+NYr3sU4sCMsf5/J6Y8mH5XvIhYHB/0LI/XAljEJJl4LRq5kS8TBoL9RW2daYovPUAE6jFw
XtxBicAi5zcWhiv6F64gw9IMntyzf5NRJN3a+PgjvMe6sjXZndwm+1BpG4GhgVk9+0v44CaFTZ9W
e8/mJK6EtGGuG7TfFbDEIec0OQrMrY47WU2+YdAqQR4r6Df6GFo9BTMEMxhaeq2B9x7tVTCUhN+p
rKfN8CWSfszVIDYWC8jSVqxK/ZDiNSWITr0MDIMg0A97cSy2BMCP3EwAoZo4jA0BwO9hjXQdDD/T
pQkk6TFU3op0cWzZo80GCwKOYM+p3TBBXkYadMghmifcheQuTKJuU6JybBYS7yS2V0YCpjmRxrqx
tEBXiwxtWI8SPB79QzhJgCk5nsfDkMBWy3s2t7QErUpg+A9+pUTCtJaVjfo7POdWoTvYjoB+24Sw
2cb4v+Vtkq2Ts6u2XNcEueVInfodGGZEehiO49o5LOvkhY+BDuOcqoQ3blXl5j0FJwE1aFGG20MC
Hv5X+ctjHo6RC7BBnV4HHfoUzbD3gWh8kk4oqNVOIPPhOqn1Cz1T7f4LxAP6GoUZ+MDDTX4Rh6d6
ia2TNRFJxd73ZzaFZ+ASodFXE+RqfJgg2f9STOHYL6Jiwx+FNUykcXooHrxHzTfi3VGJ2qsw766g
WXNCi9NsH/WXlxJx3CPj9FWeBsPsiZKaLZFQ9+II1nyL03MmHz0ijdGEZLxdn0gKA+OnpXljnH91
XsligRqD2KvyQjwLtD3w8vf6FL42PvTmRXQx/I7s8xCuxb7CkzQdSujpElp9jTqf0SHkPE/XwiGH
Osod3OqDrQ1kzR5bA6n8IpRkiYVVAbRPotUjOYwnR3Io0RI6eYoOKaQrsBYbFr/KBVgsKsqjn690
lC1USu57LhjafHT0fj//p20AjbUoErZq4aHmDyexirai9W5eYtRezizCWCqa111mMrRvns6pWYvn
D/XLHweFW+MU2s21wo+X4ubYC4VZbNUQykKIXbxoWmK7OAhL64SOnUEsrmo/tlG4qZXhmc0JKj97
3KZM9TRLbrFmtWBBMDXDotCato8Fo409xWzRXbnQhBSxiEAP0IVTzdIsrG81rJ77ZkgHXTmk119V
O/pg68Y6AYC/AN60HkrqSs4SjmMO2PcN21TYPHjJ/3kR2602bB7qTROJ0DalG9oZciPXEHWkHvdh
eeOzbezIOyrS/mGaIt7yzwHNKMEw6ssfjWlillqCJKLApgsD5oPXSoobUveCkLEJ2UEXmnzvEVgJ
nYXu/+xJdqYmxQKkNnU70c2pOFT1iUyOLxAZ6mZgiBuMU+nR2huxOkV9+aDo8l7WnUo7t+UhCmnD
NzUVR6rPleHMGsy2b/1SU+Rfrix5siA9uVpiDdznsD2cJz62tpeFKrJsx5TBvDm3sHR5hc5Dw9h5
IOscqsxTIcUFTgPgmBw2GAsxcl9zBm55VrVX8d1++VTuzY1PLF97c5SHgbKupOV7VG/qO/rN9olR
GP5mxaMZRujFmIYRXIDROkF/2SzISKH/nkZAV2PnOGXmMWpjUriqya/MRvwWuNC5x2rRSeY9ZRTW
HzLKnlgJ9EC/2bUnhoG/nxvoMeRlG/Rzkxk0qkb9PCtVp0lTpB8XJg25TKCzXPPq8Sp3LnWMo6QF
VRyR2E2cDlyNZJHgk07L3li9roZ/F6oCK3ucsEOBtgaHdnbRZqWAZIaaGquqQ++NW4EQ/wYcwak3
tK2Ap55l3eC3bbBaooqm2k0Ovs20KOJi802gXZCEvjAUfs6aJD23X5srDFlJFOoWWAhauGYMLuUi
MaTqzhkUYCVr6WYFGnQWiDNmVJXolqG1WpbQ4TIlV7ZY2SoL+PaYWAMzwwNAJ/Re2qIlWBXbDhgL
K+ID/olyxFitvCCi0wpLr6yhT5D07MwcmWdNjbHJBBFLaBzmjZ03H/ERyQGWFFMJ8Nf3bZV3uscr
YF/6462s6AO/Tj8XeMx63ZQb/wqbTb9Dgfke5Ku5zQYi8SDPcPM2A4+Zzqbt/BWOdTHByf0k9z0a
+nDsLItmQPOy974044fuCZOgFtocPoWLmy+Qv5Zg5tGUGfNhLPYkNr56doiMBm1AIqhaWDn1EIZL
5go+UnD0OJ4WfHIJQngA+aWryIstLrdhuQWSmzk7nnO5KlQYa4BDVSwEj6BB+mCtKPbj/CZpXfg6
d+LDTtGqhrUOfytqyuU6HI7T2c2AlZ62GbBgwkpBMjTLDn0K9F+JUWfFiwcmPm4x0wClYdE4KLWQ
K4H8GRPXEaFw0PaL/MfW96OtYDmM8GC03wIqZDLlDOS9KiH6cEva7MukRDP7WaNM/yc51KRxgGa1
DMYc/ge5rEVnSvyLt7aYA2Rk71kGm4ReTdw/QfE5Cy6JqjCwItNJlV0yaJtTHFt62eaEdNdRAibc
kqNZeqOMufIvkwavsro/dYsv47JQymJC44dHKsAHzkEuuEn7JEDh8UZQuyjTRyGKF3pe9fdce06p
ohx4okqI4MaPlIcizjfU06uxBxILPcCUAQw6/hkc5UwdDt/xtsP9HyMoIyrHyN3mX+yPh87OyfjB
xriD+kDUYDzp7vyQQaBuuI0r8GxeWVJt90C/bpdYF6s+QDRj41WMeSLckirTxEQGvueGjoOdFuYe
+dDrP54DMiY4lCYM75M6WsVUj4S+3wO7bqEK8nFEYxanjs+dEUyxFM6dmouvwhds92w0lwNsEDXI
4dHcggXGeHO+14+CXpbSPc5mJDRgOjnYj1zuoiYP3f83joMy/zSKwdlSsE+ZQx7ab6cVPqPATD3C
NewwFb+b1VhBRTNKXM4wK/Hw6xI5/pFgMgRw1bxI6RDbhd1HMRuS/Y6VNkqynRXVIv8qN45GbwGW
dAHdrGGJldpsFrewUlbmKoJjeHfrKgjxbDS8Tm4FPhmizzlJ/2HnoP+v6Y8UjD3TUlerSl4jF/LF
0MS+DhCtL9s6huN/xSpY+W2zglFZ1XTBv38VoEHprsQGZG1g6+vMT0sNg1duXaNziLQu63LIO3Fo
7co/FNz4CUMRaQpeyyFaBbdIrrmZNbRA3IWoEFzw5FjPJCvhVSR/1aBQefdn/ROulZHo96H3pWTS
ucyIDt72HkD4l+NwUakDXRlewNFrbXkFDFjIgD+4HqPbBxUf+C/PNiI4npo3/dzIoG2u2lQmr0QM
msaiummJ1Od3rZssAiQfBn58xlkM274cNcySYL71n0CdTtyPM6hTegau8NkcWGK5B6Y2UOeves8J
MDTwYNkteE/3f3Ghh5Zj8VUUPqLWDaWR125NpUa40cdzOpXvOnn6gpwFTmWZsZPL2FdYjv6GcM6x
LY0tdsr9YtA722xCOz/m1nVOv1kt6HUIq7lkylP0ffGzurk1HbYa+kMf3C4725qyteHqN6HNKdUb
nmRx54rAzw9mZnrD5gWizuk/YIehP0aHV75FOZvkn9iwHmjNACR8gHCFNZZNZObykm73CbaRJPfE
tCEwKfh4eJpu4DsYx+obOGJP7gP0F+kIKuQqA8jCdSbd85L9PUyya/7CTraUywEWwb4grdpjVhly
+8QdAbl1s+3XYWxpO2tGksTiyaNzltR98vXAx6jksDqfSXt9qn4SqDZqUN0dH5667LphOY92pAzl
ZEn4OL+ZcRQG7CWWOceSBLQsWtugw6laPOfcLSTu5/VHgqQtEXFPxqHWKmgagJfVzCb5lCpwC+yi
oyQQk0r5U1LcXp6+esB8BeEkeX3zNgDOlTXoOoWfib5q4pOlMNrGUyidZNW32zHwvpW9pV+Cd4sj
YBRxB9LYRevdqSRHHufeNkyW7u7uSp62XwtzNbtTlCGrq9hugq6Htwh7lXT3Pie2vLRYnN8yPMr+
mXT4/fgnPB117K8tgG5IY/it8VnOkY2h8IWebdvN5iC1nWmigoCSFyjCOCR7zGZJvJctpqAPxeV0
EsseB97kft+4L3qZvI06wWXVhqkQWSFrQTP9OFWBpNMcegqqe3HDmXLNZheSr/jjBdQN9Zwju7fn
7BZuaPXxQ3pL0uOxZCuHtXqZYgkqersU7/Ccjd07q1XUbiHJY4HTQdGHWoVMS7sYJm0txNZZPSf+
SfremJcjKsx67rBdWcbS/iCslSUCYLOz0E+4IBtavJtKvnBv1Kzclc+r8jlkK8ej3GMwVdWmD4bg
JM5Rdc9sn6BFRrB/aDaaUEFG23LBCyddG+9B8nj66anfRyw2BuOT+qaIN8jabVuvyHoDEDXs7vG5
6zuLbSwdrekz/WTOoLO5iYu4VBiy/K33NtadfMk4uqVnfk5esxTvncAw9IIXU1j4Uk9N4AvsfCyM
QFDK7fbpC9A6cvWNHanDU90PK//6KTaNViISXL+DAXtu9KlPhsobvrgHUoCpdUFxfYhHT/k5kptX
Z8oquV/UdO0YulH03WbEI4kepvRJ2/HPnqJatLnaFyOJy2HhHwokhk4deLG/BqaSpbXHla76RSPp
WrB2xZWjdU6jvDkTzHXwnCHecGWg3JzrW7Pdlk9vhSd1L9LhCsQBJa9zIhfSNgIAI2EOYq/+Vsnq
4JmQN2/6OY7wgoJOjZ/c2NeZnVVw/eqAGkxaeHi4VzGWYO693IqfMgRTZcFL9ZvyjYWQD/pdFcdy
7336hHHig2dKBGwP5fUX2IRhNDnQy7pEdCREsmssQom7FaMI1xPs+9kBOZtzsAWw8AAsdHK4sSLS
8HCQauaBGu1XrBR4tvjOd2BMifpdLPgurJPC8qztSQufG9Wxw2mfC5ZCdU0EeAEpTuCQ/4+tAb0q
r0ssjkPUgrVeGwLWgoEo7ID6Uxc92ZFx4+6dM3+6hrcI+7YjhO12oEiEYSOkCafZ8lnn5Onf/UXT
fN7YQq1Fs6jZ+LitSMRIXSbXRHdHsIKA573u6tCYhovIGIaH0RdR+pAiij16HcGmMxQQIWst/hHe
O6D7CTwrnK3ovaZVXqMm7mNqETmXU1bbbckFJtioGSuj/gj32RKPtaRfj6f8XxFeDUs5P9auQ03A
yEf9vugVo8x6Yq0tE9YPhiUOk43oJTjhDYm04hEYLPzG29ene9GpbNWZCJpCW4Y4cHK2NgODDTm7
h6MFxq/j+LesNGVauidVmGb13+s/ZlTXLcRtL/NAkWzYko7DSnQQ6w0RCBcOoNAdK9HpfSFVCG54
G1zFCulj6QF4VHYZdGYTFnzxytzKP+PVr6Y2E0asRNuF4f8rlp4UzWO4aTxYWgrLC6/2leafNINH
gbYZ/zOGsor6AZf70YMUCJPyf23TQtb0P9wbmRYNZhKlQSS0WJBtdH7hKBz0nL69lKeugMrjvz0o
JDWYjLoIffTZ3i7j7wFkVJopShHNHSpuboUJP4tPOjOyuB13BqgjedvLuaqu7ma+q3KnBAr+1sRQ
aDhpuR5GMfu6++MMOlntGKoqAgBvusmFa5vbxr1SFaV2zEEu1QphfyAWyz+ygwbpqlm38cTP35pk
UCZgJgVr002isQx6DBIK1XiWHrMKsig7fBkl/B5Afw0scNTfLerWT4DkU2CeN5li8p8tnm43S4Mp
q0PMo7BfLDS4hnm8o+lt5D94vlvDLpIRH+xM4KLQjuys+t/Ruv3kAxphv4QJkpW42ibadaHYib4w
P9ONm6TmDGxlK4Z5hZv8xuXuQh/KGV0oG50Ugecum/UAZr0X5BdsG5aj0bU32TqfGLM1pJ86S02S
oNLoJvH/AtJHZeWO1E6MipSmFBR+XzA8Mq6W385EDoalkeTNXLzOLiu2i3INdoFKE0OLqTPXgpeB
+3XZvn/bNBxE5KV1rrCGV6cOO6/ECyD67KibjPa9mNH37RNRP2eYF6qLisyZwyUqCKzZfDtanvOi
oAl8ZAx45SAlZZxyQSiBfI3tji47npcsM+CsSNgAvbrw553zFm7K4QpijJ5XyivmA6jsqrHoD7Gr
1vQDpBaCEVvMLwjJ/stBOpIiUxr3n3ahEqkhx787Wvf3PGhyp7GukP3P5qSNUFjL4AlEtObrcZuM
ozSjNSHwJbHaHYqCxNuIFybQI8hy9vUZ4PHh8TeKBRrocBlYrzGmsV2AvCGg5pxoY9HZ7oUCxTwt
KO80baGjr4lnVy2dsFE6UGnaEdrg3oKboEin8gyFxC2Wni7rq+R4ITqCUROWyN/hripXz8eNexhY
OvtiZFLuRAf74Mof9Frkgp8TAV6CBnnA7kIKJcTITJg1hSP0R3X0/LnRyDSovJHYQsMFhwzONkqA
esZSNwvcnO/pfH1L6Yvq2vE4YzygG7CaHMl7A9JT8R92/QBkWY/IpR4JYQ+z6ebAaWf6+FNS+ABU
yR+Pr/6qOCsS7yIu5GfRSLI+56AGNKtyNgLSddNjObBJ/fze6dg+zlnhoZENUavnFhVc3duMr+PU
U+vaLlDkOIHtdGpOYpbaLiAZLmvrjyyu1X5cOc0JWBObKUxhQJPNoOzm4CXmBDjgMFY6ruCPOzG3
i3+dgCZA59ZwgOpNqroUfwrS63SI3zGFLFfThcncvMQ+lS6SK4d1NlCrW0BB9SCRzafDbvY6pwdM
ZquCJ2ZmtujrA3rdR3CgH5EJ6yG5MIZ/Nl2uzK478V5HNA500QZilfN70C2V7einYL2agX8FZvcM
LUmmreNr1YgjUUWiXBfR5zZUPKi2zgg/O0hAdCYiwr17R5SkgAP9m+KuB5I0owyRpHmPnmoZPT8u
U2iGCxz88nOhBUV9nSIqC4ZpF11YBZjLbGh3MoyVRBNdeLHMh6VpUXTis1VTIRcX3iz5AOSsswA0
iNJspk5/BuhDbKIYvubQB/dYGBbqkWP+/DBykiparobRgpbv+OLR9onXXorlJ+DGr9fThfdM/Mwa
p0PG/kWUfvnEHt+GTJgm9qFQzKqhVW8BVwYYuE0NKGTHH2oQuZXjGiocBIJB84dG4dtpM23VEqJr
anvqAbYPMaf1RPf4zP+nKkiBQSL4WjPqKyxhUxWfjHh2UKjR5tq+yduBcZpYPZbPqVVLDLG57vms
bCU8Aw3T+kPeDSex/5GKRzYnPFAdXUZWJqwlXUr7tjWK756ldp60JlR7tzpPSdqrxBEh8qUcWPO4
1Q9rcgSKpPbvxPE+cM7X8Chr9Jmqdp6Mj7+zfV7h30aanXkq2wya2h63LWolzs95C4Ytbuhx10zJ
AK9VIU2XLpuV4wKd8xJtJIPtS5BPMMCF/zrumxuhPviQKu7oYtsb4tZelIqMSfe6cRiDwvZyjGmq
w1gaB3CBRb49PRcSaf68VZXxVeJMicYp1EaxQA0ddKaeBxk1vWHfxzbpXiiSpZe4FX5VLqfpCKLz
6iaQG9mzqIJQhQWzEcbJg5H5O4M+qGHKdKFcUfajRm+Dc6slyuJlYn2DanqdzswSpM33IvXbLDeb
4zkqqmSHZ/yhKMoh6BtcWvlwZSvnscJU8+7iIk3c4uQ/M+EYcpBYS5Tb1VjKSwsKkJVUTxFZxWCK
SIJ33yAozAN/MmVU6CmOVs+n3hXVNLaCuTt00vapQjvawJVrb9nuXXfmN/BOA1xl1IYK8+n9uRAs
bigzs7X1HqGfgsT7o+mOYd/P5tyxKB6pARbi33XPSn6CgU5I4WWvmo5xb88K9yHv0McG8Ybr2Xr6
zc1McR0xw0goo6cAhIQfu6gEW6q0vC2CedSnf0EMQ3VBTpaoR5goR0i880WLuRLdMPSbef+K1B8w
gSEwcGdd2SwJskRXv35KY1osDLaRFTAU/WBKuA/t1MIptR2PGLTP+uHCEcxhBMO3znyyrH5NWnL5
LflL+riSAkSQIP2S8zxGLC+LID9ZO7fh9V9xpokjcR8z/BG0GVQMs43daapmutgY86Afk+K5rlvh
TEEBapI39tmFoRderDJf8qSzIZgxGhrc6L1NvtaouS7kNj5sL4Al5IEy3wMyjBWoxXEYYqtc75Vm
FK6Bs7AY+Jo3KH17fxIyje0OWDyYgV7BNf+6hveyiqadT7m8oxwMNx2qyhEAKQ3qh1KOM4xg0QiI
a1t+MZIOiDrRLsP+c3I5OU8ln896g/rGSwlQp1qvh6yMuyqy0tKmg75WQKWFCEdwdp0u1vsNR3An
bJ+vHLHgQE0JaC2lnMFoBGOZ5rdY5OedFtlwKlUmeA3/YIReqfWM2vrdV/e/hiKhAE2bDXlEuhaW
bAqtv3I0rPWyK9EVc2aEz9m5ESg9q85cOWL0CZXAhUTAL1yUe/S1/mjKBsFV8Bp8xcLslwIehGtD
O7T+pflrqe6xlZVkfPcLP4j7gfzYb4bENrbkhvl1ZL79NQ9LFnNv/etXoyBhm8GnJxjesce08jAl
tErkcQ11OvUXEkSRVl98fqS9QHD1c6cafKnosLh4QmFDAGQLetv+7vHzvT4osVkfzQck1aiMAEsO
w+X5PSo60eq/qaKxrmiDM3ePSF/GDmhp4TKFAlB8wLNRI9tOdnNNVi8tLVodDPAAQaPOjrs/lgAR
9E0ku+03UtkNkUqeMO2yI5cuHmvTZujuH53WBSVbXfJvPhxkGyDyKm4mfqm0d9BH5v4zYDJTSlSB
jE56F79ab/kIR0xMPdDYTBFbEseCqvYphtF0owGt14ifKkeYj53wwfhO1605vGZK14h90e9mJVCc
1QuUyGHFYQr0M42oECNhx9Qg0E6M7tLDRKujB4yarOgiKjY0QzhR4PMeyPYk5YX+AzW36Rr2NW7m
C5fckQLD4CAjhi5fK6YbvGwMWZqRrmjkDrbTA9H89EMG3t/C2YEccpQDu65kK07aiXlrh/mCnBV1
ddH3sDSUBOnquSd213OWNmr/guQgHigA9XM21PWngV+U6wi7lOxCd6IwHg0LyiERuDVjJfqvgAzi
ar/kBFmt9qoPJmakAVEYlkS5S2ucrLTDrVEWsPUZ0VSkSbwZ3Q5R0ug+rqdP0TZUGtzX0EMlq5Ms
SEFGWpF1wL5ZRm+9wBSAv8QfE6XXVsOxcYBcFtR7Gumt1pxzNNpSbD80BwJJMOKmfHEZ0jdWa4kR
DWU/tU18TDL9wDVvlJR8BymdwMrV3Ny/x7CsWnS4yY6iTdz04qOiU8UuYprBkTIWZsah3V9ANVDs
N2RoDVomzJNpnjkqYcDK8npP6metqBqyWEn+6FPQW8dnB1Qi1tJIQD3i1uwhwMwkd3G8kaPPlaq8
H/LYV1CX+Wh9YN7H8vcGtPyPIUrwvEwA6UnkoQRih0wssV6ptL3UqnBpjMtAmyOIsBsTjyzTTBlc
u0XoXolMqsdnC5mHIzlnFUenA5ERhawHrPHVZmZHCewwFTLX2XUXYZibxES7iCa6TTW67QIprEoU
XaHF/iN7KbN9rDQTsbG65rkW8Ls0iRebRUhCI1Y4OJG1YFuRTCNcuwh2zbZJwJbSSzmt82cWUSMG
Hlnx6rmoYBFTYlc9hpgNEpCzPxzjFN0mxWjcYrsXB5gbga4Kw9jIZscqAs7YhA5iBySRZzlij5PH
kNTScaJAs9DKY9mmV75S4b5fTvnw0X1JeduOo9m//qVHAswNLp7PZubqY+RyOpwMvlVniWGJCrAj
vxiUY5Ly/g/On0lVFSMHY+jVkLlQaMgUvtUDzuzK3Y3QHFAFwqKHssJhhMx9cUKrT+D9pEDTLKs0
ZorvdZrQrXbiYNYV/AEYdECH24T76+QlvKutF/7RyE0bcVaPFt14sJXnEv9NvxbHtbJmqsIod0dn
PL/HMVW1peAdYf/CFFei+S0UxvvTKOnme06BayVyQuOmDUCfrmXiYm+8jYW+NSaOd5kFGYVUmw1o
OkJ000/dyCYjh15eC/6oIufV3Sk3adQdv2l+PCbB/oK1qNwf6QMljMEe9jTlcDrA/n8DBlITdwmZ
0oCEErul8B3GFmBEx/RedtUm1Jf1DeKq7GzpWvZiuGDyNECsNryxyO/N/S9HLq8mVxnV8w0S8UdJ
b2+ELJQeYr2mKhjwOuRacXqi9V1mf3NKmO6YJLhcqF1wmKs6k3aNSdUppvDykBI15PHYKlNU2Z4m
HaK7svLYA5EIEnbZHSkYiRY7I/ckYy032ReY0kzuBfIdX1jH6tFXIjMxjRcV+dCPy3BbV4HbTmN8
EUk2RrXywZaWaMUaWlUAt1SHLt5O4563CNhGomwfk0Ij1vl5WYzNH8DaIF1ksVRUZCEGNDhVcguV
aiwEukYMFBDLMn3BAR9FQIpoHAvLN9qVHwVkRRA5H1J9UXBfaWCJZsr76TYm84CUDXBYcMMItW/i
0FK7zAkzopXNrU5vU/El1JAKbs5Yb+ohBvWWRrAkcZKtDMItSAp3fWCjxI1YDsUbH5KiSx5vTK6S
AXQGH0R/p8oyr/f/zPr8PyYdT9XC80+6hl/4wSo6v9TwcJqq6J9bQa3VcNcy1tthCj4fIJjhsYuj
AzwqRNdNUlV9Y/h5FXUW45JzFVicU8A0aaBVH+6tsm9o1E5zgMAfwooW4cCWafoQwsRwuYFaAnKb
rLWSPVu3Ay3n+fSDeUe7mDR639/ugIXhmXnH5iB/H/6n/nYFmuvvEEBPSfmXUZN2/YjlEO6F5Lp1
fkVNd0MT0uptfZv0nUyd9pwHs88r3ZKBI8tScCbPyDWJVfTytH0tkb1vqSm826l++Bjkf18ziKAX
jWQXmPe62ilJfgaGu0hCxHtv0+6yoU/rLBXkgT4TDPeahsYs3KvveUAXW5PMAuVoebF6TvbDALQl
0Mc7WNnf6VxnZcqRhc3SlE2A0NRzLjcM4FfZRI3P6TorIYQOXHg+rHaBgkymkA2qKqptXyKE/6Mc
9FD9EtgJUa0nHgEdyRz1DgfrwIZoAv+DCrA7XQ/xH83PO+kbHiCZJQVeO3N5+WZMc8eQ4+nc+TFg
3AhP7b7LRVB4Stx+GH1KifH0ZS8c5O6/ee/j0jzjfMeRVPzcUbasm9SWDOkO9ry1orWK8aEDM4s6
A/Xuyu9pyYKdKqkQ6rCmnQ+rXdVNML0ubN0h6u5l3N4wAVw8vT2pj6R17BAYj37R7RwpHiuuIWWo
he8cCydVFO5jcVcC6wrrERK5Kbt85o520gCUtyh9ZtUFrpoQa1fxatMmkNR2b1SlW2AgT4FRk+Jl
P2X40OYAckeHJX245F/O5VphgeSOBAeIe8RFsAY0SfcLpJ4tywiGYjSlJtmYYzvJSGGK75I50TYD
RBtB9/5gCo4fFyodPMlXAGzSc2seCaBZ7rXhvKKYTDzSHyZL/RyhzFnmswo55UCfZxOsWMtoLWJH
yNsYCCmGuCCMX96UepZx9LNIVx0bKtMEq7Gu8mmFl85eL4Ztt1qYu5BND+BJ7YCWIttYfP8qN6wf
3hwcMD4BTNk0TewWtQzuTqJEot48/O6GCXHNCRdRnKtKc3esGG85g8njYpUoNhwqopHOysFtgj9t
Enp1vKNLIx6aMYCgIXE40yfpq//yT7so/vQMT+p0pjgf5EWxDOO57o/E9fGN6wXy5MapTGMya7C9
BCoq0bSfKZ6oGBbGOQuvLudRtmRyWbOW0l/GiUU8M1buy8iX53cWn6qqT+RUoXuuz0g8ynNCd9e1
DO72VJt0EyM4gkXaH7XwiCKEZ+Ci0TwvtPIUkXpg0le4sXwJj/NIjgssLcbdJBJgrNX9HRdKBoBo
EwHqPM/D2lE8Ff/5VDRGH+WJdmSvvoVUFZVzZAnvjugZL2YrAXVOqObo8hk5kme1YsnxLjcz0tRo
NVKyq5OI5RBZ4YY5afVCcoBNyPugT2q4CP8vMEOTDTpp8xryX7nQ8hendfrDbZM5L0BGT6MkfauQ
oyniwe9rhIr15uAc/HSIgQieZb7fQi4rm5bqgUKi9Fosgue9/42ThmYy90vN5vxNjQP2jP+rsWCz
0eMeIohaLv1hvNkVH3jeno373vAIrofSUgD8R6iRUahbI49Z8F5ARk4hKE2Ug+/Y1VQ7Y/xy1xry
myf3KTL0jvDHBScE4Hpr+3lQAysJg/IzXolf2LhN9Xy2ZzZmu0BRcN6/pynQcj2TQiWF5wpcnkxy
pw6hv9ZjqpNzkB/9iiUbg3EDXdMfoVprZ9X5O76z9PPAsU6jivp+P3XhAp6B5ZZ8so6hX29otrK4
x5ykVAhJcOlwvTCLjHT/0CXF6dbr9V0JGfvkNGH8rJ01lSFDdQnnv2J9mR21Xd0sIXyvWgamON6I
5/lgjdq4E9+PBnCZPiNnc/pP3ekfrJhNyJmDYivy09T7f9DjhTui6cX707QLmuhvC6KYU+4Rq6mp
Uj+l+f9b1hphOxyrbhLMh6QbRxm6hQSziiz8MN3RagiMx3blwYPW2jE+3QTcA30+wSjlR56QdkHo
2Zy8SG5mvp3eRQ11gPLlHObgUgYjwxDiMvPZj1LSSnjtKlsr7FZBxgO4qX2Q4Wo3SvInR/FilEgj
b3bHWS/Xp/r8qEkkypoi6F6qyDNOdlr87bAmGRANZbDDRCJwurIscZVoQCYni/YmofRiNrzboBrj
xjGU5QFbHvnC2Y5Ix0pTRchQSv3ATt6y5ZC5exk7GdSZDIKVrir+1rRgODD5MOF+tdsz46Q+K8S2
kvx9oar2bleeC6zQAq7LyZdTF2Sm5cYE32bPvVKafZRmJU8eFd/rTpbZJe/O+MVYgNMYuvnmp+B7
aTLQpyXABKxSlT8flw/LC6hIvGDnYrio/AcQJgBNw3MGtyXqwqWqSsnCRMS6TWVZET5vFmHXMhZt
7ySdm6sYpYFKPayrDlDuK8oWwu/ylKapvD8nSKlX96oVvfu9eiLr2ic2ZM6K4O0gLquQT/l6XSme
wGz7KezdXMiRSjATmp88giopJ0aqGhh0KmbKzeGLai4wHPOrELzEsUlyF99WIpKbyBrvmZauOcxh
NWXsVcnlDkxJQGa9P4Ux1iPR5SJ7e9s1uGIORp3sOdrONXCXl3EwcECbouAS7y/Lo1x472OUHV3Z
D+sA4LfYCqcxaX57ihZ1ZBP/GdOH+OIa2eRCNULgjZxkDe9J3Bdv8khUc+GMoPBwfe/EGizrIQur
Ub1Tj5X4MQbSuqcQGN2fTGOxOc2ONuZPVfakXAPDRsKVVDm9+mGD2f091buyL3e5F+kRzJ6Nt/sS
Lw5xH5QVRXvI1fayjg8EWzAx3FSCGZIBW9ZnYfCac5H0+8snYCpU0H2gmjxvP7vBoUK1xK1dXvnj
qQSrk48ytBP+oR6qHcSyRhn+pPruuzlBk7KtXiiJHKSV2SEKzcc7nhCpibS0hERwjmAvOJvMDDpG
U01lioe45/r03xCrmCaoqjaUqsf20yH0Ir61L7JNjBp/4z8du5Y6CCvQxFz+JkpdUbjw8gf7uRGJ
3U0TJXThu3c6a2nmbIaFpBu6DzHcZ55smNghYJdmjjOxgoAWp/3GbvsNYsNK4QXPgi6MiA2lgfkl
tIq9CuBL1FzTRKGG9xRjKwrARPBC4Xer+y4znkZ4pYZl2QnrKAyeGrtHTEsMm3TkWs7yxnfrM1dB
0izCDu2Euyz74Go9AGGj91qIwV3SXd2J9ZPstBH+ROc+3XFQXR06/AZgTXJPxgTqqIukwsBfdn1l
zP6w84D49KLbswis5Gm3XDcbo3fSPBolgWuuMv4/uX61bfTIxx9ZETyL8pS3PrXs46UiZIU1Z63Y
JdM5t+BBw21j4lOvOlDbFLFBtQre/CMDQBScnNFTXXgkN1jSYg0OZvLq2EYihNNoFdDNLEy9vNd3
4jv00ZO3qq7nem/PZNagz7nrN3vN9EP8Vh4GjimjNiJliqX48I7v5QuTre2qiDlY28AiqScD6kz3
FbeJuQ91oOb7f/VPM6D/ZVEPQ7Fh1e87Ltrfp/wkamZBdZzH2kRrdqSx73iqjqa210JPROP2/nGi
ezTS+e9vS9MyoOdtHiyx1dLtfguMAgLU8errk0c1SByh+Ctrt7AKQNc0fh6PkvYldT9yCujShJHs
QMUtwFmGEaz7snpi/3VYhvB6TtW4VpRLsAQReUulM9OToymDkL0cjMEtJcc67cXxybhRsD99ptR0
iAuQIhu9fTGOHYfCdDwxS5teDSTIFL/iv2P6eltmiyEb6r0Lfg3eJRq1ubdhD8a+f6bKAwMAIxrh
JOSlH3UkFfz+qkdwrmOk3RJhFpoktl0s2MyW+KS6gzzbg9SqdxA2owIV7DsrqFTippmVR5ozdSU7
A2B6xVnk3ML+GKh1mTpNHcqXyBIc1pTTi+Bm17ikSuabrSOVT2lTr89RCkGTwoLSTJrHiWGYihpA
Kl6p/eP14eNRnpe+vv4uLF9FOBD100ErkbSeuOHHWODShFRrTB6pKtg3usRKb8o3Pqwhprtf0Aow
gSJHAWSFzO9iwU0ej6XwvWypDNbhKf66EuK8R3bj49LCPRObqGcavE8xPqs9DC+lcn90Upu3kLkh
yL1qulmtLcu+apzvI+QVseQ1RRMy53Y5a84ixFXJUIjnsX4pLGX0VWLvVhlnwcWtuLnngeQAIyZX
D3KaCUwSBNzkzho5buHLd6S/kRvf2jqhaQjffR9LreAIih3b+FTz8zUhrBOTXR6O6UTUt2Tzdq6h
4D57DR/pcXg2cccmrx6FktHUj37tUeuikvyZj0fFNzG8fYyI+TL+O0kWhXJMFWdb1GzPDlftLQoo
C1FxkwG6uMEhITkrjHMusqky/NEvbemwiqDFJPYfeK7GjDD6Dq9My8P2Ladkymo1J/i4xkVFuDOy
/H8lSsOAijj3thMMnncWV9l2Pix/RxCCIjKhOPJgeU0/Dv9h13wCoA+nfchNxrAXjvdmJfkKRNDs
i9CbgDxzYZipITpJUQpNJ7ZeLQVqwPvsfOxaWTTwDdYQXPdRbD5RLRqngqhh5Qc2RdeJC1EMapi8
S0WFESg14jH2hWcGYUsuaI8WL2fdMURMM31IRia2OJz561WWXq1EVKRKIbVAfdlTG3OxTHrorBLn
GJewImwm9kOtKNNUE8RB/QYojZnb/lOOmkkjKsf5Qh31lEwaVm3l41XcypqZJMm4c315/7tnOAF6
5LHi443s8sBG2Zt5Un3HB7O0HV04maZ4U928FkBGLQYDyIgF7N1hQABe6TdauC/m5kHMnQaFDCz9
VDPHkHEVH9nL7sVwfc8EeUGO1+yS5f9yKP9wThNr9qHKDKeGsvAG8krL+Dn95Ur3VatlQ/8Swtur
K4tV+sXh5sSNLvTXCv3wSm7OwBzsMM/3EyVGTjfNP3hTCpFMKTHqlMBsXmdU/X/ptw/8HqUwbqdJ
RBdC99vcUZOZud2ydVJCBllaD4+UB/hML3TECJVU4ANxW3jfnosNyh/0pGH4L8vcdiROie69nEYN
8jk3JsbnEdwzx/mCh93ChyWe3mLTrz/VFvUzCPjKE5tZUBcmnZ0y7pI2s1b+vdVJQhBM5WJ2AqFY
e6zQB/03IbCQCN59rx4hBnhpvDqHRvyrS/os2KmY0d0PwqFL+N5orW9sg0rATmfpCztU7XcJh6a7
nlcffNZa8FdTaWlRRh5E312Ff5NJT28Ycf3WSD26MAlR6EDS+jtkFwU3aKQMPYlSijxIMyCKnbBK
jvlKfM2OvISNfR1+cT9joyFrwQiWfjjqn04PqkKLqYoM2auFXqHtm3DOvomTfIwNDd0lFXtX5czG
uFlWYv7mHUgB9kljcRmwiAahvdF8qQX8swCBHcD2/D4Kwbq6PMm4w+YRA2sqi9Y/K6d1H5MiJUny
QxqCs59VsRUp96MKu2qio7jCxbv/6gLebtW+It+ZtnfYMjOwzI9eW0YgZv5fjx/mvWqyyr00VyBV
RKgbv4gVpV54g9bgvihBcsS8RAumPiBekcz2lth9TSNkDCevRaUnVKYPxA0E1EX7GbLGfTL8DgFj
SJiXpQtrIrNQGbkdo3vz3jGRG49iZfSYc0PMWC15fpgUdbnn4NcAJNldD1XxtEson8TqbgZzh4RU
dMJrCBwgKyOVgANENZl7l3GnxbqhQlkPBSwl4y+s5oiw9VfpNSkrdFHNmtL2TXE2UE4GGQIZy5a5
nhUJ08OyPNnnYNQlfF9dwAWkHIOFPty7t54LFFQhdEjWpOFouCg9sfo4RIwOHguQ8H9BSSxi7eN+
cz5K2GIaOzB7fy4KhA5Cxw39soPzyxOlyTEVQSZYSFFYQk0bplnlWHqdrhmTaO5GJfhWLjTbYwnE
xV71o/X4PI/p3VJHFOnk8WfAf9fDyFgL4a6v1C0OMTUui2mYSqEu93mCnz1Eobm+uacmvtsHmcm9
7zj/pRjAVG22dwiJIAKOhYzdCeSUpbdzKpnvwKsVwUwp/lqv15yZC5CLb5xlFljCQvGAiJ3ToemJ
mHH/8EqTqJhGhpeBJQ4Y5Nf1Y4IoZXAfHqjGZeynMFNnmUHLCowK1KGsn7gdnKBO5BsY2gsNMR8M
rZJlgVp+KO3GIMgkvSdFWqc+mKuRe4HM9cg7fbtORHMilDgcF2Ii9cgLhg8ybbStCV5iGOF0PfsA
rgg0cZZY9JQUyct+8dHejfu/rFo7vm5j6nvZp52q8XkZZV+WemWjsKqwaqd/vWBK98kxo1RBcykX
LO9DiQR1YnyswE78tL5RUX7/RlDGbk9bypNTSSe8kIvo3EsUlV4sjesrCy4V2HoxGS+12nWLJycO
RvC1wyl1lIn98uhH/oyE6SPi7snrZ9vyRT76QOUucolBjeHIG0DuJ7Stb3JBakDg/RzEKY5Lqrzz
Xn5uWKrL6CEoYqC5a4pgKg4eDz4OVgaVoNYa+8JboD6MaVjrkEsGBe/ur0b/FTwnTatnWFT7zKeT
9eSHcB1QnizlBhd4TbXuz5q+ZF5d0NRu8TO/D9BItNO9dJD60ZaSGL7KaUrKz1zfMbEx6/dMb6Dk
mDPDuFhVOE3DVTGR6CAlQTgxFRxAaRyVRzMuGEsOmfDlbahR77hWnvdt75Ho/UyHyCKUMgC+NeKy
aa7iG/XUAn+IDPQ4coZ8SOq6S8wzcOU5MER/jNxlI6jhvJ6soENsIdf56j/TLhKH/1xu/L8DODm8
/FKmi1R2zzv5RPA+khJYMZjlhnrXaSiqqzoAwpfgni1G3Iy8G9u02KyTYA4xmasqbI0NQ2c42rue
PasPgRR2jRU4tcroabrMpJquYJ03uqhgRZ03pwU5pCLyK+oIrFC3YvXsn4EGi5wItzTITtOPUEA0
eHHcpNScvwjT6unyR9nyVGiklsQkJRRwU7NdSKrs39zAVvdcNhvbU8e7sH0LAjsEJIm/OjkeKZfS
rOrc1PXlFI6nzd5FqohH1k9WsbYO3mxkyKiKvLpohAEr1urpmkb/YaiebQIwTC/DdRPyEFPNHilF
U1x1iigqScDKB/pmYTaJbo4OBZ7Sv3iEgm4GOAdY4QBZXaf1lRI7w+8qWOcMuaLGstAl16F/pwE/
GCvFVrNtVh6qhxWK96D6Pgv2Do0pD4Kpp48ulLuiMWkKrvUH18SeJ2PO+9TjeCGnlPQwnZPb2e0s
u8c+13rZlGnMQ7S4VojfHAZvMiSEN9M6HdZx1/kDBy2djNieK1IKPm5SX1rqsFOIotjXvUXEWak0
iX8KRaz3J2F4ZUwacPDl7kmVselW52MpWsCxPRTks1iho/i6sx6OoJpEF6l+mVmQE8cMw0qZXBFB
zXyZ9cPoyL7oAOBCXGymtv2nG7lf/Ww35qmqBhg7Kjs7zbvuJpKuprr4eehY8Y6B+MwBHbJtKs3a
7019IybW90/f9z0w5VccVxssY8OiYVMe+JhlSJA0ZY3uBgMFh0v0IkhJapjeA53a6p3PX8YPzmih
0z0D+wbbcmPIPTGIXOqTFXcGvtw9qyLGXqd+FEa+7k93YoL6TobrrJP2iv4dn4KFMYWL8He0cEbu
hXhUj+UBWhjCHYs/4lddhs+PJHobzXhH946g3Uf3jF8/CXSr2+VlQ3txB+9zj0jrDzygbSpZxwJL
/hHdg28Uy6t8f3zjZd2L2y8ez2GW+i5Ib95tDfFsxTO+cdLlWz/0aQKZzs9qWl2bgH37ZOxs3Kvn
4DzdvggdtaSedjMQ1+TDU+0QplNcXzByB4nrTotFaGPA8y60AZduu21ZuZKPzLlOn0yQ6ddZCP3w
Nl2nt/Q35YyVUbQvLW3cQEGag5Ntzc+yeweTyJxsd7ApsRnH+jDZuimwVT5nU2LtMd0FWfls/ddM
Rp7PQSCAwKUg6QA9bHj+PHkRZi+9grE8IP2X1OqIS05jWOzbS41qbzLaAMIpZLGktiW4S3Bkxdj2
F0E0y+zEOkzxtggyK/Qjdxb971+8eUP+GSrtTJXHjWIE5K7i09YT26VNal0aG5mbW84KfUV/BupJ
y0+4fpAP5qWhEUGX9nULQtCS8tILLGin4Fef+ZhZeq1J2TpJLPFkkdM5liHXu31qaj8xJe05u/Np
Z9lkrnPYOs/ofiyLc7Gx3yF9uackrphSiY2fNb06S/wgAQbIuzyUABIaPBmdUyC7zHlzzZjHuVGh
JqmA21rXxLPYqtJFIUbfUbFOOGv2kW1MfvEjZL4GyCkmvMAskYOiYk594jdH2JQfQWRmEOB3Ad9l
Z0U1BVPqQIcKA+RDyo8ujZava4P9svIG5VTFU/hRtg51nONJ05KlXg7Ce/bNXC0wfOitKD77YzAi
J1DDJI+0b/lgnmUkYgylhypZGqU3/g7zTlmLAk+j/gsHkO1GiOiXtEWtEV0JdBJO1e4dG5eSr6Aq
vj9ooXGSzKGPeRCK93nWHgms/dwd7X9t8aHQ1vXWdknbgvmpQ5ykvPxkFEhEXa8OoaA0d4z4Nm1+
8WZa6+ohC6/XaOVLy6hCQykjTF0TUK1zIaWeiWKYaZ+hIjYzMlDQLccD1MmnLTgz3IhAeHpoTM41
XjiVqa9i77mz9l0BR/jNCg9r3rRTozcgWynwy6gld/C929sDV4rmABuC3OylwWuctTSsHE/N01kh
nkDz2IFS7Q9pfiA1AwUXQozz/ZttoyfFWf5pLGEeaiaVHTzmznYn0bioxmqTeU1C6MDyhQrT7qL5
YxzrfGkn1Eskn1B9993MjT2JvWvxybQ9NBqOC1t2uP/I1rBWh2Zv0hk+QWeeOC644IbNy2N4NsZa
SHlWtUqwushHIGm8cUL6jkiSQz96uGPHg6SJVa77SZwrwT0PGUurf5VMp+XcQZRO5kUJlMFmDvmB
x+HrewQKFPpow9WvMbN6V2Z/y5/3c/GTf5ephmgi7OfoHxUlemNAh3aMYL/dTn3XHuxMltkAO+eq
K9BkAv24sT6czc7sCO6+Zn62W+QYhXAkKQpu0gFtvkIeBbHQHo3ORYBdJ6B5yz9T4lmV6iAt91lP
cWOGecJKdFUiwMCuzQbYJzocWrrZrTDbvXvFWEBFBM/t6TW40ED5c0s82E2aBef8EuqTwBWeR29n
MeHj6cT1nf8sz48xyTDcocgDiNKZPMF6pMngEd1clbxnQh+zu7jpPMdRGuthA/OnFSyOg+A5yRYR
A0+sBJ1vcUwM6x7cDMxRYJsG8k8dNP9LYcV50nNg4Ln4w/vTPGuvnQzsgASPhjTLBbNqLCUsRF2E
N/Ac+XjxGcineAtRwxTlLVCmEzRBR7uK8rBsXTKFrBpDGp2ft0sMs4l8w5LjN7l50oWKnnqsvPBX
0XwqFykfbfhFCKpP5bkZIqkiHNVfQNCk+DgymupEK2w7y/FUcbgfnMup0gefOvThwdqwDa4r4zo8
FE+h6lAPCOWo/m1qHkmzPtl3MCP5JhoZT9AGz7TEpaV1Zu6OX+y0J9EAYfHrWZMhOIgWZXKInvHV
ODz/Nc3vRIRXlN5hVvF1bKUf4Uwiuyg+4ALDrQPM3aDZ5KwIxR4k9xSARkZEJi2CxW97X0MuMYb2
QLMyzUI2IRjar6KapCIrLoSV9IYCM6huFxwboijgco1V1S5nsUgwkZoEbvYeUUVGF2ZWxuexjP+4
ttmXZsgOhEsb/HRR3aypKC+HzoXUs6JLZvQIOmLwTA3cr7FsenrArF+SFBPC91aWSAxeTrPM1T6K
H/h8aXXc6XAJqDrRxJad/xIn8w4451UcecZyPxepYXlfGShwiM5e/20NBFUcAYoKM5jDPL+U8MY2
dVa5IcEm2k9F9UN5CwADdymvlhPOvydDPMKOgLhM/K2izruvcirPkwpCncIM0d3S+dM+CVKfApN1
gWPpHtEv0WmyUv6XaIFudxtEfWo4Ge8p9v0SuBKRk+gOBJ7QfkGUNvZs0KmgCjpuMp4OL9Il2OEB
4la1gGTl7D9mkxNa9FESfI1QjdPwvK73TBGv5JQB95E5j8aHfsToEJ9BVCKR7PWwLbM6fkQS/Eyx
GjHwy5L7qqPNCUh++fNd/Xub7ViQbnWOEzLl7LuWbnfXXUKJVaLrrU16m8JMaT5LGIsp2jwt2qsi
nq7VpIlAGwGv5lICo7XsNCkfxOztaZdw9mTlD/YYHnBzm5uGfwiKlOcd7bAndEH/iWRGA8Y8ljzN
YVJWo5+p0hXRp7F7qeJ3iXzl02Y1y9xOAmSCgbdh0dq1C+s15+C009YFewOssP38+DtnXH8UG5hG
wyAZsTQb5GxcK8Gb5SKBhUA4PAmTlR36RkcK4YwhLXZMf0oPvmj9VYbeIt59/IKHffvF8rUP2cAZ
eva1sEAs2nepTfiHkoHk6dldMJy+y6G48PwqMFEnJPHb+zZm+bIbcGEUDwcRgaN0U0z3UL6rrL7A
Xd/Cv70HLdLwHsvzeroqxnB+TUU8TDn9Dm6/KtS5Hx4BDM4GYEvROgIILDci3CD9IvkERAjSJ2dA
TEdtA2YE5SolhHQeM3LKY6oEFRMwsNFq/ZH7LAd+WgwQnHOIR09tnGcUqFfvMRzikd+YMnp8mpKe
kioP3XK1N488PnbLIyF/qFzAGgYFqza/h+ekRdp2ZoxtFieanlpLu5rHZ0wfZP8+AYipQKqPUrkk
UNpoKil6pC/L5D/B5qcCz0gCKvjCb9CkWZb5i2R+f5QbcNNmPwewqXNOSuJkDbVtsnvKKEi1TfdP
bReYGK8Ft4eQL4mc2ptX9rUDLXNCQ4ADTuKXP7Eu92Dp9a1ACL09gYUzTYwx4bzTUecDitbfN4Fh
vR0nnbF2J7+pjKMAwzS/T/XXgfM1ozHibbGkU0ShxGXmJrRttPERIUZyn9qXzQMEqtcGqxuLvZSR
4loJoX/RvAa9sb4yysNFHYav5PO9AXYfakV33fmNaLx/SH7wUxDrYbAyP83YHNOumo2jW3mwB1N6
B0I4hSwzXLhSCUudg60zqKQjNnHifl/bTb8asDFT7LWIvzxloXFShLXYPhlxsGt597tpgbjeqAfK
oP7FrSGVS60NLoJFwJ42nlOno3InbHbaR9mOfqAsSEvEcWc31uu4fAApr6V5SglWZy62Jl0BDdqh
7OhKXHqso7rN93ECdIS/mLWmyajr9+N08jNtwYtek+7pnMqPC0gka8NXX6CAV1Bu72/WaV2PCjcX
AChCaWVELPidPEfhagTgw8JA16smcqROKiu7wpjFBX+FKOW5/MEVawTn6k9hFljvowTYsc0IOFRq
4YAmPl+CxueR+qeHb1yLu4GWRsTM018+EZUWys1Olen2EA5B5wIrtZGlLnepq8aEUg/8U6HGOT2D
QhW8Y7xPJJJFhstBpcdiL5g0vErSGwvgFoDCg0Z3XiLHM1aLr46XhJDmh7hja300aq7SVGy6VJki
5SsygsuhXNlputBuoSUTQ2vO0XrSORHbntGBy5MpmXDpT8k026GcgcI4QBat8oQtaa8QjFGiGIJf
UeKengfSzvKc2IzjA8RNCIdIGW0xEQ9MGy3aTmICXlDtDouSaxJxs9ovbDyExksRIS9eMVZ7OMo/
leCkmU3nJnI0Ha7znTsJTkelIX7WWszz9Pe15oq8NoDLV1uKSZJoFEZPikhsu2FBNYQRea+BK3H6
9xmkgU09Dq48wZfTVuG8CsWK1ZScosG3KC9KXicsYkuRG7QenvY16cI3RaqJCFPxaZmFCQMwjRnj
a/U3rHarLveyi3NvUwg7oOwrPlo6EX+3h8WxBmAbm9YYKwj+b3P0R258SjrIDCfIFI+9LEzmHerF
7jAmaLPzbEpiCLYazIvTU9eZVsgLBuHpPNE3TwHqMh+Hm/Vvn/0nUStoMq1RV4yV7c2thwPsN6N6
qedJAOkGhYMSiJsdpSrtz/sDIyHUhJoKV/bdlLtsTMGZdidNFz+p79ihvXDoDV5nQ3bYetJa+23g
m9xgg9xjpqs5O/Rly8Kf5fTrcTVKv4vF/YZkjddZx1z03B/7JDTeRrC/WaAOu9+B6j/EDEwcW1dl
WlnuGybLUmnhSU31lvt2QKAHeSYsa9NHtsvs9G27mBcOOGEVefQGygj26Ta7jnKXMKiIu56EHbcN
HwsWZz1njprzk8RvC2/HtEqNP6y3qZznjBv52GqescqcUgHIJ/GHiXlBhH7nUmV7rvZmv9414GXR
UqhBhLMaRhWzzxxLY0W0RTmIFNnATu6MD1oye3DRBzaT4T9pQ2hILCCZFpvBd3nx99TpWtQVkCiZ
PYwplsOj20CYqzg15h5ghXSpmmFMV8Y8lxa7PtpW/X2+YPDqL5TPC4/8h2BLC54XSC4E66i/yzgt
PMbwbOuwRuTBhjrPuuch0s9uWkICSnAdNZeJZQvQN0Zv+MEo98CvCGvxyK1ACeJYXPRbTDqUx/du
ZUhkBn1eGLTMmId7bWpnZhE3wHc3hJx7d/gNXxFeYNxG30bWpYI1NcyZqHoFhegyVm/vMQwSultN
fPerGr5RBCr4T6yDQu4RfTsehgbzdoMKKn0QZ/8uT7FX/dKevpm6OsyJeTOsQJ0jW4tvQ6w4iJQZ
54pZUeMIJbp9W706OW95r6nqkUq4gUxavuICQ9DDGC51LqVjV/9MY9mrrJzV6eBXVEvBHGSaB1Na
8minmBo200s0+dVigxyatjZbZQZipLU55pLJPp27mvTzCgBi4sjhvaUwQ2t45MCjMzuSUhjtm1/6
lN1xzcGktLggMSuIoSll/tXijISG21iu0ZWxl33Dt4Kn4G6LH1yatS6M0kgg8hX8lIZZG6YHNP2d
OR4h6w1tnuCHaVCWdqx0lkzBZJs+NfJfpdLSBbuOPIFtS28TmTfVNNN7BKSE40w9iPJmNyqcj/di
sV/kmanzuIclos6tAy82Ue1S6jzDtRsIIDw7ydoWz8p2odoIMOwxg0PxXe3J779SLQX1lBhsrC/t
qZ1gR8Awc1f1oIK63Dps0nsHT53ZlAk55Ix633do70WkRkBJYg1oskUh0H4Ia4S4tfY2Xx2q5Ele
xKb/N9FatLw4VKbO0lsyGAx+UJUTAOQIsx3NS6VulKuQuTgK6xj6/off5oATNDcCZma6qOZfXP7C
3jINJA/vrzw9ozQyp2VTRFno2E8QB/vJPUBqupso2f8UH3xSx7Qdug4bXkIzWhF3zkBwpWsmSd/Z
ITiWAWrFuUcmCd2c34gkd/w9fFq0Ghtw27wVFecbNVQmyDyiNGqxbN61cvb3ZwnBUqm3FOovuF18
VzDAEMEMhI5zcwvcSVwDI9kgZrJd1Mdpc7AEbWX+HXglmPZkSdTcUrhDJvpe9feZi7IECgk/OyFa
AiS5RbZLcoHDDzZoXyWWcGh171nsaPHtVO4f4h281x2f0lB9vtDEWuk/kCrswjGHHMNpXzp3zCHP
/Rj/AIvRS8d21klzSWPKDJiBOUi06X2AvRhbn7+xr6OoiXNZn55T1ieGW15e/zwpnAugEU1Foq89
UyFpfchu/dXlDsNqGhC19RTfqhj+cfoqYcS3m8nZJRo42OfJ4Ifj5V8JwtYmM9d8JV1PScO6e1T7
UOcPEWwT7QJuQUPmhtmbQ0xPVzkxTnreWZFZzdtkT5GEC3TdlPoSl2dn7PPJkBICc+R4j3PsyjBd
iu37g1jCnCByklwc3WjTWeR2anwmBiBz1PGoP70MdStcHsuQMPM4fp+Ap5kQcfkpItuoLhz1J4tl
v7ho+BnAjM/XoDAOFmXvlG2CbTbX7BQg0daGWlgPuVOO7l+5LhHd75LzortyWvsei++Huc4DXgiC
vF4gXv7YZgZASkMmiX5oqf65OgFJEHT1BRoWc42cZdNSy2d+h6whYTmBi1Ywj3Ng7nZ8JgNq3enJ
WbvS+zMkFDkfcN+HNyRqXqujoJWkHgTE2GyjgOT/GPpQHNYkzi/dVhkvl49CbMYxXFN2JC/rjxCG
tgM0jLjx0Xr0PQ9jl7h7bpt+8sdlBKx4YoiZ8EB5QEmAPIWMznHaZCo3xuHsW6fvMiW5jFvu8WhX
PR+7Kt2u2o+EqE8pujbOUgQc22AyNT3yNbFtpMJ481QePFxD/yxVlzLKHZqg1fPHW3pZ3uPpDQIG
9Fvu6axVwdWQ74Vo0Mhv0QYg/Sre70z6kAWzciCVJ2jv9sQFgDxpyhTDpcZ0mLHg2bwMJQGM6+H0
AGRBjX802chbMWu6/GCAv9qDJXMRzLDx3hp6a4BzNjcclIiWBtyjErmzMhvBRTpAt1vDgALw7PdT
M22edi/jLzHJu7v7x83HOhxAhjHStgOn6XXxlmbmdbhV4KP1eIgCybg4VJLJDuXgncPxBiqHx9Q7
hGQLWDFK5BRQVIHl+agqVgHhX3Hu+YAiOSbF5TNTuAuqkDeDf0uLcQdAZlNSiVEIn6bdXha1wr/6
urUa5N8FvSnCyE63qtjLImAFLg3WfLg8ZAK3alfbjDldDC2r2eGpOFJmQ+t0w9QZRseV73JxqWIP
ML/FGT1CVOpwi3UTIolrospIAlnPDw2UpNSrFixYE9OUzxE5kGqXBnfLwmeNEAmQ4u3QsW4hd/0h
zXf5OGv5NFsjhyCOimsPXPvBcor6afcyb3zMWAO9AmiHJvySIojIzbzRWEhhwYxJ/4Ic1T4ssJiq
kyl55D+kpNlbEm4cfnRtKXgR7CcmuQcjE4Xmb0ErpThnvoG6V7qJrXxAe1hzRP8qHcOxHLxgyNld
OPatptP3UaDSZLRO5FAGrx/m/47kbQCgBYDqiYF9uy61kUdzVCI8xnu0pO78KkI3ZZgJbHKh8DHO
wr5ur/aECAi847Nm7Q44Lfcl7PSijNJ021g0GhMkE/jSb87QQmTmWmG8w93iysxLTCdVeK0e1qKN
AOEhNSJazf+y2f5Cuef5FcXWXgAC0vI4xM4MQAXGgCWVF8sdNRNf6hi9gyVTgutlKUJ2gIN/KL2X
RSaJgeWG81nHwX/wyoNbK2PSFRkwVgG9TwK5kKcgsdG4kyHMJp7JQxfYmZ8gctnfTQb9BxiNrmBI
aLYszJSZNW4ojtXjcrUCLvrCzoids4nuT883CL5ccWu7Hl4jSG8ci2rREc+ILHrtJ8gCykMXCkPD
DuiZBwKbtdjd7X8gikKbkzYIZs5Fq8B8wH8xwFAguPO+QMN83FChaljnh9dseTz3+ADoCrGr0bQJ
BaxuzkUipPbO+jTvXE+xufQ6fDLx+vyz9AE/qgHq8aDHB2aE22fDl8hlwwYt9nz30SCZ+hUC+9V5
8MG/u6gI3gyOShPdSc3WZpSkGdRPEybSLrsLf87qLmUi0XsRCPxzvLR134AkJ7rThOA+8Rj+AxAw
joFxdWAPN1P/LVdRMj3Ja6tuxaTDbTFSR4NED8hTwQGTKQIzKGmKcoJIJEu09Kh4RuBb6Ca4mqMT
4/znciSyDyEZLCqyQUHUMV08vSl1Eppln/viNT+SxUWnQtg+2BwyLDREU8CqvLiQVuG3Z0cinLpF
Qj49hIkZpDzJ2/zDIAshIGyOXswe1lGD7TNw+/5Gd2w9qG2PJm9ZGf6mJpfZjnde1M6N+m2KggM4
lsEQKrYu81WDKrFFDDPVxKL/oSm9qEV4LGJEYwgu1l6orC7nW/uAbCiYbG/fACDvBmqdTRsAYaTc
qk71aiub4qzgzCsXJXiRzoilN3mvqioAHM02FOl+/0+ADQNcFCQj+6fRQnCShj/d18kd6dhSvFNw
npA5hXwW3yECENaXi14YMRLbJPZVrDlD9pk7gwY3Faxyv6rTIY+mwWmtLrM9/9/QSxsF/z8wRznv
WFHn3/W2S/1Vc/GLHq9fyqw8k5edrBA06kbEgwJZt4jRbiKwRyDm3WaOaLiML+ueuI/v7P2t7TwM
l8hsoo+nU0zKUx28lLdPfgNEi2Vq3mum2DJaMXfwqnudVduCpIRTywxkNJIwBFdDSj/6tacqw+0F
KYJQtt/qQC6WEZuFV9UXlaPGoLszgrCTouHU9ETuPcFuVUAS4kXO7PMWnHSocyLPMRcf3wjBdlYk
d2SjdeyFn0yyMfwoL2KAk/0T9SuN1qVFLbZRHlZYYCwSQxNNtdBGubAgVTic31v3y6rhjid5qET0
LcSHZgm7K/q7ZVcb6GPetiIr7jLtMm5gxfkf8BK6I5DvNer8KTSClVXHCxk9faHNrkhwPAYMcQSU
kRRYuLAqTY+oKhXTs5S6gHHp7oKQhdJMqGcYLx02LzNgj7Go0S7yI5iCJFeogUjePpjkDi35YVoL
K1QIAu8EMIOL//4bmdewGUs1xZwKJtOw5EKCgC/v8xty5hHh4JjwwEuGBKz/J2hOCyicDfKDZJO+
H9unAfFVf6WlGgpTbzOpxXf7ZIsb6NTjmCcm2fqLioYP2ab8/LnwDrzfs/ki/kFMp4808y4Oi4Yl
zJafgjFWT0fIhS3UeEdGsq11T2vP0RHTJQvedFjnqeCnBbUj98kSDNfndjBhIwitRJWfGDykKr5E
ew+HFpWQ3FzkVJAvxKycAXtQZCnMS1159EwjLRCKK6DLg/07milCXWRLwnuUWbPv7j+bNqMmdFEA
1Ut++SsRs5955cwMZrC5/jIDDjgsN5ajp88QteSjjwTbsz3N7EY5b+9P1NT/oxj/8SFAqraWotjl
YAE8p3p+g3R1pEZjbrfdzaWKZ+N6PWfXDUfiu4TXQe4hjkuBmRM9vx03hDV27PyIIMCOf/roU5Oy
s9USHTI6EbQh0DG2YiCG0hXyDBuqZuWrSR6Y9UcgadlnEE+LsP1MPxOQwPaTfg1GQAOAe9vmPJBI
93amghTJepzrd6RP5foVuLG42jeLJcCMi7E2oYfR5BZtaUPbTL1tWtYsR0bR9+4CjBiB9crig36d
1Vrvw9gemt2NKjBFniyMRTE0J4UPn4jg72hwLgL+Vx6a4jGWFfNOWGmLy+R39+iRv1me2leU4URh
TTpF6qS5TgPib/XA/bc3evhuY2MH7Dq6jLb1qIOZ487yddGPWIuf+Z237bJBv3W2TI175wugnF3S
gTNMqFF8Xdi/f/2OnGvQ8IFM+Ha/WwQQevpqJdDS8BaYP/SLnGlVonT/CDDnsAI9KaT5UMsZn811
UiLHF4nkAFk3lSU62gI+zIREWVCL7s3FXWtyi6rHuIqi9ucpGFJ7pnr3HGztBppe3hAw4Q38Fix9
SdVeRB6pdiFx0WJp8HYDKCdsqGvIO/2sCsr0S2yHLQIG0SYFQC4zCKoznFz+tas56ICDfrgvufC9
fqLXIe+SJJTo4I1AzQKab0KJWsU6ARyM0yNHOmn5c6hueqLJJWn6t0yku7ebDp9dihRtOpL6o8bk
PDk1aLnxNGp5hCiviV9IM71IRewIj+DNA81bhQTq/nk2qh1yj7pCUBxkggGU1K1AuDGivpYAKTlx
XNiuXh+LAc2I46oGLnDF+xKMNepOMDWJ/ww4+n3MnA6XMQsEHB2uHneZ0Rv939UYHRVWU5WcHftb
sDzH0ou7Sj9WWX9IzGztWEgXd1mmYSu52Vfsptz8oEWoSECqPHyXYIRUPc7oMbUmgQ9qZcHMkC6L
0oxXAuXP9UOJKoM3aHvKJlE8s9e8Av5z8GP6P3YLqWeTo4aaAcVGYjz8ZVPVfSgT/hHMwrSiwV62
VYV4coyR/5RUNHgkwqSFdH5JMSdNcjIKEVYOt8Esd5OOYie2a8oHSVwffPqiqtSOBQNSCrXEN9FX
SFZ0XbGxeZMGqxcdK9+we9YaTdiUFgh02r/Cu8qXdkobY5V4CVlhZFeAhbwYGTroPMLvNBqE+KgY
mYbPl3p1QEaMOpOryc/XrMmS8cNFJ2gcSplDd+1qriyX8dRwZwzhVYPw4ra3Ba+poW0SOhSpbE1E
WupIIKB51H1fBj51K4K0FdUVexlVoyS16vlbD29Ccsc1WqAT04ePlKmtWSakW20oZ8nK1lv3cwJe
QQ69il4BcI9xjrnhDbllWw1N7190LNVXpzhqdmpYZbzfiJq3ijfRMouX8cix4JxIJk13rsA+Q2QO
u6JSIyBvrekvMWQ8J2sb4y0pIQi32x8kF7ukC6xMUm/Fot+5hgTUmgbwoWVeaSWu69PvITAyok52
inllgufUy6X3g7ZC88/V9DFz8MSS+ADR2mvy6Rv0wqOhCtiYKIf4TCqQF1d4Yxo11EoAdiVt4/v3
8a4kcMH8y4TmvCIX7aRDagu+wDe+rLtsbuZTqk8cO+LhcD2YpazeArWik3t6xsuGA2dIazgNQGBu
7VgVpROPMm3oRO+pkLm44VuYzuJDOF4GDm5SPhrkKTHTGMzLANhZiAGfc7uov0u/Yq8mUYaVYByu
y8WN+8f7WX8zc1ExQY4qje8bGwKXoUdQHuj1Bm+pcv6T7qvV+gygpQuVDOu29PpcwL78lV4AKJvC
3TPnUIGpuei+U7ztZXTF3cbQDnyRB3WYjNcu8DbSwyLvX+nq4T6NGLTaCwAl6JTqGmrRtUC7CWjc
/4XTQr+VLeX8nF7zB3bYRMYLbYylvnekve2Al3LTWA0PlXewMclluYp87RiEYDwZYaX5hMjDArcF
gN6DWdAqhsYLi19Mub2wWtInW719uyC8AwntQA9+VH9kb88brU25vSd+5f7ARjxmhDPifMLK8yTU
jHHtZxdyNowcksF22Ul15IsMtIGgG+F2Z+WUif7Gb4tY7IpR0wNA6LEidmT7qkumCxhvRdvP+m7W
GuOdf5fGeCr3rsDQpjdDJyaHGe844/1h5EYS/CP+fWA1EW0VWJgcMXmHKuXquNKALqFcRd0VDkGz
pOLGmLjt8leOedyWE27+yzhVLPfWbOtb1Jffy3ucqKKMHQnlFFnLxGh43tqPbwaS59ntipfBeWoM
kIzSXo6OUfl8TCoy05olURsedgIwBzIl+paNsi5jAFny8N5p9saSZAL8NXYDdJ5fHbgqmcdPXXn1
xgIH8G1Fwb24U6qNg0AYKFazjY4GK3RYfHaPvvwhvJy6Wvv2Uhq3NAP4xR0miOB4psYsk84im+0M
mxtfIdzj2m+M67H8At1tYW+6U1fT5HexLyX1M9L+UV6rMQ9JaahI57v+wFu2fG/PsLm1a6SvQlek
wDK/Lp+X6lwbRA5KmrE7H51T0xsAGc+eU7l/t00OSirl1ONGUOHeTWyAijyAOC4LC23LTwCssyC/
FzjD7EOttiUDr+IvLKePOmUQYHCLcByhaz48Q/xMl/dBDsnXrEjuq41b9UxpwT20gQM56DlkYutL
2oCadEdTLX/0f8xKzqZWwnhopNXjAqpJZdPIPXfFL8+liNDerVbGYv1hM8amAg5T2t8ZFwir/Qmn
L3JZOdA6qQKJGeeeZwnvhsOZX2ddPCC3cb/blhOfSjfyYHeSmmh7rT0RXjFansZS44Db9g+eRu6e
h7mVeGBMwTJLNhGrlfbmXXmH0YjTWKZJtnfymAAOc2jKTXmf8z6cP+Sb4KELYZcQaqT54FsIe1/L
Zyjyjqd7Bg3T+O0ZW1Sg/glCRtGzBdckBmLrNpKXZTsQBCHq2z/cX2xFPc5W9BUYIK6PV5EdcQe6
6BcB7rZSWtJThSCRHKIZFnOdLJy7GmKF3+Yh9vPQ9DiQpO9c941rfkIF5Ay4VVVIxIqbLB0Jz6/9
6LAnPyIMIVVjHjTXPdt0xtnj9iI6rtvHpT9wAMySDRw1hF+iW2DUHdRW7Lwbw45bfg8SOU7rp/bY
5GZqP8ePfJ3ZFPEBhH3oUtxV3CTi2uQwL1FUKY4QBo159rSDV4/zJJxOwv1LnMgXi6hjFT+jqRx+
v2q83C9boY5vuPf9njuq72fkPYP3SI6zh8ISmoYG/eUEiWbdFI7GLjhtfKPhfbai4OFM9BmgRYv0
8A9bDG2Gp++ijJEPIpkzwgQjLSkNZjXtFUKfrtrHurlujQ/hvRrjGfdu86yk/90enT/GG+Xoritv
ylZjBzhEAKrN1yxKpcU1mylVCSWML2mMJtGQtT5UBQV+HuK3kiIQJfnwLljZT4ZyvlDGFDx+9iTJ
/kC7jjlEk2fc75tW1c0PYkI71xwSjvxx/oFYvkG9iXCSRt/FdCX6aURe8wS5cX+8TGbRFg9agOzL
YRTUhRa3doZxh1AkDrnjSB7AceOpNInwmymRZm18DBlpbJsaLQ5Txrkrz3RAvtqWZJB15Lzv2MyA
8gfEX8rLxhYNbUhxUqK4jfzXI8Nq0++koSJnmMzGT5OnuxqShMXEtmQDhTgYGGlxbRjVsOuDIHdn
GESKk16KOocVpehYTCH9Jap2hoNgHv+rOB9bzjjvxU+qz3HiUUjrBh5k7xlFDCsvcospWTJa1rLI
VDWXT/rtyj68SeRC60B/5Qn7JkbRGF4OjXU5UNhNYLDh8771jQNncDCFB3oAK6qSUH5hMmpzi4IJ
aLAVEN78apLsDC2BCqrYSPOJQaW5HbmEluhs5p17n4DUX95QHi71kUleA7nEoZX3Ovi8JFqljs68
VHpwRkWuwdnbT7PPWimPShNIOoRiEM/m6A6NCTrEnUvsarQKP4IHkhADxLbT1qJCOhVt6L00MJEf
UC8D+dOC4RToz1e3VHot1jXorRGlwwBGtT+8BbHIY4pxKfuDRG5lfAfPPVHfDSpF/aBzBTWASc6G
nCKGCWcPkZnMRkchkW3VaZTAufYi0w91oOafeUazu9Hti/DjB+4WbgY5WQK7954OmX1frwTaJKcn
SQS5u/uSP6xs9Y0OHuAAxSyX3U9MUjKzhcCqCIZgGj1uuVvoUNM+mSD1DZcEeJzIDWcAWXvhCSNa
RWb/t5t2yHj3Pfo6cXOQxyykgMzUq4IuqR09dcRLNuiX7uiXhsuEKnhi1zQ4DWdsHTa7RcpvNQD6
4nXX+47YtzWfPLxzl0eA347SFzx/CR/jDMH9F+qbFp5N2CfhLLkwd005tUiRa805NwQdUF+LVwz8
mepiDtCfaxIsc9/6uXVnqakPOwnGaCmLBaneJ2av1qt25DVgsMchI5vkkvakhXhQyVUeG3UWbcVf
KFDbRa4tBVI+3dGpDh/392xQupr9aJp2hJwI1j9eeMtxj0KovxI1HCaWHJNjorQT0gtNvuLIZabU
aa5gHLk3TkI3OBg3jpsrbA9MztR/JO8vaadgEvpH8iKD4tC5Pyu+46gmdDcpB5UdhHNFsxIiFBeU
7wep45MQXdgxwNiF8f6JDcoR05Ujfr0JCSXKJn6H17VgLFOgFMHCUI3IeaqEVv1zOFWsp9KGZdlA
CotNw0KkPE64McGv/BZTn6kCLonEFCTN9Y43dKoHT2KCD11WUkROGrDRginv3T24VmUd7MfyYkeZ
kNbXvLODqlRpIbhVNbhmFZuJM9TgDyl+0dN5reqiVVkeANIiIAA8120m0W1syZVeh8DIZihNy2t4
Yuj8kY7nfhY2SP7DnC/4bT1lZDsTQNHBVnnIfk2Y8jWyjfVfuQSplpmBIUNFuxrACY9Zc6davlYF
OoyWkQGTi1xFWvVj9NpHqpsyzHLN8SBu5mobl27a2eMPQAlNllYlex/Lc4JWNF4u3sDEuOHgwT+a
Sn+rAZaoQQiBHSwoXna+y0yxPZgycEV8Y3ddHAQO0YQ3eitwmDk8xbAJvvetXH3J1bIjzloOCT2/
31w0rQt3Y5zzE1F3fa6OaBz/KIl0aGY/I67coGy2NS6fj0/g+pjnU0mWygp4c3h6uQrQk0TXqk/T
c2TZBBecXSCGx4TUkTgL8zcqVrB++HIAzZ11HmKOe5z96On8eopn9TlgWSD+snRjTEyySB3UPjs9
X7XV/hyUfbAvhffiOY+6CQVU67FGOVG39cB1WX37JGw17AUfitaiNCJC91fq1Y9AGx//Z1L7R0Dr
bDQxDaCN+90h5Och2dIvgUdx59vshEAiufTxj81xTaTvXuJ7BG5zJ0XhIqmJav0K3KOHyH6wCV1u
5gSKQfEOwuLBKenOwZ1ZTuiME6/HW1lMJwscq2BSqWPqYwxE13K92PD/mpv+Nivqy0W1ypPfw2yv
XTJ7glFEYHCvTAq2neRo0xa6LpSOtj8KD0QnccvwOAPKTkbq5DSAEc1Lw52L6tG7MuGysCF1+Esk
LWZOZYpRnLEPGm4qlQmBe5hvLshNPnx37GDKi22aR56MtzkifiTwzB4DGFFpXpqWGIN1lpF1uav7
gVEviGcA719PfAwm/y3YklvIo89YHmVR8DPaLDrzHAd16kaCBnoxaWjopGc7zJQmSTZmuzYvHTPH
XLVDoCjq74DuPNiwg35x/gq3TGhlLXZT4PHww1+zV3aXNYsuFB8/78i+7/xokEJZ1dUly0ZucvBZ
IzH3BpM/CJWt+8SLPTxR61a2mSv/9fuwm07QVt5zkSU5NOhOYkBCuoSPzCySEMh58cZmOdaqKoCy
pWozd4u+XfjOnp4rtLOBArovSOrcIK4WSlRc5EYPrgHHgbHDHJkssJ07qOhw/9lhS2mC2NCaU7Jl
x9ZlKK2rd689GD92AYcj2rL/FDhtwra9m45LaUi1yqdzgzM4QMDVsLFsF9v7luulA4iVLJoR4Gu7
PmExs5Bmq2DCnfmNqCWFisH6aASrmQ+pAlSwKAClhwe7n4rtYxF7sqPOM7s722pVklc2duoAKLjq
t+9pdCxKVcHJeiCS8uDIiYGI3+qPHZo/8ShFW5EZJrICVJpyCCzI4G1AWvfOp2OArguOx4pk9LoU
eshmrN4dHIDnVssvYvZswcWl8Rgw7dTazY9a7IH7nfKVkQRVrUv5dpQsRCrk7zbjduptkIVA4keT
VJhcjacOWh2St0q7eH0QR0gWmh0i/zq6x28a57JpxrxlWQy5Nto9ERvKztdtxzyKZFZ603r4w/gW
PWVWSPdagUOS7YSfw43lLnBkh5Z54zT1HAf1MygBiYZYbAYahxhZ44HiatZGipl9JhSwURexP/ZP
L3rDYKw+HQpwGj8a7ajYMF8M9hX2O8S3uqftSsUB+68jfAeoTkM8Qbi0GG30bdJQht4aD3LzrvbF
5tlbNSHVnMK2fPxQ7Q2/i98BsF/xpaKH4bZFRgorV/UUU5U6BNDOJFTwWYFvDK/GTqGpgcKfmeYv
XTbMFNCjULQ2JQmANdos2tYzfDLNRIExHza02UufBHeq0HaWOTyb+4jPj74aod2p0+7bAHBbv982
zA5dw6rraIPBGgtEGXhQ4jaYsvNlGMUrY95pEo9ya6w9CshxzGtV1EVym/wQbpT88IQQlTWr6nin
GiajRgqaKOMCTt4huSI4KRvW73bDjC4C8ogFMCwhNcobbzfhmJ8reeyOc/h25McS0GPNo2lsPWoH
fDDmIralQ2fH+46CR3axCkPjDLPcWiJ9Vdbp+BGbBKnzBlexlUBNh/94NgI2vfeLU1ggxURWcFVJ
bqtoYOGzaizZEbBY9z0QO9+b3l0zMT4vRhnYeg6ndp5ayq0XeneL4BQ4pqmjrrSxLgmNdnCxld6X
V9BfYPw9FhRgUxxi1C/6XZKRXh95KH5lvPrkAIwctmvFbz1oWR6fukPumNeIlNe7z0upYXgYGvpJ
nx0VOHgXv3CjaZdhh0Q0aia5e+YU9eXtgwWYvOLxrrPF4sLUJLaBVYetzAUd200qhOeqOLoRZuXO
iZjzD5FWaAo9Dqg6H0hNj9/I4zhhjiBW7PzXbv1CEx3pCJXq73exB+/lW68YCwr+/nxDxgboIpy6
5j7/5patQFqGPl/e16SDDCXAnQQuvWeLbetSDKuhB/tU8Io0fd9kGkrugNF8a4YmjatJ31XTZQEp
Ex3IF9qc8zfa1myGqWa+Yxqw1QF+VYOO9fGbWCn8CmwtaB/7cro+ea1g/6op8E1dYAHrlTMaRrI7
hlQHwbOGuruu5Uhq/ln8an26RtH0enLSXWJYhy1t4JZ9ivsDdjcScapcWQL6eRyowT4RDR3i0mzy
DLGlxL9pTdIpdElKLLZR6Rxuw6wO7Dwitf5oRHmkNwfys60ryTh5ZVnEGW0cDMncfJefDyKw1HXC
BZJxVo+J+28Bwk5SC2MJySysth3WWVWnTIpFE+tKKLDh6lcTh5agFz2QTnd0SsHcGSY+3+TPxkoO
2fBQXX6tDJXxrBVvUXj/NDkgSFqG++KCUfuVRA402CJ82BSLPGUk3YjCHhtaOt+zENHqiZbU5fnD
6U3qzONn7b7YmiaPsy2NFHfigVEnChoRaJJxbkHznHjvmt9nXUgKtx8m3BI9v+UrBUGLKwVU6V/f
sjVFhx1WC57JIINmF67EzOoHxb98yblSZAouW6HjUTlOLmcdKIUWh7oAaVDavNls1x10NaneTuS8
8gTOOpxI64C3DtF4zTNeQOrKpnwoXIfp+CiInkbsRTYYEXAEKg/wevqkMUR4mCYyYoQ5+GPRhBAd
TFOg7/bFmlkZpl0ZdfOCy+qtYaxdZbULW1gSJ+WOwwcfqq6i/XBdPpuBmDWlHPeR69yxA21DsjLF
Auc9IzI2FlpFydbfcGCasHXIm7KApz9FAwdUO25jAYwFrG7nV5fOtCbo5/OX7BAdsbvnqGiSzpBW
95R32cNSvAGgyJfhgEmSFVrPmen5L7HQYUiVxTftEBgHAFzXeHEat9CO3J2JNWeFLP+BzkODHhuq
ddKMp8/pbC1RXH5KTWtKZmewOpt0C6TxPIiUkf16ByFFUsbHWgg0lrw9oMmTU+dXP3t2iilNOdfm
EERpMhKLdrH/nXpWKKC1mqBK3+lpO1DJwQ73oI5UeTkilJQmt1PpqiDMWmh8riw78XnVJ8XnXhUE
lF66iqnZew5InZ7Ul2YhM//o9+b9JFkWkN8/hvmY3/JLLUSxeSbKGcXpOLQJlgFqfLB1A3x2Nwl3
7h43LU8cPZsJHr/5sVDetBia+HmYeQs2US1IH8QfvXubiVEg1K04veya3ETpFTyq8Qps88CbKJVo
RlCkZYWW4YhijpxaYwoExdJy5DV1UGwJbdOBoWJszROHHQpN9OVxkvQcA89BiwEUkR8UY9esTG3o
/9U9OfhANBCk5UizdN+MRPLHQZgm0+y/OagZBgekr837Eeg7r5SexiawN5KmlwvB295GTmIohQbL
8tqCnMvfm+3a9mfjXVFj/jI/4SHra8sIjeb1l4ti5ut2KUs22FhJ0MOglS1dFzUAGKiYSL5fo2rZ
bHlAu/DZgFk9zbLw/+CQtkw2d/6RFcLu03b86N83DqCuTSHgtwNvdqELzYiBkYXjP/KSVGRjagxL
2lC8FcYPiJGxH9yq0DB399JSgsE18OI1UYxnMucwNEx4fDHDLIhm8J4IoYu0fAJ9apPdWyC7T1GM
WbDPFqIHgYJr5GRNmdbEvo1zQiOSTh7Z8owcJuFgPh2SYT9AWeFTRGYYLrI8PbWfotdGRNEinTM8
C706HLYopQ/M1JIBQB75wsRmCL1jBMEJzcrM/5+hQ9/2HL47mQcd7WjyxjR8DgHw3MNVJxn7Znac
NquQ5gJFNK6fh95Yh1Vpcf9MCDHi7/cCJfuKCtJC794sTZcLNRg9u5/YpXtbK1f2kvg3ibMztV9i
f28QYd/y8SdMTEk+2a32f6ilh6e0PaWgY73CjEkGePbg20u4jnWrVWEtPr9pgmFyOu45EHIAWDq/
trCa3bKU8rW8vQtFAfjzLm5/6jlMKj60uBEWuHqI2T3KyZg3n9P15q0a6g4v5b/Fun89b0Iy611F
wcoCEpmm/bkdJiklWH61ulmMzVBrkU3v4BTacFLAcjYnzN9Hc9fSKSf8jvSJB5trqY5EFCyb+uMp
4AE3cQ3puTFhhLDLa2+uxfXGH5rILnta3fnCdvSG7o8djQg20C2ks240i13jM3R9C7Ou4URdeLDY
2xG6t4G1O2M1L3aJ2SsSqgC8SV2r+NSXC5/3x8pfO75YkSUPsoGEO2MUeTmPzdCwv/aGZpZOmquW
E8utDtYmR9fqIo28JkpLXPRdsfvJsbrbb9B7BCmOAi2OK+8hjvhIqbL8qej6+2xBZx1mrXd32VgR
l7pOXFrWVu8MYB/ldzUkFWdm29ozpUg0z4PFWkuONrQJT0cakdZDOzfsHye/Xt3tTUR39/coFEMc
37hsV0FO5JNO5Rx6YGogvVavIWCf57ZH2vgH/mPg9SnkApNfVmtT90QDiy9MHo8stxSSkzKUbP0J
WpcpjKSCO/rOv5xa6+ixNrmeWNNercFaTsh/aeq1JWkauBRwfbXjwQ4EapgP64rVSicHXO4KkQSH
BwChwtWAH2sW4i8N3PYnvFsFmylY2ge5YY7iO+SkcI6sCjS6y2zIykw2B+wqe6b0dRLrK0Gjgs6J
4QveuHos/k66o++ylJsUlRm63bqEJ59RcqqQaPKHtyKyT7y3Eb2SNRgl0riHT0x/p331D5w90GJN
W9/Tc52wC1FO5/6TjS0RSEbvFLr/7dGSnZZ9yQDbdPXjBc52zr47Uzoh2shxojjNwJfi/ldEtw0m
5S3jt8pP0pTMwF15COhUu5U96kOsB2k763fcwG0wHh5bwC7L+NBcyPvAnkXTYe/yimYkypU+aSlW
I02hzhnng9LkSK8KO79utnFSwXBzakKRFtZcl6d4bocDf40XWTfExsyqkCuxCr+nb1+FOoDgLvFV
jTbJCwm5iKYCNU8spMx4BwwicjnRaJXOsYyp1h2C5Rg7C6P3zwKocBU1KGzzUFn68NXG2qiPnaIg
RScEh20isVZPnHxw4QsyuPuFRlXZQwt2pPga75kMUXfbiWs0BufB+WmMlQJADkQo7V8OzJWWqU30
hmieHLqCZn+gcmFra6E5Xq5lvgjR6JkZ554W+gYiQYo4WrXkgIqas1SwDOYpFrhz3NTswCaRWwxI
9nWZ3VQvHd9uPHdCbGxbz9BxeZdj6GAgZAZKxkbg2mvx1+PJgWmEhuirJBeA+c36VVAUQWhPoewC
okeEFp+qVFN4OVHuhWmSfMkQgq1qNDmKvAPgLHptYmx9ABHuqxJLV/ldD5qny1obX2KwyXw48Jy1
U7AVpuKcKlHlHxo0gzFhRsk8BdDaYOuBpgvq85LvcBCPiuS0s/cBr5h68pUswyHmKvd9FN9OndWo
d7Cjl2wr6j9QHZ/g0aA4zixtEQ5r1pkzss5TmMfC4SlFbcLizo1s4K0D8ISCiXlWH9JmXZbP7sA0
DOKQBr4jNyPYSXw19B9XXjeoyEiB9ahqljDQqrTwBdnddRrzAR0ghNf1DwDeOsXtOMMNdWa6BpCA
Mgh5c9Uszpr3QpOqWpDsIJhdfGe0PW7qQWvIDS+Xj40pC+r5OHjj00WCokNrJXyp7T08mystyViR
AYHO3MZdx0PmvPKCY9vZPTx8DmBrPUeyUY9kKfyEJIpLx+JKEb+LrvvJxDJa61O4iQZx5ov9fXri
LAKXOeAaoDDwP68blPnP5zUXekRbi5h7Ei6rVotLoy+AK3lnEpeQf4AUFaj1MZVvYy6amRMhrT9K
Ks0NECUpVz/q7v74SS93FIUP74o//o+pNY3nnen6Qqk9HuLGtXgMBJd93UUUxPwoACkHRkM6npmJ
zF79LnenttXicBhFju9l3uhhmGcZ24O7dOwfQ1aBU6rY+kOejdMVtPor9xO2BVlj2BfxsCCoNrFr
8z3filpO8eslg9FlOplGeJaQr7ah7CMcHgr9Lp0OrYqcD2RAz+4iq8dD1msvTj19Fyz4UWlFcQRz
+6i8wEwPvz/NvEgqj1nEdITjCpHacUmGuY+ZkXoa4z7MdqlvXlkJcdMXFrf9PlPVjkiyomAKiDRt
9u/lZO85Ldz9Cy6nlsM/wycYviMjq+ySEMCJ5fcBn0tEyxu06EPdR5Gu7OeaD1Ue6GnpC98PCBup
rV7x9LJY1S4yBtrK9Dvdy0yAd5xyQ7ty6mK4zSXfxwXXgMZB//JcjlzW/MyPhln/2rtSl8Ez71Pw
C3CcGyUG6oWjZeulowaRLda2In6fJGCwQRvOEIQvbeaDghwzncJGS1mjo0ydFfMgTXWM/q/B3QGT
nyK0Hlj0CWXlCg1zkcTmrZe0swVqUCZLlmYTtYeGH95shD1JYd2unkHqAOAFFBZkFO4MVyVHJR3F
8PhngO3PsTNyv6/p4tBN/jV1nkYFVc3NNelgTn2Acd0/FoUY2lq9MJQhF7DHly8gSu0rudYLMQ0Y
RTtnpWmNSqA7zYz1QNF4Y4w8KW5+Xhm0LdhbXWyrM6jJDYr36gSvoL+PSeNqz8s3BXXj//xHT/xp
ClVuIf6UQFA8G2L92+gEv5hTah3vy9Gia602ASNMJJhlMwGaiItA0iAan91AoQ5IMn8/IVUlgHzH
Ft+Y3UY30pljipWbD16eAfoX9DMSUI9rT+Lcoa/t2NLvh5P+fhChDlD/oFcWmcPoQpp5P2waeRrJ
5X+iAnCnjXQxut+dm6Koj7JVU5tKBnc8/50OQgmR0mItZtkC+AtfrfcpA58ayrea4QfpdkZ2wIl/
MS12trqp9EQ/RdcntwgdMmiP7GcQRCte6DtJc1Ht7b65n0FW/RnReNjLYNWrGoL8d5W+jOC8AC7L
bidlWhd4FSJ1JjGBOmmL3aKCIJK9+gS2k9GQJ47G2i+u5XUroTHOfVLg+Te/9ULG0UZwyu86Mo3R
RHfmB+M6ZcFWjvt2ZcwED9uZQXZRNOb4ebaT8UteeVfeT6WtZEGGUvSVcOQpL/xMtoG5TID4yOyL
kxVPr+1T3x/mfgH6v7K2fLUmoVBpsTA47k8wuWx3Q2/1xah2L6lTgjnpxsHlC3VRgpCJ+NPkTzRn
oH0w99TN23wjIshU7OeAxxsk4I2rrOfcjQorcSusamPSIMhv0fK4P31VyZ8ROM+eiKtEEiKwWX2U
bn6qYkdXfr7TylLfSiDzu+OUVkjld1R8v6m9MhGDYfGQsA12gUzCUma9kPWLycsrf2t2jyi8nA0v
pFjxIGoy/+bKoD5dPP71v1+g7h8e00k3yt7UhYxTOjPXPLxHeRAGCFp/A/b6Qh0rMAbAuJHyHPqG
H0d9P0iKVm1KwPcVEGb3mRkA3wM6ysN23H50qVg8PXyvYqCRsVMB1+dpTylZyS+hHaydZx3ZWm7P
N759H8g1G23G1pKhtR/XRA9DZlyhU7Xk5EFdjF/txMwd93z4PGzNPmLyVXxoEhOtXZ8plxs7TbMx
cz0S5URWXLtH4f4qOJb5YeUxSZzq2Xobd9d/TLA6QRkp3edNTc17KCbY2laqjs4BQ/G88VkK8BkL
mo+2/29z2C6nI791DNDU5CejqWdy7I7oW4WA7uDMAd1vqTMJf/6OhrhdA13a2TnVu/2fAjuVlmyK
9rFN1R/4aL9/JwPK24fgsgJp5gPkYZB7AU2ziwXAaXNuQ30OtmfP1ISVO15XwwM488aC9K/8TMcb
9NgdW5vtuy6Yjs9rK/W93A3vfo9fnF92BTGsztQTwkaLMa/iOZVazXbUG/RV+iGE2SmwGctEP6EC
h60iH5cLjLZnmDA6A+DfGoTzzbUH3sLChxugoxc3kZ6ipfAnCg8FUrl7y+CT5tpcXm5gEBmWjwau
GbRcayQHrPeWf/dLQ8QxWKxjx4Cl/d4t62pYPpI4jRvVm60z9rfb52WdFm0hozK36YeISVPjtizl
Y89FWMKTZ4kEmBfSBYu6jFCnkEuoET9ERuzKyFRd9zoH79NL552wkw3d1k9ppxzR5w2oDVf9a7Xx
QEuhIPbCrJlcVwDYWS2FdXdyPmJ3cuT3Zywpq+NQ7F6/fGOvbyajWZ2wQIqBTNL99Mbn4XgMSgXS
oGKxFwo322748svt+1GkudUDYwTsAyoSgKihPz9Vsyp56T2gQ+4Y4cVmR3zRCNyxKl/BqkMvtu5/
+NyeDQIH2thwelaLrtCDTlJpaMcqKXSpHEhskfcAav+ZVa6pO1JdloabAa9vfiXQq8PN9f0Vyxqh
scf92MTe6nRxFJOsFLhWU+p3Hr5CTMOmxtP+mfctnt4YbnzdjsgyaPDH/3EKgghSyY7WxYoYbOoe
pAD+sFv10hggx7R/f1Kugfb+b40glcE7vRkJBaYfXAk95CVnhX018OvzqLMi041uUZBLqOcg+DfR
6bhIXiH7NkACNXI1xA+glELg+RCWPg39GVoD3LVIT3wv2HObLTIdk2tbuiIJ7PmFlK0OvFkEDfDY
qdbGvyXeStFpN8KfSDZR+djMuBAcp/AfWfd54tHl1i9DmZKVyVfNyHwjvjCsklo4NDGUqAiBsAXe
WZmU+Em+O5fg6TOt5sdtGO8vEShYlI63Jo8+Pal8nuOuga/jwD9MX8aOk1BNE+7wshvIS8SceE7Q
KdD637ShA2WDiPccJPZUXAsWmGppvl4esJ8DNc40vzwTv+fndV0H2g/oO+HiwD2rkWTMlp1cqU3X
UfN7xFzmXvc/fIstXyusRQCmISceMCJeHFoDcV6q1gCYO/+YojIb57O8ydooO1jdgVBIOr6JlLnD
a4XBzyHRhErTBaa5aNisObikCPzp+J9+4rCHc3zX3NatEEjJkxLvxrZXJ8Mu/mO85m0lxUvkLB/s
HZ6+fPOX0r8npSoMdjOwme1gl45NL7+Ck/+fC7Ah9cLXvYSfUYXImAvalE/yBa2wrHxAeHyXV5NM
li8qHm4tVRrKTzpZ+gYeJGhTsUUTqBkFA8bRihtzBaMV4RlZpXfAQFPuOUEW6x1r3f/qb2jI2Cqo
qoKXkLoWgJzHta0ijKCQD48TJ55crV35N21KNN9/aGvtldgzsD/7onbpiSC+1TDzUBIt4yB/u6l8
7HfaiowerzUKnpyrlGaHsay7D6GYkTtHDqYmbyUHVraGFA/oCV106dKXKWET5gicvWhYYLPchrmX
O9iO+nYCm3r8PWZUMsWfoMfzQ6Gpz7Lga4UZ8p1wEOffw6BUUNLlBP8/aLBgS32Vz3w8IUoJrKq0
yKyHoxxzm01wkAeuYMSFbqDq3auMPJCDCh2sYIPb7OOXEA4ARHTzYozk/EEGehRIqoRbfV0E6WZr
/dVAzJm8SiDB58NwaGGN9UCFLEjgPbeIAwgiCxXeuq7/+n5vY88L/EY30/PII+JyMvyP/AGp4ehA
vpYU8+NerNOMC1c62IHLW1jUkPUVKRQ57nLWwaoduflAIOYZBHyfla4Aau1exE5UTfZuC5IF88pn
gVnzw2pF/Qzon3mvC84v/0UJddSCjay6kPJ05QvBaT1yFJ8cRuAr9Ued50WpdTVbL2tKEmlE4hLo
D+1EjZLLlat3YF59lsqKKQvt+EZqoyif8nVltLW7+EI/X6MAciEvXBkKgQ1iavtuaPj27q1xYe/M
RVCbGnXhaboIYPV4/8dvMJWNtaytw4kRs4zMqWSSggQUvD4Fpdw3hdZJtUBISfXnJR8NY6Gewci5
/KGP69bboEcXbIC6JWrvP/cKPS/KrLDOwl03gFZNTsVkdOLYqhALc5KwUNpyea86M2WzyTBsdWhx
Ummcu0g8jSCo8NnOOAvwmSOf1qF3Wu4tkLI7aSyqvcCfjjmQxUZRr4sbPa00pEqt2xROjAFhAvhM
TY4TBSMNAGXYN6yxaMvg2EQRe8ZLBm40njPAS1yAmdtYakV+eBlRfsSRUx0tewu1CGT/AbFd2ChW
2uqPYHcX9ATz4lWHSfCptemkgWB/UJhFaObIA5KTBA5awy6OXI/Hmlr5pOXSIlQ/tPEcTMqtkc/6
chnQqIY/qQvvHZ5lDq20pZRYxPydmJBkBdVjvc5GUd9wAAWOpHw+9gqz5MqAynIHue46afjWtDJm
uo99ojkSvD53JOxVPDnbIgFLME9zE+HgORb7Pun7K1jbe+L1E7Mjcxnuuwg6K9qjLoagUIIqIcjt
B9kJVx2r1/D39ExPSdcaNJx+Gsn5PD+UCjrm64wLf3cuKm4snUkBn3BBLdJs8ZQyk/mN7jZvEtjI
eKV+J/7/582DbQ31FVaFnT9WRk6XvHCN9XcIxtIg0o2C9COY3kwVT+sHdBI6fgOl7oAZKk7rF5TQ
MfB6SrIeb1JeS7afnLPjjFFTGTHOUqlAQ1HvZn32/Iiu8RKsF2iVsZAjXCcZ1UXrVcjc32QnpeBI
Y2rWPos59OLEYFUoMR0268qfasheVrjzPY1xC0l7bpFMxvlCAAvLm+3AvDIwhrFQxut5Z5IYiF5g
s4b7lbrNT3vSwUnuqCPAny6Z+RUmbInzQRZe+chwGtuBRr+sqTNCx3SGrddLkqelU6F7c1Ize1id
M0K1X2hfq5quDFSVrzkl/N6+nRuORwaJceit+truw/N/k7WlJSU6WRIJgeEHAsfWdJGVwWnJBUaP
xD66eilRTOZ6U8HXp5Os3adXO2wiKq4lWtR4Mv65fLiSCnLiQxQb5bQGj+9fKaThQkAUK2tq7IJo
eC5ouE0Y56cd8N57w9LV06uCfh0w81J9d3aBiA2drhLC9gVPFu1eh4qCtvg4fCKlcYAk9f2Ox99M
OFf+GlMU3oc/6pAp/i8GJZVwqHtzwlyTaR29i3lLWtBLz0CIV9WmjynumCWPc3i9TuBhN5mPdWkT
4xxCK0Ngy8xSdYSdtPp/4BssXbsTm8cNtNBim9yc0y15rWMQmoAdxleJOBXw7y3a4QP8TBEF5EJk
Azlpho7eMcT+wJaCPM79oPGxHlclbeVmTKW5j29BIBVO4JE9sxdu/9YCAMhbWA7K2Xgg18hYCJmx
NmQB2Zi6V2v7n/tgVq0IHqBagL5S603ZjFDKUZKeZujWJ8SVM0UbC+aQkatllxT+opJrZKCDA9iB
Iv1MyG9fEMJGykXAY9zGJmS8ClGINxC+T5so7IS8ReCcCmIFR8CvyoYeIJE7I0GlM5DEVVnHUF1M
V5faQsPgwzAKZpXNhsZh07c1YeXlNtq+gD0Br7LfLJRd/Fwbk7+Aws6onNbXekhNLMMx7Xn9pFQw
uw34ME5R89+siT7LGcH2EYPIh3aw2EOpsVPu4TpmiNXhXz1+9z4iuIy5ysfk0EI3w7PKskYHdOQa
mUfvlM2liwu58FtSW+KG6Bm/lvpXJPio1IGAMm3kdIfNu3QhT1HkUFO2QMHLiHiykGAm9aQPKoss
ZRv0XlxM9KAs4toj2X9HuJykeAiNywD1WCCDqVZRivOHpUoFDAUfpGKildFB1E3bt7BH+N03DDRf
GDo10uEFeTgjPtdZ01OHUhdAA9SEjiBl3Gj+1lDD9jZ1ctnZXzEVNIInTvvRHbznEnlJBHbOkXcZ
EVrv+OifBAQ1YJhiV8D6xJ12DBvWjT8tYvNhG9ZwNzKynYnUdElJ2kEPNo5AIQsgRRs4YqLgOZdh
czGB9OCB3reMKKoBB01wTmjNwyRYhjlGVUFVzNYnO9CEmfAet+W3zdvrszVOUn3DYO9lgoNw17m1
vsVpIkC45IfxDz5B9QiveItvPHXkWfxypW6S2svgVvw9JoB6J9Td9ZlJvjhCnKcFuiFAoWp+VtrU
VDwmi8sN5PxdKTLh+t6VbBY5Zz1Qp3JMxCOsdQsduHS2wBc+60Xv6ML6ne30MayRhHgdAfwHBIji
81wU2Vi7JOcjEMLZEjsLOWhPktc1HqSTbWvzhqaUQVuJLuDWKQWWigH48xpl3n9itUNnX8pZ+66/
UDtPL71ZFMxaF1UMHFNvPpjCROqFsXRYfP0fBb2BIkIBmW7G6o85wTun8kC5/L55/XVOWGYlTzv0
sbCsvJT80bmgTJKmpZvyX9iDMFMAex/pb9UbMebElkQCZLhJdqekvyMCMeNUPh77uIwLcCtOm0MB
+q7BfXr8O/wbB+vW+AJTeCFh9hlQVvNIrEg/8JiY2hgT1aixDYBFMUfHp/eR8XOzFT2TzvSMM2PK
MTLkb1iMdBRiBMaIEHkbTQuRhRX0wKRLhDiam9mXFEJwBPzqTwXnO93YCHQBs84e8SU3RqqEy+p9
MezY+Elhwj4LJW/0gEvjRIL/CY60JQBRSXxeemv22obhQnWxFfIv9weTeJWTUInGAuSOJKLevdB4
ClWKrFnHVBxJmLvnLsYQHNo+CWGAr49MzUUlsQyQ7Ps41vdHLtFyKyo3d11yxD6E511Z0EXbJ+Pj
MUJERJQUFn42HtEbHh5+FoXszU4myvMnXjNSKIj31vfEJjaaS5GUEbR12ucR2viQMvNsaFgFb67Q
azHuclBW8Ln6Khek1dAD/vr5g0gAgzWimzu0dfCvI6Prnpv6oFfWJYtdkUMik+ttcniAaU1NuEPP
3EPU4gDjAHnCwsrkfLEUkp5IWS5dInrknREBD02jxi4QC8kFiWNQQ8vwUztfzaE+kvZuAoFgxL6e
L2Clx3zNj8YpycIrSorGsRrxzwkYOGWk512ebQY2y4vw+8KvZRjnQQDUAVll8SNOhR8b2dg+iVUE
gn1O24nXnls1loSr4Shfnxp+TQy66V2+DacxVrZPJKD4v7HOKMUX/gS2eo1MQz6IaXGJVhgNvbes
kwgVQYc7DyOpabRT8gKuaMEPzuOThtiK461Uou4mOB1upBdP+LBs3aNoJOoAEuYDHc3RXm/+1X3W
WAliATxAqCwEV2OjsJxEHF3mfrhZX2wGGu9huXrfW/xq0dRMQiJEH0XxEur8qwdD3Xr2S1748Oqe
V0i3qY12mGnF/ta2WT9ksxx8gQs8mAqF+YCOw4RFoSr3TEK3sLZCg2IJM+TERFsloaF1tfoxWBJv
nOL9acusAFHozyAYyy6ZRlGRPmg+kal2q7o9GyeyKJMmb5hR7SjDKX36W9MG1oliRxZb6r6UWLj4
L1aPbFyj9nJZjSKqouwDE/Va/0WzPMza79sCzYMhtj41xEmaANHd3oQMTaaG+u4az0fG0g63Flqz
sltgQTX8/ZOQIdyuLf1ke3npIUWrFXuB7jhsCmQJQYlpebefr4jZAdgdpcjTlO3u8tbYeCD+6j3A
4Z8ETT1PlgehetvRLiJ7NlyPfGp1qklasQPxWa87ODlYFjTbGfHRtYx/5dPMSfPgVvud/TjDjmYw
fRONJhcdIoX86pNaiEnJVULeIPQry24HpJwu3y0M+Xbot46m8GXdN/+Rki2TpHimHlIO8Ic8Mppg
qbGu7YiXy9PNe96yJBi0DSwbB7c+5LuFcR7gEnBtMGkwdvdhD1e4OMoEZb0yyq3qaHaCch4LFF/P
gphzAafn0yYYsI4PlI+nix4PSB+sbLPWJPN1coCoclARy0ODsdE4MaJsF/VF+ihX/RXgbPer/XkA
s+cbEMXG9xBw6g8q0ctlzLdE/3MmC5WRuZDh3dRu3YrC5BtPuV+o4exvXVdt+xlyCX5pRE06u8QL
y4/5BNJ/R3cvdjA8hHaTCnFOPVqNb8S1b7e9kft/vdRDsiA//L8Z0a50LtOYufTajLYw+7m4NkzH
KAgeUyo4QVT02URnH53SMme9JxSJKidHVsWJZWVAmZt4SobVhR32auEGUg0YLYwyKN3j2TK3wmf8
xzUFoLKh49wDB8NYI3zpH6KIoZdGHzvKcxLn5eZ+FtpczuaNGkVJZ7maXoQw1BsJ0aXOGGZMGI3n
pdwHakFxlDqxvRac0GqFBxgQwmfxhgUHMNRviV15Y0SooXmHiSnhmtJ+Mr7EzvzWA6TeFrqxA3rn
S9/qzAv6sLsso+5Rc7MNzGSYCnYQA3Fo6jqxYZo8OmdsKUDGulMoWX3H/OjA1JLe24Bt3V1sumZN
pQgi0zQkrLvrY06k07UX0CXt9ItrZheJKpo2elkxEsTtvfaPQ1ccl0fT6AzhBbrDmzN143Uuky2u
WEHIvMZN3p/dUC9ZecAoH8cAHyekRxfBaBFWgiImTQlV4NiUEr4RRDdSRDLiYCvzzkUQgu+pvEZx
XPvwXiIV6O64CV1S2RgKbKooMgfiQyvNTxUgf60RlDcKxPA/MktwoGhFsTDQLKZx6k5M8dPsACij
fXCmHrIgyp9gY8IyfGYwwyvQ9cpv7FaFzyfk8ftQzQ2U5t9VeOu3SxwiXAwiM9432lU1PiDldvNj
JubuFivXHJXpiR8C1haajZ4Z1WpGv7QMljz+TnscPrLwurspJhUyhsSLOBbnM4wWoG5VIL8Lflyg
q0pVOm9aqLqA9YCfbD8k7hosm9ePt2DyRtTULIWVydU+8iJHznUv6qL7nLNv1PWPoTZfSUQVIUM+
YXfdQ1meupR9KnxB+uFMCy3p0UfhDusc2WlGpb8IwrI0/1b2IJ3AxEupccrmESXv5SmMWoYWJ1Fq
jrTQ4YbFczGd9adVEAmsdfR3FMHjqJR04x8RpuFQkzBQ4BskD5dmqiL17pDTC6N/2ncxqpPeEL4b
r2uBDhoh4Br6cHXYpM4YHhQGgoPuQPCEps/egZoYM+DZSzuGxj0QYRBQCHL49iXPdoj6uFfV285g
Y8isiCGZD+GNw+b7f9+//WUTzRYTyQJxLdHstS+bezlurHOZSUwNSZm8BOzgHXAfSTzsdE40/Deb
2oDcl9ozwVS8VlVYN1CrSlZkgeJ9wlOVEQBgWthMun/N1GfdblfouuEmKHVHKK4ARVmcoL4LpHIL
j1HjwpZ4NEqzn5vAv7twNddHiRynCUIvCiAfQa8Hz64ynOpffry1cVfgNI0BG0ByZSEtVtJgB2/r
OKdg9VNBtGh04fHv/nND6DXz0y7x+eZZwqECrDb6hT5+JKx/lVXVlS8TlG1Rv+g93nzCjeAfsbqd
//tOT756yS64wHta6P8R9N/DlMyEL5TbL+MvcegPQA8uCYIwfNIL0ZiEz6c8sQrtvlbl27ZdWLin
TtaLKip1OcXyBQPhsLsDZfrwIAF0nNXNZSmZdbmnn9LxWoCde/CPMfv/9howqIi+faICV1BQebKK
XoBkO0sjo+O8eTSGNvMjAriFsSoe9Di+FBZnDWaiI69WT3Zz4j45dfE9Fuy4adPJj/xcrkxuGfIW
Wem7V54HWd2JgW3G/aGbqHQ2P5q5M9/b8rf3ejcmijqPopOvg+U7ZVq0mrNM21M9x5MEzMtTu2NJ
Wd2pod8SM5xtAXPO2x9pZUIoIvCpbcCSBvmX2F2y/vkSgHeb6F47B05kxHkVhYRnntxbg56af8Jv
lPZAsSS721oTlVy7vci8u5gY2234RpZuULnX9O/mPk2MBWe0CvEXlx/cwa+pFl8IEDjTvtxfHr/K
tl8otZQGbVVtikrWCmBfnUMGVktP6JiIP3kFjcpj1Fxyw5o7V8UV6jLED8dMuRxbhmhNNqXMauA8
XpmKstrlkV2INrSEoTFKwjKr0gT8ovBbXPZBxBWd+dYQ+FaWuhLGRdceEUPa1M1fcVgjZqm2DgOG
eqKPD8PsbBhPxgZlUGpwl9ERCAhy/9EOAcRrCE78VAGx8zIzbLXlp5UG36cSUIBtvpDqiOAZ0CBu
GvRY7NNeD2dusD4XQgs4tVhT12D8pkSn6oUMAktqiFOuDLs/iTxgxXUYkI9LsnY/AUYlGQY41DHK
Byb8Ndz3HHapLWcFimVGK0QnpWiiyjCVoI6NtwcLkKwY0bMgF36UpSNfR1BRxci1xVpLtE8TjRCB
y4zTx3cqKLKllRElmQGsNb+REpW4uskzwZNGt7EnGpDJVX1IfknF8cJWkbYUHMeAppHpS7AIEgTK
LT49W63c/UjyCM5nw2bUBSfpt13I52dB8kWH/ssIiik0caWmX9LJ9N+I6cdBxqd+cTJJhac6AfUr
6VrpxobZkh19KitEviyLVlJgFgWv0MBeZ3JPILUhhY6kqXaDQm9F2YGXYr/FHDaAnN+ceIdsDPem
f6PsFcfeA5N9rCs4gmtAfbiYFavta76wLgbPjE+8xTSS0vc7WkxUA3KpWt90dZKJ1OMVX2ifv0JN
SfYpfb1j3VOqIUvMul0bVXFqWNe0Z0FUxQkUNZBcL+N5Zz5c54J07BnNdFk1iQilO1NgieXE7VQK
PB4gBhzsF3qzPSwDBUYEU1wIEZywTjJ2GuZMtls3Wwm+FX5yUVIUNOS7acCRa4LuFxu/gGNUIyU8
7XpnY4p+vYWZc9zcOoVLeFfT4PzpvT9IyXjxJ6pNlpFooQhvCDW2NitMg0STtF11rvEuA8+fXOaf
7yIgaEG2/pU2Q9LRdKMXjnCPTZ77cKoFVH4gjtHj+XSYM+mHPDndaToDGuS7Keam4ZLdZ4mJh/y+
Q8Qb0nMS8DIy87Q9wUUuwSoLf6mAKJmyqhKSKKOrGNBMyInsALm7OOe2++3dzco8PxgHlOUjLy4r
Cfox0xjIBldgSqLX7ik3yUabXutjsyUVKC5MtTJpDILI84DXSHmOywD1eQRMFTOzcsTMGMcsQGRK
eUcbiSo9KlOwI3CydeTkqzYNTA7O7cdqA9u7Dncvlo4ATPvu76TVC1JLXWf+Hwi/VY670aLINhY8
cnPBG5g5mviaRTBCKUTyD31sciO3dW6qKN5h0MI3XZQUQXpRDt4l27ALVRIZ6CG1fmw7eE5S0bAR
G5OXhBPVMsbjPG9Ql58OdTcs3PNNh0GZolbFmHCz+PjJcXfpcmWnKgtbNHpdkpu/P8rWjc6XCMkM
ohY4wRkoaJjpCl45G/RX992dvaQ3yRp310noIMP1Z+O1tPRzhVNMyJpc7OOzuGg2fUNyStrNICJc
U3OvhZuwqJRyM4YkGYbCBd1D+MX/fW25oCav7dew8y1LPv15WavrmiNimZRNiRd/RU4ArjvFkyV7
ab7U7Qw5mL+g7tkVMABT4/okmpjXD+7y9eWS4ZeVXWkCFgU17mGHSUUC7FHlGEfhhKc+xs0h2lc6
78xeaNZYREalDglcH6vcEw4DOAGhy83uypeQejtra/RNUgomy02nEzUvg9RHt2PwVkNuwK1mRXz/
tmwz7DEb0Fg3/BJvO+DJJ1uT/H5SuKmKjpkkZYZowXs4fSKJTlr++mXEzhMbhIUZwMRb9nPJnVJZ
95fshVotUTZ+r7y+ENmGxLTos52/ubltZwjFzSnUCeGxmh0zhSw9Lsgn457KGV6m/fxP+jxQyfFF
FIbDxGAO1aQW/25OvYWjvlHHD5+0qvUXxu2l+ayOKM9JYTARbjsyM996GDh1eSybfcf2UjKQiX6G
Mw1zC1SgQAMzPConJ2uMx3juhVcSuqQu9KNcKMMN8K4NTZCwK8x/8DwgPWrMqCTKqutJISeEUWwu
iuPUc5zGraQU72G3SbqN1VlpeUmLrKu0jfJaeNnYlkHDWKSYCUNXDzGfLgjuZlV1GWePnjP1Yzot
R28MmzrUr7AyIp8r/NKU72VUy+4NhFWEsoXzKpM50jIDgU9zTMF0jqNAww7vOhngqyTuKfSluy0i
RZAscDNlaqenkfJo36NbQW8eWosfJZ8dR1nbKMiiQdlpY9P0V5Hji941WvkcS7fc1VQ858QKAu2u
BhFl0ndDAzPzsaYblEEiazIeA5PPhKrLsDsq7JgtgdLiaKGJjBnlf1AGXl1EIZJERA2QGW8a7LA/
HyA1/3aeQCDGVImnb36CAsm8D1m0v7CvRJ5suZi2n9frmZcTVyoeU1PpiyfqMew66ykaUVZxEOH/
S63KkUB1NKBxrSD0KuzD4SpmtZg4ISu0Fdlx5WMW/kWnuzPyuAHf4duGH9WRk7S/5v7CzuNDowHO
iHpdXygwr81GFuuE6U+f4ctnIN3rDtSRG5eNcHNOhEzMBhUuNN5WQPq5UCkxXXNBkSjZYDvleqKv
/OT9xsqcMnVAGE10YgZ3NU9BkBSGcnE5dFfeovgSZTwjDGPdfJykS9xslpLhdyH/msuyDK+f71WA
Dp5EkGylzCkHJHbMCT2hTs9P67pPHIDLeGJT75zISwKOfopI6+QhLPeTfNOPgRiq1uiBK7jeu58g
yWxz69qYUuH98DgclzwQ05hxhT9cMA8RzKRM0UdoQttcPAc7Hdgor1o3oMtqGeiVrxUGsjRl4v97
bjcIrCvOvgrITCSx1rtivauJH+qZupjp7hSuNMbJ9lmToB5iF5lhhSyQqfk5JP7kS1qX3HkCW4yi
ynQtJu9tAAmqu42gSwdBI8VChQpqwrwPOPOEyAozU8zaETTrzfZ5r1Af2/XDHNaZ8lfvfAYoMX00
vGIUuZwbFrBaA+VRjalevUyT1VXLQApzTQ+8QGPFXOsFor/dGPDRnxvDqAsvA9m/ewyIxxRy7SY6
KPWvaNUqEFJOogizuGAzrxnTgf6a/dxT46O7Q4wiNPS6KDce6MOAa7wb4JxW+cH8iKX0Tx3pe+Co
t0gpBtMYZvZz73uIIPAaUzY5mcJ+uIGnY7aptyKJbFaaAlgaaBYQIAVYRZa6uA4Sxg3riUlf4/Lw
s6EaIYyJCXuka7jH5NrdNu8we1RV9SPnSGmN5H2H+p3GZ+8hYFrRFKcY9nDa/zWKnKDdRlf2gMhY
PnwYNLIiW5yGBHVMPRVe8/5uUm77wCZf6sKOaQSPdeZEoay59gzP72qh6Iq2kmZZ1ixHIFYgczqi
IdJl4pzuTTOOsjvc8SN+KAOFyvLcUpphrQ6aqRI0FUVyAwDDwsjfkE8B6jPPEx9aUkb6gHkdzko0
mhUIZj0yKdJZJ2+xI1rDMBJ/fkMAYXwE0X9/ON8hL0csN/uPIC3VpHC1fd2FDeVksQx4Z0UaUmWU
swzb+3h5QZmQOg2TevYZRyxN3PtVrbKmo62kgpjwRD2/ZqRl+RtVcmi0vzc28e7vmptHZ2TozMb+
M6wnhumHt2rybvXymm7Nal9JkAsIliiRrWLJveH5CjZ6t2XKZkhebPv08+f/57jG+L4lT7m7GJVJ
DKgKDvttVmTFyhxoUSD4BNKBAkawE0CTm6NNmQIEVOI2SVfVkNb1sLoB395bibmUsyLyWGQYEt4B
15wpVic/+5CBKUKdIXTbKlUn7f4qO1cDORBL1qPnHAH+3pn55OSP2MJU0uDaenjljYvRbdWAs9GK
0YSfx9fY3JCsG/ZARek0NfH6YrAOd1GnRa+5yMj/U+2GwG0eGIWQBs8MgH/4kuXRgCUNsCFh6iUb
4AFNqBy/QnRignMDIJYqmo5vhSh61joS4wGEFD4A38CtOIWXR25QSTPeH8nJQiu6+fdgH85obaDn
s8Z8/TtnjhyknTrqccRN94ue1HEqHt2gpS7x7sS9XZY3u2HpAQnWyMGSDxDn1tiYmlHk4q4FqauR
exKViEcqYOGMFUwxQgSMESMtJcj5LOFpj4UwPZ4kKdMj22RgK1Q/JSqZcicLzCrTPVOXnDWcDLDT
kzr1f6KbxeueTyLgv5t3RPQWsfdqqOdXktOrbsWqgMxgmL5lLhy0VYsCMinp/dAiDqjjk6/NopeY
DktLu3kyvdrSE3TojsQpVJrCNbFAjHd9bDAAsOZ/8Mlvja1EkMmZozTA5kC0Al0PUnMPZPRf8g6m
1fvlHuNDSrvSUvXqpLcehW4cNB5mTim6ExytYAI43Q9I41g65LPqf/C3Xty3YDcStkoU42JpRFVB
vMw/eNYTtyevC2YjOrd5G9T/PFTKmGUtIjp8s/yW20+o4eWj1DLtpkEWxDfYNnNh/G2vrIFRjgNv
/ZdrvamLhaly2MGlAnjq1Bjkt70x1MDpZhX8mfYQl7AQzBFFbHXvseJv54Ddgcy2yjENrFyw55s7
Dse9hPssnxU/ShaOTBkqJXapOlDwZHrZJDlL7LxPR5+f8Nrga+yhM+HDz9/2jri2LNuGiMf+QXWS
VCZW4BIXM5mQ+YdhesKlQX3wLYZyLGkk7vQIySNXnSzTUe8VtVwBQxu8gBFqM1EhVMVckxermK/d
4bZxiFSt+dfXH3ZY3WQCdzb2wfFHRvbrTu0DXlofVzkeRGk8zY61sGUkK9Y+qRpzdEe66rp8Kns3
7oUIzduJsqRugRM1+zsXHv6zFDwIZqZ1kuJE+qB8gfPpLNHjDNLdf3VNbxgWQ0oOqgGb0ptMCOPU
Jje4wDKjwSySHb8b7yERdmoB8oQBI8375+QcTuorD6mdRlj3EZp8xBv4P0synPjOqZ4iUjL7HAJg
O1djdoa/j60MNWTzHcuEQbmJmk9wegewJCV8AA/S+FsL226YNtj2tSiLKcItwx/8icUcAwLPMSJG
g6wnEpf6sFLRzxNz02j/pBt3cuge/5o4uLNuiZnVTmZYjdFEJhXIfq45WffR5tO9UraCv4PNIM9H
7zFl8+EB7MySQveWDWF65Tur079whMPdBQtPPT1vhqL1y5fjQ0PkTxOonPKa3SL+qiKGtLhe2KmQ
hHuMSLA1WNydXmogVVcYPEhfRY3TcgJnVX3U7WttvjZl0CZyuv009R/sC35a8GYyTEvEU17fnKlr
lhP9CrhHtAUEOSQ1BMnSQlvoG/nXPskqJo2ggCZm19IwnodogoUNr7Tk525dxNHRRYEXzkhC6xMK
MicDsTrnMI8SisckCRqBQSiq4BzC90yIfnWX00gO6YFeEWXm24Tp+HldUuBG0LsYjOanpPD7bx4D
rTyip03gjuSTQ/kaVTBBN7WI/3R4kOMwoMZTPXOnz7thqhbWHsdSRwqeaQStnTLZNAgrO4Hesq69
2psvPmz/UF9mk3N2doyDvXAReVFbTWAR5MZXK9cTgBpl7yfl27LYfWv6+2VN6KvnKOoNWOVaWd0B
uyxPHTdFHk/qFIoyEXXGAScWGS6PJfQnWxvuYrIcuYyIIehi5jbmLytMIRM55+ICQp8i+DF3lt+L
qkcO040ezrqpiJdBHsPIwOCWXQ2taiD5riG3YirMhIvBv0dCyEWa+astJ+t+bE1wY9Jj5z+NnZ9D
3at2aVwj3ORFNBfKpR0vdkZbS/Th8tw/Yr03is9/UIOKcr0oK1HVOoLe9p5jMa84VUR5w+D/YtRT
yI0Vr0qQnHOstojqc6sJuzH5I3FD1axA35GQqgPoIzmwflsMJFRZMamNjhbCKOSmaDaNbtZfhdRV
1eoxH7ZEya9f8V2GqKtDMDmqZKheNEYz6yx0FpYGEbrkfCFh4J7FNEInU030CPZnwv/6eo5Usmu+
bNHHTyhV8kYsHVDc0XR7S0+8XTylHxi2yJAy99F38uhVEeV879foR/916taolSPolvEGfGzvOLbf
LJ5OPT1lDDpUZxAD3onI1lI3KHT7RUFAodmuay8WU1Y/ui0nSFgyIjfaxyHV2IkPQAq3pMqCaco7
tNGMSX0nYRqbaB0YFhJvf0q/HAplPcSZWflyorB9rQ8e+uHOvfyej1iVo37dxKGIFeGOsAllVi0x
VM6gHPvYZjMGyWfSkgSgZf3E8qOxWePBxUo8ZM1uE406P1XTmWbmBC3y1t9UnHfjDhEh3ap0+Yxz
4mkB+/xkgvERZ5Fpb+ZC7sCIHnMKGt/RiIthEr/jUjsk9KVokLCZea8g93sLyghy8HDynin1y6Tk
I9D6TCsmmcY36Jmeq+H5O5Z0wO6Vc4Rj11UFZ3cqHUxqZmjFRfkInhS3FfJ16N5S4DrdCdLOKGA6
JCGKK1HiFYAGhpsFl5aW/0xJVYf6PzbG5dcwoQFJKTKi5pxzoAh3qQ6FVRdb11SRy74AB+KloOPE
xLemrCKcujXuUMTIW/vI3zFJssNAbGouSHcDP5J+F8pRg0xYMglO9DuA0X1DVd0KUGskCXGT2DN7
qoYWdc7O7qkh/t4et9wUA+AH//5t/JWHWXIzKe25ZUzXeTts+UPGGGNpxzcz3cD7tcCTdF6u5OU0
wil8xYjUZG9lqjwd3l7KIV4sAhukGPhWePQGB7FRCIYRSr0S+Jo3/AU43U4Q216g11RyDke90d4y
fqdvrn52O4dHE2Nwv73/BVR9Yxpbp6VtwcmmF8Copug15ieW/LPOMXwDkpK7tWxWi+rXk8617G3i
WBo0kK9kf1o2F8Pk3Hv3CvdyRBm2G51AEXZNgfKqQS0Kk0XSur2DWGvyewo91XG3zGtEJHipvRRn
e8tV0+13c1o5q7O9euCaY4r+YvsPmPgwmxkUvD4eVYcGD8NFePb0M4m7ymbSzw2JA8YJMI0He0wl
MDC5bgXPNI7ALnUNZrarH8r3VcOpfCg214VT63cXATtZKB4jE48lB5FtHpLrBTA58dTV5lBLPqln
CzlXuFhL1QYnzh69Y52E06F6nEgVifCHuBMdf5+tccsr78UXdhrFiL0UqAxwGLuqJCBs+pJlbtpf
FpHWWNQ+X6hshMBsM+fuAr3Kklyqq6ZjTtJ2iQAmfXF/jQLyxgLvAQRze0P3b+AZanqDHqFPbyrM
8HlSiGQaKwSrT+lolIy8ZXF2VmzjuDlcf9PW1QTCnrWCv4A0yClzW/GbxAxbCzdajtE5MPXOcYMK
Jh+A0SwKYbc0FeDpXOrB/kF7kqfGEjyr5ZGGQrhn21rO4xlNN/WD6urz21TSFQeLgTLviXSISvF6
VXufRtAPUm54C+Y8KUEKklANgM9x37Po1eIkAvP1V5/pc1kdxKS/bapd5zJF8Ztp/Ak/CB0Wv255
6yZwIDmWQatM8/YuVdIH4/G7M4dx/yQCzuGqQEVjRIaCY6qex8R7l9b5tvzaxFk9Lwz/TrteUbO9
3EnBGXwuFwzKMh6p6fgmsy84Fj1DSWujv518x7zd3vp6W79D3DIAiBP3eeuueX5GzpnLlNZcO7gB
jz6TEkKeHpJ8G7hbvm4TDtQBxyX7yXyZiUnWKl8j4uuilHAETvcfE9uFqLCCEqh+5Q9+oHsjwKys
5L0jqtbiNem+fMm1hMgauj+P33JzK3uHY0fqszFlLbYTHvHOKdT/fZH9/FEyVChVcNHHHIQLk40Y
xfAmVCh+NIZjnScfDPcjlzrKAPH6Szsyf/roxFR+3SdHCLh6ov622TS2g3KfWiRQ312YKxzHloWN
7cmzyTjIurNY9HVJtJ7YJas/hjHKC0QoN5+l4vjYVXsz0tip8JW8pblcA7ThVnpYQG2ZF1wAt8+w
LgC1CM6x/DAJHkO3vnYGZEr9WefSyG8ElvqYp6VmahYD4axoY+SOow0LqmTczxKkqKuyJ9hhPk0p
g/nNzeyOx5XvS22UjBhHwEyMi17M/CWmwR5tMGBEhPJ0LRdLe3sUWT/LugUn8gaExL2B61JRTg74
uTZMqrNgFeSnppnRCqvAYXe90EmSeG87MXnWbtsgyfd63OWPZfTZF/SJJFpCVJKimHll2RFvrLke
JTOfmwo2Gk0pJQoKWIyI5RougpV3/R6vYVl4q3iWt4VdgwvUpo+GWCJLkhg8Q0qWOI6rp/Mdedlp
+uP7ZJgrtZUiN1fnybpdOCv5kULSHMATYRrDtsOqMTB5xv07FoAyW5awD3Q3WG5DQ42WUbWLxhYH
6qObp0IH8xtpZ4jUoSSbK1a9mfXJfE3QMcC5DuQUbIdLSDl6ngVD8IztuuOb6PKW01ysL2dOlcGs
tzZWS7WTqzYUQ1r11TQQQL/hFPsVmV1FQfrcLxi6Lm+VTTLkMGt/F7AloTeJ5EOXMPKvSQOn0VKf
91rOaJ9kfGc2CA3/+C+GNA/s8Jh2CedBCubtgS55LKBHehfbtnOlFng2H6hS4emjMyV/29i+pmXV
r/ni5VZJJN4/Olsn14kogVCBRUF+7/fydoGCvuZYEX2WDR9JrdlVkLqwGWmEHl6vVLjRUHjCKbjZ
YXNllRYDRd14Cts3/pOAppolX9Kgvee3fQ1AB9h4+LxKgNFw3tZpeDDtc/wQNCAcyzwxMChhTjSH
ZyJg4Idt9q259Yc2s/iQWQ78TPyqSRRd+Mtu13uJ6oFDyEiA532OaLBGGJdliEJPf4eukCpC7N/X
GGF7d2rK8uOgAZOfynIJzZIKFZnTnh418/qh7V0Rb07S2Xf8AGRNX1cT3NMTkckrGdWbe5yvSlA+
nlGwHJoYk9+rUSZ9RBBIFNLT96bOQauZzW+TT/Sq2JMdg/BwxFhCK0l0Yi9DmAtnsolmQup0o3bv
hBkaTnLtSF3d320b9neV6CDnQSlgRl8NE2lcLnnT1CgNUUW02lxhyGy+Nw8U4f+UpVcGUmndA503
MBcn1jRs2uMqBjh/P5AafbyfIr7IHvmrCyLW2axOrHq0eLHcPOXm4CD1YjEVXx80zGRdrmHGxMUY
qMmvA8Ouenk7w2A/x6Nmrf4KMohDXhZ5jNYyth4QiwHlAx0vst+/GpEFXbInd+JUC6teMG6Ucrsx
jLq62xe18GauvH+s0UpDBu/pssiBQwuZ1x2fnRN9Kyry3hpguzNQdZAzJi09ZZy3QeilAg2q1D9e
0SMpDUlRSK0nNe1T9T7iimZYcFei3O9vLDDZZkU/NSBRCI9sRzC8n6bF1HhG+zpKofY38xIDTChf
gHW4QmKtd3RSWP+FWDsFEV1Gl9PbuIClAn7qMFE5eR8NOTx3qkPkuPvgs+40ZYkCx6arW2NBnH3W
U+OCLebRZxxrOoWHP7OFAPy4vGkA+Gea/MOqd2olT7BQ/GD5t1aTK+yPj53y/0JZr1Tt9957xPus
vpJXmrKP3i7sQonQ4EMncxih+SqB+SMDHZUIp3gCKAwx7l69chrSHKkzmcNtA9NtGI5W/BFDKvVy
bn3EVaLwwjgiRfbGpT/wX9kTNn77nqBRtk+gwHIABwoClYi6QNI9NUnv+fze4pSOUJ3HH+DgAVwA
0GeyZAROOuyWj8b90b5PUMOjtjzT/BRWdrWqO0elwWR5Av7oilScWo6h0y97y4VgjtgeJKqoCEXq
yc8B3/a879quP8svA+gTSqd6+kT7ZVsSvZV9PDhzwo8bADiZ9UZNCHRT/jUEtFvymK/89cV1Qau2
De0EprqGKfecKTLoi2WFaSk0MvO9cS6ph13v0Ylcr9r7dslJxT3HTSRsl0oI9hjZ7NX6GIPJwxAD
gZv80ZOUun936HZUPzgu9qdQ0hDNc30sRuRTtPuQRMt9UPF4KzTDJv7u3FeaoKIf6H/FqPwnXden
T4WuavcgmLx60qumZucKR+5CvVppoMyAVpzhQc/GEOIVMeyNzBe8l1zVc8+SkD5AJf/kUqOaE7rU
5UYPkNxxfI1FRGbs/NUPfb94E1qm4mZfw760cz5GvS4OT6jOcrg5cmzPfMXn1lsjBNILRzUr9/Gf
jf5s9papeJHCRgraG12lJvekWNz0c62UxS6nwfcmYl83tQZ+t87Vnw/z9iop4+oRcueLgQ6j1ach
tN9sj5PwZG1oglU5CHzeEIaq4qMDuW+ksh7bvQhI25mjM6MRI3DjqjBp1fZeM+ju0DfS2Y0ih6OD
glXCs+9oTtsYjzemoPWuN38FHEAs1FHdLgNbxmmhnIWtx0YljLynD6VyzFrKbnyqI//EqhtMTGIj
GQTkdG38kZFUpFO/cwq0KqC3vS/CL22651gKSbm0J5HXS9FXDgPdyLPBI56a5DnfhEnVeNDXTiLo
PiXZBqyFsyDw9bfPoTOflt3kElEjE2Gw/SD+pUgyQEuQ2+QQZe97PqTfie23C3WtS076/3/yNq27
kTF9khePV0rlEV6OC3Yl7Ci77FdCxB2BRWRJzVAkuj31t0cXwHh011DJ8TOli8T19RAmKpWZI2Q+
tz2FUPJEPgaAcmX4Ruwbpo0wFufMmH7qR0O0C8oKrhWu3uMxaJ0400Ru0EveJceqsV/4aJ6WV9MU
Pg52ARCP+s0Np57byMVCAWGqUderjT/MMar9s9yTOn8BMflxBLqrnav9uMEY4pxmZSu1jq7cb1vG
lTV3E2uT6DyGV3Zh7u4j6Lj+2Lrn8nXWYgkoOssYc5vXbefPA8S3k7EH+p4W0Zh3RXblhDK0FD44
+yhpxPlY60a0qy1/fjc9DzrgRZSoynViDRiIMYm98Z0tTsexjZjZD4tuVYIj+NEva49iWF69CDIx
OSUBN1zcwwwUdnHvJmtt7G0tJFsU2JElh2ITxomzUSvA0lpgGPyoTH8EshCMlcw+AwYVBf/DC1fO
Xb41zadJqmBrPLDbbhGy43LIn+rlFjCZg2LUoLvnIyjsGeuF+nR4b+f6IKEwjGS0DJaK4llFuWta
qF+pBsvVyRRLhshFsaUqfT5xpnckZbo61xBEh9a4gW351RpDPS1XEDGeJJzkYnaCCCe5ZopP+7tp
1fxYE1363cTQxQKWgWwZjjZjjKwMd7cnjG8c7LzivC9CWYIlPPZb/Qwek0dxlgL3v/Wc1+dtghFy
wWPbEv74HeMrvayll7/q3djEDyDQXMyYTacln1TUW+g/OJNxd7/83+hsKXptT4sez/vMXeWwqASh
q5hw3k1nROp38iDSXoR6aU1MAhnfIkZ5LFBhD5h0J29mRcyWUv4HxRopKgomQwAfB13AcAG2L9E9
ceSKqz1Cx8kAFJwVV8nEasKyoabUZsHoZSMtFO5iigKERQTrgfx/Vj95RftlVm8YcsEU2+OkEHo+
qIowp2OaBV3QeQnS+wCQiGMavrZexL/JR0808CowzfVQVLFkiimEQ8OvAjC87Q0jIFztitEZjcB9
uNU6rQklpX1OpNoZYmzawQQOBBPXeu3m3w9p4lLWHu4LA/uyBXS759IR+GVeox4y3f/hkvjvZjUk
QDpGYXfko5g36lgNxSPbKG0Oy4SRUSLJV2+DcmvapjbTcxleCsJyfFIYFImp7dMPzd6Y87n4hUqf
/eI5mwv5+KmkDJYyWgRRDcNBhcLxH4Y+gFAlD9ys1w/kzReyP1tHPDgMHEQOfG6fRTsfnID8UOhx
YzgrYbl1nOgwKK6DrUHYIT0zwbpYWbcGITBUiBR2W16wwkWDtFPoB/p4lXmOqDtiPyEDsPtXiPzl
XX3lK1Rw0q9p2ZqdzIy40lZtVjUbXAtp31bj/GRzIsp+QjlvPTIINeXl97cETj6by6IW5y1CIoQI
P2Etkyv3/OjI1yuy7GkFbinexPZVaucvdOOmDZHI8EozE+8Sn+6fz/5U0uYlAPG+pIZymfWxgcIm
E5pxObhxxeL0JDvTaObnSN1XHu8CJVkSE55GtSmznHs0WPzRMDy9hl9OAHWY98SP88Un4a9zS1XU
w4dJCbN0jgsPcmblMpQTBm0eohNVByZQsnkoIKPF5WHXlARQctDamgxtFcedP/i2s6XMuBb6suVZ
sTWGKj+yIdmlzi7t47r3HP3jKTwhPxVXmLsNESwzn5WqFqAHeB8Prf717Rg+Ybs8yhCpM5AooO4e
01Gvx06/y9x4+/ejMzpRoXg9VkkF3Lo0K//ThutsHpKNJ6h2OarAxet4/ISjqUy0iDJPJ3VeraP9
oKfxaEi+Udt4+ckdEDGw5/sFv6Fu/JWXnuv/h5PV3YDLZQJcTdU1UeLQwOF8fy08h+MBGvvWQmXC
WLkBkF79/5bXtOxsOI6xmHUA9VM2K1AcAGFT/P+uaO5ZQbWm+hO0sU5S2IEbZjEuo7K9oOcgrwOP
h0XnH7GzD3RJ7BZ22aIlwBWhFd1A8DP0H72HzGLNcwemxge3bPcMZ5RPtfNuMDrFk7FcV9c9ptur
P0KSDjB+/RVneGDWQuMGrdhj4XqsjdGUtOuH6RLjwXOBgcxlf9TUS8fWgSpXFDJTrBG9rkm7lU7n
kmq5LpPBNifmmw7nbjOGjv0DhqjFPOf8irj4Zm45RV8OhTbmPXbyopTL+wprO6IThOj9uJDC0m5e
yoeSs1EQjGNLxr5JdZ7NMjI6CfDS7GWxIIxK2LafnEEjTDM2/iKE4owj0wEKxn7ifoPRvqxkuRYO
RHAX1FBg7UOkU9+8u6JHofeWSzgDnvThSMNtmZypPDdy7grZFZSXN5zK2Fvs4T9AWz92ef27QX9a
wi+5kJMbYpYdGC0TUqpMzsY6TpStjsdOKPlHBd6WaWgrcCr6cU4DrNZdTF/dP46GvBwY+IoWmqdq
k8nS8AYNkhBvSuqPladqJ+PLMXNrjv/4ZqLGTHiv29PurWuE2v4KexD6C4TZJsA7eqLuQSxdYKHq
jK6xvHPTnIu04u95uhtiWShfVAHEhKa5gbRDVMCj06/ETli2RwNM2naBcIvS66ok6WVFPJM19mUL
3BoVmpVsQlQkHcoZDN+kwptjY50ScGmNmby/KxI67/A7pxMa+Q1l/y7DePxUtA+RmyDroi4ArYEn
nhFM/OhjC203y4Z4An7w8gPaWNmrhmQWOjYQe6lOBUgYtv46XCtWAJYy9B6FxgN+teqIQLK+WX/g
CHInQL5cvT3YHux9JaQE2Hxy0cYzwqNpcJSYF0WQVm0CkNCUBuMnY1U6zPsKX0BY6j/GMUwIIBfq
Jk7lQYuTQRSo0ZlmxM/cfNF1Vr0A2iTAFaK5P0gxRO00k9Y8c974RPC24tCO8RQofPBgppbZugXo
RMdhsWx5JC2tU31zcq4dnLo+e2IqNMtvGk7kZgDF2yBDsa5dURj0zl1LI+lN1xyEMwYUiSVb7cvQ
iki+vtj7noH1fu/7x1BJSHEVsSTsNcg7Wz+HyOVRxsQZlDeRi4foLc8RME7P5tH2/OVKU9EUxBnq
OAzx4iDk8PnCMe2JBnO2JQGOXYkWM3L6xyvM8IpyocNxOUmerHC7uhlSrVjdG9XfHc8n0vtL0GwO
XMb4C5tw4FhIhXbDA8NoTcKGGPK9wvn5Gx97G1IAq/6TO+n9tjv7Y4bVBThJ+9EuAbvPwvmrQcO9
KXig95XjTVPdio3Xt8znjDJm6oGyJdkOFBm6X1/OTcL5QPz1/WPY/zf5eqjjg9+XRdGDom88Qgec
5psonUiWOFiwVZif9WFdovaDcCMVE5lRN3CXdJmeBrSZe0YWgTZeuMPU0/TKWu+iLSor0ALm5KXK
rfgtbcz0wEObhxhr4gOt9hr/I4A9OvsebTsceHQBMmrQHroKPz2EjxathKwg3aP1RqHbXyYubeED
T+62FkuX7wc0tugKNAymlY13SnjQ7SgV7S5MRF+pouuwHh6aKT5ZDKGfs4wqfelMsFg6vRT92f7M
rQ4N6A8lnQnom6SXmkYEhrjK1WRBVoF63XGjwBL6wwYv9sRdKiKhttNS66ommts4Zb/2E0+1uQVY
6lvIK745duqNo3zHhwVbecUgNaNqW5PlKQ619Vp8JowfQbTMeDVQu32ewSQrjQtQVseoq79h7IKt
mPOj39lIZrrcFA2+obfEv0FD+CVQJSIuCw3S0Vo/cqh1w+nuCMT38qFyJtjJ0U0HF9MCuYBwbt1Q
ALo2fkb79pa5uMCzh+xmrvDqIub8a9XHG2/xaN5vHRrCczsx5z/cjne90udQzSKn0Q27f/5X/dGP
Q+u0s7wAKpr+lF+31YIFoGllUyOoEPIFNiyhzw7GbYY+H/YhNwgOjaiEiB4gdRgxMKdp6q+GgYLx
23ZS3/u71fJcuTukmtri+7TtDkjB92BbBYiEi1ozWphfZ8/ynAqlM59fEjpj59nvEg5LXQk/zGxB
TgcAFnHJMlH9KI4Y8dwkVoHqtHp/xSeJMGyfDGpapxXSnF/Xlf4Y3uR/8V6MRWqApAMZJqNWbtsv
9c7hSBw+nYsVN/RhTNswLGGzKWD0zWgG/MBu2cbBRphWfYTvLs0X94ZjSMq54VOHd+5+RCaAwdsr
lSHCXISa0Pa4jXlHgvFl7TBUhXJXsDr2KmI2xXdYJcbPvuNIUhkAl4/L1n6D6+f+9LMI7Wp9GlGI
XjtXjGlzpc1DAuoijnST+ASp6kDmqhm2dFyCITJ6wkHTimmSzaClYUMJADGKm05/0MQxvvfVaQLH
T/g7FsTlaeCNy0uSBq6qDGb92UJD/ZJ/dMwowr0KkjX9uhAKz4XM+7kESi81SyIGCmJCYh8gZVAc
MHKHeXwuXeiMoKS6qEor/uK2LjBv42R7NjJh/h0tvXJmj77UkqaLdrx2MVsXgaOa5YXelaKpECb3
mFmBxKi4DH9sl8Ohnk4KZFo+Tv/D0mMkFKFkcXvsFmoC5p1QQcWn9YCpNm27uhxyemoexkI6X9QW
3407JtFTzRAYJB1sbjxL+Sh+pIY94MpGdmYKd2qbHSmjij5nDXKT6PcI1orBLZ6SLw83MzLf9xTL
AxTe6TUQgcrqfoIP4TAGQVyePfkRIHPngb4z/Rw2nHS2PdPfrwzjL0gR+kEZPLST/CbGG4/iAfdj
Ob6llWlFAEA+4UuHxPoYs9fdwdAZnM3PBPk77EQy/1v4nqgSX53/ULGKbo3rF36NxCU25OrP4DS5
JgmUrTx4KhQUZyX95MPenDWONSRMWQDDDOf8Azv2ZVn6ZlEHLdWvHWqJWACxJQ2FblOmBvuQB/+w
F4CyzHw6qD12Px4hMF6e+v+bOWA/kkEVVjxiN5uN+kUKKvCACAna8F7eLafaYpyC3g+4Cx9pqH2x
FPRKq0xELqLs2WS7evg/+Jy3ejtafwTxFQkq2gKTM6W+GasP+cE7A5tjlMW1meETops/tzNAyHqP
PKKetA6eysg4FhsfqIzh6FgJnkeAUGjoyI2eFfTD25MyJF/YbJ9ZDDNF9TCQXXJI0HfjO6wajR9s
rSgUp3vF34UxFc9yduU6igySHyeSC3Cq0SPLBukyIxoOoS9axiX1ngWEy4Y1niA4F8VLfdzDASPj
TM8KDDfS6jszs4WZp5nJMPK2F9S+VKFvaYpjJk1IaAqiU+BfyGiVZ+AM1ik/iq5h/mGnxNHX370o
8xg8R1i27YSESmZPOjhPaHo3QN6kxBJCO/ljdEPc+flH58O/n6LD8RosR40ZNWeqFLoubsw+EN2C
yiSMgurDSMqDEgcEDKDV9PBkinDv7zPXI8dtpiDoAV/Ugd6HohEGOhB3QAbjR4JTLs2W/kCtHUOb
ousm9nUG8a6/FOXwlUQMMbKKXuw+h1bDM0zSHNXQasysFoiAQZDvz/1YQuowLs1Ci4dtwjrgyaLY
kl/TmG1OteJ0SSvvPer8v+oCb2dgk0RC4R7+3OcH1Ar3tgnheu/C6IVnQipfqR/4afpPafGzcoW/
yNB3WG4nBTg3TcHaC1fpnEOdh9qBKON/+kf+F+f/Pz9CE+yFd+IifR3goQZNy1uZezFb5i6Lhk+N
Akjh7QKFE4qmjkYdeN99OKzsBdh7wNF/4LTXWCuCFKinjDZTRiQG85SPgsbYeqS+szRZ4hBVSj3P
5OGCgX05lra/oNqgw4yRJpCLUgtyh9S/j+UvbnRREtE4HDl9zTtzbgen65Oae4Koi4hJdgrMvWR9
peQljwtqh/j0OzK6TLlHyK5UsrpJ35LdChpAsresQCqkb/O7y7A3u5RiyLMB+/b/Luq+MXsvzQow
189RnjWgOrmoRMr1vSYhBpEoATZ4P7VTl1YyN1SQ7XVVW8c4lpwxo+nOKVqEAF/Sd839H3/73Nc4
G3gVOgh6yKWVIG5uY8+PbpBANgCmuvYIMlqKjQR5kNGTBuHVCc4zR1yqnelBGeJv/+gxQfcZMH4B
wSj6lB6yVnXV8T5AbeK2f/3qiEgnexAv9CP1ao4Z7WhAQvzoPT/iJrvQw8iJ4OXfQazt2UAo6K3e
iLWnjiWwQSY/hXN0Vzx/hCt02N4AXUKq/JTOHpu0ONxpWkiSIoloWQlwkqqzMTQXnlFItBd/dkYc
Zb9YDDxh3Mem4N0mX3lNl1pjHY6RvzYm4ugHZn0ygAHmTybaR19vIjfMPN5RbZR6VwKIMAIDUSgx
1VIOOQqNNUhCA8P3PMBtJpze4k3TrcSsuknEOlnBZNiv88p7KILAUgfUjrgb52thIKpHrVRVTFtk
RYgexKvZasMRV/pV1qbPm52txVDwyBcWpI4N4oylRlUw72nqPxs93WKViWN+7EuwplsfgcCQmhUx
KM2/JrcixZRziYCztcvwGwqzfqz7FV8tb4XQa02pzUjLwFj3KNV0fEaWs2WLbuYowdO2dn9aiccl
nRU8137xSELXcrJN/2a8xd7W/gpvNdC/y1f1VM3fWTgFBpfCAfJhsAwl+I5jayFNwE/jmGq/wuEJ
YgwMPsLGZtSenxKMkcIBXTkHhbBMpdu5BYEZP1FCAGkB0fMaiQ4PBf73FsSkembd9iqpff4Nlc/O
/y0mVOWZtGl4IcB4PRYW92leEXOyyeGCo44DLMeozaUXHTg2TEVU6xvTBd2sKj+GzqEx5tjETo8v
z+Nc8EEffKDCWzSg9x5MyOTlWaM7EZFleW2cUVb19OV2StninpN69pd7kGVqMdZK32tyXLRwQ8Ls
DO5ZBVC8UMvxmQgoWIl9V+QWNaxxnSk9PTRYQCSr7JkTsHLO1riw7L0OZnqooCg4SpEly9ai0rBt
lR05MQKUtE3ME9+HalnRCC3Fm2raCOBOjA5RTDqQc3jT62hnFyXGlIGVS8w7Z+D02MjKsRk6bekT
QF5rhD07oMH/LKWi+JQ7PWPEGuXF7iJw1ORwNc2HCHxFGluld7YUYhd6PesEZvmtI5IU9D0KBu0H
SF446OBeiYjb2DtjEKT4blWn+f1FeLmdDQCq5cIX7MPrE1AhrCb2ppHB23xz7Bj4bEKEhudSyZQZ
jegn3uTrvptbEI7c0kRTRMXF8QQsXmafvIpKY41LhYTpd5yGlCribPEPFUk68xP0Ll1U/XTRJ0dZ
frSD8afIR0fRiTezAnU9faqyqQxN4zO/sHcv3VKe15N+IjujgBgfO9uNNLOK9PQNVNA/a7QX41mD
njn99RqJY9oF5lhLEndA33ICNkGeHdVdoWGt8xzH86HGJo+JIN1Gs8tgvu2oV+jR8EfLD3C3dofs
8QdV1tooJaS/QGT3InDuVFB4uZwK2jXSVB5Eop62vVFLKUSPNHOBJrl6CB0z1RovXzE/Ee2xp7Dq
tnbV4BkHw20MaUw+oewn9Ln1+B6lQEh+fasxj2zVdmMdDfNkKfyF8KU1z/v171Hb87CxVz8f/9IR
ev2WK83QUmTs1KSYets4r3PQMZb3trsoNoD+GVa6I9NNDSRJ0MvreBHBIARDY0z6zV5XjoKYsedz
X5clWoS6qme8TJ3QU1v4TFeXNSUcEDfCtJoDAgF1iGuRlh5vnHPhjjsfeXJGRfvt/hmJqzJAxdr6
k7alG1mtoeuPkl8RJ7MbHNUlzH0Upu59HvwDsV8xSv4syO82v86zEx7S6KnMGGNBWDugVg+3nwYe
uFVGfEz7LXoCLKbnKZY3lFAUMVFaXPvdagYCyWBicsrEFgdYd8MpFmuSn6aehbJiCvrDPyqe8osi
OqM1TwsPw2umtDI1ZtmgECiSAwWcaGVY/UhX6vuSN6ufCh45hAD3mWiav2nxPseWQPsREo2hCS0u
gaOoE6UxlSQQLkDjI22Oemwq7D8cl27DEVPVsY2prsgS4e2sDacFdD7nurZ44VYi66rme1Joxuqq
Phq3CDPrpiPPqhAElx0PTSoHjB7V+8OU2EMRpW0ZRRYdwWgA7Y9xxDcCWrIQKh2Czzl9s4vKwyHU
JCnG8CWVDgN5CG+jzpsx9Rh+VsxMebUiS3repa6+m4l9ZtW76vvBlLpccRSNnYVuQ22jHxRJrJlE
FuWPCInXQnmFy4ZSXp3FYyKamx+TdcWgbRKDXJIYfgXQ+XyQioKSeSdD5SoGgeAW4B9qfGNmL+zd
irDKAY/tOEqdDEqZyNcHAopUl0U4UoSljpV7V9igZz9tymg8+7+uzUg/Y/vN4tUniTjqCPgDjxpj
5xtl7YqkImGOUcV8rTarl0ZjM6nWWaMndA8o9hb+18oPgE4xrAHg//K4Vr89TRn4D87KEwiY7GQc
mnm+Egm2PPJEFXXX5aWg3RCVfUTaWe92vP4kumjkNLKEPQIHOG2Fxi676txnRIHvEXtfkrM0kc9x
JWUbxdBUKMXJN9JSSJwFgFZcOLgsI+WOIg1mE3TeLzDvXBhy0FcTZOwZ1rM/ZoEP6FMuoi29Icmu
BbqF9OBK9lYuU54H+ZIiy5sVKMogPi4WyQykFMwN91j7HWKjmCtWS5mQ1bJDvaPXs6OmfAk+kHBk
WZ+BXmx8Bv3x7NJ/bnWlZTRNGv06oLhdVpH61XUVi5sspd7YCw+/UZBdZVV53BslvPKfMC2DPiFw
MKA4aK0XLj1dIwWS+zlQh2nA9wfNeQDgPWpI85jjMeXEgaHiTBBoG0QTLhhcxnSoDiChMNy6+MGj
O5IrK+ckOrca/sG5sZsQF34YYVkKUqKTVjZZtZk9IkeWt96JI3sfIfiqqq8oNHNavOR0/7Rni4Yw
l5vvOldhMSUgQL4qdqyjcz6jEIjkYrNAhTA0MrXVX3iMIdRaJLRERcPyuzoZzVa5n1l0PNuSGd1a
/gJ4jIKzfkcB9CXGlS8uHMd96UKLvagV6rYczUq4DoXxOPZU+W+0lj6W3gBLkRCifEENzkR4FEWf
x9TdQe2/friAPL/kDnCr7cW9h6VjpTalYPEpnLKGCtChSFbz6nYq8j+MZcxkQ+k3OhoibKDkbB6h
mohGg7ZeULwphh8O9nUlgTfP4uTRaX+/XFUdPNAmeIqiwduC9VaCmMB63hToe9Yo4bT8ErBF5VnW
LKXpH6I0RyKXUTlFV4Dt1nlvoQQjztTk8afmoP4vsdJcV0g3Tth8dtC+alRryy+JbMWcYHehNVaw
XeObeczzcOLA1F2F0DPAtBNykCoLgOo2bA9gWx81pgbz7BlZur95ZtieIBgfQE9aimxLq9k0btd6
xiyenXYpB77n5OxMOmbFYtX/iQS+G9Ii3WOSjHLp6O49+ObdHPE2vXdluskAE8+3XZdZtJ9lRYmU
k6MOzhtIB4+wwMjSSyaTLQtMfq86zYcSaWjv7vhgKvtqkDlhIDHP+QfZNoC5VzILtomcKXs+5igb
E6ORvXoApUAQvuaIv6w7khAh1qbcZE6NczHqOtjrfWTurb0LaVamcDCl/nHD2tMa81F/htz7QslZ
G5ftNE2GhNQ93cyH0yDSwdtiy7lr2rslFozXBpaK7v3xUg/n0Ha6TWuKJ/opD6lrSe5JfEvJG6BZ
J5J58qvmjzpTMaUyA8E3hBNGH5hTeSB70Ytk7QJJN9Ws6POJJHa613Ht1MIBJ/1wNdKZtGfelDYV
E7RGLEvvh3iZp3zZwc05BnK/g7njVN/4AXTZp3rKldOMsXAcTy/DvoA6EnLD2Iv+7651O0wmX+OI
fDrAIK6TjOTpCBOEtwM4BcmXsvBN6cWr8AfDF0Cesimi9QFNzUb2pKwKDjNpQMV+EfKNbvRzai98
fYsND9yEN1yG0LpMNR/Agq1Tz5LorX3pBpZlVw1qdWQtnOFHwNmg+0UYY9oQQ8QyiQp+IvQ2BONw
DeMO6/kxWR8j2tPA+2QPKY3i865oAbxRBwYDFpDkFyMJBE9yZlRHIl6RuuE4WgIgMs1XQeP7C6I7
LbrAgzokT0iCQfCPo3zuA9aSkRemVNxldPFvhj+Bs/P2WfCgG/kSxxikbxNwH47+D9Q+BA2xtfXs
kL9PByZwRC+VE5wJpyxvmY6v3qI+5KHFZDP+GIiGfi0ChKY20e706KswzNLwAQXZtsSospJMi9Jk
gMIghSe8wlXefd/EOakukKdv/U22PeUU2qmpWwkkLIgWz53s4m5VM2G8olBu65tmZbRh94WCwvGL
/iA6Ndq7VuvGdFRcs8z90OtVj3WvRQC87QpKSYmhtE0rxdrEcurgbV5qZ/1GgbfZ4W17Z/V3Mpeu
UtzPjqgHt3AunNtXLCNw+ixWvJO8vB62Dd/1Ub6b0P1vwc87eMOdaO+IoMQ4b+iyKphWb7JwsaZT
vf+eK9FT9+ZnBlx61jtpvk4ni677gM3Zajvv1GfuFVWz7xm8YlgJEXVNqm6zYgSRQ6S4mjnaPiAt
FI4VzhxlHcLk8vwI6b0bR7rvL+6CaIyq8o5Cy/AZS8Mcvsm4NQezwpfkCu/U0NBVohI0c9yGJ/P7
HpYwrNWRKeXGighxjjoXrPkox4F10RbbdmBV+J8jVj/+1TghuhHNDZXbvV17ow0rAS5mJX2aZiIW
dUqSCNiPj29+NStSTpWRv+2m16gvdmckFeCrP6nIXjv2KKZ2vEREWHshDtaWn6+B8Ug6rvmj7pR4
QLj9hAdhTIE9g4L9BwkcepJHXB94QEg3GI/rYKvwIv4Iz5hdEowqzVEuzCs8fjtFaUIyzMVoIpL2
TwWgeEGzCmi+OTWRwDDMrqkyl+X3w8lee5RqiSje3k9JtU0DZh9ktIXqynCrQsHoGYDPY8lq9G9C
77uM7KYSZHh2rPXlD/Oj4RktPr9LJmZkNFoyrxqlRmNtniA9fazwRLjUS+PqYMP1mRO/e3G9oUHF
cAnXG+CLD/rgDa3CEhrfG4PLVwtekfIxab9cphnimkwiiF2m4dYcvVqgpI4zERQgvXHs7TikzePh
H7kAQXbklovUtHsCmaZYgMk1SH0hBOzXXOxRbXRnMoEdsY5pYtpsZY9Hqb2p6lP6zjIGQZzYzDqe
qEzdfAjKxNrhbGoc6D90fHZP3l5iYYd1R8q6j/MbuPnrk+tmrejgKoGE67OUMfQMHspVv4tvxjjx
BcgDYNdwkO/tDUHgzzhm4vBLDPdhx635kSGsyfO5FSj/ZCHl/G45x0h6T8cLNdAvMoejMM96IjPP
wWVTeYnwDM18EJfUfoPn9P4IqtJow2tNzokcC6vrdS0hlmfU2ta91TlfkYezhiT17LJ/U96AZZSX
lV5L5/jamtCk4hnS6n0Xm8uEQhqTjqz+K8q/5lDcWGCTcf+va8y6IV036sYecTRQZm71c4lEUtfK
v7vcz8shUwss4KI0EqW1EPKJcdAuWSB88Ui88iNNwgoB0XucD2B3UiTgX9RYj5wrLSb8k2X+/IUe
CWJathqgSklEY+hWwF7gI0YpWaSbYEHfmy1zA34KEhJ5tSjojuSLnEGWtOzlRysu+NTaM4tKfrWz
jvZs4xlHGcd9fsh4Mt0LL7PTJukAIv/h14icWlIVbtPcoiRAp+rdYyTdQKiOMlPhGmdts0Fs5aEP
gynwl2v5s+w8vy25+aATIjYU8H0TBmvB9C667Q0BQntedpItn42o6vcvO5aE8yqBRSuJYI7v0w43
P/F/j7bAm/hijwGIFVd1RnL3OyiV6NYb+TGADeR/Ro1DL850khzskbs3Ik0+dxuiFdeosWcpqYCK
CCA9C5PSrTCqfxJHB9Hsm/UTBOeZuf6bOkGfJuylaWHh/eLwtNE2CJmMKE12yoHsBGr1FXBpcBgl
VQB9eHcSM5zlBqh2KSIO8vG3dsR71QEzEWTXM7dswSwswBuIYTPtALs9OKLthaqr6bJVmIvZnng9
GOF1l1CWZmV896O9XVYZvWBFvdjZYBoq2Nz4HMdhwbPGmMPG+vy0/Y85vgcPKxf0+mlwadPWfk4j
i4TDSSMfHtRdERIBVUIVkocRqaVNt4Up6hJ0EEaEqSSCFkhyyJTN86LMDcLKBTXDskgGbGK/rt5e
uGo/VlWHChYzfnqth5uHl3UanLnINNsZLZCZmj2kAIOokf8F3IcOywys29uxjENZsstqKu96LiKR
7Ybi8WAY9cKUSFAf5nZrGBBj1mu4whAVAT9Xa9axYWFudjJEYTH1Zdmy8fSQiRLAWWpMOTpKJVqg
ky/qNZS2EAHg9ZpFlzM3n/r6qW+k10Oe84PLGb2elR99LQZaowUTAB2M04RVIG/OPvV+IJxIyEON
SaJDryo8lHpykCAkRhlPQzWOwlSfOpcDot0DBeyhjCd7y142hfCMYF2ktiehvntFSf75wdbjbO6U
zlYp4SSjFz+d90RFcSDq0tZFZLKekpl0XoOLerfAPNhtYq4tx3rFSJf5wLuSGHJ/QX/dQLd34kaT
hcnge6Yzjg4TeH46B4NoLBnUEU6jFgHKH9echS37hLolPudj2s9HIDKI+lHSQvOGMdTecqjtL3DW
IAZKsUge2T+K6zzn+47KCuyHdbXJSfSzf1/8ymi6yiegTZpoPxtlyrUzT+Ry3KpJPX1UQ06tOcnu
nivyqjBvWJq4fL8nt66HwKyJ37Gq62N3p9OHnsqMLWT/wljtJ67J3bdQh3jof9B6X47ZM9zJ1kD7
wBbwPWn2x6XUdq4V7xppjfZPRGpPxaQpUusy1IUmsTNe7kD8h+bBkLLoXQTbBFUKzlzNBwlKYJUf
Wg6izfkJxIcS5WwmAQjLI96Wo+/dgdbdH9l5Ts1De2/bztCg9sqcQRWUgrQN2yAq2wDeWB613RCI
qy4424zDZMo5W5I4PKT34lHuM4ov4vxN4VVg/O2CB5QBzb1rJ90j0oK9b/vhWf6QUjR0Dgbywolq
dtb1ziJtB4a16IzubyYy7xLxGFzukvjUqlc11XBF0/oxTbcyoK9jby1TXw12BLbb9j8WaQjBq7SZ
cD8JHPPJZGumidVt03VOxuN4cvRpl7R+6rueQ/CkajT4sQPb+5CqP3/Tb83JDDrrl07yWErh++Q9
+pLxic/mmRP60a+VxUvHT2MYiGJnC4HF2NKlxy4Kisf6LHFMlc1V/QIOdjwjlVcwn11ELE83sxgA
La0T8pRMN/44Pvpi6BDoXUHont4WN7vwtMF1iBx8p89gZgmx/OCh5RNw6l1/IY2eYAA0PrYm1QSr
KgjWlm0Ugz/3UyANPZlt/L4ZyfbDWwOaZu+c5akY7spbdt3OqY2s8Xy8pm9lCVNYhni5QRIwW2Ot
2gXFVtxt4S1mkFeYG0AER8PeXh79YPYS0UOdPiAmu4YAi0C7N6KPJhZn1oD4RBmIm0ck0yJbJBXh
3p8vaG7zO2D1KVsH4z4T7U/6mFCUMi3r0Z5akBsU8YZjF8CuyDIgWo2ykgFSls/UnfmCgFg8RQay
Va9xhv0HH8mWKvikJA8xYAKxym1VzsV4qTIkoGmT7Z7piwMJMA7tLnSGQvMMVzZQA0tqrBScSIUD
rp/DAEuQPDZWtBhcuhDVJTSImaEoDsdpTIYO+8Wy7Migj7L6HmaRPlcTZL8oESuXjZr56cfMR7GZ
UQSUWAfGpYMtm8Zla1KdywmRAnu1nfokBRa6oHBnZG8X/p4TNa7F/12hEb16q16kqHCbKebbLPr5
21ZB30pdv691XOg2+BJ8lU2Iz5b44VGZBsdr0DO4d5LxvvRWfZlPsRZRSmI7NXptwmZzC/9dvG04
r6b5eeO+dAH+LqAUkV0BzoEXlHgmF4bXVzDTWf9vyrjJorXLo40KObW6WM5QiXIj5EXaNtkwu2cS
VFbhImI/npTMkrqlV8FM+VQe6Htht19044Kgy5MFzGFqvx3xd4+n9S/HqXqel0RmQYkVFBH/FjNL
KmkqXcvW3r6LPMs8HBrrXP/5MXVRgHrGPRw60dboXmbdVXD44hrmLjEh6dNhVwdNgrnCuFeatcXF
QmQtA68LIcxuyxRGS23mK868hCg2kOfucmT1Jp6kZgGjJA/LTuEenAN5bL2Zm51ZKqoXIjHH1kC3
ZLIm/m4pQlgjBiEpW5BEAnzqXWbC05GKf+Quq3N8QVYzz36ppS5srVQoFxeS65RytLxFecAa14yV
YWyKrMjAooPBkXrxmC+u0WROyOU3AOGUaD5xAe65ojYYWyk2S3ntNT14qKStVMpneKGp06WF0Bo8
yoXk5zYVZMQz/z9Awzo7wwIxkqP28Oxm6A4Wq78s5fzTYvr0FsaE4yUCZCY431q8jpBIEsFBDsiW
WzJ8LukUkP1tGQlNHJbRFJ8EeTHOT09JPDZnp17OrVeNW86P+snZBViXeTaRNovn9Qkfiac/kiHm
aHMvzMoLa5LlT87NTnkzXgWls47hSOaEr2t4LAGAZ5SjAbfyLp6p4ExNX8s94X6SeraIdoLyKzey
Adxf7bBqjtdBJQtHRCp8rN3yUxvu+YkQ9EqykdlOjfxnme/4xKiw3/vPdxI9rSZ/ZEYSulnE6Yj9
PCtnOnZlgqxYPoMrET355cOEfJ1cR08Bwc35iq4guwlJOmTvKlLRKj6kohSc/V4qUQrMkg06alwI
dTaZISaKn2RYzaptQcEsuyQU6SZEF9SAwlir9pxBDwTRzpH3OHeDQAgXyASqjfNmPKnJoatruJhU
ETB9NC0qEadaELBDfceM6jlat8jfpXZQsVRHj9X8Xyf7J73L/ARR8tGU9ZLQ9mBrys7DhiQCVCsM
tBmKVzM2OlBHT6bZU3scWJrDTWHrpsT6yTYTDMjQIrf1pEwgPGolC4ZiddyF83z3yrb9aCdTOfs1
8uRFn3lwPpuLF2XPprxqGuT2MxJW+uTTkIHViSaXnBFloBF7w3pB9ab+YfphYXh6weFNNQK7qtdH
O2z9u/xk08HDEdR5Gvzwx5LUYQp+Um98z8OoBnsoz6Hg/dRziRZO/r6zyzUu2V3YqhYORx0VOhJw
yYT9UZm0omQPjb8Ehpj6uzkZ8UR/PH3w8mXr1b4EUUvEXO09CceJ9e6sRwn6ZqWcnPxtJrdDfR/i
TrfNuJQEssLbRTQ00R/g4ykfx58rBnQxSgzYsG4gIDKBJbD2/Swb3te4/umqMrYHdcgs0Ma282As
XDgTGa4SN+ZMFglA/CCygJFUeiZoyRhut8xw2H2oaGu20ZNmbReAwoswCRC2zr4JFQ9S92kpz39b
ik6Y+Bmbv69SE+rv9+Gq+NznP5kzEJOEGyq7/6BeiEwNigvm0H1F9/pHoWHV/OgEGVrqogvyW/KV
httQ1M9SAvaULyXQWzTc+dHE41VqhxHKKU8s9BoYGUxC6lZv3H+eKrYPqhC7LzuWnj9ixOspMxRf
0rAhDFxU9Sqiy7fDwzjd+upyQfeiGb4VbBJyP/4m4QAkCmy2FRxoDONE9eClYAcsAI8zR+GkrnVc
euuZ+tuLGQJamHQj1M9wR6aRFynHzFKAuyqI1aXxfvPzTq1NOF6qflxsc3/KUHN0h8bFepZrKmeH
O5Wx4EUQKKIhrxgWtefIn6asQeKv8Gptqy2jxMF+uXK0m3N3IyMX5uDxRTLtnTyxseNpF4Y3H82o
2vTd5Lrpp1x7rpp2pdct+KzcLBSYEwhoFy4cNZzwdzz34uJWykOrvXzryK6wL28JaklEau+RiWyR
8m04k3GGOlWlYkCSY5m4dmohu0Ig4y/tCQWQ5cQ4pmUN1J0zsOZUdIF7sDMsv1o69il+J7w3+h3y
TnEMVVFDaRNEiMgQqe+HIR/v591OrrH1M4kDLs/T/OlwkkTFhjC1maC3RIQgVs+vjmr2uAEageII
jc++H5fBryC2zbJx9VDBr80cVnBslKFdkcCgOPjjflGUkyaUsiqigrOdEW564cVNgJV9AopSsR79
eTrMsKh+qVJxLM3fM9086RXZkNZirVHfANYdJFC/TRawaqfhUbBb0By63F7ylXmHZvsX2LwIVQPk
cGHoFLQFCCwkGGcaL6+9yoFjMmce8wIov1kz46g6By3IMCJ5xPZbacf05P4HMt3IR0CM7gOVCoYp
WoPCx/KUNscjI6VodDlziQGDVcenLT5kXH78DSgorxAYEJY+Ucd/bfLea+bTa7t4PgmRTjBZ0KCI
Ud+b7vKSxZW+i+plGHiq4BSDK8s8d6NZCHtjLkqEQH8DQJb6zUGPbZTbFTNZm5uzzJCgtveI0Oay
YZEt7Gg/Pv0m+asMkX0kWwSLzpK5zOnkkkOCPQMDky5NyCJxZAgLgA1zdvH4ZERMLmlWTFVJs/yj
L/smNWeckqQqdgqqP6tDFrz9cMVNmgLDuyHO0N1RYrVr8gZ8vy/Q2w3u6cfSCGVrMR8ziYdpPBUu
6hiWg6qljIoKA44rdGkLnh4AIHMXYy3SiuetjuvtIIAJJs22Bpwl4BXSz10ruYyDkVBWQ77nVEhK
m2mZkREHgAg7zvTILFxE4YesXXnY0cja0AWdHdXOF3gu1nubYJhKX438RM4cA3yDbWG17/r5BT6N
vOIDBzyHL5QOafkyRbLoi0QZdiriK7YjA+A+rziPQ3h1eFuw4uuhTPcE7eb6CIbUj4Z/LQYUqQZo
fBpMTSoSlUWaW23FZxdtnYP3JHkyvovCC2JoIaF7Fxy4ASqlDCM3jI6W/FpIm4ci7ZQMKNnZIicg
947mWOLL/+UbeZvGGs2gwew8J9Ko5xKGFLfdN5TI7dhgNEMU7PEioeNKXVIiKrxnhvlQusy3+07n
7YXSe58/FQNSJk0OUF5SBSmpnqocmwKXR6hcaUmD4gc0mWDmrIg2QQ0qu3cE34O720AhxjGU9vql
rREe24Dfb1xQG59eLEYBBx1A8nyhfPr8jXA2gYC4cNT8U5i5Athua9Z80J8xNZlhhdTbjPZPWX8w
DBnXj5/7ONagIFBIw45zyWC7XZJW0WCYgeEObrdho0jZEYcNsvyBTPiCHyDyu//YFl/+mZ6aewWw
T7Zbx8IZaKZYDbNv1ORPmuD66JJHVOexALTwQIbDOl2zbFgK3GfkiAEDLnsbwU6z78murlAQnR4M
vB8Xve2opndIjwSAFWWTQMyqu1iOXDHXDwRnLZUU30UsLV8TsHlAJACaHj2fTazqf0K3J99iNm/k
arOC7x4ECX6ezzqHU7MY/Bp6sbVOvj1/2GtAC9iQm8wOC7IbReCOvqcVBrJbsjVuBE985WU1XJdS
fLwRjp+c/ERuhlW4Ou0EhU08IW92bXZ+DvQxTmqwmCuub9jmpyXu/QQWfJQvtYib9BdSS+lj9G64
JV57qRNcD1sN05hE5ZmUtF9amlLqkIR2N7uYXivhkrH+4uZxvnSWNZrz5YTaPccnaBvoXtxh5T5T
NP5QRwV9mgKqlIw03kCZ5SNcb4R0R+4Z0r98YFb5li2gAxeI1/WkP7J1SXCifT1zMTDMzsf4M9aX
BGkwq09NJ4nY+fKOEssmaa3KquaEJtcEjmhJwigpDhXsNycOomtvZzufW0WIcX6ZPgp2wxXqXX09
o7WXQbag0sgkKMCWQ1Ey7WyFkzSvNf7X+sNzbKwmhi5ZtsP72fnjcMURWAmlL1wpe1QnAp6xmHCy
ETMuK6l4tuENunDu4xqpUHLEp8hYNLQ8+nca1x0yen5YyOnDTOctWHaUsUQOhTAwzwsdDuoZNEJj
tGg4roZ1/AOHLTx5Bm68ns+xSYSyddCZ87U+d0NkuLCg9Dhd/L/NotJpSt9jKDnQZZeizYEFeOWD
Rhe16xuG61L0Y/s2y2Gnby6JvcWKkHU/14Dh8K337Jb5+r+jxxlhgfwBymFwuNDdwuc5nBqlf0Lf
RMuuooqIQG20MXs3D5BevQ73YPcY60XMtVyr+wMVgjtjOzFsYMJYh0SeXwKBnLtclM21aIk+9E0J
+YRk/aYspu31awZ2OlBXPrnUwQlSlsAhLtNsX4zfJwmmkc+rr5YDesFoH7PKIffGjXtd4EyLzfnZ
OxJ0fL0cj1vtL3NqiUmF+S/i4mg3K7UJPVFuYcD9HCrtl3+T9foGcNXie+HlNfTjGcjJc+aze5e2
ScOaT9JoL3vvGQn3K7ljVK56M45zAh4UUbZ9TgdxMsCvK4jRmeVjzijC6kpUwF7GbnVxsPSqDTZP
vxkrUSeZSLQi0H9SX/l5Qgb5jI5VRRetvLwK60Z4htae1lsMrOQUFqhNYXKvUYZBsnq4TZFptA83
hCW37R9nF9y7hEhPCTT7aqQuGA9A6rOo8zosdVnQ2obKvsNF+g5Q+cOF28Qpsmconbf4DNya/yJO
TYrSxsNuiiLAucsZLYvOrd3ogFlpi540WSEmkiS0qF9qAgco2EfA9e5w4Kr2jznJRPphBwGkvNU7
htmIFcIhIDZ4/9a4xN/lMhpzm69d2nhnnWQMHiZ601U5Ryg5aQGYhKE7qqZlS4Vm8E+eGke6fq8T
IrPFfHvFSAIFsCF5zF0w9PdUYL3bbVdvvsj76wdl0KTD7oRaLjfDKZ6A1OjTDt3wIkrMOaZJgvR6
MS2mTpc2iInSNVJxwWzXBxrpZnBhxo8JpzG3BlAt0SaABEKmncw+jfRTEybkCX/CIBYgrRjv09L9
lAeR/Deg8x33KIinKR6G/HTV2YKBgB6m1uocwwVDAa0SnGfJkiyhSkKFQKxdYe302ApMaEBZDm2j
C1EL2jBvgbydZXJPAOl+DaQdAnWeQ9y56N4ncbqanwiPQMkgD2/3Pb5JQbiTLFuN39b50mE/pfRl
7/S+4hppV+mFICspmLBEThjdRzqV/Qi4WxQooMM9N/9Mg6INqzc2zr3TDdRxdmFseZ5J7SQK7Zsr
ov8/6ZYW9jdkhTOrucuxRdQgqiYJCZh8nPVzkpD70dTOVTN0MOTbNikvhXjaEUN60UzTGkJ6dKnr
0dsx26WAY9Olt3Zovo+86nVCjwCx859DszPQiLr5Dcxvp4eECUHqmoDnNlo14KvSj/yS57b4Dwve
OrKhGvLNnMt3YKN6bMjdlzFleBz7rRk8jxkZjMXF0/AIzX5HvWAbsCzAr2sjVyZadAnZ+buonSu6
7AjsVj8iJULtZyZEAkjVMEvgCYjoLzyvvwoKRZrtibXRjIlmSnCgkqW+tDmK2P/jz8tXHdIy9eVh
+QxVkgBsTMxkzZjgG+HKZiab4l0ri5TqwG3c22YbeL0/R+BkQa6bK2plES9fY/T1/D23VzPb9ZUu
CbtxHIh/xnPfwccs6gOAG3DQwv3F6yAERYjVko0QDwT4uex4kjhPy08SW/y5hXpyrInjuEPciadg
4bBTRhQmncMHVXbj+EVpIHBwlL5qc9rDX339jU/2PZodb1zg3Dnd/5kiQaMYu+SAktMSbtGtb+/c
PSBi8lUbwNFgxL4MsBySXpOcIvaiqFDbAUnhgGWYbdf66xTahNQj7QS9SeHsYDHuj/BbhKgthh/O
XRRSPQ3t9nARVpS/pmBAO1GWV5SQRYeaCkM10kRn2Ump3y1aRO0ZkbRjatrOmRrJhlm0/OGJa+AU
oETeP6Q/E/W1AJeKrtVwCkyXYA9fEwS0JoaEZPCs2DJ7U0hgU8wu4YrCG5LjXsTR3Asdvf+oIxZb
9j1xKcUbFNmeBwN3XAbJcUk7Ii0XBpPJXJ3HEPDlP7f5JueuccOVyxBuvmh6TVW0koHbAXbSoSOe
FzL8Q/Yzob3qtO2Jc5x2GKJf2pJA40yoe5PuzC7ydwmiHiMe6xhwvbqusm2upnlF7OvGsrpm8JeX
oWW78WxJ58nFc812GwWWxK3OAwWq65gH++gXcKUAaR6sYFu1UdZnc3Du5wvxOP/JEJnmW4V756AI
Q6WaTHn5bCgrHTsY63/A4PTctJtljMp3XXEpY5DH/h+T/G/wYXBy/NNUtrrKhUigF6nmUrBqIk5M
x17eoUITEop5JRt6VhvCUb4fLYK0hle0e1DWdbnS4SxawJYy+eTItA+pWp4WC89UffagnudwQjX+
DKMg7+MDs+G0vzut8cLci3qMw764BUeiXMpywzxqxGgqXD52MPlF9RZX/jYs7mE0ZV/ssYM9r7tS
5X0UXT0PZOMbHsEdcQufCyqgjICPOyBy5eLPVbnTOFgO9QeGhPpSfzRcEHshV8pKg3djpY09lj3Y
Urmn7Ydn4XEWbYVrnSVmj+XVQp2Le0Jb5iuEaXtpSye/IdBddllSU7DvGjceeSBA7CYspz6t9gX0
Jay5vAhxUwPMcYxkR/Psu4gE0WD66in6c97uVSwIHfOQXaalQnOLWxs1w7JIKPNxkeXZkBucoMGs
Px44srJEtPMtLAz/DfXS79REHF/+w6JR1NBVcDToq+3cpKMwDilvcbo3rJqN/pXfGhQturRPwcHw
VcuahJiLHwm/G1ISusbXcYSNzm/Lch3bm9iqcU3AezmsFimbmCSs/Y6qTaj5AfOPAVwJVnbGH41v
uY6Ey2otvW1ghVWN49o+hamEu0aLzkx16JHO5GixsZZ5K2Cuc7b6Q6Df/Eqxu/QBwPXhuZg+wCuV
Tu9xXncayc4qML5fbzadgbbxDycK32uVhUCkiJjjkW/GOb8RY4yHMH5iIi3k2YIe7VFoz7tKdCU8
te9Rk5wJwgJXsZTlDOJncJFHsehxh5k7BNyIZbD6F/qOGPoWJT1PPkfRKwALvmSqqmcs7vub3xB7
e3CQx1TvSrtXB7vPiT9ItgAQ7TiJApuKydDyKzMhe730J5N0xGEii7Uwi0qrl6F70sho9kLScLtj
JF+kDjCLijizAM8yTSqjNzGgWB+VKQBRkOAYM6cjg/h1VMka6oZrOY2paUHgWShjyJxw9bOnqFHd
OZsIU5mZFbEH4qQAuO1duuHrghWtNfxhy+X+aP5RE9FIotHnEEbrv4swgbTGJwHcztzbO4Y1NlL1
MhKWmwElvCS+scQA1bQdUCQkZIbcVZMzaBjhKJE63NB3tO604GTKvxwuS22MqPm4FJOwS9puymMe
jhjFFUb9Z81+jlG5mDBAPXUHFOnp8XMGhlZ3AegD12z+0zXq1YExG0kiRVs/k7gkqUe+Oez1lGOa
mFFMWFKWF+DQ2Hcw1C4sjWPZ9RPWbUAmx2Z4b8GoLeDgzgJcsO3Rl4nYfc/CQwhCknuyl/Y113HE
HMnU3Fx9VFVxHEMo0cSUplQsTUhL1aopgyzjYFb7Lnrlf/PDTU3Ho5KCSgVmK64DMuQzF+V6GZ7y
OiW9Ay8IFQJ7Za+7ejXiEUXPpkEvfldCVSnvGUqg2eljqCRqGvOmvnW02S5/E4B6PA77HWfKnrk0
Qpk7GUl05xYSXBwyjJ/et0gwboftoq0RhopI54t+hsKA7DnNjo/hZsYdaxCjn3FOPZW1neUGGeUG
qiXWWrH8gTsdnBPY4Cmt9OFeMNCsFCN/ru4/WDxHOCyCYG7Bh/+Tfe5rJVFMBtzgQEeyKDeQ0HEY
IDmErnkYCZLmXVmV7HKaRO5HSbwDgnQmLR3U6yiQc4xxLGxsh/PI1Hh9fIK5jqo2Xr0iKX+zne2V
+rb0a/V9mt+36Tppv7HKYwHpsiuk4+lerbqXl6L2cXxY8i9wzpDjJJJuDA3BfR2fe+IRxmhGXTvd
iHVmxhIfMnZ3ksXkCT45aOLoh8c1281gndLQI2CLiyRjMYqxKH/gIEa1dKfK9vOH9GYX+tA/HOKd
KKXso586sCEsXhPEByu2d0SpBjHjUvXNtayOeor2c082V8LiEmK1Ad2a1lxK49dwIK8bA7Qw8GKS
ZPoikFmI8o1R3IgKpzYA8XNtI+8cypADxmK5cJpA8cI8AfWvXjwGIngFE3lv32tJyStBEaosslc1
L8m0UYPbTjpeP+SFpzOdLbHfuZmZ0cSWE+RXDWXPSfUc5mL05s1A3Ms3fqQwDECdqmieRpE/30S/
DAaVNeFyDtVH7kYsqQaAOmT+9Rc4DhKdItmFMXOhYGtkSB5tjaXiztc9i4D0PhynxcoNuavjwDlA
PbyvDWgfGdyFFvYJRsF7wbKEn4hVXVOCOXsvoKP1n3GfWMSWle8jDCoT5Y80isEmBnOSfa7YOxre
TqV+1gBSh7XzFE8XoMlSpeerxqhyR2z16dhdXUiB+tUImUZzc3xf9jHWSSiyy77/99Ha8SLvJyHV
absa6qRR6o7biCz53AfKITo25bic2+9T+QQyt6yaQ9xnwfGOoxBp7yBCrrlDbq2zL/Xfjlynw45i
RrIwEPObfMRHo222lRn5XftvrK9yuWtzGSDsV5NivBzJmDSXeI0CpgVVy4y5ZQROvJ2vVHOLaoom
ptS/Ytl7ab751JCyvzXyA/e8ogFWmld4p1FMUAhsnI36QC/siOtZ7wLhW5JYkrUiLDGH/TXxzYmu
iDUOenCOel4TWUOSpncurFnyW3M+VFwZHJUeNC38hKLkldWqtddBPHf1t4MDs7GTNzstnmZT8HvU
wrK6VTlbZDD+yUuRQYrHu2utYC3q7qwXNCoiC5W/UEUMB/iFq6yj1pE9VpSwAd/zi7Ej7JKrHete
nIqJZeHQJ5iWoEtjVuxab/PYp0876+D6yJ/yX75eteBxW2nXKvTjfjumCPlYlFKX17J09YtwSx7F
gpdtRewXIdAqxFh9rUXouuF9sjz3n5LwS1keBJcpQlKBMJvysRO5Sfw5wPpLyCc6TEKKBShW33FT
wts++4cyBdhGtVZRy9tWPOd3gTOQgeQ2R3M3WhGwoM4WnWRUdNMNjEc3IcblHEAE25VfLNvm2Io4
bQzhcwvN9pQNTQi5vo/1EVA1g6auZ0NWc7CZDVuFiOSk8mEbMgvzGCwLbSPRwf+f0ETibQrQN95j
tRKmR992LTzwWVcujqG4BXTWPprgInHupEv+yiGU3w/8sDiP/7IEPWKeMy7KL4juTyug0H4PNjDo
5NIooQOHQmZHwrh+RV/Y07Vr5pHl6kVirrsZ4DiPv1NrJQ0Dur31pcTkgFax3u3fXNbh61gzyHO7
CeELb1SieVy2ZQVO1AiT6/Wvm9MOauwgBEFf/Tflynow2FeBZxhP4Hxcn5LOCeYSos+dgDPrDRse
jHhHh8fIzCEU91GwdHU+NDZvtOIGaB0JHmMSCmplL6L1GPQ4/GsL/BBJ+kKYxLQ8hUvQucCm7ej+
UZdflvw76Y7GJdb+Ms7Ag6ukrEjdriPYzeAlC1UKwYHHt/aOeseZftvRgzMRd/RpWbih9ojI9l33
sDTBKjn1W5Yhy2AY1B8RRtf41NNSzPXD4yVT2OjSKMKmLLhaUZlGQmW8MFbfJhoC7uMTusCm8kFK
BgAgHmVJpIbG1RkYoiT0nSLvuSRtmTthn4nr10Gyz0N4Mgk4W/WZERFjl9NrjUuWLmVd+wpVxTKI
a8E/iCo+/GIdBTlJHtbKx0pUn4T5wcdTCt5yYiS3mNy2EgtKpfeTLznOp57W6bOtwUZIT/UkHpC0
UxYbqpOTTzmovBQ2if3IkYhw1F/71Ha9kHu9YEJ/R25TJ1rhVdm7xQ33I4K4LHUxqMGoBi5iFId9
2E1BGkEs/f6xgBnizkLOkTj9zlRNDWGsHJdq+c2E21nsFCc9TYOQoHjuKlgufaQCFWBXUEWF5kW7
xs+NWWHAvpfOG9b+MWlFuDlr3FCFoUQPdWNFwF0AjgRE9qVd8a5SWls92q3FCwrjEBS6Ht8jGCJr
GFv1TOxeV6mbxBad6+ORWnZvVoCylZowdqekKV2CbNI4qSbd09sgqRodvvF0shHII4NusGKkvU1d
frcprbQOSPoGTwdShGLzxpy9eS89/2GMSdJdcdfDgvxHRLxOOLcRk7QB5nBbf1gdq0qVrEO8i4H2
KwBCHz0SD944Ofdbqscst6ghsiPLeLHSas++UGJ+TkmPGQA3yIm1TUbLUdDdFgb1cIRuiBD8bf7K
BUyoZwZceokB86bLd/q1v9BTIetXz1WZ0NL2QnfX/Nscy2E3/NR6iVeHexmPenE/Nzxn5o9Z/e8A
KPg5ZdChZlqh+r76BP03/x1+VeKmJyTV3TaLRGroQ54Jb4iIpeBiNZNTj8eHr8m/IMIk8ixUZ/ON
fl27pZpsfPP7NPQGwed8U1n8usdE/VW7U4fOI7F7lWEEadTTMlh3Zf8WnzshbgCiYKRuBfQXXzEI
oZ1+swTMXFtK19q7DSOIPQK4Mr+htPU8pBAp4NNvjZfNdTiX/UOJVlrJRZGbmsX3mAKAtlGvFvmV
4vr8IvT2VmvyuO+KacJrK/Wy4xpMmXPoyX0dk61O9cQIliJqviwlSXFQjEAlTHwd7Qgvfc9qKXDr
zB3LWPe+QAh4J6JnXRy08XS6l3qnnZ5DfvgxioKZVVtD7KG71KKH2wvXmEznRLdbaugKS6ifDBrt
VGK39FehgWTC1fStZF+rSIGjAMiXHhnhoOtgZ1wBdHM7I38CB8D1A2eu+zSAmMT712OFuZFPmnT6
C4X7mLIHIkWuxpNMZAudl1P67LfiDvdOGUWlZnyO2H2mC3msH/btYZMgB5AMzAGT/DOnK2ywG90b
pP/yHFIvKCxgeppUTIcNDS67nSuzny3wafeyPTkgVmt9a+UCKCO5CC6MqL61kkUDifuQs+VW7LLc
Ju8dkCw9hiHXHk+Qm1fPDv1AEA3Frk9GdaAYgiK4o/AdQIsKO1MdFI1EtJsX3WRcYGBkEvE549Av
bVgTZZCZT8EpGCkWRyB5lsMlB3uZFARCBh5GuRoTx5nXGc9k3QQXqmI8TYPRKpB5WJoXH+5G7KSO
v0LmQutPdF6GhTv1TaxDtkK7cLksCbIQIiTE/936XU26WHdJHXv+6bcLz9jYcxrcqTE781aSrQUK
UplH8tMw2fYPFo7gxl2E6cxQ/krJlhd1kZcBVNzel6t+LyOya+nEvMD0SQcpvoJI1OqPIzMV+Eqt
6hIUzdNYhm+FyC7ZUGILF3ETlEr1Z20TAw4QkhpPW8etmCM8ZiCHxoWeJ6PNbE6ouKNfs3ry/tXO
VRhvT90D7icyDgwxFyQqBd5gwzGY/KSy6ZS7nz894xvoJn9S0OE/Vn13w7FHPAw2gR/n0lWubQOl
z3gahzJF65I5a5r23/9WaBlfQpbHHvuG4a1nu2PQB/hSqDD/DTOfgsEJu2aE/JAfXIZpg4TKtWSb
UFaWUmHt8rB/7Kh8GpmNhEFMK7Rd0tCKjQT0s47Y5S+wTOkkpR1dTK4Dea1ZeGbrFxvnd96B2J6w
EKFG8S1TVONJ14Sa8oUjo4DI2ZDvYypDCK+zEsFn7EZ/2lICHc9tY48+cmIBGmEDyps/XBH1IVVk
UE6h8Z+SpF5mLdXX+V3Xil0/BliEeYn9+pHwqUZ7ckZPcIIjs2pGjE3JzopLFgx/cFdme4+ruurG
lC5wLXaGIOdTY/smFpX9AVb+eNtlPL1nW2XAsOSQo5rDLOHqHmRiSA/kBYZuC8kbjHaTRko3aqnM
jbZ3o8hdV8l3OMZalrYnLfGd2IGT5xGicPeBW9B2J5dF+cX/Ayearl5qyCNBf6qJKH1eMdECbdQV
/9nrHVhs/H4uZe1Z76dtoOXOVuzo6DlutEVLkPtT/jNvxoX9olW87+KE2yHp75b25fTzEfmSTuqM
Tx6KCt94VKHAn/zX+OnXeRofg4IXXvOD6+NUxi6F2sBMmqrr2hMsSzAGPvvkl7nN7OyV5iIeczwn
/NrEErs73Wk3eCFWG/KjqPAgM3Zyqoem/fzQWA588hrTsopCGo9jfDNvhVs1izUrsYQWQwhOJjgg
BVFWQF/9VefDHzKwRfYzLy8NN+9M2ldDMM8omth7Lt+9J8EJ3vIOTxZs4ri4IOVi1afG9Ajae551
LbNsVVdOuJZTXbaVMxY24C8D6AL9JwdN2Uzzhr7HnMfA7wMaBPjiWrGMFkMoktHlX4vV89FENAQT
Eqo+tU34KaoBct9tMJeYCCV0k3snJnY4x+Fn4fOfbOMZc4VCZnURXLUoLuKdo50NqmGd9obr17rB
QL7TZVAHup1qa7nmy7VpDv4MgkbSReriNDe1ucNqcI/hCXlE8+7LGhq+EHe2V6i5B6T+yIDQYlcL
SXsWMfID6gKDP6jB0YG8vu9r+ilr0Loji0fbyZ8yd+W/3xPWl/lCTifr9zVmiaR72kI3+ha4jBgd
zMRQlY/mfVVelnbkHpa/Ttse/7/4EDxJnEddXMu/6Gp5BH4yg7ZIMgTozA1/H08MrF5sMzAfWPBo
n93OBN9uBhmCnKhgqprexAGKW37aXMcfZkYKvpxRIEmqzCmOBemq9/v4UYMFMd/SCRCeeEZOeMoW
TcopD2hS3I+RlwK5DZ2FMn6jcAmhHAZ7dtF0/b6nKHpejVXLLy+6vKe7APgUXWyNcgR9ld42MIxR
gXc2VhFMSR2QQWu49RgJ/kOszcvnd6ecYC0aYgmpH3B8/lF7o3wKpxV+WdfkiaCdbjUFO4+fjVI0
Rx8FsJRWwGTYY3Do40EKJy0u6wg2LNz/yB1y0eWRNrWMsfR0ceexNc9/3leyYw9c9DcQILTyf+cm
NbsQ/2HpkrKERthLvgZN266lYauJApSDvo6q7slIH7dNpNb13F/JLQUevTLBc+SFCEmDT7US8/yH
umO2ROOA/2neSqAeano7Ky8gO3A1QCp4D5pzFabccWKwiWveRkTVpWu5H40+dnefhhQw7+tAaUCe
rxoXwVsCfIB+ISEM/e3k+8unA5y8vxoEkeFjr9jbUhwmFmbjsowrMj8ASl8UQlDAUaxuwAiSFuck
YKDVJZE+CSJtBWZE9Np+rjSec5Eump1DyMtPxh/GnOGJQ7Cgf1LZsy0v31PnjdjsqnMxeNJDnwB9
SNTnd7oI/ALSoegFyTvgHlItRLu9Bhif/eehVEH60YbOGpZqNCmbMk6EWe6QZOXLJbdx1fyMoWf5
gYDsBDG1uRlqSxbXlEVxllzJ97ccAGTy3S9Ryb9+pui/d83cM3B864cLp3SMX6ztcRbUiPO2KDL/
8oAw073Lf/Tr8pV0XbDQ6AWDzhK+UGIgzg2BrcHHSATrMwu+7HtuZTfk6zKeLQPgnSutYJNgsav4
OSOd2V4Sv+EoF/PfZmE/wtMnrhbRsae8dmUEfnVMLCQhVefD2jyBoGyQ+vz6HbpJKl3Ny86hZ4We
E4hI4Mxqzt2HU6zRMWIYNGGGNFd2rK8YSW1kBeqjJz0iooQBLvtmJaZTSxi/eCBEejnbejZ3iZxa
RXi143v67B161PgGBOnrzBYLDhhqdO8Pi+xIjdHUWKkQ5rHZ0a6ySYLF8qy8tfD4ffF062h1t8Ta
Q+/Ick41xMB69SiApPdE4Q73OX4Dv52cEq4+43CLJcOOBfr3bazHsWUPBuV2t5vWBDVd8HBuNBvO
qAj0W4P6WFz14T/MtibMKL7CcNwGQ6Dt/vHLPwMyvZXu7F/rXMvJ5N4CLtfHAu5MB4Zi58lwclwu
fp3uF6dS+Dl/dZ670YO74mnnKrqnVKMEAf0AF/Hv+C/AlxpQeBW4NCv3r8r2LUz0m6Z4YDcYDnlP
Srr/Jj0ZPWt6ys4uNwcdMR79RlAP8VZBhgGKkorbWz4K5Yjgj4TJZbgIGfuf4w8ubMr9qnciPWR4
zEvHA97/0ROMDDNdvsp4dujrAfeliFfl7aZwxH7Lp2eeRulyHIKcqsZRLKkcbS0/MJkaf7l9Ym3j
3jaa00XlzBR0sz6U511HHiGahAU3sTRIbUFP4qeFzmVyek68uy7eAVl5ml9rgp6UO4BoA07lRJo9
j4Lh2bKgKgAVflL4tQPgzh6tlA7aXzsVSwaSvf6mBVo3odpd51av2VnxH0dfKo9a4/ARN+a72W6q
TQcsnkweSQWmd2rnjwbXRXDXDYmmiKKr7Le1FDwPfqlZ8iLiZvOmHkCsguFj3Vembr26EmiajdeU
zmRk+pM4448skVnjWTtbr8IHNscusi87XvnTYk+PaBDVScgoSuf5L6wH2wOz8f/OHRMKCj4tAwCy
sUwEIid2uIonVE6W+rR7Hc34Hw14zBsXXvYcUVTJb180TUk+A7JdbsvbM5VtAALP80OhhdYDFKYN
28Dp+eCQrJNjebW21r7qZsnZCVuc1ZR64zwyA42ceymmNMTfgj/0/+xo21HQ3FH2FvjnvpzahGxf
kQinQ1dloybIx98F8jefRNuKKrWb0doLz0TTNZGB6PPYtL/R29Z5fwpcHhNW7M3Shd4UzoTYdB3u
cjiH5ZSXipsKKCIfJ5IvQu4MyF0qct6uGjqaSdFKpV1B2m6DRe+o7J+uK7wY46x07/F8F8dQF8oc
qIA3SczvplK3LTLSAqULWtCybSgdjMf3MnPGB8oxR9UigIZR4HEibDGtm/Or4L6rIPUONP+LWbBh
2IZS/5n7WAYoCvzyNN0MNs7YjAoFH+bsutHaCQ0OsdqAJwFPyBqiT7Uhzwcdp6Ukg0jv5/tmkQuF
KnfnGagM0x0O8LRc5sSijO+y8cNV37qgh+lD2nWY6lKbiAAUfpAJRfwodruJNs7vRpEpamUr1d+C
t+IlXTLoUaUzvXW0TCjk4FZ9dQQUSeTelLpzyB3EWWsxdE7hJGkKWVdDNDSvJLQsIbADwBEFvubj
USvZIqmcVCAl0OF8PSrimegncuxE9ILCu3bjd+4cYPvzy09Bxyn59amEhtQkmUqCupGEGDrQ7HUT
CU9xNR8GU03UhybA4XGn/2WWiz1WMpAhyKSJ59Lkskw0NCOQgKkqNtOdgco9VQJ4JJfSzasgrHMV
XuxmSnxkucv8j2nxHILoZ7THGQWYSjW92WJJ6rntB9kkBa+NsuDDvFhCQKt2VFNExxTCI4BZhcb4
SLlFpgRysjUGLwuEY+X9kp0cFdlHjro3V2/cdDGrKtwuA9eVN0Iq4S2z78fCs+qNu9u5/5e2Ud0B
WjrNoQuP0RQXef27Vt+n5XZtQBvOqGaRNvs7a019KWvQvcaViGPqmwSv0m+aBaEVho7mJTHOVuwx
KwySzfByjMB5fT3sd+1Uuxmh3pBhh2Mjw552orU6zvrADAqzoSzjXgPGQ1/i5nWT5hqYV5cyGGJR
Ntgp/4Qq7c7bEO/NLzL+/SM+G3vy5upIxKgxr3BdrKb2sdoAlFsYOCw8TKgy0KCH9xT7EeFxRw9o
BtNlawpigTT9QpSahx7TB6DKVPwShe9AnVkh4q2J+B6Mssj//YKFSl9nPn5in7y1upCmG9WaPqqf
9QZAPFR2joMeedHP5nyuSymvRzJ2+c8j1GV+y1bOQ+3yn5JW2syBuJ36OMiS+RB/shtj9C3NQeie
YQn7JXEq+vlEidVaG9dBk2bwlVUfP29o6yIhe3VHyobppYkBSG04N2lvRUvp9bS1hmbZbnkES4cw
7/4KHCaby0R9nDGNmWkSS9qYeiCE+FXcxvrTUajh4X1xd4EcxDPwTZKzWMkw7vhp+NzjK+rvtj3Q
2NffxmZi1yuDvH/Oi8RbnKzvsbHila2E91W7AZ4pcFd8DTCkEOOF13Omr0Sa8SGrS4p/PZoRyIll
YUJB8asSoSjaYbFOYq6v7rXe/RchMmjlGfF0VVhp+g4YHBzAinto/WAQ6NusNcNtW/lcew3Rv1Ao
FT0i2aaOZPfoIO+jM8QShX8SZm7nHhr92SNo+BRyVKYWijGz5Wc1VivLYUJ6x3upoK8VOP4AVJKZ
BhCABDfEY6IXkVSczrFJ8i36fhkw70VRgZs0s5nLyV0l9tiuFvKQxsNpmQokPGGY013PvXdtq6xm
DDsLO97FRYpl8+F7z72TOZADT8QLU+YBpzTmrCRNriuW+/FdA59tDheX4miGhc6vf3MUbZcQs/J/
+vDuWCAlOIr4QZPql1Dsz0ISwo3CicQBBpR4GsqTVBqrT6VqwQXjMxuHEwAFdts56g7GB5bjyA07
8LaAVRg/rHIY295XD48YuD0zmTR7hnoIPVYXLpIrpgexKl2NBZjXjUWrYNq2nOwzmlciIEb1IUEi
k+paMAYN4LUoV4fc9nY8w8xI/XsTqMCIrWPwrym9MdHqD+fTFt9f/Uy1KLpjHGYkWB/kd0NtOahk
uTcBBRj+LTKBUg7zbud8ehEL0eGr+sxzUb4v8GSRNH366Ydokq9q7NuhP9l7+RiRe2Sc0oLH2wEK
WUtkEQ5C0zMCvE3GgysK6MK2cg0FPxB8+nMPup3s0dy6uVP8/qIMk+lCAsTM1jEkSu/YE/kAgcZR
Q3X8AWVizotm1J8tekOmqm7vt0KDPBf3f2h31GmYsmSJ1Bh1mTiPp6FkE3k2HGPNGhhb8LzZUWYE
SB1qrTweXt4IwaPIkGRCtX0dbnkSkX4/h1UUXwbuqtaRhC0hg+FJrsH7xnr8rYRcoXv2GO0UJdMC
fwdFnJ2Vp4blEIxufWrLdHzOH6ZEzrIsPzRxB96WKXaNFYUOxS6IBQ9XU0YOt+UMK5pMhy+cujWW
39BedXZR5CTbJjUe5Uk1Dszg2RwpmZT24fO1BZkR1qqdgVz70U3P0aab3s5u/YT3nOk8NmPv8vWj
Vsgn6BLTgW7P0I2lHywwCULlwKVXKaZPleor9lXHrjKaIp0zJ9B2qcA7LgZ37t1hDISsKkcrjrkJ
3vbYjJhaPM1dbFsmtnYrO78JK5/2vr4WGBZNMT1rhH8qPnF4MoAjer6OK/lNmQauUvwYbm427o7/
EY1dLAGFHAgsgS4Fo71oAA/ucNQ6ROkEqLU0ARYnWHYjmR1N7jba9+Q6y8wVaITd1T1I9boKQ2Bb
DT43UF95+vLTSdQXHqWlhgA85+t6WTEVP1iCnDW9dPdbivty5OREoT7lbdTTTZJz83gNGyKExGNH
9EWaA2fUkpzYf92QxDZzs6jcpQ43HJ3eeLTs2NGAuQZh+4vD9lG3zo2fixG6ZyTpa1m5zOz8ghio
wmzspiVq90SoRR0hAQLKsVEcCdYsb8F76CDMqN0oG6zEWlI0q+KIr0lIJIsb2qMdW9sklOi7JW5i
xl4dQrJpmIbhLki5pC5jwWRp4gGxhujV/p0bmdhk2e+stJdyl62T5ldhl49MwNJBnIIabe1ZidN4
9rMq2vx3xBvBA6fXJN9hn36RZVBSFvftDGt2/Yp0hGUMy0VnGOVC5yGirZGF53/2leWxd/a0ElXJ
EkhUPh8DugdRINyJVO4WtQLAoXdkPyNePZSlWBu3SbjNksVEuH3YE58SDcrJ8ppnJco00abebVPH
YOvMvrJFk4ATbupzlz2Cp08EAsfr4QcelNEYDUpRAwAR0uodZdbR+9ivTnLgIOybr/zEshsU0ymu
jU/zvHAWKgUZ7g9XA/tegJtqU5Jz99XVR7k8sStDb3wX5MXCjwwDZ6H10jTvo1nxszCwZxI4GLNR
a6Efw3ZFIulrA0+OjJhJmAJwAG/03IZN3mUjv0EtonGPkJVI9VgVuetYmE30zOnIwZ9WHDISo/u/
WpdkTCFr+Vpykkhgnocl7gO7jIFrRQrnvTZ+iVbqwGVyz/GF/ZLuJ78JHmH6rj7d+astkJX7kAFL
7TWCLx5pZTIeAmG+qR9DhWskUN4OJ+bAGh4RV7uLLBi4Nyu8sWLWsNDkUNnsflaU8eeHgyo0gkgu
cRuqGAogmSyziRS0Qnc0BlVeRHCXxr9leLWdhDT3Dj4MUNLYZ5K1aJCrEIUbsOALHwjFmx6stjO4
rkvnHEIz70P7RQbk4Rlnqf/WIsSMfSk789TC0AG0E3eGA+Ed1Ug53R2TTrhu6wuGE6Z+ixZ9S6NN
MKRfX6Iraih3E/tm8siaaDJcI6vFk9xFKhJZ9nv32dU+Bc0usqJPUq1u6OWlIz7FG2hEbWj7z1Qy
0Fw+lOnHhSDF+moYD+LZ+l5HtgsQ64jBMt4RAsw+QyhqCxRi95WY/H3TS7183E+l6APJaaITUl5X
+KaQ4MwbCwpzRFatpXaBbVb8s59E9vvA4Q19wsZaZp09+fwX/p7Wd4zA2o2Z1kOY6azVvpMtCO4I
ug3EBWlq2hTR1BsWtsRx00EPxw0JQQEAROc2ydktG4+h/iaBF56N/rNY12YME1U1yjiHavGAukkM
ZT50aMcMgCuOLY+HQqudXTq7ap+uGlNaniLUN5qBY7a0CLUHYve3S7/dFwDPMOMYFFb/h36OSYB2
18pkmwPws241kklVoSOB4DM8ZQm+1aR0+sGxdrui+6BmMEtxJ8g5ai/W2j3X9LxN8mSFhBBr6JnQ
MlbLOo1CsM2fj/EuVingr6f95kuQUeMabJElWYPLxb1bb1ctmiKQVJC3IjBBC6VI7RS7Qa8Bqk9i
gk4jk5kQzwefBfqBu3cBNWRXuNsLI1uhNZdOt5n+d/ZcUN57qllRLfn9j4iRI1gVXdMRX/HijWAl
7tDMygYn4b1tdRFXw8YZWIlWVBAFNSUyVSpG3NdIBrOeB2MqXzbOAmtayiuDa1YlH4iLFnQL6G4A
XfSpe2d2HAeOWZennR7Beaei4mGwQHiIpJ9GJbrd6RJWwkqaEbhljZiskeQillLatUQIn/8QkqsY
gjWkX8IsYb221rm2Px/eGHRIWP1R8xYARvDprsj7F68HlVJ8qfELlyT/4UXRfWel10Z84ti2RnBi
HK+T2ooPcLPBuprudMqTel43B29W153XZM9UmS9Fs0hRop/Zq+c04PBjOiEB1UKmjnDxhkyeGmuj
ttGYZ4GfYynDeT5DzvLVII2woXU97vhbJql7g2d1mIbZ8Ydu9Z4YHBHkJg9BLUdBgumYMzEiOiMK
qclZUQopxBrm2ZOMwEqco9vDeaitJu09pVGsrjnij73eOhFTOHyA3+oIumriquTnOoxIhk1a5Y+9
+Jtne9ZRqgf+ucrCBNhXp3xA+6LWC7ZR+NKJMxQE6ihaL5URimuXXSbm7bIgkElnQUEPqgkfE8w/
79ZT1ab8DoiKiDfKyyfSTv3VfT81hFR+uwRRAyoXUD5k9fhxi/EOLvb4L8awc/QhyImSnfI1kfBO
6QlOMqjEWBnZE9mxbLjvcWnIwRridfcL7SmjQX1D0NWfQf1D5f3KNC7YoUr+/dWFGrsg/b2QEIB9
YFeD7CFJWa8jtID7B72Xu1Dq9x38g0eUhYh5mTj+nMtmOufhppkNThn8e40hRo/PDCjaHDQHduzm
Qfj+GEkhLKppHAypxCJ3GRWX+25OubLgUaN90X0hNK4Ti3QC+cFsUFeuh8qqraqHn95My6yKqaP8
/KeQtbhuoSwyIOGMlxwWfqZWzBMuP/Ca8ErUVxWijM2O4UhYQ2006F0unrw60WSpHC/n0j0BWESe
qyfEfyunNWTsyPiDEY84xIHnXJ9UUGJpdZXcl5TdGuSO11p6zgTai3cDOaOwkgxVkQtZHRWRnyoB
UY8M3y3xuvVfKwvFGo6wu3DpfGF7PvUGLW4RB4L+uvRQTbKwEwjwBarzygzbt9SmYd6oVtSSnK/T
+IFWNnPNvZJKzm6bsg4jnI+f14DsMwyB5pc4NkM/8sXKUX/74ODd4e/ocSBHUT/dkIIiXbqF+GHM
rku+l4INqum91U4K54MlII4nSRZShXUkQ8hG6MMRxim03jIn1ptPoXHUbeW2dEItA9NmGyh4xUQ4
Rn7aiXv9pVPlMLEJ70+An0HZT4Cnj++QkRYe5X+UFRaG5PVVQoSMJQ0zn8QZXuLkcYzIXCaKF2FH
8Z5SnT0DxG0HQQTmJPaKPCwA4VeI5YlO7SVVUIMSFk6Kv9UN7Jsvl9C4vFTqEgNf7gam66QslAUJ
HhUPBOd176Ku6fvou4+PIVTjE3dVCt4W5StSi+VN8uFJ+S7ooDDVyxXybYkwB3hbFI71B6Yky4Ws
piDcpUCv+PHfA0IJZ3ydOy4CC7R6loofCMEZqSDxC76U+D9QrP8N3WjegEvs5vuKz3ydoX9fSPvl
EOFpIHg1fXQh48tAhssm1gbYffz0TuJK+mIuSWKUbfNjAoZnhmIy23bKdttpuPwEBmTZ/q7zwCNY
Fp832Fotj/dskOKsVVd9OIKRbz9fl9viN9yIcNNGLeEVuDBSHAEdFZZlzfUgOxfkOP1Rbkz2Y928
/wagIgFnJnkI2O2CP1Pzt01FA6ifQXRL5B7W05TViBORcL4u1R4b4SowMtrXpLbl5LL+A3FB1wwI
UTTU5kRHWOjfL2QIQLh8NipbzcOABLwIbIXAp/k/fHYrcVrqOV8GAKzyIc97up/4Ru/TSmgeERUO
Twkaw9cvFWqXKI0PyL7oxhmoWIvGkeWaa1hfCdVauc+ieeglKVrq8VhL96GKeamsxNOx+G3yTDaH
stZe9kaO40h17OUedf3tF6IjgY4NoA+gdNnJtD6TBAEeOn4LTrwf/NYC6kN2xzdYRtXfBxILpD0b
xE1HuuU17DLY6aTQ36Zni6E2rmkrRAOXP34wC3dtoNrZQla7ytzf37KVEcKld76v6GvYzZyYBjjm
fd/6R5wjKPkp68AXNm7GJBKEKTNPmzT1zWcfkcWgkIyp/c47Ln4jSUMkynkMfic1SiO8GGz6p784
nIZiTrQi5IsTHyIIaBbBsePqkrv22s1cKCbWAoNskHsAY+ha2gN+fasrZsusZez9Gtq56bbNTiIO
x0TFtxHVljjoapK5MwnARyw4c8r2oGchiVqqH49m4hLhPordbPpwufeyHfGed+3wVVhevyWIZmkR
BdUGFt2/06N4/wy50GQXiUkzUIDrepzavsFvyymP7vB3HJqg/6CtmAdN6ZXCuEzh2GDpMdqHNquT
Cx8Rx8oEFZ1xRct57LyfF7xQO+8QOukpjYM0+U3wEkDthz3BQqqnWvYAr2GOUEbRvMiMjnjy+FCF
WED3L1en9tdYFGtzizPe7fC2kxhDBcvSMWyCOqRm+QzUh7YNc7lAELvAt0ohDL6axZMkZ25fCVZ5
jsuHXYk9vWspXV7wMmaf4jYJXgowMt+iP8rOzEuNWFVZlMeQegwV5dhkpbAf0JttQOW9NsIRqy/y
VCj7Sfj+yoBqVrIY6HbbFERW0b6Y/A9LkQ/8vlidlBxSUdXf4nVZf1yjybKiq+Qe+PWnT7uL5Nrt
O1xiCG98wV7P6YJ+TMoIbsThveI3L9iAAgDQmNcCv74FluALpyfSxLJwOcvTW4ivkgJE+JrfhBSZ
55h1nLoshovAcRnh6hCuAaluDdzj4vk738M4bQ3zhUy1cB3NmKMeovJcxo2iVOd6MtGuF91kvciM
pwTP3O3xgdqSU5VgO17Xh/NM0cjSevfjzQbdQ+Fjt38L+Q4FbEDyc/hHKsE3o4gVc6wRhcgShwS8
PhOOIoJyXJe99nQ7zCFhHmZ9DzSqXoxpjd8ODLOYyf6K04ijUAn0qZW64kO/dRTRuZDLtFs9d2eP
doXMU2rGuQGRDsgqonH4TFZYUjU3hgBbaN3jVQZPjLzE4NirbdOmc1SvUNZ8ZRqpNQDa61zDALhc
o6QaLmRxjBrVEBzfvAWEtKxXDyEwoqcht15QGCzP2o2ZkHdIlb1GSsbmse9rythCJwnzJKwOtlGC
ttc9vzOg+6KFdm5L5rMyahGZ02nPEImP3loC7uqB8byWKotXQl4sYhuA2RZS0SJj7XtJIhO8R0MI
SSbmt9J5r5496y2Z0Z5KBoGM30TSe4Z2a7sUjNrFCutnXkGu77FEoDKubz9If1+xwZxIm7HM9/Q9
nC9VbqKehQND4tsQhdEXurt8stni5O41lpLje8p1UKy9yCz8znfH8FHX4BB5WAuCCYs6KhIRjuHZ
xYczYxSQi2TdqjIvPHoMYXTXZn4MzHHoGAQSl4jZHMhHY5jzJadNUr0/v3OpjO/2xijNSGSA7j2T
w3EUYwiclX9RVRRaCgPmddpvOSBLwgQXR4hNvPhmg7sKrcg1hqUTDBP9bcnw8tBOoh8mm0gh+55V
Z/Opwp5pUfLBUrL1qBOn/eQIzdAXFHPUQOmvEEEzY0XmeOIFFoNUdGtVtLNB3GppLu6Sn00p75+p
FeddKN1fxsvhnyJuSfp9BU/g2S62o6wU+8IytVD9sTnNzTJDiX+4l1uBIhEsCQuLOa+UOnefbMdT
qqeYjxcqf6mCRQIushvTTijXlNjVsuyx0xn/1yVhD/fpQEngmpx6dHl/+mDmC087SABZtfiSCvrh
0aTaFBdpz11EUoVGNix+3FfpqBy21DB0Ofjl/L88++q5+1Qc3kYMYLltPbiu9DL1VmQNU/Q47wdJ
p4XoS+vDGqALy84soKhYMOq20QhYRcwRTDnEg6CCi/vAQ9mCtq5XYo/WkKqP4hLpmItBIG/GSTMF
qGpj5S10wwXuGbwm16dEM/hkmHXeeDJuPDUjfrg1BZNik+a1kvpwA1E6qLraeej7CgskokpN6iC/
RpslLPTi8w6UqsFGIRysrskaRJdd4VNZ1Md6L70BWGBz7j8BZoy+fl/IMa+TD1LVsjPqZ87eFCCx
W1ddUgdffucn9/WELapzrgv2f2J/LAZCZdIRyjs3df9F98k66NC2LIVw/Kd6B1yf0GvFKeYSvPqy
xKHbJ0iXvMEb1ot8t/bk4+v4ut7q3D3hOyjO3aYtW+yWdr7FGGxV9Qlq/vN9SBsBQ17Ii3qi4Nzw
A2pevPlYiMvShm96DjcbAEMC5DOqoszKkLYR61GBwoPFD5aYMvFxXPIczLypwt24imOg1GV6sXId
8EcpRe+ToyXy3TzT49K/mGG1hTlHLtqOtH7EHBHyvNuPmdrZfZ8rcw+tXi7LkORZs4kQOBcvT+yn
eyR1AIluGNpcGvvoqL/GPCQ44wt03QZdZiUu49ap1x1JEmcAtyectBFUnJ0XHygQsFBS5Jko2j4y
p1Yd6gIrNLzKHKuCvrq9jJqpzkj2Mf2/YcS7UuKpFfa5komkMJkHAtmD2LEPODvtprxSjH2Q0TVl
SNrjmm9KGgSk9Cb1SdbX4imOyB8lBdH/mRj599fAzYcjZ31g82fgHKynLXE7ftFoEa3D9mNLpK2F
oqHlM8znP+k4CHJeMwJXgQLsg29PSA703rGsk2mneFK36Vud1xA/K2BQqWAocN/P3HOi0EJbIMWc
kA083/orRliB5lyUQ1NcinBndQNDZZpp8kiyvGO5klqCQyJefoz+Tau/zmo4x0cxuafBZZbjHiz7
qX+8vl10de1qJYK12Trh2D3NiKP7ZHEh5nPrxwUa9pdM2r7scDx9ZOKOKl7L1anV8ZrsOjkeXQ52
h2MdbJGsrPZH94WLpX6kGhUcOO7iElKh3uZ4Mrnk+nKld5S5m5V4PZxI5Ii5j1J3wEiHl3uxrolh
6ji6Jag08sm/d3hVnLahUcnZxuz1lfeiI8+UZJlSiXf9PIBm+KVTpIwGHewZ4W0RNHd9c3GtGP9k
4B7Ck+bYJ0SAJ0WBNbgCJ1KSvUccJN7nvhiZuw/dsxxXHQu9Rv1jbDidzNF2S5nB2oN0vdEoFKf4
LryUEOhU984K3MdBO9c9XRRyIpESn+lS/tqNcaw0vx867vQyJ7Z2bquFIxDAhRjgBRDjTU/lCzFS
t7T5ufAqns0r5i3lsXjwH1Lv9Gk1taVoYXCXwCmP836Sm8Cgyi51MjmV/Xg9BeL3oh9rWkB+VATS
lfP7vQI3oHi0GlK9f4w+nR44+5Q/P1mp786VjxmS8YReet7fDoUABxpcDDDD1gH889pMKfVmKaPD
9qbCtsxb81fNNxHcOr5uPI6pYISVLhxvOCEtieKQt6mMvMP9PCOKWg65D7Kp9IY+sQx1/Y+nNZWU
TeVg93i08jdp5DowoM7eUEEdSCEVH4DhQZce2mMvFZ1Se1aiph7EDcz5Cqgqs7x9TgcHdX8EOpoX
kpYgjdq4oQhDO6wirVzujeHhQyswa0gHA87OTNVuN8ZL8U8gzZSWbX1lcDRQVAu5kedIP16AR+GE
S4x5xtBdC9rik9HBbPiZLZ3kDI1h+Ppf2cUjiv8Wdj+JQ08Py/iyK/mzM0LmtbpcMZfCKl8lNmz6
A8lNyl00e3K1EUOR58BtWXIr+xBCHRHR7NfGkv+OWD78+USOV/O2hXsZS9AmJxpnOZ+eriCtEsyv
Ob8+VP+or+kNBwEGle1dDRj5zJbwcWv5BmUotq1wmZktL297BxgwCFK6v+/25XS51cx0Ivr4rxn6
Gzl+3m5naX8mXLNDc9K1hzRAKU32K1TIlmAonCM9JobFxMTqnUZK7hE2YQ6iU4vbPjRO5l6PcESz
8LabBh2YobhNlT96PxJlEMwhpvFw56kjBAwumRktlKWmbnmoEHgDHDvOceR53NetoB55M4iDo+vs
B88BGdw5eN1C5VIASg4dKv1UxEg4PUrdt6Cccm+JcAega0J3F8EjyxojAq04oZuOSHx/rHr0klon
MgW1kAyjWq9VnpF9JfsIh/YbykpAVRDuuKh+7CSOMNYUxpON/h43HluWQ0+f1fpgLnnA9w0IDtfH
JO4PIIt+7IZAcLjps2/NfAnonK3mF38EVnQtzD3W5lmDMxLDQeFJrIxEoRpkaThmiK2XiWnDU1R9
/p6GFsUrg6iK5n0SfHlCMmLO0FucJYrC1YzNPofO5ppOLoJ493GVIRbVONf1OsDPEfV5DpD86Ten
CdMyN8JTtEnG6lcz44XIN877+guTU98s95so4v+ksni17SrFj/HTlmnPwiw4S5emkXKBMqMU9xFP
qkJDl/ASORfjcbYTThPoK6kUhlVybfQUPfyKwCa/jydfs3sRNneDilPJjvDLuyNOBdq1npy9o0ed
jx9ffHwrBXQ4Eb8ZhtefbFEHkpljjRnfOe/OnC9l1y3FXM03PFONa843JwnTHZejGwbMmqsWE87A
N21oAgXP3DqwggrIiipgN74Sgqjr4yByr4WPmYpa6VNpk9L/E6STs9QTXI8E2Sz6zkhNvZqu2WDX
5/rj+jH6T8vx6anCOF3aFkuhMDuRr+99T/6ti19wgqw++TlHaMbKKNpFBz056lt1NcaHyyCxPd7W
cV2LKPcw7vSziwm6YZDwTVk5nc5CgbN2/WTjkJy3VTg2xXAYujAwtb8NPuGNA3yu8UhR1IMqfJU4
M+ubfCfY/WPG1UpGLNl3KEbLh+ODwAUD4bNXvIRj5tvIOVmXsqDrGbyKAUHWXqeMBDuTAfVJigid
b14G1M/6/OR++KiYfQmAWdz4ZRL9vtqaser2BUaTwmJBt6ZZznCfGDt808m/y0muzix00+e9clMr
fCTyQMShTlH8y0pIjFrjTeJbtitCtdC1YbMIIIGH6i/GSq2sgvHd18otyry+E23xxPRmNzVeTDVw
wXOqrgIWk9n0jRLZONhbU42oL7wX/B4AnXF4JTdH9pPYbpBRxLFW02LMPzooRQzdBbSW6i62E5BK
Xlsbho1TjRnVPnCz5hRdKAaJvWtsFSxnTidzqloZOZFoyhNk6TlWbRRMR1slArPkFs9YeLPAcd4o
zT+r+gf/s8u6yUp+TR00p0ErjBcEdV832/uKpn73cOuLFnq3ak8s6JAOXfJRih8Kg8OvN24ZauTn
JDoOxQ+1yAa5zxgGIlf9tS/vKc192Zuu8boSOtNMBx+zD4xLtSOx38xWpTJl0OnzAirjFZbtJ+ZS
bejaicz4GM7q04ESJvnpPr2kPYXvtajKrSRQARCjbSRAw4C3GZ+84r+B985U1s4fqAs8Iw4974xN
7iGPUOViaMT7pYg79LnB/ORUNJ+t4zHIHbafAVurcztga89qbDXKOOym7Ye7b16vT/xY8ufDaEVw
Nv09l2EIsTLvbuWapMqrLc7VMSTHKZxzk+G0SA4Lz2lML+xLT/W5Q2eCSNyxCdBvs/mJveDJOiYe
xHX3IKOM2cYSnr+37zdT3bHmoU9c6mXNjUEhwfpldKAQg5PgnTJyf+/w18FyWuaiQVkY0YyAybPv
tgh64hQeVG4WjFcK7KfCZNX3xiUQEklk2gj9WVKpPsKKjgR0hXJdF2/Q+ls+TcEGai0Au6k13lkH
7LmAypKoMy1feWMCqo6kfyqQmOPZmkCfLBIyQJ73FRafA6U/D5GWxQYqWQM5KOr+cmXEJDf8kV5F
nvLJA2IBg04HLXPB0xlwZqWlK7yl35Hryq4218FAhEx4ENQxqJS5WuVuapfl5V27UAXA0gQBzbYb
2chyar5xri54JTLLkQAL+5xyMlR+q8d8F0uTossHcdk2dsL3CpH9VaTOuww4Ku92Qnh30Szt52E5
aRmoH5TFf0m5Pkosuqx8l+ryvCy43KG78t0g49miFmgCAGX6+23Xmgk6qn0JZM36EdhrM9cztD0h
GtEWpTXerRAEjz3tvjOV9m9ITFp9YCoXSIWDV0kvRpoOmuFz1demkobn0ryhS3s45Ba9OCvLlI3X
3HwluYl7lZ8qBH6gXm6qsauhMTgMCN/jvA5oK5YdQh/XMhtU7jQM+j4iMSdA9E/dnXjqfvzQK9Qq
z219yJjmM6oB6L2KtCkOJo/zfZsZO3BzHk6zoL6Qru7v21GlvRQa6/0/JQZesftTyJ3RiG/kN/G2
9Daf2aag2YaQKZT0u4oxhuouz4jQ6pkvQn91myF/R1q59xct1eyqeS9aIKjoLOBe+MZbq7qynX+G
XpiLuF3c9IFFOa71B8SW9LhyovzKcLdeZax9x+0FHQJ1cg2y2WomGj98y9iLnTEOeH7M1AeY/q2S
J2Nxqm3ZZPrWG+OumwUNOMpZU7OrBJWH56omAlwG0viSGcNSRCFqqXY0bCVynK0i6R9BbvlR37PN
HBkQ7SHgI0pIclQ3ZL619VP2OPvDCYmMXcqXTjWT2r4Wa0K66DL9Ri5uiVWcCQw7w5aKVHSC3ghy
HM1/xQi9W+CVkkT2PNMeQPuH1GcgHCyR2c1eSqgrQoZVI1XQrDAtmfMj8cPjkyYUhOHsfepWiQTB
5mGk1tusS+Aa1HGWF+3k2c0zZY5iX19JxV/3tFZB0brJP1k41+Wji9U7R/87aesEJvRmduW9rGvO
9ZovyjrUrsP4vrbp32RvV2sQOXSexe9u4WCoBjNsl09eMFtcOExwwRWepAVrORhibxJsN58b+i0y
EtZ+Wnqnzs2tEd1Kyz8QDq4qALbCQBUdOj/vy+y0C+QeHJSvfvzN4AEcL97zFtZ9YRTy5pBn1vXx
70CKS1LovBybots2OMzN//3e1TNIPXnYlKDeWPmFALT2aTQbkRia9HxOhjgW/Cq6hPgL6OrRckI4
XukQI6yhUCZIdcx2GuKPKnbrN0WX9cVR0rgySN9NB4g1F9gYeBs8DK7L8OFWNHJTqbN5TAJgY3Bx
GhNLuUAb9dYelI5M5B65QpVso71hKjK4PJDdDy4HBgbPVCTaRGIOeyz+MJlyCOP4sT+W6I4/Rgke
dQYm0CA1X0MwT+wi37fMqoPya1+Mbvo63OOSVK2egjQKs0GULRD3TC4VKHkIWwPB7E4vid31749L
3RpCsd3ZydN62vb6MoAdp08SAbg8TOeXxZaWOyNNrYq5fLu9DcDhNyfper+nHmr26gLq4yJ69cmN
oh0auejvflNE3r7WoPhB1+8Zcen4EgJLQN6rAF6J9BxKgvCO1xE2WWPKrv4ohizxqSSLaP5h/wfv
EAZCEqSFjk6HQfTTih2ZzztfU/uUnBkKBWBu8fWUO1GmffcG63WJKu8SvgfxtoB8PbAViFQqFpM/
wAWjZzTfEJjRqSz1XWB0r5aPZJBjuF+fiUofORfcyejWXFa+KSCq6Ce06SBS52vDimpsyzBghm7t
tDSsjNcWqv2n1eNjXrkPlLPiUbwMLBRLBsmSRxOdXyKdDIgnOCWSy5cSjmKaMCj7cgVe6q6t0Dm4
NjvvR87cCAF4yZMC1TTYxeks7g11+nHjxErF8r9AlmVOndMd/yEcuoRAcrvqdHhZUHmXxMpFuQXL
XID+jXMyu3LmGbkOKl3MvldR1Sx8igaiOQds0De4HnX2dvsLndy8jkUY/7OXye2Efjy7E22jNuVY
ULB+dAl6NkRn0ZAHZv8hpjHjtDKUDEKujem9Tnc7KYNumjBOjlhwxqeBZstiMdIbGZKCCSgqh0fg
Pdc4oLs+O0x0sn3vI1TwVvWpRBQdZA/j8u9x4VeC7rc5qO4QXeKEp3rgGIDAtYO3lXW/WP/0M3RM
kVSnxay62C5b1BvC5yvjz9KrIyE6ZO632dUhn9iDIMsfU7mtoQdg9nKA6lFYqxFkGWma8sD/M1wV
v2nWI8510phMVaCQsBZEnwMMfnhGEUOk+bos5FkwrODge+PcrmViGL8xNFOH20pFs50c5+L/LyAC
CoKMUah7PtnPvh16xfNCiBUnmr9D9dLqW+lHiZ0mJl0Oyc0s6zLuXYZ5knuesD363Zo8VV0IPiBN
jVZFtjJMbm6RiVNozmlhsTVoVaABklzurOsBMKPAvLbQx1Oc2a1lFt0jhM64CB94axl412OinO93
ysgRBe/6f7gFRJPUSALtKSCTXCoXpXkxzsf94mzjIDQd1P9NWKhHvXR3p2GoXvHpZ2xXDsDP6Uaw
z8Oel1Bth4ukGDRdPAYZrbIxhI2/odXexUA7pM7gAS7X4DoIUG3FvmvBB8Cm1IJ3lREOdd/Btjz9
5HhqmOsjC6xRTINvNd9sFKmVI7o922LCJPdFkUiWvCVp7fP5g1HMMxjYwlSi9sgoDGcxBYOckhb9
pa+9Ez8mQ2cWnUdNvwE8k+JxOWdU+dsAI02mAQmZpxpvcYZblaPod6GZeUnlYenK2j2/SZlTJi3g
sGyI1f6V79/xwr7Cot/9FmpYK0Z5r33REhP/JbgGsZGG2qwHRxvIq2rhXkMYd7oNl2gTf8R/fg3/
JT7LY3X4OEDev5MlijyYZugOpsX/8eTMx4yc/sc5CL5x77I/v6MwAAOEWJ3aDkU1wCgLD9tCfyDG
3/50Kq6UGdetpWs7u6xB96reN9Qv7lFkEsK6EXNT65YjxtkJjYk2Sli3o79X2m8yVEYNsMVDn+3v
PG/YldRNbE9h2jZwyPw1JVOy6pH7BkcwhVKe15nxWMAaiMvA7fLcyPNhWEFFH6rlBxfhgrQecjcB
eSkpueD3PySjv3iVF4QgQwxK7SEiTRzIKXHoEheQW20/WPIeNVv9MKsc0wSL6RJo552KnkQijViH
NclJRfU+hirmqqVyuQ7HZjTVpsJ9qgRBd1qeIqVU1cYeqXowu2YM7ejdqkRrnNmFqXUWmm7FkR9V
cTVYl3SZ/tHT1SDAepQlopd49SBQ6pr/WMrrIOR8BWsSQiDqjsRShEOwdrLchToEkvfrgRvGNBVy
r0PZRy5D8fZUxt3dNebB3CJwfBuWoHn+qiIfwGDggx/Z7RJikxvITi6giuvVr3KIyuLR65uuWs19
7A/+dmcZbsuImfaS2DYW37puur3+IXCUa3yCMudvQiIVANSRn1BXcJhexAlTkdEoVgN2TQI4Mm5t
fnCXVcghkbXyhP6cxJJf/Q4ZC/ZtJDSZBZmlcZ/NQKVQSuSDXgoYYyX5bW9/him/B/812BJ5CoHl
kbrUUEiZ9211WEgIw27Z6sZg7Zc2SrEzZ4Ocay1QV+fGjWW8hjOQE41Bmtd5BFRl+w2jwQ0q3OL+
sk1VBsOGBcdSoQxjogYmKTDHvaSGqFWVA6/NTjRY6S+WXMAs7dt8NaSmTx77hXO0zTAd1HuBpbZq
JSvPwmzZswXVbcqlIz4zErLoL5Sx5kO8s0pV54SrI+OGTwrTVThNfaYawESxBjU0If3AXcNsmVsD
tuRAVM++zhVUy3qNX+eaeaEFAxQsw5o2evJVeVTqqqTvaPtWXUiwvxtq1qDuxHIpiFS4aTnce7EZ
xWAhAPIjhcZdNanX3p0Cx+/wNd/GvGPxXVerUFIQdD8HNNrWOtoLxlPrKIyTLWZ6X7LFX9d3Lv41
4wbKODi4RMh8HR/GjrVeHPro0jpGaoFNB5LsW/3tEG/ZRGiAOGCxEP8lCF9YlR5mqwu6LVltcPO9
5Hm1BjrLOIL10n7QL2bSJBQvJzeNRynQ7RsSyAFzU+D3NS9e4OP6xt9MEHZv9DqwBovq2KR/qElT
VW51Z7lpqZ84lym91+/nzsiyL7mSNxLlEmRVoFmwcs10V7CsIenMT+GKiMDDg7uOOghSTqxNkb3+
Jd+4QOlR3j+lxipmMlWjnGQqebpGthka5gLU5B+m7AXgplSGlzAh3q7ZqhIY3SJA2OSoAyOTDDKE
JC8NjhpwFxI/vl20eO5JLY8H0wsAGd+Ah6ws0/LOHmDMckKe1FeIYLf48nYlLpzWgBuggm0mh3CN
W9/srNbvYYf4DPO0LtbIu6mzmy9ziPsWAbCqIVdFyezK1+YjroUaDv3PJQlHLSNA9RjXEtC3G9xZ
IlKWoTzM+l9WgNfbxOaL68SaM+9gawzwDmTGk1gyb1uZi4WNQwz0Br6nxvxUWy0vNFbcRGZI/luu
Sbh91brGUW/2tVUI93CTZ7iDWn5pDu/XtWDOO1nes+gNnH/eRz5VmHg9tI59S+sgyraKG3FgJ2Et
2lnQ8PdPPXS7xJzfVsaecuhDjFfpLxhmu44lisHIUJkCUyBiU/vrBoRCxNfJkg83tuHLiNQkgf/T
XUJUPIh+05AalyfKFEmM1hn+QPAZQaa6OALqu53L2fyE3QbV4h+qMrm2ed2/EuJsKIwqJEP1oygo
xAtQXoFWnYvTI28ifO2v/V5s+wVfIKYlwV0+KDNuW/snyGkmMO4yld7aCYIXWgaayGVEVRD9ipf5
ZeAT+ecGIAdDmn9hxUY4yKD5ELb/82S2QAArXsj4DJ5XZOsHK4doD0y/hoYXqZ5rnhD6eVGuDoNR
+oIUr3rWNpveAp5T2owTqGOZgA/hTDtMiSaEYXcRmsGjZGf8jy/XiLz8pWDkYUX1PA0znSNI2f3b
Chkoh1WBx6iceFa/NLaCGYkIf+xRvD9ej22biiwY75p5Hl2WTNeh8VtwummEc4258eq0FktmbjBN
CJjlseZ6UV+VFxoCdcmPHARAmFokUT6i3z33CiYmqsqN+WUetJkCRugoSuYi0qZwm+slqQxYDyuz
x28u8XeAT64LbT2ziZEf5Wl9yy4yC7epH0+Qq91L2U5NauFNrx60uD8dxzh2q5/93/mKjfHfkgiU
6lr+msVSVz/MCXnFHHGNGAV2OZNe0k3pmk5CXgZjv7B+JKhDWhOMSaBuAX6dV7s/YvAp/CYjAi7o
Fn1xsJxrZGsLHYlguartxO2Juw/dCfoEMEPhk7nIBQKTD/D5c13hjwohVPkNL4tLIJ+/wlPWq8gE
Qm+D3zwhhBJajFXfDMxoK2Kf20veP4074FKHXKWlQbl/staj/Py4V3I63r068nScd2BxdQYUsTpW
Zo0ofRfV9CyCPWaUKvyU5TLsBmlbGInIo1CBGdYhhvUeERQBNT6mFjzhFsgCKX0XfcGkHZV3o5eY
rXKiV99K8EdYPKhEkyImoeXRjj6/WK/m3M5lf3WNniXGsamKDzH7samLHfjqg5YPv7OC0dDR0qzb
mF2u40Co+OIKAk4f/Hndr3BbtpZGZ/0vrq2N3cpqMbZyxirEo6iZ/nznxybe6etOCyLPVfLggZJc
b63TfdNHBeOIvafOH7vKo3zqjs6l7xYWTCQBv2ofPJ4EMsJkfx0E/GJhxBqMOkiHuVogM/QTpX65
oxK7jVV0Wm83+jEXPfbNKQNOOZP6h/MtWKg2ch0mt2iMhZjxa4pmhSebYkyA9eNrwc588uT77b7X
tWY8nuN5x2RETiMiHDynXxZ1AmJThz/Dj3d6BeWVxRL9HwmUQnlmnO01JR3QIACU1yKwIzGArR4N
jF9wPNe24jipRmlLhFE2ugr1eYM6wuTC6YjuzO0aUAUhCw/vVdJriz23r9s8lzWI2//HSqZQTbE9
uUu1PVWQjlVMiQ/2zDzZkXvBEMj7HyhjXrtM1GiP9EAkxpJUX4vp6Uv4LF0xddgZ61GoyODVU4Y1
ACkP0ogHgL0LBMqRDFwDvw5I31zuV9sLOW4u8BP2rQHsgm/YCwsliVzVJdPG7hSrADT2JE0lR+1s
bgmTSoxUNIutOdjIUFQ1auqLVsMGf81ve2+UA4deSI71S9/RSypCoVzNjO2mv4tNAgi6WHCrtbtK
xmnm5/Alat5AaD+MLmd/+z6crw/ojXQgwXuBGwj1qwfBWKhtYbcflJwQFEPdkZnIKobCNxwNqlRf
Q9FnqdOsvXRLUHXXUe2+gnbfZ+OTkoGfu2RWVaXTrBj6qsTwTkyEgCeVaFrWapnyRnn5CMmVxgbO
0fff/GuJnlzAJtoGMHKOjDbDdopOBJyxQbmoSx7H+olrLj45raNyXuTfyjI8Y5ZYH588C0QZuqK5
dMKa2Zrh0UEcsxUf4AnkVEHPvI+epOczbeYtgm42L5F2Y61fPOr8P+lK8NgxG0utQMdz52GnkAP4
UCIHTR7dA+pjEOUZN1E///FaTa2BHx5jU54AcynmbVOccNtlEl9UZd/W+HPkwdUhljIaKRaURLJQ
kZhCYWLNK3RNpXJFehaA6xbu0uNVark5/bbW0yE6o68wWyIud5xQFrcuhnNIMy+lmT4JqXv4FaIj
IFkgnHXwc5eIp3q2JVfyZkWGpDIhMbGzTBXcM6D7ic8OzMGt8SYiOPDhojthmMO/eijfYOoOhzBW
hGcyeF3zq9jFEwoFWMKJ9bPgC9VQUNeoPOtuYKhGrM85YLgNsBgn4oCtOlkGwUgElg/lBbynZf1l
BXbCaEFVW14+Ubu05imqh/Vpr/UxXEOh4vtLjpWFdTUXxpqizCJ3XzcHsxv4N+bgBXePofdhMKsz
tbdG5Q+IEWzwd3RrdNSVixw0Way1Ur7U/CPERo2vbXlzeXsdeJdIK9eloFU/608G/K1Jhw1ThXdi
znKDp5Z7O1jB2Q24qLbIGaxGf/+DUwDuBXhfCkgTjjugIdF80TyXkFuWihOuI8fjYV6WO0wGDF4u
XsRKCpwfXkJq3P+z0xTYtSxzOOoIt+KZrjBFN94mPorS5LtGRrBkE/b4EOGoe1PdhmxxClXTFX5L
DP6Sm9YMobh807aZL/TrFRCYKjz5OfpC8N6oWpW8rSaCI4f/LVvSW+sVn9mItO11yDK2FvjZY5yE
+M65Qa/AKQDJrjLFzZlh51wUxAWGWB0YCi7HUIfWdSo/8iT4E5HCM5Gl7dPrnXQVp2B5+SvU6yvE
X9SggD5SG0vAu4t4CcAvA42seCmBPFeilSmtfpHIpu/3hWz9pgptFeMRrnKNLdtYlEaqgIQmRpL9
SX82uOw90T9YBKtQ9G/kLp/bN0mSAkf14ksI5pDok9U5uszM0gOIU9NFbhQ8B2ZYvW8aODFKZvZU
M04icmIxcUocBKo40oYjySdv1nsn7M71E6lef92Ptb2P0eyxrr/tp3FpjD6vOimmmWb2p/Au9/NE
A17ykbtaSFTopnEN4w1iMCiYRvr9dqu0zpBNK80RLJTTwNjZKVlTnKb7aUK9i4/F+22HEwUbSWD9
lzaK845ugDhPclOmvlw5jn2DFAqCXvPqYPse7ejkalwBdDJDHfaaK+kVeXiNc/sZdX33VC3oOZf6
SAPf15bXKLbUPbxhjRpioVnD2GK+geher5psUVw4KAmT5hVVf/dlQQUx8voFn8TiaBnIRAQyY/BI
hldAr1+tC76gtzgqPGRilNK8ak3Sup/ZXTmjk1YgeRSG7qtYXHMUUI8iBcGN11nNAY0ZA0PqmZHS
7FKOjoqTmSkmNYpcwt8CNQ6O5TJmUeKWSedkQzbrIa4z+B6GtPxwcG2LEll57BV6X46KIiQIT43k
1FXXhfR9GpqRUTb6ARECFR0cZ34n8djmZGN3SRCMLO3YDWfNOZBcVc0Vcu04jH/366OTaGBV5c0X
x7CbZWIrU9lp3rNIaR624uQ/9xZiimMEaqsYdG5KAD9qfacirHszdmLl+h/23PZXjK1LCd7wxUZ2
lhi2xcRke4V04xZ+4vefvq0fgHJJmTDxqzXndkAAtgveRDwtJuPCS86Lyq3ccVyE7LCSBwmk3tpf
iUI9yhz8/YmkAAM/4GKHDjUFMUFNXdvmTFcvzvZxOtuQQw04mu7nD0+JO7C1YP2naHSIM3fqcM6L
FQt46JQoD8ga0ECo2Oen1b3HgOdVZhPI5RyC3UROemC0W30Bv8/IHcrVVOm18eImYU95j4rf80b5
SV8soY7KvGdrD+KcW1ZvfU+ai+0cJ4wol2rCeGHt1HRuLqbNaZkV57OdPfTLLmU7fJlgTSehBqA6
UULAy+kH3Swf1k8Xo5z0IZH03jHNP+D8qv480rYEjed35teqV4zS3PG89yWGV6hFxlk9CrcB8eql
h9uoZUYXlLl4bGsCBgsbqDuEVEmX4xg0Dws7BdlzYeNJAcOh1dpogoul/jZrq3rFQbNbihWLz7NA
qLY/XeRpWaR7Mdeo2JQ/FWxyuy7w+D5psiCaTmUpXk7NgWm+y3pTvgbnoV4bbFBJU3ss00jyk6lO
vG3QCbl85r4VOWBt7OjIrTuq0o2TyZf1x9KUaN7GhB1VaihLxMKMjodMOzpJ+33BSZrFqJ62Zdy9
R+W7ZaDb4D7VdRyKn9fCecKfi22CUljiVmsvxiv9joqrQtMYuOeR064mmB+MGZOfH65sVtljOp5c
OpHeULZ8RTQ9SYrfYtbBxUUxOgPOxRNMJVsJwJqEOr8E/5Y0gnlIU0uaaYOePbvp5+Q0emQultWq
zBi1WYqWHcwYDeNKDpQNC51lt1O9Mysd7yjeAMt0A0EGv3By4XeKFeB3YI/wVhFhB0ZschojcZKC
5uz62kM4+VWosf6kFd9gHIHUS4+pMAH6mkIqh0FjViNGLFpMJn0nJqnIDEL3REfuj15pIix1Hkr3
4KOLeNyVNf/70m8TIiecj6lw0r3fRxuCBAzbSyKqbCHPETMhYRR2SA6bepuJ9LBNqbCovTUN0Dom
c7dw9EIlK2hf1S6pWjTC0l84UQ8IkRgMovqHwra8altcWsir0D8pe4AN69NADMoVYlMiJZn/b33o
2jjV0RxYLpg1ZR6uvHndBGZgKAZmTZNH8gQN6KiiL3WyF7/gIV4OPq3vhJwu6liiWZ6KMFkkrL52
p26OxUPZ6v31HPb9yRj+3ilVpqzqB0KN3kp+2bqB9eO+Q23t32DLpEZRT3TicSGvObmSv/zw8Vo0
eOK10sZ9yjplUoMq4NiLoTbRkBQFzDhV3IsE0pxzeDvlM+VDhljHEJrUKEqJHI0TuFqss9grm7Rr
TQbxeOEbbwDBE2iQE+Z7gGAsiIVvIRgIpHUPs6OJWs4zUWu/7uRFsYDcglBAnTrOrec3BANTKq5+
t5G3CcQXfSIDrF/V8s9THk6lpm410qq0oGIwBX+8iiMgnFKdxsbq1pTvXTdOIR84U84SHzrwopxC
3JGsO2ld9PJz8h6s2/lFZSaYmgdngmyKWGVrNp9RTi7bUdIC0s+d5gFkJoxaUkCAKhQuualZwtGK
t1VmjNjLsLE6iKlKAqrmocV5v4iVfuPPXLX2HIzof5g0vihBm5Os1Mz1kVxgePNX5b/5QDM8quQy
eMmdssv15E9XW/SjVHnK3AUvAWXZ7CgOlHTIOOp8yGp/p0j7XCva3tTtswCH0i1MI1DxrfOD5aoj
ZT2CRVSzBfowtNDgW/HC9zZ+TFlkhq9SbhjnMrLbrCxPqMqSF0XiHwfRt5chCyKwwjKw025fCeLG
LXjrpgQWdampTMSnfixhG6iy5Wgh/e9pEWhZ6LlL09DIgyvYhTWQBtTbnF+YJl2ZwjYWn0Mzsxdf
oPuIgrNKHra+CJiQTRJMt0Z5xJMwIuwuKlCkZ8qUPr/6V626Y8JQy98w3ztEEhoBRqoh+/kgaQNB
J9TXmMQR4q6sRDVbkDoom61PqR20DAsNfmFIJ/pf7rRC6fL6vwJClnUZNj5+ML6C0ESZTkJdOz1+
UwGJl0vFtReU1+4b0228bwCBjDqT8g+HmShM+HsMnJbHD9THeo1yBzvWjMZ41IJjWLryeDW7nCWT
eRuw4TIg2lLbpKQNVO9P5tiF1nZgSIrzR8OOkwjw5C/otLz1KURHNc8OXY4g0UpJXCvyCNFD4PjD
lw8e1raOGHgzHfKJ4AfYQozXTTLSqhefNIvGXTvqBHzg0hLjjyRIjMA34pRQipOJ8MifbLdDHv4L
OAkwJmVQRIFsaz3JC4gxfY+c+2KI/l1r24ayhjO0DreejvzRKrVmF5JjADLHbcVavKTPthdW7AFO
FKazC3NCVvRrZ7sh7k5GDQHdSPc1LXPKvfVWsSeEEgSZ/4FH2rvhEfPPUO2MJiBZD2MJTAfLvM9O
M8nR8ohe3pFhx9SzfLlLxAzoFr9o9CtpSqrPJqiQxWsLGAwy85ZUwbeUJMkH1pOLeqxwSP7DjcED
n/nK/n4hCuIQ4w1wlEtyblsSS8AEiz5dDg7j0LE1xAnVyvirEHhTUCaTeu6rvZZIZFObORdJ4uPR
5CGxZR8BUXVMAYXBRttRUrm8VwnN2QaFOaEgKUBKZXzqTuI3h5SOIPAR2z9jUXayK4kxnubL+bMB
hBeDOSKPPWuY/ZQu6nZTAfvTmOqkgF5FuJ9scXUs6npNXiBQhX51l13zHYvBTihEX9tpqY7mJk9H
2hHrr+sO0v1TOtqOaqeM9Mnx99MxHOVQ2n4WGMcimRqcM/+TIT3OAhSNvJZUU/gnPftpBCRmWjv3
WD0urORXvy9JRCnH/7EtkUftyc3tKh0Pf9libwJTGLZluBazeBatSDeAf80S0mnj2oeZEG7/lNfR
PtMn/d0AZ1/bHNKFPFQqkdxqC4W4cm4vRNPEaUtskLvcU35T7f35Jt1G0vYq3ToFcPbchBl57Kqn
PJU4qYwpopDdPQ5BdVNXZu/S0Ca0buQB2tPdJ0ev2VdlxKZwP+Ms6cTPpco3syI5TvyAe748SJYe
I5FwMWA0sQi16pdMOlvU50f7IXdo472EhDY4p8yYQ31Gnl190OGOeKpF/OoKI2PgR9uOdF6fdgI3
a16A4duPTSI5IjrBFQiWTf5xmSLGZhCx7EMC+cKxV2vnAmaTDC04eED41acdqXluO1mQcUOGpOB/
8sLBDGKwpOAbaqiudlcj0a5ZAYnvSS3TV4ZAH7dTDjam+fK22CUMiy3nDJRbqc7X34iuX77Bnl1O
MqZnyEPyyf9BsZyGMfm7GT47WOlExwXLFbntqJd8h9aUYSHGHlWsLucyaGkdGeK2CsNwhdF0xrF9
QXQPaFTBztmG94UTeF9+zxjFMkdiYp2SZ4C+d7/b1Vx4t58gdxt0zyhOjP6W5gctp5f0GK+7H9vC
3azfGwMC8BjYy8VEnBbPS7usIIA55/s9uptKUoHuZljYrkh+AQM/ymXxGOmiUR/FNriidghgYWYT
RXSQL5lixVpwSorm8zL5+COD0oG9p3HNpmbaEkFO3XCR4HrNJ18JiDPil/fAgOlbwT/HVw67qOLo
JkkdHytFguymPD2L1ds1Zf+oC8bguHHI47Qr6Zuqp7KEDUouIeYu4INLBsS2T6SShgyZsCzeYJSj
w0S9WMQSUSVxgeWg1cKQgal2D2F50ike7RhL+9DyCg6jbqIqFyaap4EjexeVjfPjNLsTkSwBOFy7
1wrb70cUF4CktkT0NF6NX/e25uZhbKc61GdWM4DLJMpE94e1rAi0m0t+sm3Krhd/KwAUPibFZD/7
p5OjKWlY5PLVa5xM1QAorbxkYFk1CizeI/OsZpTKnIPFT3KO/jRQyv4XJNTvWrCYkb1nw+Kfpky5
287dyX1pgqIDvsYs7DFeNb9CBMm5lcTdY2iIA73PXxz8588RLwkWavGbsolVIa+aupo9FRQ7o7y6
aQsCs8xjorjV87zS1ffJX7DSr3isqI6fakqwhQSXfYRoCoZ2qbWBBgn658sBtnGb2OZhumk0LSWQ
/yA7PV9HKsj4xGorPcZT4Jm7+yUh2fsqF5qdkTGX2WfghEIvAM9jz8ENKKuhJXPfusO9jw4UGVAj
jO5lSKy9C5ARQicbb12Oeea2Yo9T+s0m+oK20NjbWt2lsZZgDqeDj5MVZ11lm/tWeDtE2c10w6ew
poFA37look/+TH40jBH3jd4Kai9mAvfHhMBVQthc6GT5/XDpYl7Iv3/Nox/D9nVmTqr2Hct2jdg/
koFcKIJMy4Qevqzw2ynwmwD79PJsT78HLgihdD+tjKDCnoMSlF7nB0Da6Ukyws3jGvW1M5HdsZN6
Nc6JI7sS38e8t3E9oAqk08uBFm7jnhtsUDR6AIvofzmlel1+SqqSAj8TfW+lA4vkkp9c3Iz6wH8z
lH0Q0hKVLxWIfsgunQm/CF3AQqcq5KwLbVjScaju2Rh2xg+AzVh4RqpquQ4OwpGO3eHtudayo7zP
TcupPoqJX9x+rRiCt83feVGq/yLVYSC6CjttBI9CltgBW5dN3OJhCHYXESrfWk2gUG1Xw6BpaH1w
KCPO4ZGGDpsYm4blW2zsJUJ57Bjnc5aZbZl4JvjWKl/4qOjT0j7kP0FomT/HTpTYPbdCOWMDVti8
HDHfPochIZW0qvHfPfYFZNwsqkHgbHtuSkcaLgMv4BnhN+RX6B0TywSJyTRWL0ZZiHUL+98M0wzW
LTxq4NFl2F6mck4Qb579vT9g7iC9l8irOsmiSJgGymdCIj3JxuI216JWW71DHRhFSM1+vuNX+wKD
v2CaUm0a0Mu26NAI2oHt+P4j5cFru+PmQFSr144DEkOeX/JityxL/hFGzr1/Ib4PG6StixB0/39T
2fP2WQqJiON2T3+q2pvGjmP+SqH6hkipOgpkOev8txjps0Aku1OTVXXzgh4fjsk3JHSwWn3+R575
7bwB19P4sYZwWxccXkm+KMqVSg1kWHBX2WMOtdCBj7GPSj1jVH+PjK/S1YFqeU1W41U862vbAFNC
yBSqdCkPSTKYITihyM6u6je1EIj/L8URO/o+SONTM6XXp/VweYgEXqYz4KjDKWGxxWXB9nYcHp/6
Kdm3r9onFleQBSaath2UKQJVRBZVY6bubIQNiruJpNJ9SHHcgy3T/61YTS8kxxDhA0DNJpr3Mcv4
tc/Aa6qADhYawrSM3u/9wq6mQEMjYT+LjLIDjl5IdUIGvyUvZylO7myyeoIsFHV7ujRVomgB/Mo8
9wlWh5N4LSIfHLwe4URQybpRPqdJ2O/jvB24M+3PtAcSdhf2vkSZFqJSWGwJd+T29+HkpkH8YZdE
N4Hh/LMxDrsQNiGKnOomC3b9aeQyf5HUOR6R5A46fj8mNdWouAh1pNz72d5XePyWDzQy6Ja0sZZB
DPrpZ2x4zKspdaYSjbsfxKwo1cwqNxqm6lCVeFsSyTqhFMY91KoBjfhtgHlebImY9RhXtn02ebaE
vTpD4s0vTwfuxMX6z7XUc8yJEIFfjhk2gufa7Nkj/Eg8PIh3fXQa6lZXbP9439yL2PNaYrjAY9rO
3vIntUZbezCbzZiAj8X5yqtvvx3+L6TA/66t4MbGmlxwehA6IwCtvX/qkztsK46Z9RWcVapq11qZ
Q64X4XIJ/rxbhWIUUCxPLCcGE4exRGfEQafmpIWLL73p8XD7MC59dEz2bc1x704H4icaInnnLwm4
Ligku9b1DN2WNvfVovgkV6UFcVUPWnV7Zu6Q6ApbkGzPze/UZhBvyXgsfKeXeBUliWrKTAJ2erLN
sIuM7V6jgd/jVENTK57/9Lg1TTXSm90khTzPTR2pTWHni16qf3JXOdpa48Ba5DSEnoTdwfrTffns
QtSJ1/UHJ0X3ryIhiSuDZmW5SY1KsF+Ncn7kUNh8mZdlVER6ArchscgQgoB+UjXCtW6jjoOEx0k2
/0zhWCfrP3XXINZ1Z7aexQSgcy83jdBgQka++Y5Tdq/RmCzhC7UXNfR010Rh0k0jbNJMRRC/zYq+
jXIOoqmLq6jfZ22wje+o1Fff4mrA7QDfCWjseHeOogLUBegZeguR3GPfTFWCdsbEQ8MsI/Bb0Vh5
Rw1fufZmCjVP4vI9vM6ll/9xhkglRWpSVsIYT8L2A0x2cmQyl3DCpCq9YP2Z42fhFhzK3UlmMz6T
oNEzVz7SWE+cqj4xYWpMhazx4WSJVEKzhvz00Ld8eNcqVl9byS1SOPkMHO/+zwaFDMOlswSGbZUS
6v7IJp0UuvfYed0TC3A8Rpf49Q412cyo02hgAA52obbNM7xDS9e5uWFk2DOXDAWoZpEPoLuNkAuP
pGYOZCg2uD02uacXtqcCeLml3016ej8EoUDvMZqvqqkm5hjZsEAi9q0mZXS8jw/iWoszC1NMxNXI
OaIUrNzBUQ1gXSTkbVPP74dpICsxUqFIRHs8vgwUPBrRh832bWHPAyZ4dU2+hC2/d+MXkWZTz7OE
YncsFGu3FD5meICKaN3BPn6i8jngdBvCacwAtvBhmGwL6GsroESr2x9vCEfLGMh4hzBePSJze41Z
zVyrlVsT/tSLIJ1TJOWR80xEPrvUnQpuQ0pfBgisYAdiyg0Nrz710IXPTHGGkagCjQdAphO/Hs7e
bjikQDQBoqrKfBDqXcusMS0Y1xtEsje584/wsM7g+A3EEAkH9w1Hjjsne9jh0q41/ssTgZBBsOG+
5PxSInaPk7Qp+nZ9i0oHm3+ScW3kYhVbYjjtLjSDPhe9IF7RgtuLL8zbYiqxAgphKrCdQD3c8RU2
VustGTyGdBJbanJMWwLtf/AjbV+HKl9pandycsGsMBu3+oRJ2Adh6dST7w/66m5Lfk+3kconwvOn
6UBYVRbpzDyEFXsnEn24WKXSh790YGFEYnEqZyU0sDG5b3Aarljg6WzZE+agLazCI2EGi6Czwy4k
To5eWCdhhasw0W6WrYT8/K1GNqbOt3Twnc7v8vpISrqyG7mj5vFNdfR2F6rdgy7Xbq+Pk6vW39Lp
SEmtRaXhd8rStKgtDjbnCYu64kADA5DjnMaoRmd2/HUxiqNRcT0rOeWMexgOyh4SeXZ63tT44Bxu
k0eMAiPE3nf9Rzq/9oLb5OWSBj9cFeluS1N6OfDGKTPWWtb1AvR/psieyHfppczMZX3EHyC6JkB5
+KfDoWBUkJUS23E8BaRuT8XJUd/MXrf8MoFjVSmJGSTtD0OaIno91km9fgZWqwEwXamDXgq6TVz9
7EpuLbH1jcOVaJUsRRuMKqRPEbCDBhO3K+2WEq6zoqzCxhGgvFL5Tj7Bdmub7RoivFWHPWzPqx6C
hHnTpVbwC4WMmgdMXp8pilPbGZT40uUriFaaumTZet3JaoIeBcCNmG0b3HfEfzNQvZTzLTowZA8k
cnH04zJJwCf1KNhVOHRohIVHtG8pvW2pbIjYVB3asntDWc0JLUjvmKZ8k5Hsa3swbrHAyFWbe0Bg
T/FyzMYJ9h6WX2oF5amEK9k6ODr0Rimq5DK6vF1AEQUMbEN8Xzns0qdfpTPQc+CVSQYyPSol/3ja
Rj04xM2sFh/kF3t+DvpPRapLRgaiA9dowQSazwBL7QSzQNXP52teukV8UxTse9BO1QKHQJu/G+kR
TM5ATNfsxb7F3+xZogw+UaAYQyhfO+HmwglyCJlrRXeXS8sKN8DmagAnNxqLvk6Uob8VK1DALNFz
HL8oQOnMcH+c5RqMCRhOFfZ68RoUfI2FKPopLUdLNF97DrM3MA6nP7U2pCCmrKlet6cvY/F9g1za
7Zfg2VqoQVYBIQll40dHqzsb+sIU1XIZrnxXI3yNP6XiWcDC1UX5e39QJhz7VJPNqSBTHyVGG+lQ
f46JoXM4u00fzMU6Asa5dqXUIQuUaza3EynTBIl+izDOsqNu0A1g/wwLQtD7dHF/oVPj6GkR6xNx
ff+S4cZKXemVR+7XZx6X2GUOWhRFxHnl8PtTLUj4eWdC2bBWIBPOUAy8XLRfbSbs11szmFld4otw
nSYXYccqKT0jq0APW86tAnpgVz02Zmrgx7l8jmS8QUdyF+P6jY09Qb5193sHfWc183BGdYFKOX24
yf2q4+BIgILYQ5B92+fqA3ibhx3e1SvoTxswaI7+qp2dwJdqj5Be45VLRO6qZsCDY3VC1lnM7hyL
Q5Mz0L4dSDKtibIdKzevveYQK6yYqbopP9LJ3S+1g86COhKwUtTmbO9rO8d/R7uRUxnwDEPubJcg
SvrUtGrB2Fw3MG+627hfDzN6NV/c2DZRo5mEApmQyeWxo6em1FAmDIuvtuAzjYut55/VRg1iy86X
uejd9uYFa3hVeDpMjdrXE02i65FpAWR/O05unmA/qQIt+2N/phe6dbKm9KsCud+jEEI2JfEUkFa0
G7kDLyuO7VNCUALSWcS96hWZXn5IzN5Tkvl53RRliH0BgsH7yPButL1GytvJtZsn1r2zUHXpDiLc
QuN7em5gltFa04SIYN5oXkJDXmAa0k94r8FJCBqbl/38kwGbZemXPju62v1EghZ80Qa5BWkWP/KB
Xjpa+E0yRjGG3Bl5Xn/bZnrnxxFDXp7UmyCcfwnMikF79w5fKef3sz9ZqJAvAgpjv1ihs411d/30
LsLS8dpPwd3YbnI6MKJev00rJOkCZPom4ZIJeXg8EotpQHGSjYH3v6NxF0qJN/7jHiMa8vArnrJP
vofqm2vHBaSpczIsqVbF3mhMVbgaRX6x1/VWLO1YtvQ3CyfhiMSobT8uqLgpbH/zGIIeDHHlXgHQ
QsdAhgbWMnS7RRBnS7RBLPP791Zri4VYw4ymrOCx+10xH9V4OqHlYO5Jwr3+7f7ojHrmlJ7Fhu+l
M6CeSwmPktn2TbnFVnj1vlNi3o8WZxiNtWuM9b+x3qMFUZNKoeFwioRDJp9a2j5AIZbIFoqH2dS8
q0SM/V+3EzTArRv4aZfhydWNOb0HQ8VwNkKnsZAmFR/DUf5OnziTr5GExVuuvwuftPcmM42i0SCe
UoFSQdVW6dBeP+MGw2k1cTnfagIhPSH9S5kVfC+n/xvXbb0LLQpETMQ+T3RDQ0JUrYsntKImQzfN
qxCWf2zq0pAnzW4ktLSKv/DygJf/l8mhx7e2dXJQs6P3RRq7EAiJqm+Lwpp4cvfROnhn1FhoP+ht
7pMhVLgYGbb0cdA7kZu9nsrqbIEE0TWJg54Kln1tQwJgHvRBavVRAPUOdJFL94wxk/rn/fKvJHNu
utW03edZdDIMEcOcpkSBY3JOctx4HD9eUs3TqN/4/TcXGG7oVGUFXBe/yGq/Uk7rwr+hmuXlsoJZ
DQ/awzFCrVGxoTEPSkNDqG7gXH3P4bWtUDvNqvpgbThvR222AkY9AxQmmZ7YnagugK6l1ux6xj42
WzlVivC5l9X+Ik9CvZrnw534W6xAZjyX13qTYRYlWrRK0wtKeaj/BZDohR1/mTNzWUKl9hJFodS+
WndOHkjlutOWVyKPay98RFHAosQBZ/72gYeJK+n2dVhUbIkFX7nMTDGRHQYDOm6ud3T0UaL/6Nc8
pahMVww2+YIbnep9OogI63EgJH76lY/TrD+MdUxgtXPTLeePlke77sVgy/Tmqddf9BygQJT/mgsu
sT6SraoHaT+pRDxxIdHGOL/BuXfRbVxToHVGhtU8Epmo1vJ09QlMBZhhtNEx8oL/miIp4e6UZ22a
0xRhcEQYYsf5tYNmp0sEfKJktqH6h0iyT1MWj8f8Y2Lfi5r5X0/u8hRIlI2bFoMI14J/6afsBuVI
LQp1GUojsowDyF8MrqmNGnV8o3eTqkwllbIlFZQTn0eWkYSm2YGqACMLTFJAAIeWOoYqklwc4xB1
Jrgp1pXQ4WEMh/a9AJRuDeIwZxSb1uxEKs4IWNRlMbSZ0C6N/VjxOZGElaWFKgKxPGStZbzBucRw
nlaRMl60L3PgnDCzx43zWgmI2AAb6lqccSsXACWHbh3ksdh35UXJUK0+FTqNrGMIYvayJIN4pyK2
PkBMDxQmNQTXbrIx7Za65JKtq59FTpoGY50VvQnKb70YQkqLiPFPNsAtoO0KI+5y8VDvMqqfKOxU
qkP9ugceKno5Ne9L0Gp/blrCXyevzdzGMEfxqz1TohEiFCGZ2aEnkHoZlCqcmN6aaQdV8zaIrVUd
LL/S3r63Df6QohqVU/GJSxPAT5fZ+CNJZ7aSVLwUrhZZXl0ZoJqP/b0kmqlJY0JlOMecZea+rLlz
HoQGkARjbVZK3aG4OUYCK1vTgBV8BdWksZuha3//KyOxXJFC1rJYDzC1PI9k4lPtrRe7oudsyQVg
pdwaXuTFawm487zLweHCCg2z9Xxc2Ji//3llzJ7r5Y9Y0sQWFViOzHYAtz5idBtLys+NiG7ATBx+
hMbqWqdm4lA3PqbnoZRE0iEnTLA+eZW5z8DCcNIUOZq9UlQVLQBU1WvecVEIUNiMv45aykpd9hGB
0otMeC0IA9jZnbrRxGtNQsVYGQqWU/Cbq7jjWDj+GtrlWY8eVIwmpZL8oxYKpPKWXFqVvhM2deRc
DbJoTMgRMnj859cVKEprKn/s/qcQIVrtCphsHAB9cmDWm1uGviNGcoVbMfoK9No6xStESqb2dwTx
UeNmxBjup+uh4c4zZp8DGWkxlfDAOsBJHp+TrfhY/6sL9sPd7Y+/6+aMgNX9yNRR8X5Hx488BTSz
j+tf/+cLCpjH8oJWzayBBHOYO22z9L6NaZgk58WMzxHaDZ3FScSsex+7zUFDGzkLrNnd71o44CPe
TEwUTBkz/3piLFBNIcuBoGUwAc861hqZyCU7+yAyap/FM32TDB1f9fzaMAJke8/N6/J1lBCrxAyG
7QOlSfJPoshty5nznnhSn868BbO/ZhUeZV9P7XZYHSzpLuaqpmesnx5+Z6ezoh6JgiOvtVWn72/d
dY30bL5TZtUS+4DBglPm0xoAuEvMQ+sUYL6lakyq1jaGhn035D52azqbPJh6qMpQ1/i9OhyLMAPr
vuvtBuaaU2OrOXx3CVHU0XXHnSNx/H/ZqRU7iSNb/CqwhX7FRrIPI5ESejIE/fusvEnCh+cPPh4U
f81esmEoH0zounqSkZ20DkaaXiYKGY7n/BHM2BWTZ1x5wHrmahIwbEI3+bc3GA6sIiMFQXBgYOdg
zi4j5WzvWq54pTvQs9WfaidklOe1JaOU/R9TlwS6HWAK2kGBv/csA5v7xy9Wo/X/Mx8bvT7H+uTo
8IHghpYMmHfxPwLbP7ltKE57CXv48IDUVwcg5Ww6lJe1ByKkHrth9OM3bRPd28jc1dpehR+dfX5W
XytzQC5k5hvS8KLje8EYuZykhFig6gdMNkR30RC2RbUs5EaSG7Y1BewdUnp5FoidO7PBCsyIio2j
M5FhCj4HPxDD0EkLy0dCC/nmZkMXbQJkFGV5/wPp+qGmEXBTjiglF8ZIFpAI0kHDl2Z5RhTXZC4E
LyIqhMf8JMlKfzh640iWzkI8o3VB3XB8oslGzaR4jEjS/yUJrrbfi4LeacJLeSfg3p4HAGXfMERv
DxiisGRNdrZncZ0vcaCXlSMKZ+5JEYXK6SWh4645Jq011+ZLnGE9dVUKjgtT1Xz+fTJdEo59rvnM
+X1UkGMqBxzB8Lhwy+FKPu2KFNgITtpXNhhgPF/IT794lmwyI1kLGgHRGVh88L6kRZ53UzZreur6
KBX1rIIjhVbL4LDy7U9D59sw1EzsU/c0eYWi7s8fHDb2LW1wv63DpDYK74WtQZneHITLr/0rYs24
Xd80/ZAzdAlyWfTQcXX4GDRtiFKGLufuqYdZbu6Au3AjTE9Pblj1J3K1vmPVgoH8oyr95JOU4QIe
sfm6Sx5nTKjZlWNHq+a5rNP99Uj+YR9jIg8f3udKSRrHhc0UiLKiscTSWapqowwK9kL8Aan8qS6t
4AQvervIcsIYtqzcM7K0bKD2SPfDxULkgTlZiTMuUeYHElg/DwGxpIhTKG2mQxxgIsDBVPYHUdFZ
gU7CqcVgbQukh16gLh10E1RinFGwZglL2w5xjFWUz5QrqfMvYewhBegw5oDX/lVuegS1nBsWR9se
7Qb6Qjn2SFQ+we6+WjCBFm9tKJPh4EhcoD+xCnRaASsxVm5YoAAeL4a89VwyeLlsAzRRkEvHcvLP
tj2HY0n7bxENmoOR8RjugXb44X/J9iqDPJF675mLpXq/Gxjx7vQA6ENBuSht1lmUq8vH1fYexuJZ
3ukQziNUXwQ6X7sFzHvjnA/0oXIYlVZFlzaI6fFIhKPOsEBJxdIitFMurt/RI09PaFZRRbHgN0W7
doSZtPeKpJHwWD0redJj37PYg1QwP1YvRU/YkBcVeXk27uyzopmHzi7VSYmo7hpTNUxlxcnVDa+F
JmyzWck1yQ1w6kAEo5A/dGrIGE5kw9hMF4nnrtKepy4tfEaLSrO4n8Dbnjn6T5t59zi1Ml+Djdv/
AcSrs9M6P3CdQO1CSzRxID+AnWkcN6TPEOhDHlq1Qtl7ES15eqTA3AgPUP22Q/2nQj/eSJlna5TF
5ovlBTCpGf/AAIMWDq555lUD0Ez1m1vBXiw4UXECSPP4WJSQ+j7+hq2XWGAYktt4Qu8EBSzfMKUq
ivmmU+Wp5MG51I8QMbcAgUZWvsuXB/WvLsBxDz9rcszNWD+EAGFPfQneMlibg0sYWrwi2rLWINDZ
olLpu9LrzdtnyVyfRMlJqDGw7jUuObKkzNKZzq+O6ekp6lf3gwmzgUkEJp8V9FOg0am7on68J1Yq
A7b96Uh834qtbrbCL1EXGrMB6k9noEy2+Zu7Xw7B5f5p9dd4rox4hvOUvY3L2g5WAndE2OCQQ2HA
jVli+g6FYs7ax93qbyuz+3J1B0W9tNwLWGKFn2RlAUbodFgVnjVrogGYqqKzOWpuOxSvCN5dxy/3
kcdwCdLeepLgeQ7q7QUQdm4/uNak0GaZPfoMKufYA05XMR3AdCZ1ss9c9l7KuPL4cmBpBr9ep8+E
IJ14XbuUyWupPMe2zByxSwFfgq9oYyTa+g3JGMWaRfGXpeaABTmNPuiNdVk1m2hiPGO/mzVvYFil
xSawCAjhiq+8P39h6XM1EviWAOJTBgh3TRwTvV74mbNorwcz64Y1DPnxtBj5CbgDf50QKb6SJJjt
d8xjP9Y6BTvp/QO5ot1CIF2VVSeWrqpAvocmu7skZQD2JYFY+y6acAVc3z0up8Art1dgI+r96oer
5cn8qs5WE1N4pUoDF8tjMQtEbVudifk3NF1wI/rFFpQQkVsL/syo2smbjznqhyVLZcdQZ3kFUv+u
XpCdyZ25hg8wllVmWlikuMvViw+IUq/ijN+0+kWuJFze6OyRusUm9lsSvUzu4inaq6pXn9EQ6ROn
guN8Deyi3A2rECqnX0b3q/g27JiOiLCa0catwT6OEx/jomIxKKFpxfnIVnJCk1oD1W2/EJpLUiW6
W2GU+TYDmIY6GxKCJ+jLcT5tQ2Uk7T49xrypdNJk6p+H0bzkPNnrhpujeuaBIOAoMe8KUHIJuKxq
ybr88JwyUhRqm1n7yOE8z65A8o0klPeh8gvzNxSp11dcklRILpl6D1kmDWUqeYQ4/9dCQkVsu1YX
AnCNiqO2IbXOu0a+W9DxV62HJLhX+EjKMZuxPLjwa7wcZ6slEI4ebWvvxLO3z7+OIO8VqV0h07n0
fQu9XsDdwUqt5bYd+L8cY8NTNAtWTcuRmyDPmVF4hAHBASj6dKY8znWP3h1yAe/3yeIIWu1kOyli
QErgmv2FgcY8d2Wxk5pqUVyFu7h3y8EszBw2TC3MQp3m1HJJjgt6nRZQt6cNB19/HQQaCzpD/Y6M
7zkjKN/x+rkhsnvzaL8Hb8k0kH0ybMvRxKHDSwkAs4jaKU3B55XsWm4ObcVMoDbyPaX9vaLyJ/hn
aMZEWlpwyVK3plAcBLTtCMJDz+88wtkOSyyallZnSkb0WCEmihrpBJg/MwAp5eVsc3Y4kueif4P7
ERFdiBLIi4w6ou6yJZmcCpm1vpJd96Q1+lOh/FIB1Tak66X43bQAxsSug0qVhWHPwlow+/uSFh+c
ny+kfCzpczqDG08aHjY80ndmR9x8zEh6nDYO46RDS8I5t3Jxyqw7db9/3kcD9F5cWABf0jr0UYle
y50vMfjYWshXAkJj/VhsoCGn+F81oqQtq/1PTPFhBAMaVuWeaSmenP5JdEkLLcQe6wVIAW67QO+i
U/CDEttPu4dUa0T+7Ipf3TtAPoa2zKuZ4EluRM8pWwT1SwWGwO9d0NQcNXdmcFcEqWda43pyOG7j
/AcWrrbc7Ac/F+112cIrgUE3jNaf2M5eraOhp/KVUnSZMXXsOZ1F+uMshH/WXq2x5Jw+Rb417iQT
TXUhfSy8/pzdejnayA5EHVU1WIC2qH8MFxjAjuVVFizuTa/xxVSumIFFGUT+TOnSmnCOLxqPtBGq
8nKJG9aPaWjedKnyMp+3ce9uJTZKPhlNDWWQkIval2X4Ui4FMGJOvQhtuxObh0vdf2XlOCsvZv82
wmMfsTJhGT9u1afu/BtO3vBWjtZ+ihE8grT+KZ4DrnP/vja1yA+2GoMtHFTQZQnqIqQ7P5Gmkysi
2549TBOep5kdD3lG9oV0aMVzQofKiXogaiUsO6JjHKMYfBikmEsKW8J5c0/oTMcWRpzhm7p4OQ+X
jU/v6TsDXOrUK3RUYy9+dE51MyFxkThZDU2YAsOGn3lk8N9vcXmQP1H5dCZXMiRgJd+1TTNFqvD7
uVZ+Dg9l3CFLkXMH8iMzGfYylWOz0FtXO42/U9g+VYcMHSZ9fK5i1fiRXmfhImcdmiQSDh+g9h8A
NSXZhnCHESwvi7KRETapsC6o9ciJ+CngtjvgTXWvbNPptcNcKGsk0IFSd0k/y3e5sg/zRcS9SHWM
mhKrMweE3bSOqGKYaEKmSXOEy8UDx/HqHs+sy5iX0bzFThoDyl2LfFTDHRCNcw4jR2MpeArEMNdZ
9vKKP3ehu9yftWkM0eJIr/JPp0Z7Se8TzqIl4cQLcJeDCefgD7/qLCn3kYICt6UulQk4jKT8Uvpj
8okE62HGmhZsEF/ajNIX9r2KoF0ghXr5TTnIiLtPQG58PC3vOoin6y3hc2KGVQolupy7K0O/GQVl
R2CzDeysbAgNXfGptwC8OrP2YrUABre7h/RJJLaEAXvoTzjhvcXuIzo1hLtz4E0XVNGOxL8kmb1j
CzSdgqeYgY6BIHIgNBGfvipTvtaOYis5lKX31c4O4yKhaHAmO7/PFNhaDDzk9cx8iAgZDQHNkStc
9Zwoc0FoZ1InYh+G38Jg0JtaGdWO8CxaGbccK3iKNy/hL0914SotKNRQsrLkXW/RIPp4lDZIw+Zj
UWHxWJ40byf96pDbuHaseiVpgMD+fxF//AdTasNmNHexFLuggcuDv5uw7dUTK+JgFBbQVqv4ufy8
2zGX9Xnq4HbMX9UszeB2XDv9IQoVlCGNIE0GztUNnhQAiEERr9rf/AF8jaAbZACj/M25jgArDYwK
XAFvmv1yAlVr7nF7ZZq8gOI8um1yhacY7VV26KPS6NI1GyifQofcs7k3tbAcQV5/TYsSNyKsIB6/
ZMe86oXA+5Bn9/bomvf4zbRCdfYURaOV4K8Rxfj6TRXUMqrqzMj+JuyjSdnq0N5pjUYK9R1vx3eU
YEwwOFjYSLENs4R9LPGOzxTiyh4qgD98etw4e0zIHvTAH1DqcKtIq9FXoTSZUdnJnrRnALGumlRr
NjZ2MMscoz6UXLP2Ikewls0R/Fa9N7nEzH5QZcOfwLGkjdeG7gR8yZB/2zR1y6CTLka5+z/WdUO+
PIb3Jk7xqHUF0BQpRBw14VkadT1SSNnxqTGwhTNYab+KkIkFXK+3HsqzMssoDDjoRvguRVh+QAFd
mKkI0Z9l/dW/ISFCZbCReRtwclJEE1BhBY4SHfz08inJMzqpQ4wUHqfhGq9LvryRrgmHK+vqv8Uk
jL2dwKYePWTG7Q1fvsnU9Ede5CfRivz01vV3oHxdi3/3DyrAvoYZ5rY9BgeEeaZmG2v9RBsrkifn
azhcobOXuj3hI/XUts7MZjEkTGRWZyLEpF3Z9+q8DvZwIQkZu0h2vWKruDUgiIgEbj1XeCa8e9dn
3ZuL5cQVE3ETP9wBmwNzPQKmGK5PXs36UBYy3p9fPDJ/+7nEccCZ3Cb9yg6D1bBfu8qk9qcmV00v
18BJ8p7QiHSnWt5G1RsMFkbmoFtTH2Ag/rxp8d53W1g4/1SHyvwN5htEOhS0qG9+NdsRcMxHvKsP
wO0CQ0ED44WE7Fr50oM67oAQZPRWEhpHmz2EEGeR9CgITum3lNK4gOp1xIfHdeFDsZ/oHeb4Ynko
sxQsvqAeWYcZOoOpuKZPSZgozfRewdlnRz7HskEln6i6sVeCLlm6gEQ8++lAsc9ZnM8GXvJF7Yc2
VqrhcfwcQPz2sNm0ppchjdTpjXUBs38NMee8eaxGYYTVTJFy4Rqbg1u7Mh57YTbB8LSlWAecZIPs
MWDMIsv+lOUjEiIEuicb4qshV0wK2k9I4swWx45+t72QvMUKCfN8hxIJB9VcVF8eWdN1/zjpN+0S
u6hWRjqsPwpf2brFxwh6ScjsBNJkYAHiyJVcpLFncz4VYrE+fBSeROd5g+BGdv+Zqh5iM8qoIEcC
wys8/2evWCeVTH4f/cT2EA+OjPeO5R8c1+6tGyxHBgqR3TkZ7FiGXrAXK8/MFKmByeKAl4TFyk/O
B05ml+wpc3bRSVAXQAMZjPaTW7GxjbGeEvFDeeubZHTjBky+vbgBKMiU5lEC4RQuZGVE1xTCQS1i
ivwPt5h0IhcGm2bYgJIn6OXFS5PIg6vsAxjj0w0Z9dIQUkv33HYVX8fKJ3HjmY/NrOnEsGA4Nynh
J0t07ug65qLs/flstBLMDSLZraAs+bgqIlfLisRJNb8aTB3kqLbLnjH6FwB4Imj0LnweeZN8JXm6
71pLau/rP6CmG81Ol77NKOaDCvNBu6WKNPIbH4yuZfd03h88155JfAvqn+ycuJIDPvJW3zU4GxpT
DMfh+lPlYn4cDHB7mC25jvIifdQ19JaHRYRHnCS+6VffqIjP+rRs2HQGYEKLLhGzEWlCFju8cK5R
Wl5077Jzg9csRUdE+8Foy3SWeA1ZoRZI5bDqFsYCO+U0B71uEfQYmVW7qXlGO3LWKgP6Bs6T/Go8
O0RSy8T78iCztBgSE+BgejoEKZFeu6LN5IQoUo9Ub1dbmQEWah8DYSUeK7J3+kAEd/OSLFRR+AuK
S02SNIE0nQQqZKaG5L6TnOOjBD5WqYnpvnSF3ZZ0Yktcvi4m8yhDq9ZRFocDzk+8ZG5Jq694mrgM
iB6JU5CNCZE1sCyTNQXn6R/4h4KFkhUykEdUutXlaouJOZ1lWZgOC+B0G9YwuLeOlE0rMsBMN6Br
TnPRMFw8zap2m/B0qN93PPooHJHuIl29/F9S75DF5g0x+C12bTihytxmyMwiCkxFqgil1v2HALJf
zttFvoNa0HgXBo2mQxWQ9OPb9W7lO0UrdgQbf7VQCRWYfAca4ts5qW9MBJXqyQv71arf7RWwZjaZ
U+pMW/L+J1voi5yZNfdi1+B2S+OYezy2ay3E3w+r2nZfpXfmq9rP7hB4QHhfQcSMkMZ6wnuLLlho
hQB40xKRNL1aI8UTpkpQhYfT/XOS9c/X+Q1/ymOhAD62PhzC5YJkjQBECCpklXGX3CE85F16SWy+
7iULXBWAM/wkMLzLHh+VRDmNMbGwLO4z1Pn6UTUaD09trn3YzLBKpKK1+akJDo8oF+j0F/9oo3bq
rlSavp5QXVGj3O4g7Hru/VhWwzqbDVhkIPayHUqE7OQ7M4k2Ene3pUNYoQKSvy0HJ8UTTWbPvT1d
G76HYj78gdM81RyPuCX8O2GllaRuKgTe9mUn072QbZxhryNlsf4Q6T0evggBzW3IIbuso3Icd8Wc
kGpYuBmkB3k4lTTa6bhHFcNH0+8FGFXRl2UjyYfZujO/ZjbTWXSuKUXJ5uXuGYP7gcODOFHtMu0J
jgrQtMnCQZIqEh0gNG7jyJGADiIbJ491Pl4lRH9y1rkD8VjM7fFF8t3lfI6u2x5OMMhfcQIpJMic
AKLLdg3VGXIjen3AYafCrQOH73skqduhbltO8L9qPpw8qnL7w8bWxxPaMrKANOPDgcvW9B8heHIe
ulfWlNplauUFaMsSbRuRx6V6H9LNdOZ9HB4stSbad3Sd0uBAoPJDQlQkck0+3kX1isDmp6vTzERR
bC0MV4Zyt0ES6HSLOwbvc9MnTaUIn4BSvQBepuwaQG+DQsBo1c+SnqSWBQ87aLFkXpXN0hX6CIM4
+gXot7AhqNMuZ10RcY2GjUUvsHRp3UY03D64d3kcpAc7nEBkoDOgiDSB5+GPN22OHK6MQZY2dbFV
s2YvrIkIp+IRLOmcYkM0CbLDz929sOpOFILUyksFP4N/AazEd31+tpCrLxeXdLx5DvNUDTmdrTW7
jCPIroo2+5K/QMiRL8osj+Z/YWmc96O1hqqmI3ldVLm2QpXcitviJUKQJJkF25rBdmjDf9l2pgaD
xXnHj4YBxGiuSgFh8P+mXJKVL5Z6hYK36a69WXkjGTxuyY9UUTE2uIJK+qGCie1BzcQ7I6V7Gk5c
i6O2a+8jIFME3ZXE2Lokf5DgrSNkzJ2fKHz90B3s+854jFrDuAvFsKWiNXg55ZyYiTwh1L2wVeYQ
J2MTMvAJK/ybRsI9B2qnrT6vPU+6F2uWaa3H5bx5dNQdcb4Op0mrWbEw7jGow+UhGZx1qn1eyOLw
blrZY130Dxf/TyM77oyZqOpjHdtvzGx1aThyhYdVrCQt3ZvqfDn4C+vx+2RV26evLhjVZZsGBfR9
pIpCwUk/NzyqbAmynglmfJOoNo8JXm0f/M7bvY/x8QtlUb9q9kgc8hqr96hNE8cuVMZnZa8vClC7
BOV9M6YEsgcg0kz1t3aXUYWVcI7HKgzEQmEBHR89o77eEPPjAvDMi+0UzuvSKZLxCI9VKPItzWsl
VNaubb8ThzDjgBp1yD9ChAlleJob2lFY14musl9fidfHLNSXppHIyqdyycgJ5D1wMzs/ZctwS9/P
1P2c8q3kHNeaW30iFHiV5GqzcIBkXGW5Fl4j2g3ld0N8AYzanXvQ9FU5OPNPzosynnU/554TG+E8
JTHqlvlxx7shsdaGo8GhjG5UvTN4l5JWfu+XY/VexYZ8IzRITMjXyYlqKDhjN63RWoXkuXNFMZ95
+5+QQRAWHwCBYRRh+HnqRIBa8Q4a55tlZOc2yCugq341iluInGOjmpk2G6Lnte1IAzHTB5cD1sIL
HZDicmROyVb4tSjdWNlMsUGz38N5f+K95THjlJJ25Gk9LjxeQ+ChF8btkv5u+hSoptH1uxs2DLaf
T9f89vhLkR+dls9scP6l5vG90BN68ze5c7xDRE1fvoO1YwP3s869axI+qjUvXY17Ey2EHw2WKs+r
/zmGq6hqbtpYIw7xH2MTT2Vb5Kqx1026Fej+C0fLot3lQf8rHMCgHTB6ULdnXhRS+fIE2LvhH1a2
srp/IxtNKa70ReEMtW02GmocX2II9m51o25y/M1mNLtIY25+wNVqJQVtLHnB3pEYgnJqrHPOooyv
kn5hZgQI5xaXKiKI8QqMB3yXq61vFfb94AoQwL0ECN4eEgTBx5Lrj762rLYRd4XpJvY/x6whwVtm
9HXrVefodgKubAxmzxy6OLoau7TCnWjR8XL7yq9luMyPk5OhsRR6jSNZUZT8/4n+1FIJMl0d5l1q
RXaMlYiG8x4LIUvJ5a3OzMZxMvxd1Gk555S8rTEGQm+BVVJvL6fPykPNupTxPXtrxiYi2cJ0j8/z
8bYTyZh2GexWXo6En1HaDc0lDhJJZ3tAu45+BWAIc/jg6D8SPW+iJku/4w58iDCZFsl4Gm8rAwnj
y0ZurixsCPB/wL0FQTY8jnUN2tqbEd/xvO4dgGQoOWruy49Y1FKMneyZdpUxW1X+zDSsntaAkhxS
ntCIRyVwEYWSdsmH1KYBOOVCin0XT+9sg3LTkLNpl2gQhVU8Qf5eJSvp/87DfVQtGzlUqY1l72hG
04nwxHF08U8n36u883b7iJdKvHm5oWE5skJXJ2Zkif9YidC8PH03vVqPWs+F2INXHYDG20ZcJpYj
3ERcBY3R07Isp7puJp5K/3bJBSOCPEtA4Cuc6g4G0VsiZRORixJRxmMTuN9AyqiVl+j1m7PM4y0R
OwAyFZAwWPeUhCrM4aKXCbmRkdxX4V5XNiKlkXaZs1iFrBIui4BGIBho/oUL1onbkI426OZNldbO
3nTh7R/N1buT6g/8QuNjY57YJU58UJVe73ThobwQWie1s+KyMij6HZrhZV7yzXUQQ0EiVIyjlY1X
mfl1wpGa/59xS8m8TXtW8O/xWvg4SHNyirxY+L2MmkNMV8/fk+HdO70sOIGfoz9/qCc3/CSahYQw
G5iLv7Hc9F6MaMQzwzJ7ziGbqmQJ2V13AceL00ODS8Mb3T5c7oxv9GMTEm4WM7aHmpPjPDi7eMF6
WYgfuTXUOXJYzHcZh0i7+VgSFpbMv45jFBOSfOCS88uroEkvjCAaPEjmA1SkgqDNcshLTYeIa2gz
/yQLnBzqEQDMjAVlPTviAn9t93Hq040qbL5Hwoe+CPTID16f7ZaqlUm5hHDkgpVO4m35bbWJ5A2g
FhcY08pCBpZnYikpsiO9c9gsic+sxzdBAZgJ7KPUkqJWUuDvEQoxbhw81/XaXKgNJVssTpv18bP0
VXbddMKpvbZWqrmDnIeAk29NPOAxt3J9k3XnzpflZ1Hgdhu7OW5fwv4hkKeTMJtSdyYq37v9IG1J
4PSW3DDpMHlhdNZ8tEM2EYDJ1fTaqewHqbUdSQYI3rUMwtbcdZXmDbHcLOTLKcRitCm+RtBT4Opj
4/GdnWiWJeOTpJ+4blqM+NwO/o2GoOHdkft/bbWEJk/XP5yyBVXYCezM65r7RlXhgJC1NBu45+KD
MP+557D6ArGE1Lcg+ocPuq9HwFQgCdfAshBozE5PRXF+TOxVy0dllMwn0RMOcUJfAuC7M3Bb0fI3
tSl4K4tb+48wEkpIKtDTICnNj65gkjw6VhdryIX243WNOBkrvmNH8ctF6k3HeE/EXasKgzoDb1D1
CgNjX4Ocj4BadU3rzY6mOTHXL+k45Ts+dbl5f9vQ4rKAq6Gxe+jiLBuWsLjoSVIYt5mJLJggF2Ce
SJ1x2CEPqA1tbexBW4Yd94ShYWVDoJTK1ayC74R1GFhAVrG/H1Tyffw8VcBszO/ZWUHCvUebOR5+
ESREh7PwLpEzNYQO/ZDc5VBPNfXI4FfFa92tjkwK0kwOCVdosc7zCIa0ciJVRWzD+ijmZmP1rasI
VKYWHiKyNCrJqRblEIu/LY4WaiOZe8T1+5puKDBk5HyUitXyVN65avEfXt7UYu91OEkA90FakNp0
5lC50mg/GTm8k87gGgkn/VKxNVyhvgqywsRFv+QueeeCNA3w3eNV5raeQCC/MAvJoVieH2rpgRXR
/zNLUtIudKVUXMeNsL8lyTAAprMRrHL+kgfVlELWTomKkhwAvkReHwoLnkEAVX0l7iq5gysCQcaL
f/Y6lF6mH7uHVUncjrDJQtpD+ZtqfhbjLM/LSXv8FP8cKkL/6k3lRKAO7XVvH2Tw7JukEYgcTMX/
65NMbxCG7j7dL/tPqOtLjBDOTEUb2C5rXpUdZGa95E1+AqVgE899/p7DHoxnRuL6HrI6RL+a5ip4
R/2VvhwV4X/POcuHXOQlP69gjOhD05ZgiYKPH5YoXMozulAGEmBWiVV5j3B3D2mGVgNBUxhzsWwT
eFJJU10Hi388o0Su5kK3hcMvo7qTrcpd5yeVBqaXq8YWlWI4Mz5voDd8uAsMjVMTiW/1wg+cOSj4
FfHv+ShmE7tdiT3wy9DkZPMZM7X7cUaW1/QPZKLWGOTR5AIs+ncRYG7MmoDrZcLHl/tpSd7w3H5D
Oh2wo+8CpVwawNMVBI63ig4/Rv/H5/bhFa106WHOUe2kbxT+TV00dYRGLONplefc7sVsbBK+BeQt
DcXAOywh8KVUzKs2R79xxDosAins3fsF4N2twPui4F2vUR2YxdgUyTcT5SLuHA6/6TgZB6n9jYA4
xQH5OQ+VIJPwBsPBlwe4FOkqtlIbwv8Tsyo10KI8LXsk6laiA4NfuZVFZgpXv3a8j2/w2rXRcXrM
u55xeAX4Lu2gmECFiacN8Daf/zq4tDYtkX/0UjE9HWSJBN/xLAWE5sfpebN/RENuJUJD4sbgXd2m
j1LDi+N9oz88y9B27nxyvvYcpSWoIi7gQGMO2QzHK5yPcHXqjoN9+jPFLZJqGs03D+UWk0E5Cx/1
DoFZHf1IRiuMYSYKkZXx1YIuM78/JC9JkCF/ex/GRnwCX5MihyhyPWhrJNVC4kRNNAGZwt1cUnS7
DSgx21UekupcbJDiYPUjuLYMjG1kSdlYZotmLbs8d+nIzqaZ4lAICaAiMOxvPRr30j3IrJZe5ked
vI9DzSLT00gyvX+6Ph8KgJiBoXEdX5eNDTofHZ/NuVYAEt6DX08int7B2sVgLV9uu3Ap/pWpes2a
k0S7uYH9o6sAUyKCQIuAPBPGGpQSUDUQBbO4swdPZBA7N2EeGgPNOquXhh+Jpj5pgwfKx986A5o0
LI0sJC88AgxMbwHsNXTJUexBQXP+6TrXDTcdQmFSftRJABsAzQeRUss9Y14DJUrpMPZmVhfJMp9n
4QRQP5Nml6EKrB2FxPgniQPyJteSF+6rqJa4ECtr4osW3VPC+pb1c9jII7yuxvSTQEJrkA/32hOB
ZPVTxxQunMSI9FMoGP1mmelOGJ3NlIRFaiQvGYOzhj/Gy+MGLhXBRQ9TOQLM8S8ohyWOgcclfciR
vT+htwbz/Vd/rpdqz39S4OpvI1wQEr/nYRHj+CYsjjPxHglM8HgcW/oHvstXtQzuVWjVP8cJl3Ps
akIF2sWUoVPsbsA4XAPlyYvBtYlS5Lh7FliCIDPc4XFt9PHCvJ1+AgRYWzG/pz+TBYUoaa5AkVKf
YjANDpQyv7Vs7oYwknnqckHdwB3jH+KkYNK9BAhWAzcqc8hp0hJ94NTS0+MLMqcOA2SWiOnLZEJH
F5a/TvVYGaawi2rz8au6R21nsh/pi7fhNm1q6MIQWle0kj8DmG8wLBEf35X+gHVkJgDwnc5+Yqck
f+G8avVf1MLEithz9XE0kX9YSfSO/hAyx41M3ZjQzx6opuCjJSUuKL54srb1YZPXJLvlejG9D8s8
Lgfw3TBwLliZUOBb0f3tmrm+3+p7KQah1UFxjd2YdNN8/cWxOfbZChO1VOfUA13abysh0nin4uAb
qwTbL3bfBj4qV3TXrPiqvMl6vNVreXLLi+KaifjxCqi6kusgzELhwRTW7jNJ/Lj5oUYaa7RfdPye
22AJMj/wjPQ/cPFcf+Fy5MgVCHPP6vrhQ5JaPzQ1QWWGfzQoxczvbyj9ZF5tFgtb6QomUivyjm2Q
cquyyvqmNGAubeIDY9GUlNS5FOz8yZZlj/BivOSwMwQAcSGb31RWQEXWLc4dFiTJ2H+Mu+XBRHIv
4wVFTzgCF9GsbrF4HnEjA61aEbhfezqmFT9n6jNRarFONn8a31JJprYnB8/brhEKYjXzMGxMZ9PB
AogshXG1kVJ+vnCpFLu026znjzdtZYr7xc167Wg1Ou8h8VxvyoTbE/s7Oqhz0RjAIlBG4SFoMslq
kcpA/DPbLxBWa7aahg7iUFemwYe4hq3+j+4laNZxUKeYBBcpspVkL09nTCy4iGIp6mvJFaAJCJ8j
fWZ6e/qjsNt/deJ5fb4h+2rDR60uz7ZtLoj41/h21wCiZ6qVBG5Yr4ui968KOYjjrO0ZCHakt7Ou
y2RZCeM/sf2TkS/+S+XEXNjKiISEtZCFR1bKj2X8A1gVTbOVSfJuXygR9OW+FwUhvS3idmmUzdiX
kmzE9OEpteJL+NUTyzEgQDTVDKAFDgmqmMyxZvlWEg5sBZJWC+rHI0F+fuXmQH6I9uC7bb+V8vrC
Nf3hndYC1Rt7ednasPyIE5oYy/cWFtNhxPKeczbPOiK6Ehpb5pi5hJMyhDhlS/gE7Jji4KGKCgHr
KsqyOX78RxdSJdOv46Xvm+2/F/Lkd4M8iwghoKWpCvSKNBqcje15KbR5UuKXfOZnKA1WKURv4UGk
f6PQ4XqNDb8NCAuRkH1ArKf1spe9ohrH5een7NanJsn3d6vnVmoRuD2Yx1EO3khqKi1W/+zopOpZ
QcL0SFmkSTH9gXuoAWwh+OTxSpAI1oY+Pa15cPQOBv6A/IGXNOlpUgf9bFnji9nlOl9B/FEp6A54
T3HRDJ8d2DVOOFC/vEr5JnHane18CveDejuYz1DXLJDyfBXpETe/VnfEnobcX/EANU0xY6aaU5A8
crGbUx5p6896Pshg+1GXq4gfmdqlRgPAhczN5rwGqXc+9piTN/4JIULGgLEWeJ3byvPSDwh2xVZV
uLj7BbGTapF0ZlKjdIhdKvO6p4tu8dP0NdPoseYJ5qvDhvlV+MUmS+N6aiFtkLOSJoCdm5tL4+Zx
dNyTZXPJ26rRin+5injynaNTBefA4PC1v9Ebj60zlFUz7K6rlkgA5N/d5+fRl15v0RHTgeZk/Zmi
102dezGTwZYJ1CBSvMTDYxYjzhJgIZMkNM7/2xgJ/BEsnqWr4lUJeI2Cw31cWlWS7XXMW2/zI7k5
tG6BcivMcnWK/LsXpsO7umh/rwjoFCo8xWnNPkfNVPGmqmOc3VWuhplRiHKfHGBvka2h1ymokoKz
+93GHAcdfk7+HpRMHGY4lka0KIK+d/IhLV8qLVJcxosD2PXo1nv8vcK0DhlsR0m7EeRJEFatJReO
xLcxgcUNpj0tP6l6gdqz2kVIdtmQR5oCi+KCt+qB/9hXq4FspPHnnBWoMuwMiacbvKcNMDqQNrqf
C4+MWrPxr/ow7LoLh3y7Lc667etXUBNtS3L5e4vnZwAzgD+tOj2O18VYf1+EboXYgMpO1UWCacG/
wR7KEmZDOzFcIAfA7V1kgrNfzRTO0wZQH2DG1SCDAw0S371x1skho9VvrP/WEXFdHjfRLnlWWYyi
DosKzRjwExrD9RIyU3EoPFILX6jspYAEDvA1r6lf5JY59nb3K8sZzc+ypI9lsh1sx9IUTkLxSerg
bWA2pDlRMyOl9wvVVDNa3nkw3PLiraYsyfLMHMSDC8pEfzNBwRHJWYj7HPMwXeu+e0jI473GXMFi
A/5jnSt/Xaa8m7vQRKqyDJZG1GtBPZRhqsnjS9I8h7+rrNgjICR0vOdgqHHTBJM7RdWiQIICqgex
N3uoLFl5pulYJL0j0arOc6kLxIlzKCQn9lIyX7+AorFGd7tvMkLX9BqCUgKNcnbWjeUi/WYJevnT
411kBHHVUEc9Lz4rswLfDVLwVxnFxYddiaAiZquqWFK/Pu8r6l1Zw2/fLEoVPiAlooKFSnkLq6+v
2FZE6Ist4vRMFg6rXQlVeCEqIIC2Svn7hmTDkK1nxY0W2HK+W5h6bt52dcMJPqBk3vTs5KNp13sF
TkvpCZJ05Izjnyva6b29VP1xai8ZFh+7MB+O1BzChyVQ7tU1yHqC/223SFKIjVM+9CAbE6iOBPyw
FNDkgLM9oLYcLmJYHLnvQP+Y7Fo2V8v2HxmMgogfa+szJoo6z/IlNRYPCXfBaP/2MC2xmII63RFD
iF8TeFFLzaPHEhwZ1HnZ6e7JdhDeyJkdVEeAIZS2lf3T6V+m850M5GlQfjYnq9tccK0MkachTv/r
+RZiohbPRtAo36oc91UOHaT6zFvUs255uWKDknobnbE11pVMZBe+d8Bwngm15qubE1MQYodixCsj
iQmMH79VwJIm9cf5p00AtZaqCiSSlO8yXdmymWpqNqNKz1Vv/LhtyIWzyAXbnPUwnwJOkTov/xwB
eITqVQxZimjIzIaAGH86v3OmaOIntjsYuASssfesLT8TTpNBIhq8pBuG7ez6H9RNEdR9DUec8mbE
6jTRVH0AyBIEXaVdbVadqaaGNdW5659pvul83x6oca73uSviQB2mMQKqeKQc0nSU3UmXEIeUoHgH
Y7K3Nak8j9Dips8/pGRt+eI2xRlbOdsr/uqHr5CAcmHo3uhcBkESFEqFU5yPHRHszSs8hSG+0z79
r/ujd3sn/Vwx1uiZFgp0MnQlU8AjKzbPXBmfH5z4l8+lhE6ZYLQYU4+9Q8VnqLOF6KiW5IMv/PqB
LBcM+hGT7yt9Fvc8YttXy3PFXYSClMJ1XZ1MFAaK/tifPFRy3Q50eHk5EstEvg3nb/9tLANQ0W1F
KnsMZgRePzyFSJvhtxnaxKrRCwPSlsJ4A+tgydm/VZqMnvnbKdEzgroZvSsRFxFe4/Mhd9kbr2Od
UwEuDaM2AbeMu0zGkGjvVasKSLdeITNKh8GnRvdVR6+dmrrbTZO1BkB82P6RgwSLPBiAHM5v4Qx5
0qk7x0s35B1WvW1XCYkEpewUrtsKasv7pD4Add6e0toiSQf+OpXdWG1eed1XJMCipiNowB/cCwdy
sCMyKnlx5dI3G6HSvh7p4peC0nCpEotnO+NxaS/Yq5kPL5o5tSpkxC/YVfmF65eN0nnRZ9L1iyRI
prQQL6D0b5Pe2apziSuBBrDFeLnMjoNSvzxrRSWfv/bN/ISN/9UbROYfO857K99cvmhg5kH4JmR5
/sZL2MhZxOrxQdHimypCLp4gwyiTSdvrBBvjE3eCgNAdUNl7Q7Qc86hIiziNOsM9EsxfujRRtQTO
hCV/2si5lfi9o1Vpq3meM3HvbauOwVjwhznmTh4thNAngIJ5VcACxnHPi4w2migEMRddf7pCxTd/
vwrrO0n5Inwb7+sg3rz8oQVmwBc4V4l2q34Cd0hceWNO1/A0yMHjY0C9Y9OQv3iMKeB6Eif9BylX
YvaObGSMYXkiQUZeGvNAnGhJwSlrj7NxCyaf95kMNt6OQPo1UDRuzyqULX3Izdllqbp63kvVE9eU
AS79hA4l6B4jnRIdCSBz8ItIltKfZVhKmE8FFETswR2yQwVS4uFemUUq3c9oA9tWWFCGq0OtvFrr
07l5IsJaXos3YmSg5+PZom2SCyZVSGo2zsnHBFjeqF5QIHNSYj8C5xNE/IVWgLvsNB6j3S5cl0Sl
kjxZl/USXwcG44H/IMWAUDOpP93um/9yovWyN4+ZRVlaqnnR1xSRZV6wET+6MK63Dy5U5rnSf+AN
0EFXqVyMlPbQ9ap2g8nYRvgwzSXjbb9R+rE54fJYXcuPkOIFLVabXfgk7xfxg+4bPx30VeOSS6EH
5ISiijFgsgoj65T6G9lZkqPVQXGC5LTKwsbWAi1LXXIYpDqx12Xw7vvhymhIeM+BTwY5cDU93t/B
zpjltRkCWPwxPMLsiPKo0txJuccCHvDFqsbiRoEFXZYe/K/qiFX1IxDW29hO28p91GRL1QeBGKoC
M15U00tsGvjBiXk8ccqmg6tp6oUx3VTaJqrfNFle8IorIITvuVAPEM92NK9FYrjjpgUeVp++TgQ/
QM5oJeWwwak0e2X5jhrrlDoQUlky2cu6GGR5/ElL1U5+5seHt51rHktmnLRrCgtMjBra7N9Wbxlt
+a9PtOAPBjxeLQiUJBcfrl6OO2tKqIQJ5MZTaUtzeeKoIURz6ahoX+aSzqZ1Nw9S4nyVe0FMP255
QAEdDOYLOukzp0nGuw+Eu2pDeMhq+pSrShuBazzVyH51b0POiLzo5yBQsZp7R2qQrB2pmkohosL5
tlCb8sehzEkfe/9i9D3I5lqOjcf0ckW2c66hfURl14/Rx1LTdUu9jxDkh6BTGQFlKFHX/LGA7Rnv
+58JhOl+xLnPo/yozoTIjsTj7CeRs5akvgYj8QNOeJQrPKGiXv/pQMOVnR36NjbEGO4X0lBp21e2
wZ0diivr/9lBok9wXYVGwweUS2f9kfb02Kc++EONZlcO+f4VLn0LaOZmL2k87e+nySoqQJRIH33o
ToDykqhrkSDI7MfNoV1mmVF9X91ArT6iAjoFIhT8AH7PX6B8o7mo+LsPvp/KZKJIrYEC5PaXtjxC
tzHqAQle/XitccOzeizeVEkCyAzrbTlAyEY0jdiE/3sou3q5BSqr/8H7fdr9ZlYXjoQr/givdRkz
LYS7pIWSr3214XjXmb3DjVlJNlErXv2Ibcd0JKTiMgbXb1yMwZnAsxGIATVC+VsMPYRC1tzhIjW+
O1U+YogH6zQs8ewy/nwH3pqHOX9WhB5XwK70QAl6+QO/H4QNp6ZXTi3pXNk/BHzEqdmmPJgo6A1r
K7VerounHSnJBiNa06djlFEX7r2Dcu5Dz/KjWxgw9siyiinQ24DHQ1lsbW3jEJEQkm7rch+hn1db
HoCy0sjH6N2+Zrc2wt04Z1qt00lBsL7A6Q6EcO6X7uTtUMoT0Q/ijlzG7iD7yYw/zJTQWd6srBJJ
KanV3+PYpdtyrLF66fRjlsNFVDRTJeUqKWea/+fBwmZLvVFo2v49e2YCblTMv/h+PTBSAbLzvCY1
7ZpXKn1SUrVh0V65D2FWjdp1YBjjuNPdC9bMgoqgaT146DPEfqcdwPq9snZDM6jU888sQrpDbRF5
NwfmU9HBgyCLLirumxZoak9beHYqxyDmxdrcm+fE5K93Xqd7bDpzgQhp8ee5XPY2N9WR9ExzTyl2
vrPth+1BE/TIDue3gj23qYrFgZl4f064Opio7xCSApTWFbFmjZzod3Fw5XOB0mVhEoFSTTLe4UDb
ss4hoZu4MCxogMuLQJdyTk59KZX+0NgNN2yv5JONhD5K4tMFcs6LGtjXK0S2JHm0jRPI/PJ+TGVk
n7acI0zALA7ZstpRrpxdGirI9ZyIF2MBwTdZupPGS6XuuWC2vRXwzDvnv/ZRASSPI7cwdSphtp0t
GuYh4J+lWq4dFw32tvXjH0P292CnfuwZ4rBSzkACAuPyq0PdZnG4ZRKnWGgop2ssNWocoBbh0Mqa
wQv7wc//pIGsLPqtFiCBZeWP/N06nLqfw9C/u358hynmk7LRfoRiK783p8IETiclD6QFxFk6vef8
5lewazcLHFaUD4j9r9QVQYP4x3t8pf6fb1CnSJ8hsEYSPGEaihnnxwwKPDj3dZ/mK9SJh8tKyfQ8
wTAe130BNGtAmbPaBauFYLTqqVryfpvRifHD9cErepA1uTgHpjSnlgkZt2cr+Il+D6L8ajk+Zwr+
opBVa4wQQFA9iL41MHgsw0AUTq0xX6vYJz+iMZubeCxCIkSgLyfV29nYodhqoU1n4034CW1QFD05
72GjL9LgYi7oJYf8zp5XizwvhkvGx+O1tq3bM9cZjzqmd9hR8GQZjvQL5nvOh7Pl9wmsdblXh1tt
VxJ1u4gmJvVorkeXuIPrN4ORzu4GVdh0T49fAvO+xcDJCG3mlm2QnsgbLg5hZX1uJtcXcvPZ9te1
QrMj8zQkg1J06+53QMLHY9pPLVmfeAuDcadzG0cuBmTRCChOXaPfhRUUMQyr/RBcEpMp9fZyR8JY
9peZL2JRXkcIGq/ba/jyOVZTE3/3vr2uWkNYZICRJa1Bcphv+qATq02c6GrY9kAdKkr6xRwVneSG
1pKE3lt4qugw5vQBVkYcxeUALFe5advk8TWzlguUULgLTdRbsNFPGDo0FafJxg1PHkDszOUNjPwO
5TpI8/p32eOWk4Jetjz7RJ6XAYGTBLlzUg64G7YvACEaXscgy1EPgaEsKKA4BarLEvvWnfh9MmQc
pddyNqG334TnBRlYYd5I60Mg6w6Nk/ToH2fYRSPd7sxuSzORrU24jNUPR5LIF06gpKtIrl+ryxd6
8kCAmhEZyvCiGLXjAQ69hz3AWuLEonDpzidwSHA15uwvjcOHKYiC95KS+0NUd/CItPUHqVdPsFUp
MuA/e/RzXhren07pU979Gae9cZF3zWoxWlQAfCEmZ4wJwKWFrvDe4Nl2BDNmF08mwaFrINiGS/An
RxHuJ9RAi+bXxP30bCZj+0G7tRmhOfBKHBlMBclfqqiCnzU6MdwUZtZwDS5tyTD54WTWnr+FmVcH
+++79zUk1vJBmWyDTP5ztye9Ln1vguU/WmofbhMhve63i9AxNzyxuKwuEXizIKnPDh++J0ZwpPQL
L4T4Kn/jMAzX//FFel8xPJvDHCTasE2+JwUzVliv7iqznrLcYfeyuRSzbMJTZhWHJ9FrFqI8t6RA
Eq7YfFnuvN2zp2vWi32ejYrcgmbQ4A/lzhtdtOfHrbPGSQ/QYoDyw0z0Q2rWpb2CDJ6dGODN78NC
+5xgJGnePjcaFFQyiw7PPwGZJEW03Joxj3A7oHY2+41mfioD9Z84CWX0euaxKXfUogFTB78vEnoX
dkOVLCNOcfeb3u8eCUL3sfQp75kQPDqcvmewEH0zT8Em009Cl+jrKjrpNl9r3MyzAsNEbrYPOI6Q
uyIsPT1z1uHy3vZol2mo7dnt8nPvIjrmE0yWgZWKHpW/L4P4KObtlFl0+waeQVQrazA1mJ6WG+Rq
+/FbzQNxc+mC4QbOUBZBOQEnNgs2/lt7r6jwsaTfrQAyzKsbsu/VgFHoNcE14+2kfpkUU7StwmWy
AfKNdMEB6+tV9ghYpRZoJhAijYJR45b77Q71cW1rdkueQpgkDxjbB8Md4LjerqLj8JJSkllxfIaj
CyNh/gjoyzHPg3VnA/ywYaiGBBZD/77QDDJkousDvTy3yMPYiyCWlNdyAwEx/r0lX7d+T/+9suXw
kbwxNqiKK2QXXp7C4UzdOUGtf8MiRmQM7TJft29Me9ybFlM3NBs06n/bprEoP1IIdsatLCf4zB2n
XHn5z5+6T3QMAB+tx3VghJIRHI0HqcJDD/rrH784G+HFeDjQT4x+q/JLGx69iVkwkPSyR6zPxO/7
hEGMJ1Wk2Bj7n17KVonK5K7PE2OqIvweKl/x41BkI/lZeYdJEgmLjJLhKqjWKLNayo9EOfE5zD5B
Sw9DvZvP4Em307Ic+e8vkxGP/K0llUQIMWjQnQjWkPRHzLtlpWrNG0quz6rAhxmO6HXoUs5aF5rf
H++cpcEbqCM3ujPLmDTfGb06g76736E+iHYxqcwGpKquq5nZXlfirkpsbZ5fyR+xD5FScAEkk12R
ivgvCar7tpuVc8Ah0+ECr3YItTYix9P7/l0l1uZJ/kiK2KVkibpk+F1OdpT1Ybe8XHKsaIWAAfcB
poXwU4RaNXW/6ZzMIOA9Jr91PMxTQh+X/yhnq/FwqW+UZg4bZ9VJmIz9qXCyjVseJ2iI7nth+1Uw
uCt+uc4/gxHbrzRylaJJYkJfBE67ekH5YfxFL/03i8jiOlkw3oMHpEMPPFaDh/kdKYmNoYnl+8nI
VWEOMDdPUthSVCK1nOiLz821s9vuPYYIPHVj3E+Mz6g8ndjkLR6uRHM5rdh4c/B0hVDCQrKR8R6S
2/QA80B8+zGa1nikx9Ry+J1Cy0m4lycl72TV9eGw4c9zziULFFm3w3vq94K5bKsm/EC3GeMxWkKE
7gtqHCAHqSSOv/PkKY2p3AUin+kAiDkrTcL4thtHDtJgimiMch1daugBCtc2s4DKk9Tn6vQXAFK2
UJKGi4oJAGhdzMafDiYpF1dyy/z0OtIR7VdUKbDnT4N9a5yC7LH73AR5UoQ8ZFi/b9uFIPYUPhAG
+DaA/Ak6DAVmRp2zBWY1xuGB/WAuefgY4wxZvowck2haSP4JPAhvDdz9ngRfDssN4cIFnzEd3FFs
tojh32RkTfDh/ESH2shanULLlz1FtFvlQgx9dDUe2HUgr35HWYF3jnnRTE2rFVhKvbvoKwFD0/BT
whiJweqn00qTe3PWdzIqxjTJC/GkWAyoxvSDNbJ3TiAxJTA3kMSc02NLv+1jUhYFnhhiU/Yxlw9t
5wZfoxNBXRhsHDao9gRcI80SGKIPvJV+mbXPqGvQlg3UyhtyNTGoGljeVn7UnO28Q3LCUk4v8FiA
MjMaG7xXpDAH7nkehP1zkA0YuywpSlcsMGgjKlL6n5lE1FaPV9SUdA8ut47GQBI3/YUWKKY7l2Io
Cy5y0o9Iw6pb0TiU50D8kZZVUTXICexz02bLxR3U4NHOY5NeERxdZNNHgVTQ0vyw1ms4B9G4arRo
xAbGjW/YJwjCyOcIDVe87yo2+QDxYC/JsiaPRRDc5lGkV7cSGXibRyo7VnZ4xWWMWsUrtI0fEW8l
K5Wk+lC2oJdMgrwyhEIfSYljhqHBzPrbD+uQdALB/rfWGCNqVAkk1mFVLB5QBnikD+xSo5bs1TgD
2Rasv2Xol+KCAqsb8LfV5LEJDASLgrOM/K2zhq2fwv0X0BK815851boEPxeaW4+5v383Ttmk823Q
rw0CrBoiiBNq1IsyI1fGpANQye38mPswAEPk9Mw33J/6CMm+fEEAs5INk01GdFOXN62YY093mgaR
sAdYw8ZuZy8DsGME0HNdI3NfjUTHF9xJ+iB7opoOxiuhvx87rmuU4eMhXge3F23JS3fXx2s7Ytzw
qWVH1ChwlnmnsT0D9gVKCNjp6kwLyyb21nPMwBgp0MYLAtHztNgYTMbpr9I7SbbiZ6Kuckq6t2lb
DNmsBu5EW/Fy19waUR0jvcY9SEtr+WxIEy+IK0Vo1cxLsv1cXtlPCOX5mdkhe7q0DkuMsegxWxou
4oj8Jrf3I9NFt/tgbqoqtHYqG086O/mg/RTAgtCqzzX8XXOa1YjTub6uoQHM+OLeRVfVkPn0Zqge
xC2vhm3qWjRZCysLfU9jjwkC6RPsrmAQ7oFuofygFMzbRG39F4UqK2E66c/B4BZE1INtZfJw56Q0
+tWILh22Yaqsc4nuUu9ePGnkeMxD+04/fl8dyn+hXL7jMWOzM4eEF6mct+5R9xf6JmSA89AVNCs7
fm9OJmt9ryz3fHNS/ZRcbn6mccI+vKyEhrHQdWJkRZ1srk3gKaJpiXkWqM1qSQ0jwAVyov2+fSDW
gtN6vJwfQl5UGaf28tTzcymgG5FHz0JBfoFmNuIP5lQLVzCjSbuytPYtL7N2hSOv+86KAoFeRIa7
UbvJvEzcUvyMzSZ8XzNwSaPi/I7rcKkRquglWAl7Qx7KKDRoiwnTJXOg/KZKgBmwKe0+dRamD+S4
ZfytuZshlcUyWKe7MoaTg+PSsH0SfPioxqls/YkyzJ9TwWK02xssfbqewZlFcgX3d2yKEU0oH7tx
XUlmG59SGoGAU3HYHicWANbKMR/mmdffFVQquVNzrZ/CrD1WEEgWVvAa6NOwoCQHGt1fwit8nd5q
PXViXu/Gt3KyDKPb+zipfbu/V+2nJ4Lz5gKIfuwOX8kSlQ7dxjdz5NvWmHgQgPrW/7WyLHde5Ns8
eklGamOSSGuPF8kBXsmby4EbrcU7PWFAkp1rw6epDYoDf9w2bMxkTmJsWfh4r+Ee8QWkoswx7OTn
vTAmMFDJ6IjdlAC9Q2qFFncKK5RHvmNlSstvrwKROS5T8WmDiFGXw1sPY2fhllY95RZlE+jmthBG
wZJsEitVns8KYVSmjxGTbwiRzwjPdU/vhTL2CwVljkCueKA+xD+79MBEdLJgpuph0IiYkawF2hcv
CaP/N37rjDjZRS8UeOpVHFkoNggrQ4GafGlZUdWgXgoP+dJuyiUtFPVzQpYjuQG7k5DMELfNdlbv
YLoIgP+zvWPs60r895d7XavHSI0jC6fojqQ1cRcXpUPNMtok4OUkqnzcMjLDILD5MjvMlBmkJS4m
x7cz4n1hzjHPwK1JtuPfT2FJcz8RZspq19EpiAqQdWsbqqfSA5V9ZVo/QUw7qTvh6hOQmhRFhDiE
QgY2ISnIWsb1w4ZoigpusLLGbocbug7aZ6L8WYQcCo/gjORMw/9ZO4Iy8cg0mxb1BjswYsMNA7KS
yujo6VGJf4obXWnBP8YZsCFhJWGBBwZBpXxtvbhOgokV1ZP4Z1lDmT2Ktdt9uFcnYpgg6+vqmzyN
rLhcgAQYprueB6Miu8f5+/V97c6/1IHMpko3vtFdfafrjzHiDFTlXmg+sAtJHi9k0eS6bOBInouY
w/2eEczNOyU949CdPst15mfzT9huCKbRu31XGnbjIP5iBYysMXYLXAItHy9z1xeiAsQORm2iUFsk
AeCSGfLsW9rdHapdHDV8R4ElPYNUaYxCO/q7bh3+AM4NNJlSzLc4m4u+Mlau5cPLCAf/FMhpNhtN
w5V4ysREEhTwH1zFCRMZXrgtphKx0qNSI0O6a+qfeCJQseylylPYQ+gdyt95pw7GQiPH09RAdC1v
o3su6xpw7PUhKvc9hj8bcM45U+ToqUXzplvuXyz1oX2jrHE3ieIOnoGN2rYMO7KJ/QymjwG+FH8G
XoNRZk9GbFSe/QWwTDdqK1BabzpWMOE9peeac6Y7zwQb97lnpArugWFM7is+ffsw3DQJ9oLpM+q8
yfed9+3W3V/7OmvYTNgyfD6/PedChYEF2J7DkK8kiMiKUchVz/RHbHZpTgt7uja0lIbBxV01iOsY
HF61t3UEeb6c3Mv5w3KxfuYUF/iKezxKRMUKpI40Js3rKzzS/TDXEHj5+svlNTD+jENnlmpPIXrf
pG4zadlxWjLbFsfRPh1M2dkcT/4Em5BALenAvbkJnHbNyqUXiAfhPLq1xDkhd+ry1z+QiL/6aD+m
K12GpO51J9e9sNNzI8/e010yZkcRPkydTT1X2AtC4wwk6AJ4FdoyAy9954h3x9wAAX0Bsw15nA1a
bAr8W2Ozt8fkA9PtXlGkQMkidYNjdD7IQOMGjy3tptb0J1U9pU49e9PuYXJX2JtYFvHn8x3EQIU4
F8qQY0lfSDaf0w1LkMy5A68H0zUoLRjlCiPj2JYctYqoFotG6h6q/evPEOCxbNLvlJycQUZ3whLG
hBnh+eHyXzfkxUok3xWEPB40OzBJn0GzVUfguTnv4Y9nwSm4D9TnFIrgWmqgLyYKcBvnpwh9W568
7d4S2s/mnUonsWIp4qZ2ZGeYORQsg6UCSEfwgIQBwuRNU5Md29ReTcAkR6jTcz2SU+v0vSSm+VIg
lIBENp1/THR8onDDlGoiK6naxqjSqbhApEdPpk56gB5GUqhQVTR9Zi1OCGmLIuBXTst6P/nqv0CW
GCvV+4EYoOrVyhCHXD3uXB0KGyUWD8Du3ADUueCSzwZIo7WU8IO2V796TN7zRSem/6SUHPcyGwHG
hhaP9YiZMiGbxrmp+hVq4Aaa6GkmaV/+jFQeDb6U6vk721nIDYlo8HJdMTYgodrlPXZP+sdllW9Z
ak1ImYIR9jVo/hf6LAj/D5/TdNMS/XEvcraFts0FSUrg9s4Xgo7l6quvPbJrje0mVOYElEDAFB4l
2XX9E+Q59e4bw5QlXDnSMRpr111tF1D9juBu0ewWHVeM8YhrbmclwGDOOgXav4ofNcXKA2iBlfFB
kqtGBWhF3OPDifyU97xRclzDdYt9E1db01BDnEGmRi3bqK1Vka9iZkFIqtp0uM1N8AagrTkhEFbK
NbhlXdTz690Ob8/DotQIVyPGhVY7q+8mKx/VHRH6PO15ql5UawSMvjVQJ0q0fmYysuXBEpaT4fSh
IVCkyzI0MjwZ3ICHcKC6f/fMcd2JmknTrnYBwYMT+vrSDbmGHeyNgZxmt3PFel+1yIn+auF6tOnP
cXGI+IEZAi7Nv+H4W49Fs/XG1pCbV7HOlAvLXfBUmH0VBcg36585cHbNDe4yxhCa39BAiy4S/666
vKLT0IAHozklkXBPJGx+/IjXGe+ktKAHoIxF39ycQ2cgxGZ/mFyk+lf0DWMR0gzMfED2OfUsXtKE
rFzzaeTtJEAWlxJS6eJpjaUv7T/DMA5L9X9zbFo7s0Hx3HyDBYkO0XJK7SCe17oNW+BHAYSYmUyS
x4ar5b7xuRweWZ0rdZ5/J/9RMoWqtKobRET/aALNgY/hQXvcF95hf1lCTo/KfaxMP5nvBDmbEiyr
ZoyaAAVjUEgXzJtklU4th1piNlc++6TWF4sOtokmCk7ANawlblArmzed9Eqs/V6H6V1hkmPv+UNH
FWdTc9LRZFvZEhyL7GH7cvlknGGzBrLVu/nCzXo35Foj/erFixfXdThDQfUdxb2N4IKQwFMXbTnm
SsDgBXj8juJaJedNqtWFgU/RXCmUtFJCUE6Zvvh5d7RTimF/uAKYBc7uwb85fNmHMumCtgFn8MtJ
oGYk7T7iaecQkBIqBEZcHab8b/fRMXYQtDBzAIoRfbOvvUx1EoZfjq16R0a8anZpvI+q3P+RY9Lk
zbQecylIHOzBLt6VVYddnu4UK+svqdA9xQz/MnyQljLe7o+wEzMMvfHVmTdePIItpWuzaUhnCb84
tHceHj0SN6ZY68Xl29kFqSuAld4cmEZiLVprWRPcfQ+lQFHDzQz9V+TlfGp6TjqH0IEoSdqjXgyp
jYmvnsY+4xpCFA+Tkl39PskPDzXORdUJ8Y0eW3RG07/fLNcSJut1aZLtrpAsVLlhVLHvmjMwucbd
4XSDjQG6Xz61uRZ1Ez/9VacvH+/Ad+122yW3BD6jG6y2cAWq4gOuwZ7oLb1q8H+ETv9Kz1yV6MqY
wv/D36MIEYbPr+jBusHxdcIp62J2axS8C/pG/MDv0lyhnPDXNdr+WT84AKpyinquO4b8Wz3/wMMx
B5EG2+rWKye0jPMrNE7PJoVCY7Z+F8CEqZwq/4CaqJ2QvOq+eviqG7ju/4aVSWIMSAlyVfrG3r+t
fdSyacfT2XBomXnubMbAiNEpgXeGKFHhbLVFI4J7Ocfd+JbO9Ptapp6hG5yGI2GiUt7KKQkWEr0I
zVR3ieRYqTsO+SQdZ02dxZJJ5CSlQS6rBM7d4vTB3Zaa3vFaY1yhW0fiWq6GNGTp+QBgz/1YDF4X
0l5+Rl0deeBwz8Ti5TNYm23IT+/ZlDPRFK8VxRNsoRusrhME8fFsAiWb3NbSNJHEGEm/PvHBDXYC
d9WiD0AhtmLUHmkKMBCHY6dglthfHEln9vrTz8L2qG4H15N84iVMkLmDiKQFPcDeSguR43mOLlm3
V68DDZVzT1znh1L4IxmIgG0L+5Xz95AHhOeLf6K/7UKnpCVbor27z2vSbg+trwn3WTRcczjppB42
GPhqvGrCGt5KuVSU61EgO+cWbLLqWB6pWZl8360kg9Q41Ik+O/G2IeCIxX77oc+vvYxJrmN6fE0k
HCFdgPebr8wAg8ZDlQXr1LpjMlh6snYiP9pe5ZudKFWMgfHvFU3Hae61pLtaH9bzhbhbnRaTwxkS
Y1COHl4AswkQvsY0ASGIrdIcIXQH4FFAzM4pYjOeOnN9Sv2xd4fb5NzQj3VMYXVN0EAZyv49VERP
7gnOr+3oGPWyGQwafH5mEnMeiuKoQNXJXrLu1dwpTB/EwXYA1DlO/wjK9vvlEfDfg2QzXZiIWFMZ
VjvnNN3ikd8HCI8DBmywUDN/j27b9+tgWZ3Hjp38hzpuSOI4+y8nHtz00SzlJW8cRW0E/pEsKVZs
rL239zTjjMd1gt6aRcaH9RQY3k4L3o9qSrnPgXi382Z3R+pd+kaAtIzPy2eK5+Eqg4oE9hVYBnjf
iVw6cmGVsEIawJAT+efWsB0LQs6lOUy5h8RuZZReF3upxWBG6kWZzMCSOpVcYzb7y51zzbWotlEn
v8OTBCC7MMb/TSXNNuSU5zAKuQXDXvFhfDEfFWWBteopeMO8AMDn9Zexcw7IUvSKVRzg1IaOCaka
iFc+nOksx8hjO/p7TmN0gHkXinpKjBLfM1akLvZPsMra4qI46yKSBVbyFFavWo7QqbYfoD22w24s
tYR44a1mLqAtHtJVvDYH5iPaGFdNGZVTpv7QKC8CT09OPjOqY9CQ05SBy++gAvbdUmXilkQUYmY6
tGygjrY9Uk7SD7eEyJDTitaHcWgVAy7R2/GK3gG2+qLeJ/Z2NBHye0OtSbohOhGys5v+eOsadifv
n8Qv3g7MeXDW4yqAbfUXtKtFtgtI5D2iRY818b/gGadH3bGQ9neuCJsPWXZx/Hf1K5rDljdA0oEL
AisJP95HNTheFCCa9zoXkEkmCIYKsYOGL7AwONLrw/v7DE1UbADUSpAhgkIOJ3YfDuLHdVoRn+n3
cAcWOa3zzqdd1lM0wCKaLY6vq5osApvw7fxwljSWhD5eFAltoYoCt4V+nVKnGtGDReFH7hc+ChfJ
LIaPitBFYd/CgB7W95OQLuXPMdSm2YoJfnQAq5TklPqqxdUokv7JkDvYwvMPfX+RMlNB+V7sEHH+
xRtY6AFSvkpNxB5tMMXKtuP1ESTebVlMrcdCmqYSbYMOZR/v/dXrJyfXTPH0rFdEDk2pOOOBgcof
F50duaGM//MQc5dMd7VHFMEwFoufMMrbfkBRx8pKgjJKaKk/nV0xCNwwTPB1oqCTt/0etYiwVYO0
goZyN9Ifk7gC+N+3/PDQAdVL//vPU9QFd9SWUPWAcYRhF6sd3LL231Hrcnyhj1UiyBdz7FcC28fa
lM16UlU4iPDG6R+Onqfp03Z7pfMsE52PlOestoCv/V2is4GQh/y/cfIHv/6z/avZKkupUEFtfMnb
g0LHvLKWkT43DhrIUnh4SrmqD7KFsNrU5kdl3DEz+Sgm6aa5nctMzyegIXOkN/bebb/fXpeLOFbr
y34hzCLXzEpbQcSshFUZCKFKTZnOmAnNjcn9hgapIrjt+LSMoiH3FtA3C+wAQyvlPLx/U8bVlp0N
WUT5vBi49tamru/HcLM6q6I3o4V/DDdVAsZOWgeJ89bHFYTMmy4BenxlmEbnm7LCzNWNVHXzvCQC
ouC6veaIcnPfvq+pT35XVpkvpIO7QfJA920nsjPpsC8YmhLjl90AaPWoaqvmYYKIjNu0lq6zgKED
qpKUAWXiHKJeJjORqNRL4NlfB3KS07wjnuan6tHfbmSFCMBq1gsYSuyZE00xvcV26WDF45XiGg2l
5SUbM7Pza24oXDZXBOJKw3LwVXTdrgfxGrRJqm0gguoXRUpA/HtKNv6QIrtm3lH0X/zZqMd9qnz+
zMEx+y/4QISIrpXKtViB0Wy+l9n9qrBZ3Sz6+G1Y5SY+HFWSFlCVPHBBX+gQDyPGCQQmX3+kq0b8
CVIfrwvMl5wBD5JooNXha8zwKc/DG85OQKiFJrbXsdlWli/y50ljPa6/EukNjTKjh9LjJG+0eJ32
PeNoIuieHn1HgEQf1vzriMScVrF8D3dimS4G3lOBdbuM8p7GGxLvytMbKYhBB17gCtKuRApMjVtM
2efQgHgzt06oq2wcT66J8v/qS5iO47ieyqqbWhDGLzlXftrp/Ee0AWBY9hBy8mld3SDJIwFtbgFt
Qc79hi/ZouiTo5lX5ab7RU2ZZdKRo9YDnYfV9u7tnqipn/60NKAyVmeesGgZobT1THyjMv/Y+exM
lZr6LMKXnTOF8VnJqguyAG9372MiW0HdW0X4zxw3xE1XQXs28cH6smn4RJtg78c0fndMjtrowf/0
4XEDUbtOJzr9zw751NKjXWbDZuxe5T9Npc6Vw5uSXd0FUKEgJtB7nk7IRKnC9Mkre82/XmSLEzUv
NP9RPKXb6StQ5wuXjB+3gu3aaU1bm+odJKDVaZwYWJ3N8MHxyUp5nVGHVWzLbHeAouo78vOjYzc+
lKrNIHZCo7mlIGeKLUtRL4lch/nBqj6VZ9sO9EjR5yfaoocxJeHp2bsbMnN7xDfnsZ0Lqa+cnPaD
1TnG8sQ1vnidTpSouFIeYB7su2ROyOY9b6jGyiPe6hwcALai7plaow7jVpSeyouTsh63td/8BRX3
G/3Jih4u5a7LvTEhDtKWEmaeCk70XlWZ5Q33hWsGtFrXxr7hPDdCdBUafZdoPcLm6DcOTDcrPnVt
YVv+bBOmBn5QFMPoSXnS41XGQe6u2QvScyqldk7jzDNBazGFMSiJKN1NB0r0XIshXTWL3lXIkCjZ
VYqgIlsH4XlTgmm0PktSwZUzq1VAmH/SoldyleeF97KSZWG7arv0kibMsRgiLL8Ovd9aVCZTMhzW
H+5K4I+KtKBtvdBnYw5kn/THSAJ6Jr4pWlyCV4nn/vGnlaho28m8YnnUnCe9tSK12AByQyTo94aB
PgKlxtazmGyV35bbChwXaaTWjpVhWmGIwsz9Kgh1SZa6o9WlIBw7ITnWgh9Exv0TKiEd5zoaL5S8
jd94zoPjpcSRJJ1CrGf97LCrDUXtdnYXkoBQcmSgf5cGeCbVIoM01txdg2z9Ht1juiJbNpYHIUFE
r0IDPRCEqYPpVoFWPhHQJZoI6MnlsXko/W9RHZIAXyUKbEA86Jmx/VdmilPK5QADaNc6d/RrDsPM
SwABBvd89uw7vdjFPqVeHAqinzBjfnRkq3nZwQtbkCvlbzZ/CKCsEk7f14iWbC14MyUCNZiSien4
1yxudGFEc+Pnu+kb6Iiitt17+RkGJ5mDH+S7c2rHYX5R1xDx+Nf6Vguts5drr7W74q5Zg25jjAIj
+jYYrU07LXsXtBwOgITdIDwaBnJDssnb5FsUFFDJAGp7RpZAAUrQypFg1Udd5hRi0Q/Y2Ntr46fg
kBOBwpHddb63bSI8FAQ5BGlJlgdqA41tzqWC4Pl4GWR6dn8VJWzjWnlDC7Htec8IA9Lc2ZIqhTo/
yh22aicO+9rb/vbDhKYXDvYyiLfKTwzEWV0QdqTSlkVQml8Q6NRLJakKxaU0QN8AAwWm31GECRyb
sOOhbbhI/4MBywgJts07bjFSz5prGAs2UzMq1W34l7ywPZc7pKK0Zm7M9hpFDoMT18ljWFcAMwD5
SEfvjaCvnG+xT38gXGPwEwLFm+Si8clLBy+TFTO+AHW9Q8r8WoeCENRwFHcSX6kFkyvrWbE40B45
Qayu5Mqcrmf0jgFjERbifRWlQP/n9xzGFnEurrCkVuchrs4XpNPLSEtBK25XX9GKbcEGmN/xkF68
WUWubm3Xkn91eGu0bqUkLfpLqI/3nzHUTYWXHGbyTo7qplS0OoCdErsOSp2fmfQd84gg+r+xOD7X
4cSFVPd2HMRuMOSvz4dFw5Jt9dcGwnhFk+blPhrZV2AV1V/ixSTEfYdsbVVn+YUQ7jolK93zO7PJ
Vzi4cjFma5BDQmrnp67I6ffBgFDKW8U7DapXWnUbd6jAukY4CckOTf7+SR1XWKml6vLemujTCKoN
nsI/X8QLl/8OTMZnUqJ6LYFu0ocL3j2XlLMVsutIuy6rJM+kzh6jy6UMULUafpFzXCNdlmmMjL17
DRUgUuQcyFOWz5fQXJi/06w7CvX/7byA9xAtHPZYLP46yuqjCl5+Cz+0pqRQifM3uG4Vd3J4KDLY
zebNVDDZda6oEWS2MnrmNJ0ibmA3159j0HjdniSGmkaNzuYmXwEnZdakyiz8b1zbe8b4t2M6zCAa
RZtNEVAmd9UoluhXXF8Lfj7BObxNWbIJ540Ld4M93Yq0bYV23WTVCLYF05ONga9rjhOWeVwhcOMe
KExDfwSTKvtwSrQeJpvnd7eaE3FLln4xxDjXSvwtBxJ1xWKXaK1tvVADBSSRmsAppBcZ89fQ1+k2
mc30x7vy0a4dgPNs+T7nkSpoP0Q/xMGv5MvViil1Khn3z2XBEcChlLUPYcbPxXOkyt7s+q4aQpad
z3pkt/NOTVO+kOK73MBCMKgid0JT2FrzckQSdqXXlvLOovUnvWBPrKKfATVgwp4g6SWxiV6y3/Kz
oVhVndNnf7szMPWcqDQTgQ9uQ9FzKMNU8tHsf3gQ2IhA/KGtJo7ncI3owsypg9fPjHCmuP+fr7Pq
XETVxF9K2ZJrcpTjR2P/mJNhPJd7G+Cvr28IDLydPcOvCYH0fOFEkYe6I4DRNGzOKrL4Hycjjt7O
0qNdiQyrNJ6hmAhacZHaj72D/LYldBpHxNjKdpKcM40JE5epukT7cK8NsYvlClTok9fydkpNoBuW
eOTzw8/byRkbzzPN0alvvjcHrFec/aDADBPwMj5OnSLEjmr3TA1p1pP2ssSRnr2uCo5wJp/w2t9c
fQ4bapESTKy5+7Ohof9vEGaiRiQUnVvygrCK28uE7c0oSLUZV63XKTAB9n30Fe4qcTEdzr1OLrz2
FlWehfEvdTfSpYrYgjKxvNyLDzw3WQvBnsJ02MpKvHQhh2TecMJU0bGLKgFmJQ3I2qBTy5NBxreI
MO+iyNorRlFakN69hl0ZPvrsGcL2mXO1Pr1u3z5MyjH6v38jDbBNara+tpoGN9xV9o8DFRp94cfF
5SNzYHqW3rCiovsRnzu31lvPjfAr5N/R8x4ONSVZI5iewkTMQVqSHjW17PS9/vmA7tCkJNn7uiMq
+aHPANvRtnX5FhnLEik44zDzC83Zv8H6cZCk9QhOCk90Zn8lE0CMEGDZlLshFaC4948QFhUajlKL
Qbvwe2BiYKKmY/APjLRM5xhRAJwAlTzvJJavm1Jj0TaPfGgWIjXxmG3ymuZrCnEuRgWKOd5yrxwG
wpmsqGBwBcSFr1Du5KZKWf9mLp59HjkLBTC7fbO0xJO0UUd53Ly6oa5LYHEIO2KqKVtC+pbuuPc4
/fY/ezkyyPdkfv8hq6jzz3uQorytYTrHr8K03j6AP24TpdEPYolLwBNyGo5iDKQyZEYChmHyulnU
PBD23arN2LwL1sJAhQNujKuwMg2pW/AaT56j4i5DpbWhCa/4Y9TRCboAUe7qI3EL0xtQD9Q2l4xJ
dOiqnKr1QkLkxnnfZAa5yyRt6C8TQtiufxj7/FkJCcj88+9FaMElYYXoXI2mKT4chvhoa5a6MRCv
rLkCKqxUKect1qNq4gb5Q5uxnxUgb2YtT/28LV3ycDg/ZU9HuLtPZmVgR8jxhFUe5IjoHKU6jDoE
vYHj3AuA1jMA3eQjluPsLFNXgFi5Gi3+VvzZrfpGpkviUzchqT5FjeZkxHWkD9BZ9Gjcg1NpoNt5
9LrDz5szeuJF3HeJDAGtiByj9zsC/OL5VXQu3P6VW6mGv35akWeq5olnXriacdvhlw3KK7fY5BRK
BCzku4Jhzfxw6U4IAmf600t/4fzGn0hitdzeYkbQ/uCNr2xgZ7CMg/9cW1NiN0/oDkV/AQDQL8Wj
zVEe4PqKlQKbyfMCgS8yLdhXGRBcOq2GGEwfBaPz13E4/4m3O5uAcBy6tWMN7ss2KZ4XOdMu0TI7
yCby+FTg4RwKakS31BShsJuMv8wlrN9OtUtUOVDH5uaThpYCgAgqdID2fn9W2wL4PF1M/MJ91DWg
wXXY3q/Wuc/BqqiqIhxjLH73AfGgfUCW0fHcO5doDvrYcMGxmrOKRphGc7Dh9NImceNXFHMAGcO9
3eXLhdyFsasnQLyJQZUK/iPR7k7WuKiD8jm8ijkprFEGTK4VlwuBuHVzGjq6hV3l3u7TVFUnxBDP
2nxhZUl/IXWlBVWcL38Mazr9nONd6K5GgcVjyQ19Kq3yg6LULXMd7hy/aGfpToNovzYQGfdRjSr0
LaasekXM146JaZgJ9avkb8z7JKi51KMdp0esrPCoe7Dd/D2MQmOR+Cy2eBvEVDZxCdbfbZIi5Ef0
QDZODwPwtH5GSngPRJK7axP0+YfGsHRy6Lge+LPrNfDsShIGcdvEdXJ4zbSPFea05HdOGrOS3QDF
I5H97VmrlEwRgKIO9gb1Du17JO+TgkGMVyLoNW1UJPcaSuUFO5gvhc7Lo1geoAHgze/DpTd3mVaN
6K7w/TRg5WB8gNqtqkva7TnGktmiLPkE8WfeUG7hff7TY8EXzj4Y6Az2xPXT8ye5JUJuwOnmC/Cz
xnLurpIa7c+fqRz9Z/w78AlAom8S81KYORkAnu226+RcftsTdt0lyomC9PStUN8dTYcQxUpk113K
dmrslprxx0OOmAlucVp0ZHVW1kMHghteDL3IkPe5bIQRFxirYCLt89KHd6SexTXyS7LQsO/LnaFN
k1DgMTIZDKz65etJ7gciok392fBKW6tlvjLyyhRLLWUwWsTLHnxJPCLdv9EQUI30GeeHxxXrBD1W
S5ChrrLheMpFdJQIPdYYm3ybDUY/ElBw+YbCZkfitzw7gHYmmo3mYYQpCBKrWbses4vG0QDwVoub
4WEiHe2cmGy0l9fjRb5BeJf5gn9teOoHQoBow6PPh8qUjTj3u5a2ub4WbipnTbylqXg68WNiUJru
LMEB6dafdQYGgB+doJ89SIGXr58CKteYxjxk4+j5rX3vNv4VdawaoqYEtqceLzEFjGZLJvlZYCqU
xydJfJo13O+Lg+B9y3kq5Hp0rR9pul7v65V32JoA4dI0GF+jcTOwypT7G6Qo9ilzNyxgwsUuv4BB
TvGrysbI4l9lQHSP76KqDyKORs8CuIP75kY4TgUZLwkIhmUlFqmPEm3jZwmmlrW5FsX7NF+DxqBm
N+bkoya7xNH8K6LNMwljCdX8Aj1H+k0iUwDZ7ne+njCZReKHzXgfusNq7/zhDfy79RInxt2PxpK2
LNFxDJETjC4HnTjKPm4k9YGdL1qiXIAGJ9QxjHSdoNY8rkjnMxv92L51/HyysuTch8nPi2Gg1a5t
zeriBhGrmLa15V+QeQ/0wzvvaXeHsyv+t1J3NJqyPNBZjPD9bnKYa7mB4gWOxqAbSuWA3jiHNOQD
tXokt2PJDji+xIavMtMY2Em5IFCYGAHdfnHMxDXPIGvsjv1d0iZEBB4HcgLzJ0qQYf7PUJRraMEw
qcslJpZHLWS0QV4SocbKi/65kr/gHhHUe5FmYNrev+m3vLc57zxJiMQ4MyDwJXh0BUFQMkr0P9TH
ghwjJYZO9eVVliYVV98b5jP+EaZejyjB+tRAYNucECloEASNuAnGm0jZDWfLWTTdVJqM33e1Ax5g
8X60OiYUgCjRcSx8Cs0md478QkwZVQYJSXtGFw8iswteU4IrETqOQC8RzxjcLfsX+CeveQOprBmA
wrpr6j8cw+LQDG60JJgTol72tyODLYFgM0pWbVg8hpW8XV13C03r5yBAueMwlbUboCTVJ2j24d12
7QIALUpgHZRSU1hYNboQHk07UVo+HBBqLc0tWWhWn8h2hdRwfLS7wTvyRgyuwhrIOtW8hTQtQvGd
OqQ9RAVKyoDzMQ9n9+1Qbr5UCdLBWjy4t4OmFXTXr9Q8iv9WuKw67FtFwHItCfh5MkGuJlvNY5su
tBCqkmXmudqrKfSYTwNc+tKxnRWmasOy+45Na5RusmUEcSi72ZZV8xPcSuq+hIvclb15skom/lG4
PwNxNKaiKUeBvNmsi/i7k0CinGsP0prv8kLdKcPZK9Ak1T3OfanHuRavJtDJ1GuH9Ry7KgARNian
ylNAunvUpFAQ9dK+Tw5ItD0jGZ1tnyvDtKDXEEbT4yhxwFIv+0zw5xLnbtcPMKEgAgBeiS4kNA6s
uQi6VNazYJ+Dj8IYCynnWLkyB5kt5BeMmgEo3e0zNbcCRi14X5SpfdtHUVoAgj0Daxdsqi8o8Ua9
irVU9Y0JvyZL/Z31uL+TqqMbcekh0myPVUFN2CEtJujbTVQ2tLk4fVMgIXdGw2094rzCebkOL+io
cPnThs3PSmt4P63OMy71jHvdKvutDBneKzg7dFTklvPL69GhgcID/IZsjJtCgGAU7TQkEJcw7P69
xeHiNFa6SgI+j3S5MGb7798a5GCE9KSCWKsOiT8ssA4h7TpWarshkidyEtLlwee+9ivWzjyRGJrP
Simf4oENbPnI4H9YyfjmaETz6j+CDSO8+lEnLItXbdJNVL09hU9t64rB3L83sMRwomLIMZ3Rs7qA
Ko2vwe4iJY8QWARpRV1l3S8lZETwuQbI3Z1Op2+6eylY14SFICKPVFnu8V6IUQZs2DTc/aoCxEJF
y5/I5pvM0QQ1Ubkg6UU4x6XsO1kJFc7a1Wa4/Bawd/af+4MugScJujpuI9m6MGT7uMYm7+uVDYQr
zBqluHKN/zwne60flwEK7YsEwFKmk8ZVFoPB3XTFAu/kkLtLRlLWXf1fJoa78gLENA5YyViXPTZg
R6JWGINGIlHIMFuZowvqBPuhJkPEYsoD2bmQMfd+0CnY+t2xCFJD9S8amAt+flYcLYMA1PSctWae
G643nXUCqbPCU18fq1r7PzCzGWPMYrCOyGyjlkLuEPgm/mDiKGIfQDdpiYCayPZK8M3Lj9Yi3pZr
JHExWzQQYoS1O4F4Q4gaAUKuwAhKP0ihVO4WOoheDnvvQg31amN9SSc8QjO4sM9Y6LH15VtXw0eF
en/+JNygH60cXRQZEwMQ4Hjnbv5znx4a7g4FXVnDKCXTlntXuH7k5u0TKPhLJTwCjn7qpaJEE1WY
PHAbJk71mFdWuwj2fkhJFRGwtHQKe02AY1+4v32Oxk/T2xaZFxB/xj+OT+iDIV1RSZAYe/nLJ2Dw
dmII9BE9wNGqTtSEMNOPZjcsT8++5WiZbWwzgRmsL/r4MiIDnu58OVv2T+wO9uZsOj9shJLFi7Cg
Vk3VulhZU4jjCtEkFFEXTIEWd2YknhSCXF8Hc3CG/9Lf0fjLCWVD5uyvjaXtS7oyLLwFefogFYAC
CivBabtLB3x9/ty/oN/40/S+AMU7QSEQJwxjcWFW1bFUpjpiBL/x6xOZomSAqeM8wIOdAk/pMP+t
rNeGTVTflua+O/OwP2HcYhazUvn0/XYboGe7T4Tg8Tn70Ys7KUD+d/S7Rdd/gFX5b8fZ6G/AQLLt
ys9YtAmBpmMTOcXj74+P++A+cGt0XxL6b3Z2lgQoUM606jNbMwZ9GdzTaOLNBD6OfVWZKK4Wl7Bq
D6zYlgEaINyYNdkVC3x9pfmPU6IYngS3vswpETKllURcMRcdBVZ3IMVRGROcx6z4v7jHhQAyN1sa
yh9K5BApVrNwGGTAHbCb+doWDy7NAo+VqH9Gyyp2VdVUYM1+fZLz8wHoUjXwEKNtPsS5VPotJxGz
KQgyz4ctLnFt3KONOfnMTMtSHnAfRbR+m+hUiBmTqxA9jtnoBPjaAPnoOVXKMpssDSpBpT8x0/Qr
3tL56Qxl39YmqRITbuLcHIR/jbEhRYyHddCHEoB/yXlKFG8QBSMA3UOhmad+1bK6eClYptOO4dUj
NKHZGJ/8MjwEab96MphcX97LDHEFvwyq1zDNlc5NlH52oesKQfCuC8l9KeVdtDPqKUtzkcPxwWgK
9MoPabCb99HnBRMoe+xv44ZSixYTPXSbby2gtUdVOfeuzIRXvazn1xTijLf1DowFXL5+pUvhIq7U
LpK9e3viTb9eW/O5laDRZhZaKTs27bhDyZXw+ZnS98h1Ri/sMwTHnQUIshioj9r0YxuIfC/O9gfo
UeNMZZUHh6yrJN6vRSZZntn54IQAXQrI3jGzAO1vyQnM8/1KZIAQfTiQ3XXsFU8OJVDKSO/cKOck
FnIx+TjrocffdUJ0mViE01f1i7x4XJ5D84hs55vf3sfMd7n7MAfO1Wnz6xK25rI6pwtIDUpxUBbu
PU/nU9GstUqwb+pLIlc+426LiCsy/fHdPjDzWhyuJGWDsqpzqRgxmsyC0vC7peG7oPWH23tV3A2e
GUl+Ukj3+qacd6oXYfCDLyCnBJvGKhwQwWZdJOpzPOfn6FRIrV50YXWq0ZePd00XEs0GaHBiWu8V
CaXq4toE7PuJ/eipNPLbaxJTr1ecUCTT7JhZRTfY09enZPf2G7uvFOmFOsq0+T4ZV95cgMj2hL41
t1HDdvTGWQ0n8HcF0hvT/0etP/g2XlOWXCheHvckqY94EX7Yl70qEBpUVBrut018eBGBVQtlgWs6
XXG9KomKyR7UGcmgBBaJA/+HRt50Vr++OTsfjbXkp+Q74fM8zb6jxLYwQVxD4x08JmCAh32MBMW8
5Agwg7FgI1I+EJ8d/2iq+u7bDRGU5JLJDJd03F09CRIGHRSTjIZ8m/LiBP0ANPIbxJMtFNFw536J
yVZRejAMsX3xcm+R0S4FE/CzLb6sOauT1K3hvD4CVR/CQdjCPFofg2RXAuTt3uM1M8t6mwpD6MQa
mZO0fXRK1WkusYRjfeyw0P4DR23nd9SbWFvqavyCJD8vCqi3Kl3vJ6Gkkac9Hu6uY2Kf2cgY0mj2
6WBtF0N2NWpSPrlxId3y6xJRftsW2eoQ+jE+8pbB0m0hvBoJyLQOe86mEHTY1+LOOIqLgAnvxhE8
5g80MY/I4s+tdrbthKkMavaSayQvDaaxsTFOnB8iH2tUQeDhan4udM1IKRSZYWqlCdh1PfGhko4C
ooqmPbBvWcmvLTs4HiY1Ydr28VhygRsSdyF0lirJ21KT3y5cgb3MA5k7NnmUasDFSonO1bfKiBp4
tF/rjUcMGxoaWdBwCWZWQeGdHqS3Bovgw5IAkFRUNZKdJWDVBjlzD2Zzeixjuf5NWSMbmADfUUN1
gCK6gZPQLZFdH3APuGkFPTPG9k2dUhlQvynAYzChxqmBIahamWh7vjXgWASGZmYapVe3kMnGSPgM
FVATVANwU0i0LxV0R0o3IXzLBjYHLMTNeBFTFs6pFMnEhhrVITa0CIt9/QLr++iEkYhxk/O4jMsG
aqUvKt4QPuT0B8raRGLS8HeNbpO164zTZob8hVdWHzbXJ2//rQRHyHqJ7PNTu/GQU7mqzmb7gxXZ
cfd54ZyZ2ZDL3bQCpE8qmjmUaSbB6qJf+sYXyvIPxraWj75pnAUXgW5rFJ/RYi5pPtSrYZEL2pQc
dZR2jsIpssh2Dl6sdS2U/DilKzesUKyVJ0M3WRp5MsGKDjc17gyz1//dehAPFjNSkzRhKew8Gkkx
SRM8nDZ919HwLgovR5bOyOuGigjgzHbmnrnZ/C3psGhtjUQhU6JJVagOQagc+9j36QmrHWBIznBE
RzDlvtJXqUG2CPOnBNK4MMZ2oqiy1LnydgwyZFXci/1Us1OV/Rdl9pTuyN+XqBlm1cgWVEVLA98z
TaG7nbF8P+4H8gh5uFGQW5uukb3+7gaEM+guL/RprHvaf+0pCDnR9icH5JARpXIdiyQkdfhKrXj9
gJuAuc+yQGggJyZNm63f3bKhUpseZjYKKM+BiO9dRc1K1CIIXF47j0mBZ4TOxAM6MyWzabAnqfBv
Jewe08n5EjNNuMOUGY6JhtQHwbU8iHCPCKaiEQSyN1PDA51bEUtiyTo6BbBh4AP1uNnwf9GrfCf4
qWMxhM+5I8jcEKkMo70p+oVSYPbmgdN0PoUuzOBczuZo8VlTDvMwyI/n4KdG7uoj6BeNLLnoH+bh
Myq2m7u1mkwS2Zw4mrjjyLHPnCA3w+PifJa67rMK+NutEoa+89m588rWsOfuffhgPTNGwefSGj7n
0tlBFgDum40KPCdlM2VuosUHT3N2AAWtY4f/aF93xmwAPHepRww2woDEUZGc6kJLc5NSa+zBFOsC
tC4zvd8C5x+dBvdERqd9z5rAHE/9WFnPZA2ZGtHbeqEOqNxYL/J/j5v2+H/A7TaVeF4O5iXPKjVk
LjjV/ILtAZrWHuyDGk2B5wXw3VlzISXsTETWF1kofDVCgP6t5BIhhWAzyCAttO5K3aSxxORrURRS
ZoQadqf+o7Z7mI7f6+xvtQaHXvGUX7HxPyMeFAHxkgktYKz5dYE9ayNSvKKm8JD1DoToQ927Kz6Y
IYw2JpPIhQPdy3ujltVY6hfN52zQiIfubHivAzwTMDzgGgKd8uKNniLRY6+f3aSGfnefQWulhcrX
RsbeJ9p/yafP7RWuHnkO9G7SDfYsBL4+5FTbPVDTIfqnwac8yTEL8G/Cm4ZyOFaMtO03qCWKH1ED
3fiSymsSdjusGpCKtduL4DMTTBQ/tkA2bHJ3JgIPJOmyrEwaZTYkMR3aPbsBEH50bjuXEzFK17xi
C0MnBteUDytclUQ035ite5cdaGOPeCO3+s2pRaAKCNkpXvwinos+Oe1hfmZfmbutQ1gpFupNXODm
Y0bKzu0vz5xaQD9Pcc34LDXmZPQv7Ee1xyiVH3jGoAQIzvgM1vbYha1J8ZNUVWu/LPOXiC4rNc5O
AUuN/EmBg6BnGuy+
`protect end_protected
