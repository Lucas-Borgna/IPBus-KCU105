

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
SFpyA3WDAkH/h6gENMNzEC70V+GWX/AuJRjC9uuhJRzuSJx7LjCfMePfd14YnV5eJpUmzZ71W3kb
9tnOI6KXTg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FappTG7uNGFdZRwaHkH1xaFvi8BC2aKkPLd6PQ4xkTkeceiv05HkyC3+B1zcjatywH/Tgp5My5jL
RzYpXDHCiS+WLEnVqDpcElLtP6A/XLl3ajXqKvZhmMUVZsEI6d4wI3wE8drV6caY5dK99YnGiCxy
c/wD5JKxsx7IEFSu4qs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LRNAkwpKrud10Lp0Eq/NqP5B49JnJU8WkULh5UDIksixm1tOfz3iui+8sx8gHS1R0x2iJMsSndD1
7xzPuxZn4a1eVkZa4n4EghKA1iQCL4jIUagjOF/A226osIvTkxPBVZ56YpbMiMwMMgRLER5z0xet
LPBfedO96PfexivUiLv1asz99hmC5fi5UUap1VwJdrnsIHsC0bEW3N+9FFvOSldno8glOl5txGSe
hOwrv3syYadhoBtySSxq9fjTH5UTCT6nikZqZkVb5yhHF7eaz/U8CnmNnm4+vrB5n+GG7KIVkI6G
7PqaCstXyxVZ0I0FOvUz/cqAZvJcffVN4NdFGA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u1B6Vk0Eso+5EvY7kmrlz1476LggIIsaO8lHvFGJ+HKHly0lYN/LsIll2vy/lYtCwxTSlrDsJgNk
NtsXioC5DfcQQ4kEDu1f339J7HYisXvM7Lhemt1gBNgHhAmdUioIYx0fpzcnzuhwqs4zH51jdAXH
PU3S8K0B/J5Gty8ttFjVJwRIoxIqhWdYqBDiUuGzr/SoWf0A03jx+7IJtD5tY/voAJ5g3LhC8YQt
AWy8nfe7i7XNQN6Y3WxajBwMrXsrAH821hCM6aadbQ0v9Rva24HNcIHmfKUDspzFekOzU9yGfpW0
fWulISNFKBsu0+/BoJRhSZ+oJMcibfGGrXXNCQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ufS+qjgKdn2oE3oh7EcYzivo13DkHjOXZdvg+7gUZzbjFQGb+M3QU6lNcH0LrOEXll22KbI2ohfG
TzYR0mnCNIzsPfjq3uw6taFIWJM74+oLYtSXEeuY6ANmuCGlqaVPg2smc7PFDAPdH082wsWirRmd
5thR9q4u83J5L0asBhDI9ZTgri+q5MwrlbJ05yQiFPUliJgl6amNWt26C09sTCAwIMPW69iBKeeW
4vt5DSJ6XyglFS9MDI6DvF+Cy8vysZSNzc8P7lm9H64JZqo1p7yTgGY0TjifISAPXC1fHwrwfQXY
BsZz6suWdJqjyzpfb60JVTQ+/k5D70Xj1MXLQA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TI2B3m1FrAeKaU6k30ykyHfDnWZXVLw3GYVFmPwE7PU79Tu2R5dzZ8wRPsdfoPSTye6ipaIAsPtr
CwCMHFOrInoC4tES+00nqn8BAlNtkgIns4JutCAsylfO0tbo1jdQM1s3ZfLRmzO8TErqp7qh34cJ
cDScSpPoqwYzQG0FgIs=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pRy8ixMxliZyP9cGiEmLhkLpE8BPUs0NUJLS9EUfKEgqPIYh3TC0iGkIkNMUl3FvP77e0IxaktFA
/jqS+a9b+rZb/lQQUSJMP1pPdZyeKNO5EYTlJkeq4M/QPt/jHeYrB9fa/fTRWFaLSO4suMctHSMB
vZbG6s1wo4stlPecixWiLDS8vMBqt9xY7MLA6d9rFSok/TUkwwve+vf4FZtQpUFEhypIh+/V1Yj2
bwgtk5lfZpX3tS8eSCYcpYqNluL129jpVqEYjJIDkcuxvvuRJPiKMpRwiViOhJULCVRU7pAOu9+4
kiLxod5VBhsHJGbgGwc1XTZvGawHjedADbu7Tg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 124208)
`protect data_block
BdDPRRtvSzwYWfGSxnubswSuuS6tvYxOofcilQz8x65cz3G8BIh2R6YAbMUCvR6427zxSZ77LuIP
ULN0CKPX7KgM9S3ydzEbVtuLoWlmhob1ouikP3r/TjuFnA7dUspak4D6ZB/fS2NudeW5w0Kuwfrs
GPhKAHaWk1X0yj250MCv+a7U4xu7GSaulvfutN+c6ZP+0KHiyGl9Pw8nLWfP7hAtnz5vM8/PfpJZ
8+qXuvUCwUAhL6CPc/OYn9Z0cwynZS6PlYuvS/Wu+5kBmPyhkNC/ADtCGE7gKvJkpUa5xK0ZniCe
o5RBWWJX5NZQ7JIewVxqB6B5YZLI0x4H5ZeUG/FBc9+9mR5qlzd14/uo3ctqbJaQOngEaGXYHvpZ
MpEqSH0MOlzR1iXm4opLttyx8OKN/YG51uVqhsVyJ9w5fyrwCdPE5IoYYy+corrP4y+flwFdk4sh
oY2bhrkNG2diK5aQLqxVyaqmx0CIz3bZSqcebNRCXx/BpYgPNZzHILCC7x9oNXZ9tWu1AWpniWtG
ldw/K5N+5W1pc2plnS0qVYW19FTDs8LTDA0rFY5AVfLzPAL8qrAfv+Lll6+XUpmAHTdb2frfqERD
JsrdVTaZ0wwtVbSBWVXhM5K/aWmX99OykVJCxUM6ArLz3UDVDkvU1iwTuGg7FrSerXAkhwLod5w3
zx3UPd1//uIlPMm6EqSmNeK0mltq723saIlhDGMCe/52GatCHi4Rfh/chxEKc+q7bSgxe7OaCsgW
N+bzqMOCiU9g6rM0aMUubgmOf013BrjXck2oQL8D/bBFdYt9GwhpNjBk7XWdvx5qpLBYFQJrPPBi
7Q/ltYIs6bk8xe0dJhRmK+mCWepLielhIDM7+QifUYf/3FqNP57lVdUF5BE9VUS24IXeIUQY/bPV
Go02o5J1vai8TY5aVGeVMZAETvm4J383pobTgWF98+hyoajSQo+2EltPBiuLMqRTEQVMhoUEyp7Q
fbW4Eqyv/qrv360awU+YTWrrtZzXJiM8FXN2BTDk+3gLyocNkIizHhCTvIT0Nh3mb0o/dQlfRgBs
85UcNzaWAZTHGluKUzXzuuZg+Z6J1JI0g1ADBwkMkygUzopZvCr/BRzJaJofOXtwhNzbccglPusp
dFS/YFxypq5crMm0ixcASbmZhBLtUUrBGqIaQ6+bMPKPM0e6dLS/lci9xLvp0Ae5+UifAuWjI5Z9
f04qZq4RnRnQeG8zbtmkosDb+Ix8OyiCb6eDMkHX8bNPMLBAix41qdtSfDMtI0dvQed0rUexzBhA
k3Kfb6fgSGM4a+ajtmUCLFYUZmd+5mOhEw+8JzNl/pBuOlA+QB4HMhD3ySspJwIgy/mSnINcWfep
VAiT+JxQNhOE3CeEu2u4mLLsJSTDWreWjS2xYaz0TL/iSNfSAy6GhsGIEehQWBtlAg8BXVviy0lz
Fvh9hAIiSWvTzbp/m1toJ4yfjCg+uhPf9w5McX1EBvk+vbLydQNmaEsP7U+KEnPJ7PwEHBTsVv7l
cCkiaB6DB0PHr8WUdvHVfKD7O+hfaJST445QnTSKcDSaJP8iJzOyLz0sA7DvFzIuOW96v77ujsrJ
VfZlqmN8jL4UnQHhsHLhAFu/xBXAyVKMvdJyXvck3qI6KG4Qe4gmtKUgb7wysNoPzBR2U0E59Ue+
djE4MXXyarjaXHKz/LSi8DBalwwYdEFQSbvEWEmN0o9K57qx3gmuFr+YPf9Js4UkTH0M+sa99GVM
YJfa7XboWSn2xnZv6ktJ6FXzhTNtKQlW+M7HCiDUdm0/K713TWtuSywzHpxi/sArzMeaYdsg7xW+
1KN4HLwiVxU4MljDfR503SDla3CrmVGVQ9It2+RFWs45QF07b2tVE5RcWkJcFHs7bmaXhCOyVLhW
Mw+Iud9ZwaIWy+XQ2wlAofD3Hs9hoAeeqIXWufFC9eScqNfLO8ya4QYIHWpqqgm4X6ILwb17RrSO
Gt3MeQ8RpMQp6RiS0ed7DEIljxagLKo4KAaD9HbvXDDOAZpcL9+Oo7D8U/Casn6CWp3Tq9hTCSLm
T+jlYlr31FGdRxfN4NOf/tJ0JhxfWbweuDdpUQE/Lex8V8TMlGnJdN7h9TXWpNNDKHcD5RyzH3tq
tI+y5NIcAkwKY4hc1aWWUXWHKPA6PtWbnPt8VMS47lnnlVQb74758KLqzn1Zay4m//UeAJn3G2Hf
QjAjJljRucGoT9nXvgy0yWiKsOUVUvTfFYtVRs8/YJLuZv1fP0FCpEhktUxhq9q3QheoXxM1JUv0
OUdLLIGWocjWO8M7gd6kpeEkXJrdiJROmoYGlQX1zkGlPU4D2CVrgkb8o6UyrMq/NmYC6DNBYg/N
Ze9bclDB8sJGdBx6w7IY3hGQDnFmwAKLErniG7hOpby4BjB2ah+PS4ICZ2OZazWn6VbQKc5U7Obc
y/fKNGYUKwnDe7Eqcj98/X9SdK7WNnV8wneEA7oAzA4ybgQtJ5c/vx6vMQPmLApMSJn43QVsQp/g
8P+M8V7xpdhUhsRcLgMxUUud7cq/8vx/GxKQ7FyCbNSs8Yvl0jUEaz98R+MdZQNeHYOS3qhG7nCB
Ge4VpyJVBlE2XST/xo9uAdo3V2Ewkz6tHcUZTulS5LvgCStXkEwtW24ZoKNqySg5wbpxCAsLzpJ3
83wdGSfXLQBecpMhduxMRPT/yBdSOnR8Fv4ogLvQGERvsItOjIvMViTj6c/PkQbRtvRaOETmA4qR
yGhguHdtdSgYE3FA2bD66cAoZZpPwAxkQTy5nzStY/83xA5EhBKIsjGh0sMiTW3GEySsUub+BmLc
ld000oRNzc7Q/plEoFy9IVe6kGAZqXafQ238umGvhqisDoUTn8VgedwiMJO7bnLAZmLf+95jmUGY
fWbMZYT63m2WZRO+fPK5CHS54rBVatVTsDYwP1A/4U5KtDqKEAf2Nvp+FxNZ2nQu89g3iQ35MotM
F5b3bacEuUIBPuzsHgt4ZRhKCA34o2iDs0KFf/zE48KPC+uYbcehAnohDnz0CZpj8F097qCf60P8
NCOK2NdVSfbWBO7vwBVk6cb2OZx4sItD4VMH+KajIAU2QQcO69jqg+pTCaDVAvCj8TkiiYJDVVRl
Maxp7W82I3RJ+I63i90j1yppNRSPhi/o8xeeGoR0wNbfZZKCBI3Bul74AFoh7nvWcTnPOOgM87kj
l68Cr16YzmIxryyd3nT8oR/OuTXUwN1uJpAsyQmwn4e351wYdfkdY0xpwsaPrKH/kzD7bLaKSPkV
p3Ox088C6KDb6XL7vy2tEvgzdkcSzf42rTzey2tNOgmOMfGQh+SMQX6RyhiZJGNHdbAn0NgYob1l
zya9v1V+SVMWrmrRFgSyFhf5BvROSnN0zZJO2N6NvKlbR6yFfT2DDnhWVBk1QAvzfLfEZ+1j8wWx
QcIyhSpi6uSIY3RfJ3pwUQTA34lIvav/Fk42q8gTxt+eayn6s5tiEkZtWIBxSjF0+eMmQ9NYH4y5
UNQJZPEGBXR88muvD90HR3oCgopS8K6MWhNdQ0yioA/+ghYFnXq3SbbyhX7knrmReRIEpOuLXPqF
TurfO9Ryh9+vgDSpwR0ZmYDo6N2HAp5MDYOjiGD1k/2EOLI4OTzY2OdwSAcNQ6MrOOmV8nJ6nXh1
UYpun8sWZqvhYPVo9qXMdyntkM0hafxylXKfMPklAl6W38Dpy/zo1xyNJ/KHyxt1oktPwQSseH/l
vFkYAGd3tmXe3s2tRz1oEB4Oi5pcDVYpb1wUtCvVPTEhclB4cx1/7iQVizPDEuh84yKwezGPxryj
h45eFyipcsTt8NT8VEcwLhdZ4OZFiwSe178qZH51r5sJw8wBN2vWNgQ4duv6vXEsP0iUOhAm0NWw
LoV4+sZSE4fjPA2I3U/WGFyj7HdJmFYxnnGG/o9i2kdAMD5LjRraw59B4rp8ECt5fnoZbf8e1Uc+
GhaSdA7u8AC/0gChradtnz/9ka7UZzzvHGXM5KcgMWcGqHbdQqqEj1Hh7u5ADEaBAtgdKFyAEWE4
l/4HyiAkWOcbLK2+Mc3CdgxREQvWL4lwV1pWDR5BiVPaekfiqB5gu4FdcpJtFNo479zG1wyL5u9v
xo2gMvktxM6rNHAGDgkFIgg/yc7WiD3aFox2UN4bhfrQI58QD9FDuTCamoCMu2eLnB6zLrRrGBMv
Ra1IyejCoZr0dnI4rN0z3Aeba8NaaRPIRG7A1BdizAhua/qGK0hFQKDZdrx3zVV9HzDAuHlogLmy
6jvhALY1OOqm5eF/Ev7D2pnff0hDiHasrHrioCMTHK2CAsRfVfs4xKv3RN6U9hADfD+DYN7LRA9h
xnyvbpmqhIoGWyqJPGxebFgy0yIAa6HFoYGID5pV0X/5iEBFuYqZveNGM0ylWS4wUI2tQb9nGmDo
CASYe07m8zo7o/EUPdjEwBHep+AefFg6TFYIuIfIpUIhQ/tv8FOIjDOHlf4t9eWUemwtdGEmtJ/q
bfRxk+b4/3lR1WxW60L7XuahClLA7WEJxe0baQIoppwCtkdvWTNLfR/heuSjLIQNEvQixCP4iput
qAplWbY/YyMPfuPF7hZko1kzOalfAh/xBZu0c0G53vIUKfgr6ZoudGm4z6NcM4l9/nlkIjbIADDv
JM+76QiKacB1AhV+TVkcGv3S1uT/pkVHZGnNMFMnSwxoH/C/I1owy4Wtcu/0qksGF/zJgj+Mp/sh
AzTpqCmxeRPHvuO43QD/MGPhcgqUc/JWGhlxmD/Zf8fzPG5IMn5denTxi3BiAmdx2gDQZ5XI34Lf
4HZrkWamVl/RKOGlgJ9FGoKxAr6dsccHyaTwsZuaxNV8mO6TU2s7XpcFFSUei8dVKgHF0zUMr5T2
Mpjw6PrucU+HS+0R3VnXtcOofsiwl6d6CN8mrz71vfSy4wdAk+CN8J47K8ue4Jy1aYiWJG0a+Efv
pIE4kwZZw3ZDNouuLU63PedEk5tvwkldry6wb6o5hXpXwjPDJPAEsADKn+axSQa5cXbRptRzrRKQ
N5kNMR48T6+sqaqVjzZ9m7tEnNUksn+1y9RpiExFWHbRk/XiNQmt82t1gpRw//Pq5AQc9iIxDUiC
vEG5f8G9UArJVvtb4yqnGA27KojX1+cpN/dd81A/LnVf5KtwUYO5uVJtamX9B63Fl8sTxUZONpCG
4rsA8vlLwj+nc39Adgr9gI/RIJNhf6yaoRE9+BMFZzR1oi67y3Z+qhQ1lFEPqGNYKu7N6b0CCrVu
TuFxQBUACey0ANhipR/1Hn2KXJ2/I//s0EfXE3gfAv3iW6pNVPQRyDnhGopIDqWaZVeq2mfXxS/R
ca3I9wQqDX1x5AiHx0z63EIOKcwn1XX2vM2u1jo7/vb1WC1/LZpPw0eApJ6MXlIeDLq4vz9arp+b
tiMhlIbJAK0pGNHaG3VfHbt6pjlKjDDTutXDMYyDpqCJiATYR9U+hY/ZXOpmZ0YCaeTRviqFr9qI
Z6XExBB85i4te3ApKl9L3mkPhxW/WHrD1XteRIX1qaaly0EcYzljpFFq1I62tAqWuG2Xqr4imTGA
LUKZieltbxAk+U+ITRf6bKEEqZbhFdxYU8Oq4rEKTur+IDlmmO4xxlOhAOc5+QS52pDS3/kZc+l6
2hWx3zwxJdT1IUKSmpWrftwyFJAwvs6ca05OGbKCOv77g+qCR6yPgj3z9JOazo/tJMrhOjD9XYdq
r/U2wr22phND9MKqsqY0Ku8w+8fvY2lDPbn5N53R5z1iqJtlwFPNx1mHUDnSk4iKJKcXVGpzJL8J
H8WwZn3FVJKEqf9pRDq2R0ny7DGEh3DC6fnCTuaydPk5B90J6wmpoZjPHPCOunRRyIgT/Zj41s3E
w4sXfiv0Lr+gc3AmiHh1S5rICeD7A9xJnjZoUAyd8fQJHI0jmMJg/lIPfA4IsaHgEqV2KHOVrdCS
tN7QdQvwvSSn9SNhPdot2R9LJer5kvhYnbv7oSy1AAgUlA8BKvYUMU4k6LA8jiKyD2MO1WiomMEZ
e95t1e4EybRSqSJrNB+RtB+N2JMW5c717VrmmhAHPsy3Q+y89bnu9IW/s5fic6aEiGBpJUJJK4T6
nuzFO/to+8oAFuqr4HInbv3pRV8V2f3J30LbMaCOkjq0dzwGxc96nKN0hfvmZNGwGsfHSUhrFR7p
3CdCkzF+SfgwxfKzhJxA7QTZXf/UqI6Iba+h8pJs+4KKfsAFPDdiSNDtymWNUSlDOC3eHLUxyaSm
9GRu2G+pCR29wbdWeod4mraMGZn/4jgvu5RvXkhb9PcpWEJZNZBqpzZtscYM183g+LKhfYLf5V6/
Kj2FbIHNrV5vjFHKDZMu16bCnfFnlzmCBd9TwrwOosztHPOv+ARmC1PBRZgcfDH2MWNbuM1UaQ9h
Bp87QgJW5GlqyqCJtHS0dT37VwWualAvsrUvgmdyCTGwmz07maRma4q7FS886tIEcfevoGzRer11
V02vWgIawpBY6peNLGM80//qIwAabTs6SIbH/en9nEjHPd4okTmL12Tmq9tPrhUcjj67WDALHsaw
FrRiPtWPMnQi2IWwraP8h6tP9v16KcIujqeRLlLCtf1wMwlTCrJTX2PFV+HDhkOxpyk/D1Zh99Hk
BCV27ywbI5MVTYnsoP/s3ey8REINichVltJuooLKl05XPXq/PdxGSISNOwusaLcAiT0Qt61UjFXb
tktsl7yc/pueUWWlT+ovhCLvB1ebzjSR4cEn2l+SpwHEd80iFD1yiZsg8pMjRakIalJxOYyrO6H1
ki9kkAIyFYbVRAeh0FIthwBSE4PFd8HFvu/+5tTFyMuoJFf2iW8mPdzWB+aAEgebODJyb19WVMI/
Z2d2UVEy0sPSqCrNLQffFcMarL0Gt4KcSf3xYmxAUnVCgfgLqb6iOrrBvRVjmSNM28K5iP1TnwPW
UMzzOD1iBrJxZpzpdmTm+ikcX/eqI/CNrB/eD+NBZXuw5vs75HNF6JGTJfT1rTyXeJFLCyejLWo/
FoR2XS8+jAAUs6OSWBHvtWMFsoh2YaecxxkwpuR5hO0qPvInldk8C9DugYtRllkFG12X2WPfdMTW
q7ieClyuV13VaRazuBQhs8rv2FOHseP94oOJkzY/Az/isxJ/C/YqQ7hmFCUJ5kgTbartFmLvrGXA
WAc/PWPoSo8udP7+iZyANylGQw7mQSigJzxkc0+EpUJGuA5y/ZCEbO/bn7b24LBRuyn0ytz1Zj/I
5O4bTQkTimAkthJSc84zgvONUKxH0ZNPTOYcQV2a/Xo1VQQ5IRY28dLVGYbEAlg3OMZKjxa5AsJJ
Qs8/t8WnSLLgB5DXkbKFml1mv3lfxJbK+MmxEEUng3PpNJzIImied/wYZZFmFjataNZycfpMiMir
BJHQlb8Naw4Ci3jXnzhUpA2i+YrITiJC0milkOSocKIGHz5vZ9G0ZLVG5+k/22FuxLQCJOj1kjE5
1puGZcrXRUgN6aq8Pf20ptqJrvVDCqmL+GXTT5etNhawEg9MzrTRT+WkBKecR+8Pxcwtlkig61+5
x19ySId+wQvvHGJiEThcgMr2DRoCxmWR2S3u9p4SwNUK45sJNgLHAT9gpU5A9qPpRlno6/3sjAB2
qRj6XECjipQd3zWJc1i9KdTLZihDtJII5yogOBDdPg/pt47yeYi2H80uIB47PZaVIsg3akbyLVxh
+rdc/NbEQydLyh24gaPr6UtQ7P2qtiOlS2T1IX55DwQ1/3FYXpgn74ijnA0mNqQGta2AJzWoGmOL
zF8rb46xo2TAb5RdoVg3cQ/YBiNsH6sVHtUd/q6UyANP4LCEmOpVkY6IZiTJQaRNIGZpr/ZpMLcX
A89Zd3rkRW7QPVm7bG+XNO5CCVDTReJxT/jBF/JZrcH5zI4zeyyrcv0FqB4NFFvQKTacTXj/2vyR
zNq+Am7gw/DNBoN6midVjYmeTwFMIM6CXGDl9eI5e3yjefJbu7ayTqwnTwX9yYSLu21PQuyoihah
2tfYOjj6Qq7bx0jPaRdeEAIq3GM67JJVukdIWBr9VqiYsGrY1Uea00Vp1y5em/rUDlolz+XbreYB
2H6Lz/rLQTjOFYhGctk+YuCsTnYcjmHe7ydwoEMFxYmhyFxonBwFWNZDk9b/uIaXl5sfYiv2XbBz
f470UVqJF2B59J5h+uZBQSQs9+5SyP4b/7vcbtzenGLEOXDizTDTETeN74pCo7ziouuBiyt/NGp0
q+HDAtE1emBIz8qPUPOeyXXolbXObuKbiPNfwdzjnNqIsJSBp/PvlUQxhRAghVixZ9g/JFaxls0W
AZrsvfrvgZIVpQfTPf43ZtC6laY1Zef9AFOprSBXA4+kUHd2CPJnGuve3cnBdQSnO53OSx2tHabf
9ymhJuHai2KHBmOiOrn2Quq1lV3nbgtXQ2i7jcKYzofWCXCuJ9f5STao/bMCz0ZqafQ6xeJfvsN2
e/sPZz7Wfz6PuLw5JaLnp94njJBQOgcVtlECRhJcFuT2TYkTJ0MwcSN3rU9R4rA8AK70t21rdlZ4
18xMBuG+wcgD8lsVZTw3zzEz/cyoN1Fte11ISH1dLS7LM7DZE62UmUL10QbyhlQ4Mrx+Zkv6ut5V
GjGcBCeMaaAo0zejDFYiEUzAY9dRlkzAJOqLkXoLFSNo+EGLPpGv0F5bOySkin+cX8DLinsBIOV1
XwYd+ipY8mUTCVvd/cpNkG5mdnAED7Q9d0kYUudzyp/ZDYDcNU1adkgPIDI8F2PqXbOFkusjiZix
t9PM427KUsc6l5c0RENd5wQDE5KYnNhp38RgkK9QqCIpjxF6lqULFrQ90b1FXR+7Shyydh10wDCy
DYr5h8/lv4oIw2BQR7unGwHUyyfCDVSN4guFTnCZHSyLEO9IzNAobbeS8S6AkeaE71fhQUavLXUX
nO0qzgTE1emFiHBciBXLo5C2f4ceVZHm5dVO8+sMPlBxcCrI2pvfcfHhweUZJjBQHwA0E4aFvlKW
OU65k0kQccJnoKGgOE0VfZZ3QJ8In1/IE92qjh1REFKCfl9ReH+8pa0IG0gFLt/PYFH0YvVwp/r1
wcnbCk74S3m3wiz8wenv+W3U5tMxZlnvP4LcwpbOw8aBJXFB2CXfPFVoel75Z+Kz4/61OH+7IWWn
2CP3nSGIhjcOaeTl0jLnRswC68hc366TPzvE21ZkR1lzR5Ds8+wSkE9WOupCOQ7+LepALs5n2YN4
ZtCX2AHA7yduG2ZmcrX0vBcKVqTmmsjM0zWD5uD+jBrxPX5xsb7AVldhhRNVicZKaDPUHUyIDtSU
6n2qW0ig4mPdkXf5lZhwHxpKEPq4Hd95PEKE65Q9nC/HFpQ1AaY1AKDQ3PXmDUumxEiuYn1C6hnP
cTCLwmhutwEi6X9iKLmz7K47eqphKm6l8AnwsIfJAzsnKf2nC8dxs1k9WtuFsj5wIeJk/82DwPjk
2qd+jSBlnebpkuucLCZitxiTypJCW8aAZv/A7UPQxa1K8mvfsFajOQ8rR+yLlHtWNxZg14DHbDHh
eQV5XD4eqaLnT/LMBSenfLDkCm7KZ7Jqo0hv/7TSKw73IniDMFZkHR0yOoyr1WU4HYQK9r+IhLrW
XE0/Ll/2U5PXoZEwl1f7kAh3MYi9u5ON2wNjYVfwuXl5Bwk42WGUyInpswMCxTGRqEXIEJmEfr7X
mncVgjaWvAXNcFRNgtediYxVLE/NBfBsiIOPHwFrirHIQBYmptH4Q/XS4wqT8sekQs7rjsaV4JB6
YLoYpWCdTfgzWo06t4jpGe3GGXVBQA1OkxcVY07br/X/3mBdIqd1h/0ABitrxYyD5ejxQ2XPLBi3
VN+6FbhL/RtKKrSssX9S6ZGkpUFNmrCIOINGI3pyhPGIAXgT2iJ48/KGPCX1/rlHWZm5PFQWiPoO
F2LZb9e0ZUPcBUAEFlO0dSHLXdqpts0IEcqALLCj0u2qkTR6QVeNKNyy9SlLE2XBB0tcK76vqjT5
VQ++2EydVITbqxwYIy28jCcDezGoqnK6arNYCG7pVPsRMTqb0XzPT5yJ3utNY5KlVUzkqWjgTxdy
iMUcfUWhSbW7JMIOUeQE2OPSZFuHIUIfjpWzaZMK9aUts/Soul2OCCvrRVMzaV5IicnMUNjwALlw
PZMgkP5JQ5ffphdySTpko68zBHScxidn7SAYBanYAh4aCTcA9Z2/45rOGTBQVDpTTY+WTtO9XU7x
tL25K2yaWsvJnnQArTLEFprK0vxvq5VG/WPUwTeqPT7XR8Jn5js20tlyevPvdLtk/hwSeM+tzgbd
x+ialVfqgMkpKLVl0zM2LVf9bXMLzfBEDpIhy30UY95w5oc/gNl3FT0Fo4bpKv4EnA+HCvfY/riu
9LTEIPNzerMThVcHhlneBow4mcEqTWZZL50PkWDoAvw/kzL5wwz5Ptf8DPGeSG1QeBNqioU/msD7
4LYfppV4a6y/ia2u9oTmW/y8Fj4mXwpKTbcQKKm+fPUxusC0jJa3rFLz3SIbOYeVguDz1GcAaUvt
NEmYF6VJGg3iZ7kisrya1NcraOEsTqc5bAxRimf1C5KgUMDTbwL37/7Y5KStD12ydgAUD3IyHlRW
ic/IHp5tmK035hzizybpzaju+dsCG8r4KjP2Zaj8bzZCa4I9PvX+e3OyFCMOIqdn9Uo1xNr61oYp
MvgFMk7auCK1RKLkGsXrnVez5v9MxvSNKIEC764gdwdUcgx26x4yPtce83tBYCTHgkgXHJSvzqf7
iqtPkPG+VN5J/9mKoOPPFMVoX8HD36KW3iZWa7T4VHQ3pETxWX9/2GiufuVxHfXryAR0Ckdj/ql/
1GKf7lBQeqqRPxwDWMF7M2Knxni0T+N+ojaUa5kUaHDxPJnV3A49PymVs9cWp4i6qUM2+kBtm322
g3EELu66353BJ9ExTt7077R4K37Yf3ComTPzHk1IDAISV6f1prSNj9eSA06NSmJdjkTcFs0PPj//
EZHkl/AcLWOJT8PvmHwspfNGKW5/0YsqlJcukvz22daB1sSyt6POyYsZKWElvzy/mJV06MUzYbZR
n9iLvWdvJU1Y6P5Im7hJ8Cpje1OGhj2M5PXKRM9ZFRmkAziIMSPIUkX4suehpp5OS75pzW2p4EUf
bOsvRQHlkOd4sVlNY25vPth7AavjwVAaEOk9quFnq/6qmbXjJ9Sd72FU7/c5OSU4jyGVsU5sgmLa
/Rbt9hmfG9DZOpG0/uQFOsAk6HeDqUIziVv52GhbuR4Rin7u9fUAttBmjqeKqFKQMvuwFbfeb4RN
m+B/kBJmyf3jKY9NhkcjPqaOKAu4/57Q1GXMCMCNF7XZzAluRs4pY3IUPp7xX+Yg4ae2O/Ap3eQ4
QRGrWqx08tqdaZQxiLsr0QnSyCt69jmzJ8Hot7+7GIe5eSkqY5GPui3p2hfCcKpj/5jZOTW+wLGg
8PgH3loI+EJPnU/BGkY67MxG83xVJVEML/gBOHjJQ7kHkswiHHbu7XfQBBuLqJwn6jDNvDvfdwsy
2Rd5FYYLCzEHrXo1MOHb6nOnMmKjjrLwh/UyCmYGQDM3Cl3nzdgM24hnu7MHBwmPbZDLjQEPaF7E
5xS+9SJv2+jJjYMw9/mo3fCjMkzissPb1BHaMiE7YyBKbrd2uzFMf3DP9t5o4hHJv9oBygwXia8J
0/im4/Kt3SZ+tXZWDwn8420Dh9gNfbsYqoaoG20Eld4w9CASUA6FnU6P9Qk33NNRG8crGrTZH0Bp
Z2G7d7hnRzdESDR+fbLkDOsOP3LYeecTmEMP5mEpHlApx4EAblldNU0viFoOHw7QJbfvgGIhk2ij
i6KHIqchyk07HKNd2JSrenpiyiX0eXKMZZHt3E//exR3omjx5XeT2pN1S0K2gFfXET3tmnZgWaXY
3yuf4Q67E3Qu8RHFeYdjUOJs8xwtvg2GHOyvXTCCRAo8cJR7AcZ1tghgKqC/mRGOqHmPkJ/+su6J
fw+N0FcIABl8ADm5gC9WI/ljAjh3L6EBf52Q6trel8xfidv8Ka75EfE0VroFLj+j9RJprpqdWbQx
dn8Pt2AnRQCMIagmWRxnkI2asVTB7ZMhcMxMCtav/5Ru2W/K8ZiWmoNKf4eS3YEHSdZMlNtE/Ftm
b7xW8TqbtmXhPgkN/6CLST0MbaPFlCawmzmgGJ+D8ooW4SPsrT3ezoXHMjCZgfVim+DjzIuNlhLq
X8w3wJYOCD1yMnE3Q6CSkuJS7dO8a12mOzuw9ptHEx95n6moqcNaz+bAy/tikCEuSxEVuboMSuxf
Sl5FpYTUZSGn+1eD66byeL9H3O30ZJqfHfmMJHQ7LdspNEox887VxpjZSz+Llzv07ygUlkbC5ij+
zNjwlQJenrr0rjtSbH6oRCY7VG/NP602MVy4dcnOWYrWV0zIJNUAQmyPrPPw7rEgUB4we2kSBf1j
IMSoKdIo53m1jsDCtRROQ8a188wD461uBuvSNcRlxH1/jheKQ2rkLdhaq0bPdNvE2WZYkAnLO+cU
eGtL09Q45KcYiIywC6GXGTa8uUzD4GLcr7MiITXaydgnLs1zMxvWyVs1XvRtYZVqwmvPQp3moBVj
LlMmGbuuJL35APeX1Siu9ou+FmMjiRah7C2wiALZaxVnPtbF+26dbsHNY8PQ+jJshhlatf8cuLna
c2joXPju+XM8cLtEvKPTlYeFqy5tCmScTWXEYZKN6xs74L3SQ3/YjTum2Kb/jKIiUPQDJn0UV60U
1kxitk1OjgHd3tvpAPREhx6eTWgcYN4VRj+Eai0Fr3flPyDy1aIoHJDSYHy0S0w5RrU5GB2bOE+F
RUfmHIP2OeJD6YVykFTg5WYsYGFNXFgJU/cINx97igvkXigKhdSbO13P3GTHvqv244I3ByZra8/1
E8vF26vsiiBXE3Ek715ZuWaz2H1JQYrb9X1GUgeQ4Gldz1lPTE/Snijrv9+/Y9K2LXdzU/l24NMD
g591NRKBFauyatIOBCBFqVkseR7J6GlgDhofwMgA2lUm4FNw/exKyYhmVpjb3c1X9GzgupSFf64K
wR2rrrzNtD8O6iy8KZJkV3ATBwaEGEs+ywk+QvjTzyzegYFLa5cwphvS/4Gm6xYblJTN0cTOkJBQ
NFSEvfZvqSXKbwH69pEFJ14M1J68tCY9XBsN5Rwu7ayPaEyYEsln17t4+1/Gay7I2Vx11Topxfcr
d/Xk+VkC6HdAtBuKO3YLqvfvBzeMFxjw3X/OFQzBd+49TvaUHG26tnsaaLW3F7vYdXGiUNO2H6E/
00J72qfCNOoupc/1x43QXhWsGIcOgNvjIgDF8OfZBARLm1Kb3Y5o/9QEtiEh2rTgXC+Mi/CtjRZm
z1iPQKAxDnvj0cdWyxfPqhKtsdHLgsSzkimy+fouKwQ0Jm0tYk5iDWz1OJioXks2c9pn0QdXiv2o
WIwfuLatQ5T8YGY1mUphO+/pthGRIH+d1cyLL3XjmUXccfquIO7uOSTt8Yx4rZca3FBSoUCSzRxL
tiEZ3Yq3wtT/40ykOLWA5SlcJGE+m+VLohZBQ4ncGn7zK4VJdGKKfrkdz3cq1LP8dOYh+2iy8bO5
8zpefb9Nw09lmGl2El4TFvwNOcZdDnt5If/vJw8RAAlpfsQujGQp7pAO9QHjpnZdCTwu3X+xjbl9
KZjM8WZ+5Rp1Kcldd8hH7sNpak3/aXGRVkJIs8IqiPhMCxwaT5r+KJQg6iQM8GirfeljRSDs/aYr
ukMaaydJsx5TdshVGxjzWVLYneWNERDalWMKM2Jt8BhpoISTzec+IpYbMNAdnzcjoOeSVOQtRqlD
P/R6JGnlhcJxStC9StrJGMxyQU69CoDkv2LYXhcQwF4zpl5/8w/0g+emFT7ZJ7O1jEiDYIGjQSCE
twlBFGNnBQIMM0YmG27V+IKBQWElOuA8dZaOI9S4GrLjfPBrjlV68fYuQ9nl7E4jYGD7fTIlBw0m
KYCU54+cdEX3MlFUv7bIe3J8/aw6zr2HSzDatLFwwUts1k8rBC7gAXyTRPU4RezZxfmImf8t8fTH
FzhcOi/4WnTMX09UjOX4Ic92wr6FLr49vZC0kG+VCqpRlPzeiFSB/fiHR9NCPpHXcFI/VWpYaf2l
3GWTXFDVz07lXEvP7SiBVc3owBnBXM5TwwM7TErc99ytqTuRmQ3hVcNMhwQKNG8jwEGtR4K8IdTg
Rl6MfxMqL6bHBXTZh2/Hu+1dVXKQ7Fsi7rgcynNTFlhHfPO8XKkQXlO/475fYZQdoD+SIGw6V0tD
a+K0xkjw+vxoYbAnmbjfVRUuITm7IpWWNYUvpEiDDFl61TL2GORPmVEzP4+ijqqVI8UgV5TX9dWL
kWarI8SNFy/jQXdHSyxMpUpEl6t7MuQjlDtzdA2LIvhp90tp5a0aJ2yMIcBQ3rG30cTEFr8mVjwR
K8p0gZd41Q7s9t1zqOlHo5dePobAnb2h18+P/6ffklNwLSLAUXWI9wlScV+f+pIYgtvMyYcEbSHv
GXXbMDELlFKFO3/tywi8pdbJkD/Qx4P2EfmrxGfEyjzW4y/LFGEGMzXJAwvTN7Vpogb4vIRYXedJ
CGMPoYi3o1qxmFShZ1pnxdi3Uk9RyGbg4RPSlxhz8VZrc8yAqKMi4pRXh8BvNY9GkagJDIuAVlZw
1cFQx/7Oguzrcg5QOtPavJqyqvIAdygIktvdWCaP7qugY6K0g0u4cMOe7mF8v+011ny97zFirWHa
hDa5khLCVYZvqgpnBk/ESuZr+8vCceDeXgfNUvLrY7mnR1eTj0p7+oGosrdBasZfiLKkXNSPJsJe
zejcd7h0YarvWIDY6Ed6y2y3js0Js9FhC51GyZGesueLZI5AAcE802IbHLs1d9uZwMxLznhQo8lr
a4xXcCcUS+8KJJNoS7oHs6mXiWfxuYaJRdAiFgBpZut8pTrGTxxU47z4EMBv3JtdwMGquZEwXEu0
PTtQvVDbmS2feEz2qOqHtl8sxn0KNWRkS6nt1jhE0oyMmx9Khr0zVLb/UMnralYKM+dt+Y9l1Ezj
qhS6Ox8RZ68G0eNzfRb/8p/jAbgWSJB6ZPHJecNW61tfdYQ+k+xskCDlyruIiVvKfiQGc0XCyVvk
u9nSVsloJ8O4SVy0+2wFkWE/lLfmdxtWihINSucPcsZYPxlErrpWe6K+ivu/tu2W2/+iwA4CE6d6
AfYmsjSs4ETCo/uQuZ9Nr+4D9CyBJJIwQPBAUR05/9WGDLWIV7deOfXmtAyXUGxyNdrdx2TEAjaJ
O7j81ZztnRLsFH+GymGTkHWjPVlwGy+UuoU11v5yuUr3kKwmvsYmS4Fp20X2tzTRGwpelV/Sf9JH
q5DWpbw/CgTXpWJZ5aThiuvRzhV0InNA5gU+nrvvjKtkoClHdCWtYCQL8X2S7voPAIdgJ5Nm+75g
/r4BpmkLZo9eApVeXdRTICz1PfiMzE44re3GJswKNH01oNfEXUOJu1jvUtXZREXIoHv8JOiet27b
Pw9s1XyESOuflKnKXiJk2ekxeeBivcyCQftOjoahfErE9/3FfHPBEsQObK4PO4fD5nymYmMGhNQe
4Qz+Mi040N81Vfju7tj5WTP5SjRRu+mopcniD7maeaDOyILLD+GIgLz4JjN45/XjGJBsqCgzb4lY
093rERkw8LcE9YfA6lzPMBJqRWuNP5Qm4r3CkeGg1aAjv/51weaK/Hu/QSr8+/AciLEsbQfShMwX
bLdS/6kSFJMwXmPbzO7hW3FotXjNMGyrtlu6TN1eIrx2nouQ2dEsDOK5lueWq/BDbLrpIqoItxt8
p5DZHz0waecbl5HWYPvku/uFUQzGmNnXbTGpEHUyutk2Pk7S5y5PKELS+Exn0REilF9R+ga9BmU0
dof4uXQUL4a75ZGLI2b3MSTNBOQ6pDwriu2zPgw8qjPYxS++qlO+bYUGlpgZW0I+EDMygfQziiHm
Gd82jG20e58L/nFsABm9jPNRjhvLufhH8Largm2HyrWpvVYZYZtl+TPHWjGd1/vq5Cs8+jFJdNon
6vSqd9nC3Niwg2USuKmxgXUSyosEeZ3yxC875l+s3tOkwUiXIMAnbltxk022D+xdMms+IZ1hxlhy
D3Ec1spSUzxLuEtWCK5/ac+fxyXsdAXn8LWnRUtzkQYoNpKgGsY3EbvQ4bB5zGS3QXuqj/DQuyLO
JbTelugDPEeGbUt8sS9AX5Tyn/jcqpCiuWaGIdOSxDqFkiqCHB2of9Zk0CQbRzMc9pDuv9n7mk5b
oxClxmvD2SLmrszZejhJzlSwARNP9DJXeOkk9C+q2+cmBE40altj+aalGZcHMAZ5utaBjaPMowdz
krF8cIgm9sOKw/xLWLIlOWykD5O9pRZkCxisQyl5+OLD8RTtPIP6GcZn/XDPRAsbg0fTQp7JLp77
LOOfucD4DddHHyrvqovm61CvhYD/S0iLzMQFT5591Vh0Qpr9GZ2ENxaL57zyf2pzVkgsZ918XfIg
QuWTNUtWw6S4huMKsiRaXFKxUJfQmhzW8jOPsOU0S4mvWfewtxi3WUNDeD4OMU7ScmsSvgL6cJEK
vYY+Xq6oDL5s6yA1FWAyUrwbqQUKrNNt1mnOGfu72OnczSJFrxbGGp/QQFN9HyL5cK+vkSeP3pjS
w0dWSXdsgNQAiXDbAAyVBi0QHvfLe/S29ezClXquJ3NdUYjlb/qloe7nSaFygAeFqLo/S4qhlZhA
ZiXXCEpDOjX7Nn63BguAg3rO+fit3bqL5ha7GwNk4ZFlAcIYpZDvWwff0m65TC/uFrn3VbHNTAGN
Pr8TGW+b/PS3P+GDj33nJ6RxWf4xN9x1b8nvhgcYdU0Nj8jsEbFj8x8YdbGTlks4L35XZsW+QQG9
62pfGgx3bdalY4l37c5kbI5BMCaAwxSgUMPNdBkIycL7ktRhbift7wLNoTL34/1Lhx0uk9cQaR2P
TDWVbJmM4eqF5hU6Eu4f1sF8ABX0ItWYTykwTTM3vWOZPud7T9HEYw5ZZvZtSA7CRX4aX0g82B3O
iQDy7J0T1lyhy8IfWB4Bu9qQtr/BW7qkBZXIDTvpMx1nBrF6SQR3cSYHdy3yoMkhbePy36EcInTG
isvBNiZLYZcWHqBoNaq0gYFGVNcX6XNQ7glAXc1ivsJVLteSMcCPUP/8VfLKNOPj7S6i2N3A7HE8
UynFqoqEPLIfXdSXzGNvvNpHdj0FdGeBqCS9HIH0gswlJuZTOoWcv+7+bVJvhdduC/BYUIv/v1W+
mZvoeh/FbFqYfiTKMRaA7+GcPiMKH3zAQz+L56a4IWBMeHx3SeHxYfIusVuhw5zw8kwbAfp9DvpG
pZbegHn4tbokkHmkAE0PphK1RyBa2HidpOPq4npc6xkJWT8dxydcChy5bQ3I8haccBoDfo7FV5QM
m8PMYLBZSy22W/AkVRZpsYLsdLJSqvQlrX/W04YEzX3PKv7FHvysAaPQClkrAC6M79ZsAqrUODnK
ykhNGR7AMs/i4829Bydx/NH+dzt3cW0hirlFOhKEU4c+8KL6P+d5r6ORkwnZf47lZNczXjlmXTL1
YZSolY9B4Lqm88/DIBILgVPj8gSf0AKNBPx0pcrZKTgd08afhm8xrdQIlQN3NH1nCkeMXmYLhRLo
xnLxBOWmwfleeLVAEbjGadTBQflVdS+63x7xyIc1DfFicLT9N5o7i6TNLRY/jYsR1VMjOTojw/gT
tMiiYd3EZ9+vtIfwQ9yaM3KdimnRZlyfR4hk7XhFzMbHkGf8T+2NcfYLEt0fntsIknGjCE4ZwVMU
/ExMGk0t8wLru/bhDjSaQv/nhfwhyYqnIPdzisrreHMf8zDBulp3aeHIU7HLG5PtfciSOSmcxiNG
eL3SP9vDQnpHDN6txADZMqjN7TQdVUz6PVl4zs+e/KZ5J8cTKuPRSNXTNjkL9IcKxOwRR+8WCcu3
xi1sAlcDGQSmEtEYH6L3O442Q5IdylQgq6Q6ZlDJ4gclmSSpAVfjpi1hz2BIkX2w/L2sYj/c/JVY
F89zoZQcDdLDPUrWiG/tzN4OokOyVExr/Vyy/dfNSE+JgkPV9JjCsRwuF4kyesovNuq5oT0pdKHN
PPAXnUQELbH131+ztA3mw43V4jcYdTf5ZpADsi9R5cefj3+ZcktQB+iRyVRH0wymReR72dGNkBy2
QZVzTnEzxleeQfFoq+t8OMRyZ1gkJ9G31n3SC0kF6F2VY9LT+jshc4mnK6WhqvYNwI1R4sgBBrJA
+WeGF++Hr2j/c2wrGaEJ20ZFH1XTAcINlgo/D50VZQVDdy4kr6xuLrlOIrGm5kRXHavCXCtzjJnU
gnw9Ku8c9PS+ndUAknhzqIe51jdGxlhab70wUeDgwzXBrFyD7KhlB7bVd+6/auTpjeyF+932leXN
5cLiL9JslgJKWyh608p/pCTlG/d9mW6TXtNVJlssCE2wv2SBXrJ+IaD6XMg1FGH64r+O9fcgml77
KMqAPiXLxtQkUZgFJoECjU1nmhUNM0q3x573GodNAx1HNF5tbCfV3oqsotuNVVNPNkb/k0IWzxGm
Bqtsnrzs0qgCE2cVXZHem+Bz/h91bM4nTrzzN8eBkHJpFgBztGMD9X41lIbkbqV4ocf/X76w/xsE
oCUrOS3JciMONbLNum+Ttqg7l6ZmfIIP+R5dGJHszSWAvblEzFc7cHb6BfIl5RPVtRcuuywHBd2s
wNzCO0I92z4cX2o4HnSlgzPA6S60pKvkEVa+J79LPh1cqhKaVxI5KlDFkWcBExqAP4sYohckTlKL
j64qKCGxCEX7ivyx0dElAn08AgfsGr7tFxfs8/NYp3v0k7MIOFDrmBNX1uq64ijl5Y/2lvzivq1g
BYItC3cUinyKahGIULwU5NxRoUem8n4YslXkOGB3nqG1Kpp2mhqJ4N64RQq9I5FtlXvO/mcrKhIt
i9HxPYYaMQca+DnRCoL1K/h2CfrJu+Z93UD6dPkWrnvqnhLwefjsjCp7G16DLWjb+N5dcnkz1q/e
dmCPj0eZ7TZSqNz3chEOHpHGGrZwXcsaDdf3Ui+DaDOdgPTiPwOmL5Y+evzq3Vi1HziOoqo6akOa
fH+EBzhPSOFXgF10gR45PWqNKRiqC7wvEEMHOTv4UfOHo+K6yHwazLn5VCJFrV7e8b0HaZIDr7Af
hSYmEsgLjv1seOzkS1LVd/KhlTgqvJQMuMDsrkPqaogGc/NsdEM0LLeV++XQZwfpONesR24HM92Z
tV8Awh7meCybqyE80ILjJI0r9/aChBeBoBebdMgBTxbZimzQoLoIZqFa1XRud1oPrQXEOEv0Tr4j
lSIs7oddaevc+TWMzWKIdhXz0EO8u7OZUPpg2Kb+RyYy4mCnpP24P24S8TbioDB2nKx9TvKJjNex
8VsxFC65vxqNgmcqTsPex36OjwtvgWiccIjgtcD4E2cFZDxMBoUx8CoC54rFWYtDdtlbcd0BIlxe
vEyf3kIj3QS7qEO3XQdGrO98VWPJOBLkiIEGYAXmicSr64v4ePoYkfwyxfnbGzCjRCp2aF2OLaJL
/3DhNSl5rFvhVAjZqew+eGsbJ3Bxsf132xNehfhAHsvlppRKrqHfsWJga7ooQgfRpMhop9D8/JVX
tiXHf95I5s9Kk4yZYFXD3pVd9PWsIR3uKlDBFA6lfaslYS+1vy9AK38FywIXFlW/80mWPuuTdLur
rZOoVwfsVSn1rJt8uagnYL9EPOJxIuqm27T8puAPJ++nrJLM4taJZY0kImPK9+EgkySjcGFvnzMu
nyJXiqcxOjEzrbd4C7vdSkvYMHdq2iyryjuYUPYwNM3K0+ydV8l01cSemgSvZcuTllmki0IydYbs
EEwb5QGMXJswMooNtrbxba30dAWrQpSwTsklq9yG7iiHCegW0x/6VGfYlODjB97wF3sbJPLeGaaq
mrx9B37ZlQbMHIVMwyXYPH0W31sWI4Y5I7K3KPsQN/uBpUxN/BK/1IOVMtiVDkaZ1Ausn8Im+wRy
GMO2L2g3qU/XEksjR1+NfM7LtiVD9vMdHfQTB3ovg99kotqsLR1OiBOmtkgYODYw7261FuovUpul
ZQf4fi2sh8Kns5UfEaFJrq1rfTiQgeE1GpHNdICc/3vYtpYvrOKcxrgVhchrwfkxLMFI0L/PuYP0
Tr7E1SWulqe5FbJp3Zc7Ckl+rYc9L6hBaoe1uPFYdvZTlDivNGMXXRIB7cULAjjj+lhX+KTUtfTy
tGGRp4BFTArrdTFzH5eLWbSaqCT76sTijuHcNDnj+SU7sjBs+dYFuUnnL4syLv6Sohif9nMWAW09
5tzeHFy3Ayrk/LyqqVgJn6/tPKb0SzjpDyqXiE2eD6fqZP+q6zEBcO2tVeQzqFTgeikvYWw2y6yI
2TwBw8YY4ERwi3tCp+WtS1TcscJW15SWLZdb70+0Frg3lS+ZYP4pQypQ7aPgeSIS1SHXrzo/qP5l
tq+rwXW4mWWPsrxwLZQnTO6S12K0XFXBb3l6Gn++v6zMQia4IIVAmFcGn8Wjo59PAlvNSDIgiwy5
+wWNJoh2pYXDDMW70RIv/UMCHwr/FRXkSYSgkyM87NdgMUGxIuLFbRm5nJ+arjdyGkRnw3C6rKTC
HOIfgPiPt9B8hbqJvc2wr/OigxxOVxI9sMRzbTVliq8bvhszOJlmDc+sB1jfM69NJY8qyq3GkUVP
LHn6nlhKuzJnixZujz67CjNWoEW1Yeej7lzBqOXkh/9Wd7UPOOpQw61yYUEz1yjFZ5gESq4W06NU
pPofF1GOEel2q3KNKLzv07zX9A11WBezkKeVMpOsmyBzyL3hm3/TOFEuGiWSsaGO6sXgUI3MR0h3
EwFQmtREy0RFF2CmCRW4zuJl8qaJcuksm4N2djEzqLshRNXHHkyOJNnHUdsBLFLn4k8kAr6o4okv
RHBrAzdj2Zjp8VK4G0G7S8lLjOtVJSbV7WqoBx2igoxw7AvziCaww+axcR+EHaixkxaMdknpUzLd
GKNaz3qKJdiIY9H8adABnzZc2CyDXt0nDfLyUNphHHsArUU451d4QJqlN79xbbM1OJ+FGtrTFMpA
qIGIgnECImqBejfa+VCtkmn698EZ8iRr/LJ0WSYeq6NuFP0huugHWvq60j5hhxMQOUGNSSXoamZU
Usf5UQfo+TheGUcOD3alLtXmLQ5+pQrZWQrDSiljzHXjTW0O+taAAC9g11nPHr12R03UCmFvOb6W
15apSeHuaRA+eFr1hsXN5v9ZzORN1eXBPma9Xx1peayEeuv9LL+OyWqL5ISzFuJAdVpVPDKfKLAe
UO3GbLLnO6vErPitN+cKb9adPiP2rDFkPr5Uh0n+wEHBQg+Ca5wjs0M4Icz93npZCJ1UxXyMLlyF
JQkwIXzueQq4xoqA9k8WpYNxo901cKBzQzcE+OzVg/3E2Q3m3l1no1xvBXq3Eq/T0w2fy65Fedpd
7cpnXscyE3qQyP3htaxgyyJoFBZoT13Z40xm1e/ZloMdTf1uaM4eOtJ3mcf8+UmMPM9dmuyvsnHC
UyOHFjpYuO+THXXXSRN+q1kPCfAJTjdf1qxQgSWRM6f8TceTRbg7ZtDeCknXsn+W/RFm3ZI4EHzA
u+sGI/Jrco/WPM5/JJajSKjjIct7GPeuP4RfHAvCoU5mulaRmGEBlArnrHISZ3Vbz2Xd5lQA5Sz6
6RZ+zceo+6JvP/JbmMAySIDQSLoLznJV7R7s0meocTkdXMd3Eu5XquX3FuudC3pnBmL4QhkFmN6W
/wbR3WFpv5KpzPAWb1hmKWqdqJRSzNaQu4bOMCRrdDbI1jFawmdknv7o3uagt0N7EWftUuAFfy86
EI8fWeQRFYvFfgyq21iwtrmMk85gWAFodl6aP0JIv3hR2AV79SPEUVr0f+M5xmLiyTgj3MMVEJ79
t+W1biiGM1NY3rSvRPGGuheeKW9admnwBKEZ5sYIlmKklDMt+q20ovbZPoWbgObeG421i4Npxujg
Afj77w+Du5QkRnPeGuwOzvqIU8ZRBv8mhsFm08sKcpaFf/fDCkCCEh5VYPSxYHnlLOxYw9o2+8JT
iG7+HlZfV95AcQrSVhVK+xPiCFUgroC+WFK6k7AxgnJJlIUzk2mNxDD1fAMMhukHh3wz3wnhaJ2/
EsYezvH1AbuUFZIu8ukb3yMqKTSsbqZOND+XUblGJ1IeqS5AdW3PmswVg7t2ulj54ax2gV5woe+i
/dchUwrwoIll97aG7PxUL6oFllN4LhczrKqBgzHuC1rBwa3DhJViVEnTd0qJ/6PMv3wN5Pt2XrR7
4ln7nm29aEdE9bbhpz+RsJP+Snl/rFfdp6BAc08eY2+58vRAPE7wQHbJL2NgYbucHwY4VTUW4sOk
3Q1bRGcCuZzvEdzaZB9mX7cttgfe/TiSYgAnRrA53azaeknP+JAu7KA2/iw+6pl9xWpKux34kGZZ
PWA9riLasMNakptDPlpRERz6tx4GuwCxH4RhohuSgIYWZNdNpQQVlYXGDYFmSn7SL/LlDZxO7o66
bRl+9a3YvoKPT7yPU0klgdHUjI4bTyfRbozcbz32/Nkk2cVVWE5XtjZXkvRh37oGR4guTHF9Q8Za
yrgCTxCeL/MbLzehqpQBea/NUTsicDMrsp5bhOusoCSb4KnwxkDmdeXgTQXpmc5Y7SYB2Qk1ng5I
cnJS1kzu8StzAJf/QVykouK4//bkT0C6kwTrVVSyRQlxFzstmxYgiccyE1y/TEItHr/EXIZpib3J
T6bpbO/QYKFSXXtGJ++p3RnAgEgxyS19IdjUHkAiUhtOP8yRYVxVfb777vun0Y9qmyiv1S+Nft7V
WFqhpmdHC6OQryGZQWjZaNgUDSCgCUqp0vnndks/yd63QeXznzHg6ApYw64nqu6ZutaGbaGy2sCW
nOCTYOqSFK9CgKySkdSbgbDzdxSwI9IGIM12phY41zdzGPo7yLxHS8BVO8GZ6vJXm1tgGUThxSDu
VBM6KMie+HweAANWmEAAtYl90lzwHoSbstmauGCyGwYVo6k8BKS3RYKC6xrsyxFxKKUAoIYoDK9X
RlocvqP0wZl+niqQXjdkJm+aYAXYWX3xiFpWsWh8jSJJyMnOwPpp+2NHivlLgQd5PFdBGt5y+WyE
hFEgWK3+jyU74mIVu76GNP5yj8lIg7UbXPD4MqvHYzQ97kNMDuJoJVfwzjOJ426slRs6uTYKPcvu
5r+/2nrltZdYopo0ZJWzjQCm8GFFKSjv7dUgP+MJjJQj1p92U7hlspsTcN0nQaJoKvNe1PIbtmD0
ZQLHP6gnPNxbKYN1CKhL0pz5rgZCQUtL9QNdlmuVtmBzTSNFR7TPJgAv5CX5f+Ll8etoK+ii4Jju
c4ZLUdEsacNCf4ZHDF8J48FQHY99AZYyt9UQeNviaNuJUK38mqwJbot7NJk8T6sAwxulQCsTlCQ/
G9IuFvXtg1ry72a3uar3LiaLed3E7fgQnPaNyteMn6KSEds3bcTqaZDWtM/g4hZLUHNjmq6INi0a
jiPAPuQpwNJTgP6r46lDU3u3vVOODo7WVzV2kY/iK59CF5qF9GT6RM6ODytU+afFctnS/n8iYrz8
zFMbV30o23bTn1y6GCmbcNCHynvl4ApDhLWbuqDMd0c46ICNZb7Vkgfyg0Oys4u/axll/v3KHv8z
BRm57Bgms3l/ugrKlwpmQznXefTL0e4tuoGU/olIsP/1KArfOfworW0NlSnM+czUp0WDwDeX6uR+
SfmeIlyGClsG8xjM89ybGkxBztgmdx8syDz4bOONvmAGK1HAm8Z2LYEbJldmQKzoCnr7Mpa3u2Ju
jIz/6pDc8dp3quTEJZG9lXye3dAbqyMf3575kuWYYw6FVEf9HiyXZy8v68hMJYT/98cUTe+1WOfR
vroCwg/b34yud58bwxIVxLMIj7NBKIpkbKwR7Dj6j6adw/PwIIaCf+Yqtin2DXf7WrXN5gUiv6zW
EGzKUynHWneNqhJTPSg7rEFE2N+ohwsYrCwtRLOg8cmMEpRbUGkpQATlHKgdpZKMzQlLYR01IrFh
EnSidC7IyvNIHath1/ipG+iF0XskvG/J6BOpAj7gf23OuIqXmJNyYcb1Sw1x8+B4VtdciVIFa5T2
WBl+EeFLbmBDM2ZXeeYEJpz19nv3nJbKVXzsOz0MmdGZHkoc++kZiqiuj7KKXs//OEIxNmnn85ny
oFOzffxLK1ZsdzvtwwaSOTfHrVMDxXvH7azHP5f06D9ghMuhbWrJGuCsRy3Cb2/PIx5xmlKNYloI
JLyI5lMaUIhkz2+m1mCG6w8beo50me4XzdZ++O3zSq3/ZWRUuhER8/wX4HC+vEKrSc9ozWUzCVIA
Tqik9CKB9LYSdZBWGyI+Bc/e7tx9tb5YlUDfFoaNuSJTtIisW8d+E/cWKyUwG7/TsrpyEbt+wdLT
NC6vpd7FkAMnpH/UXf8Kz+hf0W4BekPZpwTlme1Pvv7eYjGHaKyV3LbDmSUyoPIZUC84tM56bST3
AF90vWKcjqaWmwQJ3vot1/aXkFxlJ0IMdEJr/IgJchccn3dCZWfWcV9zSkcB8xpCSHFyeSZwaeW6
r5Yedtmm4a0qiJmeeGdorMw8xjEMadaVezUM2FqwqC+dUa5Izbb6prH9odHhznPcpzLp3oMNBY0g
PQo31bAt9/+1S9kVqTfKCwn5X6VQQIfJjQI6lerOEztCyXNiG0/0QLytBgQApvuyOkmNHuu1YAmO
KblgyP18+SMzjYZUtGltOf7Q25zJO5gGNYEU6BCzVnrLnhUJAjhnqxRyK9VDUG4idBvf6Nk/lrfT
9XM/4uD6/XlSU5PZ39NPk/7j1vuLgUk9j1gKvP87dqJH5iWqmsdSWdyMmP0ehvZe+eSjCEWGojuW
pFuX2v9j+STpdZXJhsgjY8pmHrTtTpywOKX7Eyt5wpzkczPWOdUCo39/sEgc/TxPyxC7zGZiwJfp
6dT3DfqvDqCZuZMDK/PH/728vyx+q5cOevisPjqBaoayOzBmOKUWz8kBIgJi2OWGceyhgr5HJgxm
GiCI+1TPWx4sm7avjVujUaAfmxwcol6SSNuZAl8RmA/qIOOT1x5mo0nXjqZU9wckGqGtMsYWlgGg
aLX/wBRecZczEA1OeGZTzX8Z1bLSg6msvjM6ETVxayeN+Sob/0GGKyToIMLkt9vGGLWNT9sx5f0l
ipMa4DSL7anJ3EdGF54a6UWkorDj5pOIgEJY+FCASgmdfK4Ev/+nO4jUo/unFoDZ61Xyzo41rai1
YEwsyC8vZNAl+7YeEmYuLAdfUs5MUNuZ9DjMsQSK7XtQWJFwVlPsJkozatJbxJTV5rcI0R1HgoED
9Quo5UvU6BzGRZxBAQ4OpfyZcjigGc3FswKaadGOCJ0MiOGbUj7Jv6G6t3/A+dZZcjbP/M11uRmv
jPXZzLWXi5OGprqu/ZQw/lQnUxWIUlffeIHRdMGrGR1HX8D6IPi5nNxz6lhgS91HFigvu4s6esUs
Xonm+OZxe+Oke5GTw1u595ta4o7tVnftWUWhvXNMQvaxYFVQwcuxqvayD5/rBQ4/7jzj01IavpQL
wacIsu241dSQ4Fc2Rb1EKaefTOfimQzLWv3lKfrVXUAND62Eg42RgHoVk1fhNoM8/4+hSuU8GK2V
uO1qMAxvhOLdSGorYZH84JtD6VGVleCeMiWHidIegW8FJCiuYo6+7iqsq0nYVnDwfDd7u8DRc/zT
ASLUBxevYzOWQQQ42UqnIdAEkXhdKCAHOswEohVXVg7JvhGKHLgIO8j34x2WxyJxPM78u5d1n4AJ
/AMAtNEnv7SsJ2ytTeCwpFEhZjIKo/7IjuNRxBq1sNOG0Wk1vzuVUP61WF+sz6F8o82yse8wg2K8
scG72euYig5pY+qJBwL+yb+Rv3xaK8c1RUevSy0F640tq3tOmaNOug49tGfaifvedzzndaQNjNHt
dVap8z3Ro6J21jHnHxzs1B+xM3qR4FtlcQ1narTYztGvqP3Y4Sga//D0kS+lfYQcAXxl7sewZVeX
Jvmp5U30XZ0r+SUjq9VEtFs3a7idQfku6VeuIxFSsujLuhHRE0ohlXtXsw7+erXL+ugd0IHlHhPM
gCcv4z4GBeoxcnrpPL6/KmhquBG5053Pdrk1zuoQYZFAW7hIEu82TZMDuxDKe6FKpjJ5q6gm/VTS
lyDHdoCNUnwJiNuhd58qaPZ4RHNsX20gdRHaeoqvo7UGmyFeTllqZvNxIgA6e/WLgRN64VyVS2dU
nfVQhaULWt6FyLU6cyU68CGi+zN/isbAEOyWlRwb1MYwdKfsII31hmWFfKB+xW++Bv4Et5DQ0Vin
l9Ow8BD1xYCDBausUW5jUjby+uiIwPv6YflEyyMrn9ThQNGHeWOBVY6/vBeDrIyQKCFBFaDFiN1x
ESEP0EVFnQuuC3U+3XVkdK1bALmjY3rX7d/HMNy65MCJMKLVSId3txh/17lDXKcxPp49W+35IQYn
Ptkgj1q28DKlARhMDRnbAnBEAgHBaztsWNoS6r2SyHhwkbj3IBFE5AEnvGeu+YHggJSXLXL2AXR4
4wutBhyAL3wpwBxx6IczjSnjB7fs98NHhF5isH1bA+JR2AXHsP7Xmivi8PVjC3Jsj6Q8qYtUgz5r
LqwKh1+t2fo8GrXaWxXmzfVR5jkQ7YEMMM9gDvTl40hQ18vNg6JE/2l4zQxI5ZdtgG0y6zvoA99Y
RtvkKJQ+2akyRRTZtS8c069Kd9NgdtLkV1UVnDNDHS8Ohj14JRAQoO8iKNQjTbWrLXTcLN0FKaV8
fwCNJhA8eIvrxNBDPyKuZ5DtkHjph/ywlepS4/+km9MjcbHpVIoEPmtTwfBtbT1sf4YLczoO6DC1
UBBQ+1TheImaNg5m+Nyr0wGwGHcVhA7ZiLJNXTz7O3fprLWF+5u9FZW1QIUISBvn/BjDFf1XYxxN
Omgcp8bghtP91dxbF0Ou2HeJKB53GLmEixn1ijHDgQS+TL+mOHBCvtwsnMRXJYKoQQPwFeGJyZKG
nPtw9ZwIr/51v1TA0x8i+D3hlq+Vw81seVMo5beOctSHyyxZmTOSflWRskS0plAkhKv2pUwacE3E
MVE1TEYHq5CJ4mYzItZy9jeO/HJMMdM21gIUaIgBpQ4PwIDs+47yZBux31zk9U365g3SDZES+7aD
eB2bmvlnFxRhFFyAckdNxNUinOpwgPAzQfnJ4u8iMTApyj+I76s52Qw3UXriFDyLU8LUhIqyC0l/
580WCtsGrDL5R780AwBN4i3jPJLkjc05R5D9djOdm3cSyuukhTEJUOEI1GdJYhl9CsNdv9z4MNEP
YD09xXfEdkJQv96pqpyY01aqK2l8KsInbEsG2SEVcfXVX/6E84r/71BE9CwqHckOCj1eT7pI+fM4
6drohBOKK1Ge/2TyBtDL5XXaLcydiTM+5zWWFAk++RLbI5izdiDq1ViQ/AEoi9sv2qZ1eBAV1dsC
hAIjgEnGTq8zF4ieNGIjnIQA0lZIfUJ2Nf7cHbp4Q4JWvCwyZ+Z0taFl5yr4Tu6Df6UW9fOnp4Bb
QhmlmYuIEUrgOADU9ztppmAe+T/jlFLABybsMDl7YyxswmyxnCViG2Don5IyI+5fhCctDglcfPtN
btvkNRgRO3+e2vJGAVEwnsTKQlwGf5KtZEwS4VuoS6EWhVUbJ1tgITJzkOp21mSfbkRtZvsbllD4
u/I/IJ1ruKMDvuMzO/EHvd0GrG9fPVetQmql1MpErmhJPvxQQmodvma+jM3Fhd7tMwBA1nFPWehd
D2miC2Ct62X0aQpCh8kQkQCLg/Wn/BQfFDPdJKp1C5/sxDJyrZe61zVjFiR8tJRRiMJYlZ40QHa6
oGThT407k89H0CCbKtqDHkTfo5Ox93nJgeh36L58fgkgWaixtoBfvZ4BM5H+amUC/bf0+EUIqcHZ
aN3o/GjwOWCJbMIl5shIzLy674yR43B1VtDKSl5ARZMs/1bMAmmKvFh2ufRaPG/mr8ve88dirm4r
NJ7podhgGO9eLGRis3D4yTlA6Odm/0mqDg3YPD+XpxqbgzGd2NdrDly8/d5H/OBdxSnve5hyc+U9
EnQxb8S8+Kw+DnPAjEtKp+uxF2rtKlADAJCvS/NJ3bq2tcW6RDkzyPfnMGL4O0s93dLzEmm/+4Pv
I4cineE9+Br/y46g91kh0wGOa5uWNjE6Iyql4hKGcT6n9kAzSaA34wohODMDT9G9U3YGI0l/G9L7
Go5f65uyyo2i8Xjpqj/k+acBm51T8M6b39x6btOKwQ3Pt4/lTMysWr+WVS+2jxnJdKHvg7/bQMK2
3oSXMjN4ed2OTtcnRmazuGu852e18iEjXIrCH5+sQ4Cj0e2/aUKw7V7RiPHSvWRKoCKYTKOD4cmZ
Wd2nlkU1NYO/BH9QviNQ7Pfbsi5nyTvBWFjpL1tJUmSaJwUbr4rjrleXif99OLkVr5vUHhdpaUue
uegJpKJuc/Rwu02X9DoKP5nnpVa76b8OoR9NAQayMwqbz3RUBLAFvRMZKiWaXbLJIqXWsNimjcGX
tVNo1GMKRhUPhIG65Fyd8qQN9JsUaTct4YXEsrRB4e3X5sXHNPOveZgF52QktsFdGsQS0cSNhZ6o
9FnyxlgH1jJ5uYKg+zXFo+Hmwb8j7UdIp3CR3PA+jAWUjEj2KmOx4OnybkyxSv0YaL+DTu7D7xk4
ikBmiXZ02mqm5TCjpsfsq4Dqwl+tB3nyBTUMbaOivCSUtK6pVpeuIaw4ONSN/G4onRO826j9pm3z
sV8TPiYz9U8/8xYqcY1M0zZzS3JwpCQAvadsPAyGXJtL1aHNZO3e0dANsn1GqtbnchAyfE4y5+Uc
qCE9uL7fL+gxhMCWVZtcqinqgFmXj+JaIIHsLaDqjw5IksZxecKBm73nJx9EYX8tkqQn01g4gMSH
lbTdLSNf8O+XhBEKzOl9au3UtiycA6EqXkWwMeuX1+fFKnP6xFUQdzkCMcN2tKut3+xd4ohVGU1e
3d3Y9cxne8NLfWTqrhGhBiran0pcUYtS383BCpp5FuFZIgwX1FNdoZrKpRulU+89FNkpcrB723hR
AdbLuv9ZfjzKuEBoTNeT8aX770qGXGc3RNz0Uskc+0pfETm78I/P0MXFq5crXbzhevYH3cT61oXE
afRST2qyCWn5fbUAarE6W2PXdLmwczePzl9JBta/ivLyD1PVeHhMTf94uAlVovGHQgaWYe1UywnN
ds8XUGt9qGWnYiG3yN/RAjhDzpuWPBx59QeYE6Gv8NiFtbgGC179KA20jXYamQGlqQXJ/5PVOd+5
Z0dLS7Y/oiIi/PFYft8CAhHAPVM7pP18RgaIOIfo589BAkxctY3vSiV6hPNvRegQojQflkVz3aBm
S9Mv9HkJb1MzsV/uki5M8unvs+Q4ipqrKFd1xS87ufWL+X4i6fibqDeIPV2Jy+ZVuZbDmQAHKn9e
gbsULX0jojEPO7yHZ8avxQyQMUO2ijca+GFc/Q1oc7sW4vhEbf9ljjdgh6cmHN8k+3gPu7OZ9A4m
TPQfyypiwFDSr9UyC1o+V1/nPjlk5EU10HZJvcAcrfizUBsIbITR/oavhnzJLUJCfQvQp3wu6eK8
tlFcIWxLzVo1kdqKOa20K4hs0GCvjG4ZCn7oFvwCMQF3i2hdwsVkRObhemwhLayY5sIyhPXRZG+t
UPHO/t0pNOGdkswx8kh9nGgOyv2Vh0FObby2QyMR4/1KGVr3g9TrbeOqlY/MQIJFqV+jAusWuLsg
0/3uL+TPj8I1veapx2if9w3k13OeReUhsiiAcvBOgmsdcbToYSjOSg/+fEdZhKc6DEPst7XfUH1P
YfC0z/kgavmd98xCM310xtfet/rLMY4OrITRuKJox17vkpvP69hcETIMAiiPVLBvtMj8GcdpUpcl
+X9X79nNyQw1uz3zmgycm/xAnRpYZ2rTD+51qKSl/2iEzggbpqZ8kyM95G51bR2tqBqOmN8ogbw7
0STNXwuY0NaMOlg0WLbNlHs2+BeTND+Kfc95FOyCMGcr/2sVLYLZrfh9r0f/Eckrghrf7OISACBJ
BRUg6Q2YcgFqUu762e4AN2XzQBolfwj2iYk4Eo+NP3jEiWgEEOHMmGF6TM8RfvoCoNFq6PBFxpQ/
GO7kmKAzZKblZDkm8Z5q2N3ezUJXjM8z1bInsKKvsE8pd5nLfTD3FPG70qzIPWaWlhLFB4e95Y/t
YaYZiLj0/3UP8wNmrbRpYDPjz/iA8QtH5EUDa8Avti9vIpCWY/Vf5C6iYsqMPdSq0WByrG9IRxiG
Vi3QzRQBHy2AD2KN47i1o6pmUCt9jWYzvLxnNZ5L8LMKvamUPXvZV2wpNNFUvYj8rPpOhgz5/5F+
CcKY4OoRoB7Xvp3AvKpDqxOHtMCsIBU+ruiEIX0QdGEgLfF8Yin3nifRLKXY0pFLrpH5UpB5SYVW
66+YLQG8OQRp+47EMAR9ao+bxEjmuB4V4P81Tk1Nr2mbSrqkMTt9jdDEV5plVGSwAv2uBBTexNS4
qtf65rWtSNJpwHqqZbwIaNmL41Siwt3DiOVGnFkLJjFCN5meWZVUfHWwYb8DIzvBQodB+JgqFPdb
2+EoCRfN7TFGVxSXFoSmVziZYoawknwTs+H3MNshjWd6hQ2yz6uJuvAoo1frXGGzxZGIb0XB36tr
RUM0zoF8i0BE6dh1f1casVxJtL+Qv2bWGO3LlvGXWO5VUWRdlePMQHy8ArudyJAnAxnmMtkb0ntX
BZqTxGVC3htHAllRBGl2G6CeXu8Wg8jjGup5E15sHMQHYlQIorcW7gXYKfcPNbtunQQeZGZ0dVsf
x3zJumKz1U+xUiDRFrGFXa4YlEW5gVAP/T3uB513puxx8irgkmRqgjJY3suLstj/3d1osUbsu7Nr
AX1ob5+lZxDNxhIZq/plenaTeLkZh/8kFLCoSIJEmY5syfcZA/MQLejGb8hCHNZNbmWleQRwKjIj
8C+AMPjfdb2vBYFSvVE/CvNaWPijFvd935r9GX2cWb7wBQGB5M60ICIe7pvjMEx5rA0y6x53lzNI
klTrb5nfZywuwbAEFto3pHDHIYTtzKyaRZoURE/0SBwXPTv2ZzVIcLWNJy5Eng6eBNQ2stiZChv+
bGGRZ2onYYf0xbuySo3+R5Fxow70xDZngOV/6R3EP03RCCXV9CI9Wo0zTwGAsMyc9EIM+HJC0AZn
Rs0kcp827GaNsluYixc3WiW1E+fKDm/wdd4r2kQ5+N1wmcJ6N/OoImYWt4KW8DoVJIgsqPX9I8sy
Y/MBcyIrecDC2g24ak+VWwNRexQtXtSaBUNKawpFhc1cUJ3npJbUP1xBrXRiSHruze8nQ29Bd9MT
auCAvpSn7DFho1qXBVLQwH0FJr+/D24w9fLBIIiaPvxdxrn/kTmWS9fr4ZKrWNceOwyRHMWf7sdi
/aJK6x5hjN4IwPiGliSSzAlPzqGrpiR0OnhkE3XF3qLTIDeJAy69yqRUra0EkjLz+lJ5uSzarugB
h4FAdlV4zbU1k2EnlAZDpB3UKGmV7eZFbSRX09biQVrUVNs/OagYiYk3aPPRbbIroEyu04qinMSb
8tud3EVWXOufoi1GWMBdxZCX0kF/L+z5PODuPwukKKFDmpj0lh8dFJJyzitVeyV8Gf6W16EW/71g
3eBwL1B0tug60zIZ7UbLJ6XChtWFFbkjv+3CZzOmgTl99mzjZe9qRoHjWcOZlyg0Kt2eKJQ0JpIU
LGZsvFVRHyJHPo4sQU0JeucX+CJ/CPSHIO1b/i9NF4PFCr/rBxJ3SflufDbLrUgbjF7644L1UKEg
2oBGjRHOZs42Q8NUz7zhPtzQhksGDVYUMgVFka0+u8Kx6X2XDBYRZ2n+8VO6sC28NiQsJa5bMOIs
r0B3/S8nNIU4cA4aryC520ivQHdR1LlqZoimC66/KBPDE+TINljdC0UHleEcHgOzAhOy5/cxUOrB
TF14PMZ2lxBVj2WRdomYo2GE352IDieIh+VfiTUzSWoMm+/pnjpH7T50t7XfhyCf4jeqBMKjOJvB
iRaKDsQswWqx7X0T5WCTj8/Su5d8Bq8G3mZC/kJQUP4t2uNQfgHoItyUiTRcblskCXz+eqP7R9z9
hv23Zmx2VHygwQSGxs4Xtw1wNKutAlrrLR6lnJz6KtXqAChxcLkoqixU5MfdYOTPZL3bOZvPymM4
3EBHkFz50ytjaMt+TihOVrm3kI0tlcCzvVlg0qWFpwfGIDZYlOtpf75J530xM//u93zIyRQlolD/
nowT5HdTIvFsDXbxmlpBPdfiabohw/ceV5sHjN5u2mc7n+VsSViIxLtZACBQsLapjZJONMFDulVM
RaT9EaizbyYxc+nHv/RM65+2DdH9Q9yr2zX6W4OyYIxaTncC8oa/IumtrOMPEc62zNFbLzklBIGQ
T37aF4P6m6+HASHIt3HLUITfG4FFHkqBxQX2kWByv+D0LtnT3a2kSaloD6NjzpSGozIdiosmte8o
qRBHHadQBc/maKY8ah4WgtoF0lwriBr6qW7/FblCa070bNWrsBqvo9H/ijojaFIAZoBzBjjHtzcl
DGx0eLonb82MFtJVei2n1rssZTvUHbA6bnt/rke4wzJ1YxGOq+t9N+axUrwblHiDElMFfdQeXTke
gy8QNM7mw6IYStn/+FsQGFVlICbJ/VNgjBZUR5LAzDwi5lMQDheCihTxmZ9DGldgJexRalh8Mk7h
5mrTIEHRIVfh28381Vpn3GO1K+fPa1Z/J7qSdMOsLLSePva7vlSdbM6U6v2RX72yadiz9O3sbBzr
Nd5LmmSYQdOBTL7MKFk2F/+Ht+kcVQ+t+ZaLt3VTR1mLPXvIpAtaWX9ygtcvo6En6DiWobOROGDg
GNb6D7c7a2z4zrBnbVz7cCNX4iaU6nJMae3kpMEbp90YNIfirL6AOJYuP+P6dSUzqzYZgmZYsnF8
sfaWzK0MhwcnY4P0tsc5gLvs7KaPxTB8x9AcgaXygeaFPSn1EO3bTv+P8/NJ26UQ5rxNoGD9ZP3C
k9T/kBIEu5FSc0tfcoPIkr3CRmkdZgjB7ssEvd51gH4pP44+bf/hDN7wIArr/OVn5qbIXQEh73Q3
/lIHiBsE900UTmv6/phJg0nU9stcLb3fA8NjsV3gkXlzuZ9bPKFPJSFEwZ7DpmTyLoCJylgX8XLQ
Mpa6S4ufhOjpW4IUbvlyfesv2TLoJhzGxX5BpsOjZUQLvtYWPjz/n7FUD+k1btzln4j9y6mkm+/S
FfQ2zQKALUWc9bBvv5FxZ+mblh+Sf8jEoPCwOg+Nv2yndpi3q545FyC1FJ3t3DSe9dG2FLSm/xrQ
nWE7EDS9bjqQzxHpdgpKLbNCq3QUlPu2kH76fUY00na3YRF8diAUqVnNlLWluSWP7bbXYldQkD9N
aJf3yHrdboLGOBo/vvJH+8+iyVSSQw+8cI8S3WcrmulWGHTaH6mgZ+Be8sjeZRlAreLZ4gEKHq71
TA5biGLm52xThgbuNrecGCPFt3paB4GkFiMigyiPuJnivNASgPSQXm+4vqv7/q0R3TDkAvRQoAs2
Fi3VTzAL3ZtViNVP/p3jCDD5rvlZbYgOZ3rr0h/colZYAaTEtsd+BFDsmEMbaO1Cnce4eaBHdOZq
ylfhsQ0WkwbBR5fi4zEyltuSgPMXs76E4qHCMgTSHi+LtW+aHfaSGqu7mkpXZCfH7LYl5zHLiWP2
pFD+L2PFtbmc9Np5IVcv81O6y97QIeoL44la0mK23BaXMXhRvAnHvb/x75O2L9KxUTue/uIiLmRZ
kcZoDiTBb/1m4xlqU4NNNnC+uW+T37JNfG3MqwRTKdnMxYBgravzNWft9xDB+NT251cpN0b7SUK8
nomZsIt1QRGZyoaXQ33Hd4jK3wMdC6vzYHKHj+NUiA6xkGiFuGAdf/pzoCehvvEzKkzFTcHke65Z
X+PKsspAVL1B8WVEPsQl80S6PpEK8ysZJcfEAqOJ7l5CYMYNsX3whmnMxsloig4Yb8sPAY3odzoH
kQ6dlE/SsALDgQAOCKk9a8Hinh151JoolIi2vsyTZ1B0+FgZWyODN9eQOWTp0Bak0Z8ddf2VYDf9
7Luiq6tusTxbv3tZxnDBc6KGtS41/hqbiV3n62D9lPc+LGfX5WPtND/ucZITBKh5jU75yXiFpw46
M6bIFpyDfsK/8CyQmIbQ6kpLsYbsWSwWj3N0RrHnsUrGINioRS472Cv+oXDHIvpetiyv0NWGshy6
38gBnWO5FGRJhr4LPx4JSqN7D5CmonqNk9G4ZcbyKutSKHr3pl004FlRpPZGewghwWQLtrPEWGpm
VRhWnElj6lVOEWt08cWAJwjQiey+VTQ4KdI1jLS6xiRmV5k/P5shjEuAoOX5Nz0c+G7MKPwxnFHl
a+btS4Z3TlS+TWp7tF4Ybtl8baPSWHRMM/lcXt4Iptpyrl0kfUpwGj26XAgqsPu++Bh+qasw+AjQ
oCarTYR+zRAUvKKjWYi+YkujyR62eg+E3DsZb+fQYWjJ79/dndRDHlB6hSh0rPd/wozz80EdP3q4
EtXqLiBtBPywCrQVET9kbj/lw43Gm4bnch+sX3m5PdQ8ji/umZDy37DzGOKPBJOoqXTYsuAyMLcM
Yb2uLnN/zlY9/Nbat/UR+nyp+l2NdOFi1YygdAH8FPffRYvxYJFiIKL6LYTPtaPb/5wKIt3AisCd
PsA48q8HO16X9J/MuQUIRnfkOdmCdmiwugwzDPMzSpIDWwh5xglMEccMZI8xr/irG8VTx8iATlbc
D/LrnidRTdrprDSsQGlRC53T5FvA/+cX3NBe+WJNryILRNc9wDeA9Z32TYWXX56ejI4fqxZfmD5V
pOyOg4yU0vAL6EpkyaVJJLcpZMxMISnRk8CoHzTKjy3XbGzIv8H+Nl1LN615SStBzwxUxcvlctiN
najkOTStbpUN+qsgVl0wIUSpixhs1AKtSPsYK7HwOryBzsklgRQNBDN7xqSbDHXoMlsEq/xmNv8y
NzSVNtfTBvrvLhO/IEbCNHMMUTxSjYrP/bgnbkvCa9jTT10VUGC4Mb1vqAHIumd62TcMqJX/dLa5
Whoni8ho/EsFqaAUW+ELRuJuZNPpsi/wca0Uv+g9+wQryRwLGPdQ43fE64O3wBW3BD4f75jNVSMs
U5r+lKvkcv1a5n2F89clKtu5Zl1Mk5lB8Bm6ozvei9BZZ70NoFGZ/0cwvZk6c0nZta2arA6oeYto
94N0o9FEcduljyovB6U314oZj7jEWnQ/tx/pnIZ9TwWotYcBrTwUCJ/jVB1CKc6hSL6lzZYsCMHU
/SFkVMmesmV6AUJYkepQfdHGS71CoaXmPXic9YM3/HbqR68x8hhieyVlW+HsNdXrdESUeECPcnt3
Bnn2dJUTgrmcnhoZLfTv1kjy6EC+4JLslZdJCyU2rjblgnFBT/awsRfMuqybJKS8e3Uffpz06e69
8/jWVsNDqNgbMX6wdgb+KI9e6AHoK09R45J9SywCVK7o89UxBDWO2uCYyzvjinCVICDB50giBTpn
OSmtTbLz3DJkLQbCCXmRgZMG+mW1ETZPYQ4w5BEWNlXzc6Wj8h+srVq3rwzQ2Z4RrvTG5orptZXs
Eao+mmSzDk0H3nQgQhHHCldBISIMwaeAzvXKFw/fTo8PNXjh8pn8E0T1794mtzPsIwY8zrbV5ppV
2ILEEpTTAlb7jltP6RaNMLNhZhO4Y0YZvgOK+8SvesrwWimuiPyR4xW7h2J9ioOo0T0ifmnMX5cJ
F7ccdismMzJgct+BzGxBm1Qg8CjoFMCbIDKySt430kRPqqPQyvG04TNd4yMYAg/omxLrUxM+Lg8T
f89TvEL3Vf7zhQsbtsBxVuN6+5uZEas0fZ7XR+UJ+fScqxYIt2V14Oy/2cUR2ENem8L6a93zFerk
0d2crLLUR024oyyyIOFqp9Tf27/XrpSbLSrxXsEorfHn1TJZE9zbutdP40kgF2ealk1ftKDtErQd
Fok0RTInsPlX9glsGdhimQN170+P9fd4JdpKC6SPBrvo0jhoG4zvcKSK+IfTEAg434+VdnKttNC2
8KxP9bstlxs4bu6huKHSd+T+8TWYMfKBzrCoBjdnloVgHXKQsWYEmDk20PBGrwmltTX/d2BRU7Sb
KXiGlWEqWAu+pad+utVmJJWG4MnXoHa09lVhLGQ/hmUZJMG5IvKF6XPRffunof5VgvnDWP3H1C5/
jiLsb7b3iWW3xIDjy9AW6E9ecoX/SCfxItoah7ItqFanHgDeK6N5OXF8lEi55Il36odeMER2TdaX
bzob4yw9ToUaxcMQAtP9uOwQ/DfWOCTUDSjD4PbIoubNhai9aHN+HKHZKQmHbRAYZQXgSrZgSZln
KDS7Tld1rvMm7eD3FhVoIc7jYFCl3TCBJh/JeQ6JedgoIPTdiHFm0H8gqI8lFwe4ZzOx375MsQ/k
ZsoB9kC6+KUN3a+VZnYh5sv/juBcWdpYD4+gTHKwOw3jdv/ywNWj+SE5UVxBtQhZqXms+I5Cg4qA
JD2xUYKGCmDZq2hGsB/Zjc/UJtra6HILdNkQNU8yXS6sj21FSVJI3g2I6XmFaSr033PMhlJOXZrx
iri3safPi2k/kvu+H2DH2tw6IIR13VndfihprQx3bBEGn/vXKogngs0Pc5CLbEJ6ebc1Lma6KEtv
0fC+2liv6SF1ZbzSlijLKomt57DZ3FlbAEhKjMW+WBQiJnfxqHVVroOyZLECZrFpXwWYBofgiUsD
i2eoyeCg66Ft1pfYoMyLFAsVoZKIMIM/IfnYraNI2mSp+5uqc1CoUz1EYpchAHUbfMt0q5OHEvv6
HE+G0GDFaEMvBa9OK6orx/Dxxen4L8HcnvEc3NLeHFUlXbSm/I5iMIY3l0eKPea01DOa6eRf2Zkx
y4V2VoSysQGOclJteRt4UTwDntsiAzf9puOv1U2QPwV/lewo1LwUzWXXG/ozseEK529FABbpOog0
vnjfkOrfIQI9IRZU1gwCb5EtBPZgO6w5O6V/BMAFfo+HmdPSHjYSVifOjUAxeVZhYS/BdHr/T9TG
qql28vbExCXDpOobUAtiexglPIzmrKWs5tN7Ym5DPg2/tp72otnE36hbfDeHYxJDe79HwVVqEpHb
Je28geerZxwcQk85Ox1hWNWGai46TCLMdSxv8P7umz7ER8gR/cTxxBinu1QuqbVMCZg/xe04HFAp
suuVi98Jk0rHsstB8J8BzbrpnwAtvd/54NhOC0HSJSnTn/vZ8okx/0BVVzLstD9NcjIDETMbjC13
DtIhNjrChwWJeRWgF3UkXmVSzrwusiH/yM3dulGYuElC/HSG+TPnqyocjI/DV5nBVSQa6U81E7GK
4ydyqZLXuksscDNo55p7PRSxv1j3o0DSdLjWwoovh/70lH4jxHI2Y71I5fGSZeLvlFnz+KDEkrrU
Lg7ccJ5fp6/MTDN4AoYv0QJQ2tgLDnVq4D/xIXfzgANY13pyYOlBuUqdJLgT7nNnhVswYsXIv/LP
dWOxHPdgoHK/iWOjq5kfFKO/+1JBhD42OM7lgUewmTt3wMRp3YaslBWfJRlZfIBWsfFHlaF5fQxt
wMApUZWjOad5GuIdEBnCJXFZbBE+FfaMIQjZHF/paG7AHf+hzgdhQ3Rfrd5KK2H3vDNDtHViVv7r
8audOC7OEh7EU8G+hkBcKzyaiJXzLIu1T0BczpfLWkAN2VZ9hU0Ey6CLqvULJ/QATOcWOmPWXshg
2+MYyD6zFlBH0dqe4AS9N94BRpLNNDDxi5fnc4itVj1doMkvxogrtOFKCNKojW1M+g2YjorvcIKB
vUpBKLDAM3QuCDgyD/Y1WAbw1HdU1OWm7PS2xRjsxegDIEfApisaUFV+FFakdHVeqn7FXCzQvQAI
l/FzVgbX7ws/1rEEcM24suUL5gbqPa4ageU48/uEAGxg2lOG3jv+lGpIsJlqXSUkJrtLrGQyv2w9
MQt8TUrUokOVEjRRUk54ZcsQ6O+gMdfOzOiMSMGtGQPj0ACClscv+tTBaVXMwMuZp5RWv6l940+6
qPM/qUXZblItpmexNAi4lDDIeeiKCDRF/91VBIMySkSo9RxfdYbfu0e+Z4ZHe4V6W042NCm2c2Uc
7QDjsvYYf0inZQ4GVbI5TTs4I/DPMQedxiLbl9Y4/g24D7ad1f7y56GMvQcW5hMO5uTqbuwNIz3o
yZi6HDPqwWQ0VSltehO7Ajyyb8Dt1aVwcvWwtThgYvbrbfCAaQN0gnlcVM4wUsHjXTAoiBcqR/el
IBsAUJNfBVij2jis82tmDErvL6Hw5EuoHseNGztLF2nDAKG3WMX4bCsWZb3BglDpFwZsNx6cMc0B
uWSP7JRQ4fZTqv5VtdsDlbqUPVCemZQ5O6v940U6sAnP5qy+5IVncFidymsvoxdrw3RM88vFhmNw
D/gjqGQ18EBmpblFIuac0aIj62XJIROtccRAsKLXGoawNMDPt2/e5HQvg/Ng6fpKYPLlMrPlKIBr
AVE357AOS/a6gMnsuxRET1/IXuT2G7ev6inJilrQEM5ye79nTSi+VqiyWS6FOohM+e/9onWyQkr8
zfcbW+bMLOCmjmC2CmxKQrSL/4YwhLTAQD+JCA0C2uLuAC+vUsVC5yLtmel+PVbPhzhvN22qJ1iU
mgR3LdKx0VMJM53pbuBZwZcg7pqp3TtjRiTLohWSznVQFnuASVSv/Lt8/fMuqy9kD3o0wzlkS0u1
BsSVxfCr17RtkWB3D5h6x7NP2GsrdRVs9pflabLUmyKmYLLL2oO014lNnttQU6z4stIwlIUeKR8h
/DShbcxlmp4wkx2rC5c53+0Wbp4X+liWVYThIW5Np9SanCWGVT09Wl5Ii+u0pe+W2TI9Wml6+4BH
UHHNP8NMzJy424UEXVpYDri1zqYhPFySKWvicXId4LMVhrD19YBO+4wyoFmOvJFP+MlNLPL+vN0c
70xtChwSzYmFEj77pnSrx+r4zUv0JkAVx/OcQMvSxbBxTEzFVbqYlrmT8hYQi33BNDTCePlCAGrV
opsBKjZZlfVqweTIZDvQ3LnJCzWJJlm4hHeSisYCBkTH0A2QHiivUlHQIOFcndsIvpaukhkGpkko
sOkByg/OJ3/TNlyRnRO0K/CPLBEKc4sxf3GnjlVYuTxjbmNpEKN2+lTh0HhfZTbCJKCT+UsocMP3
+PP6xoWQabz08VVGSSdN2A5NeiTtuhOTESO8AY7ZBF+WGYhSUxjDWnkz6g8mAun5Qqfe5qXJDqHW
xn5bCi+620qC6VDhRgeLVK+UdpZtPc1enqnm9UByH9gLSu67Q94YKMFGKA234cfp1oYpHVh4Su6T
Z/Kjk/RTYu43YKNT6I7bYxw1EWxvxwNC8s9QPnbo1Qw44cO5TS2gnsVMsGkbNjWwq6Tm69SwpIc7
X6AkX4OJnjtnEAvzbfL6OF2mf9AkFh8/M3v15W5SdCKEEzB/3DPyS9y6LAe5thgghcbxiCQFpc/l
FULSkbMiouqR20GoEZV5Wgg7is494nJcwCljZ1MZootutRIRiOug/L5V7Ob9V8s9hBbGmuAQXcR2
olDkrTU4COxinOjE5A7CeDnXaPGEIrTjNOciBLOByeURi6F+r2VrPxOOs2NWOSNEObtUvIUxxmc2
W3mcNTSSMhVRjDhT0s0vtwGmG547B8xt37279j9UKsDkDzYr//Xd36iGLTSmYdBydumOhQCE4SIH
+wBJ8Xbab8GH012gAAOPfVjlbJ/fwEtprsT7spFY9VHA+sPpuWTpBOj4c/VGU3c9q0/RFjHW1dWp
bnl1qcqnZWeq7hVPHaJoIA0vNs4Y9y3G7TeylgVIPw0kcKtSMtY5isWj3t7hLd3ZW3YvAgGrP66O
i1Bg179OP9uhqSWGhzBqK+Hw2LUWGdXBSg/tlXjv16ZX1kSscalf7SIAmko73FVtc5LcSSR3Umby
jClaMJrDgZLUTFMfnKcQX8aj0Ck+x8X67IyTX50AOKVhC2ovCuCKbFEj4moCBEa4/MBdEDHx8cl0
MxQP4FZJSCes6v1kY/5ukwjXI0lVdZ5Eequa/ThKFfMBFiVKK5HsvmKhQMx+lkNIuuze8hcrQ5f+
sbfqcU7iQBRwpqWaBRzpBjsj9+wY+AkH277S5k99lVszjxoebus7ZP8WzyndJfimdsn3lXq5XpZO
TyRquEtKdGIn8zfM7mibNKLKwLJEQcvPqz2TP3RIiEB04B/XmORjNxOcZ8dHZwS0o/nqSH+z+e41
SyS9IWj9tyqelgiwM4SLk13LTc/GK4R0VpBUAro5QQnO4FAIOZWLIfpdn2N1VVVk9S/BXoA/MkPn
rUCB9W1YZa1mWdgGfyNB9pA6pmwPyvH4HyVBU58+PUvqiij1Lne7Zm2vUWpMjIO25mB7fBSUl6+h
FqKrO9OGzmVuxIhfQzS8ePLZ4Mse6Yz3nkA5su8HRXkfxyC7xTKW01d7x8En/ecGwzSVDwE7BEra
1KCFffXpidBWQDGzipE4YL64WXLJrm4PFpVh6YrEG4Q8/cjKzSO8bjgHnSh5VBMrJJ7HK1tn2iXy
dh3fbt8qRr+3obyPD2bcgKEAY8rXg7U3LC7cn2cYLryVJ8tCuw7t0WF2OF2NIDIqkPSSESWfe0qh
/4YzrUZmVffZy0oq9Z30kM+Q3nNj/hbkrmlnY2XhV8Tk+Lp8DMJ31pqljC9wmKD5gpUiWxtcJdXd
Od9GM400Ix1U1RZem3vBbJrvoY9oBPKuvvEBqsJ+AR9BxkFYzchL4zgGvdrsnFXqU1pyURoiLsvG
4HC7HlkpYYphSXoxSeqtyV4LFjwfC1Ij0AceRySMJw7jrLNGkyjn3a54wQZnfSVo3ToXAH1t9koZ
AYSeTJpGAiEAkFLDXc04K+YWn++23fdhooDAk56CuVyuflm9SD51D804WZm51L5NM3LFn71vy/4k
eUkJqBA/A1Q+ptcO96E8E3I6SS+p5AzKIvidfmVQOsb+E4f0S6vaZ9NCvwv1+hcBV1srZ2MS7ijn
bIoyBMVwS00il7VSMrKhT/SCYu6ENXs+/n4ICSDhZM1HrHBBcLU8nOi+ScyWnaccFTqF47ok5Lhi
lOVM7oaafK2NphHYczxrGPQM2HWYArvyACywwziu56VYVmtyLHVu3rebH0LiSAclwW/7mLVdRgJQ
LY5LjwhVzapzJo/D+dwrzj/g1kiIQJyNgBv57vtFqL2+6vMt5nMFQnDWdU8ZfetXpwRLjsRgPAjq
c87qsHW21mmKk2okBBpsFxOu1yuCNa0kNXidBZl7FOIjdpNcZVZb7AHOPJdayxItirXQ/A2Einr7
cpGHtme/rI20ES8J0krrp8cK/3GB4rEOSCZ61ZmIyRrnRJMKDXzGtjSxjriQLfrdahbi9eykAVLb
wLFNa++6IebWdYlfnD/b7eEu1E1tKycjwmyy9aL95LgywWrWRP9aVNkX+mVIq+kJcIfzc14yLcrO
9FirRcq1FM0cqazLjxPx27dRpr9JWX00X4I2bQmpbvRmqkEmwnUba0TbEQdG7hduQYiUar9OtHpE
7s51dfi8utyASYe31Eh9NkB3wIjiPEKLgS6r9aryUJNhlRX/VezFeUJzKQZql8AqRSN5IQc6rcnQ
aQbMBvzX6VLoGyYtnTO6l56xjy3xVUea6kx7RPyNEr3sIEeT54JRlBQM0K3JqyGEzJB5nbPsT1KH
xXKPObNpdIMTbIe1ULFUTRZEurdl+d+r+gfKvon0Qohu6xkr0RhQ1rCYdWDwvSomfx5cF9aMd7GH
uiOZCUrteKLQLgWhz/w8XqscbTjkPBiCJILu/4h3CtZ5tCt8xBVPLadagNDYbB374W1PvsUqh4/Y
27Y4LQpwsLhtAQAKsZMs7T9Zc10MxRyFAYdSkFMkjtV/sQ96kH+yyqNsIhC2giP16SJUzNRpypQ4
pO3u03t5yeljKk3aAWcE4zLTTz5q1pRdltf68fPDFt9Q3jA/NESKKF1dKA1zJDLR/Tq6yeaQX7kD
KSzFUGA59emj+YPIBUOi5aa14pMnE0aEChrR1n9/gTcAIhnR3R9/HE5Qb/od/I3kZH36Dsx41AuB
TBjcWo3x62/sfQVLu5srkWAr1P5Akunh4ZB/NaplcnVYLZDheG4CQ/PP53vPzcIo2e29KAPYemqt
VbOXfoeUAFzWeZX2FahCzqBhosnmRG/uQyTtfBNgDdxiIu1JKoTbVLUbSZGEJzBwxL0XpFywq7xL
QnZqFOncGq4PQbwVjhefRwSQHF4tIjGJvb6ekNHNrYxUtRMFVucFHrtwyPtvKX7ZmrZItEjY43t3
shIUhxM8uCFFmlQW91J4H7AlwCLLVzWn0+icxK82fpN+VQPtOc3REJOJ/xhr4uxHp1y3sqN12FCu
XAoSnaSJ8k4ilwjp83SFzNQC5lIjFkRSWyDuG/AheNvH+nKajyQCpEWgp8gwo6D2NZNpcWMXWQS3
cVU9MJDfpwWJcIux2ylZJxSigaxyu6maX57iEENw39VzsPNmQAxgK03/iO5UwfYDlyU/C7i8IBxJ
IVmCq8qdnBiSbpi1koCRk0dMRbgVjLnOiL7fVsn8ktzdxz2r6jg5yp0OiguHwvL3+Dw9V8AFpfb0
bm8j5//ijhuKAHACb7MlyETFTnmedQpAk80CrYnl2Hj2huWJOHz91TtNatcJikeHt2QjkOL9FIvX
HedqhR6P8CbrrsHI5PmZtzvy8WbM4sBsGnpdyxquVPjGP5NznWpBzEoMF6moL4nnIva02E3saRTS
SghtG10spTzYQjd8crZP0uS5KkjFlfAkay8t0C62ln08t3+ig3ZdDVKn5IfF1tzveLbNoFkUgQxf
jp7qqbn8NqtUMW9lAItnYSVNbrvA/aTj953NJshrsV6byjJdkEpoHvVEYNKnZ9iRF+1TlLB2GcIR
bTYoyGrAdq+f9Ec01zv/qwA9xLld154VJlPYpfQXtl/Wk5JCx+lImJ+DBv2v083WcSVzOcri8XyO
xztz5FY+iJDMGWx8v9pZhNh1zsXBS5xoppIJCv+LDMinwTO3sU6dLn2b822qVS6KZoxRRQRj+rWI
F4Q9HNeylgN4fY7PoqO6hIaqqAFbLIbCdSX2lG5Gow+v5EF2FNkkkBAkOJ6PL6xJg4/AZBNGGNJZ
4DGaMBl59OTKj2yiFYlA3wK3C+/DzEwAbBAJOu6pKdo8L4HH0TISIfw+GuVlkoYSFUUM1rTgRBJP
xzGZMOB79QAW63vqnU3tcBpTLdCTWs70LpH6SRDHqBZrA2ycn+ZTiDo2YC6uUKAS/P/8QWjLtCof
ePfsOOdh7LiD+f5Uv0MKvXwpiTW5DQVJbOLj7sDfbIklxJ9gCaOk5ucyPIYbh5D/M1cOKK097pct
xJPCVp5vzCqdoKRCn8X+jh4dzqBR/OCwdXJBqk84cghiHGuVXg7ovCQ6Pg/4EWy5sIe3xeKAsQx7
Og4N7+w9wv+PFcbQRUAE4KrWMdgqLfuqpxaXA7mO55RneqtpNkz/E8sLbCXH9dV7YuSUo/pr0AA8
/GkUUh996css6oBDyyKF5RnDb51KSiMCrIHYOHUdjJWJ3/MBUDY1oxyQ/OSthMYQJXNEhYK70vEK
6yODAyyfSK3aK3EYtMjs6qg05bZZr/IezZ5hklMJWtK9+TYPC1H0WllHwW+jm/R+/hvKJC9zAAl9
BRkPBGQzhG+bWrXMwfMacFKsj4EvA6PtxBlvYqHBpcTpyqc1mWrTYkgtQyWLZWfjmLkrNHp2SJPb
EporVp4RkjRvnAMkfCnaBTcoZztiIOvo21I/mj+unT8fJ8qG4rBDDCbJeobDTYymiWH2hP7nue/d
vUA9hHAuVYiO5VsefNFJcKZhR8bnHyo501jIkE/oA0NbsvSXprBCsh8SXtVSvHdOkBGwTK92zsDl
hnbL/FqnPjbEL7XNeshdKSyK7H2NjOx7sdqO69PyJHc2/XNyxXEiX/NJzaS0PlpakxecI5zDbIwz
Matk2QbAk2Pnd9csTQtSTTOD0744SSb7SLgzsnBBQ5oVfHjkQwqbN3Tgj2gBVv2cEEeXil5aXPEx
zJtMr0T8Nexc81FG3h/dpTgIUu50XB2u1Jgl8WbAZqNmxeKq+Orssf3TUzJsNU3bRh6EpeRgo050
kYbw64KfNDkMo3WCPxhZ/qRQDiwtPzUNfpNyE9HMXxnU89izqEowLrXmi7Vskr9+f02S/80Vgy0i
MfWVnSFZVAaA74jPvy5sQZoOBIcum1UXhUgTqBrupG4gpLzUXsg79zpkQg8s3azC2WORTMoRqZEl
IOpmsL1sxvDUXXAX3S8ReV7hGXENfE7Qpy8G/xViKLmbt574K7IXN4qjZ/6mMtjCVw5jz52YbFGb
kMtTB98fcJ6n6UQmQSO/fDb61z4jz/3vdplUTth0pDc1atA/bce8fY7iq0Qf34IP4XBecfpW46Hk
vnaBPSavTXbzx20yuTLzWH5VWq4bm7kWl6gZKiHgFEt84Dxb4ZvrNQ0V15qT3CQJ+VsuHGWY1D7t
ypuHXYbLxeVMhRUeAI2oOrM5vKnTnE+RO8yKnX25OXXpntJTBc2eHdt6A9+p5mpHP/l6Ysb8b+M0
7GMzwxp04usGdaSoUkX0T/TFk2KGb85I4HMu/kVKeUqUSSrkWlUGWeRx3enG4Y+n5ForXkOXGyy0
/DhmOqlb56fuvDn0GWtJG22YLD18YfukkfIEJF7FjeN39SRLXOqSBlVsX2PB8k5otWE7OnIVuE+0
byh+IL0GKQbVoqsLLbfr1HwWMyzoC+Y6tz/POj02Ik43xxGZnljhz9BkI9IBKvQU5RxQ4PjZsnvI
mhGPzeoNzJ3YXlu2VXZPIMIGSMhnMnabiUNmlsNZ4NNKltz7dULECMgOlU0X/GT6vy2mHXTOEn48
EUT+vDpCAhOOyPzJnt7/4+9vyeGwP4/eXU2f3Z9pTTt70FLFzoi8JGf/us9WaPIp3JbeWSCZGpwK
6RdHp/ca68SawFtJ/uS7Y+Ftx6VeKLhfQavPHNTRkb4vou1pqtIuNiKpMPDNY1PaDS5YPt3FcxgG
Q1oS8TmKMgsqJsficlB105bDKQRYimYzJxJ8LDB8+lc2C6eKN9jXagfuUDAcJk8TBTz8IvPpPjKi
OggAzPsSSa4p+MM8D7Xxo1PPdFpS1jmRxIPXCYncUOITJK64Ljw/PVsfuwt6wwvjqJfGlCrdUIeO
UHgfBiVxMmlrSF7TqbYAjf/kmd0d/lhj6f7ndGxkrn41QOZwOYPAhLAT4UzpnHVcPOMfSuBhToMX
yuZ7HjBKVEh1R5G4RoARtpaCud5YXEdzQxzsMevHPVFBkx8Mwk7kqG7VWK3KxTzDwlmnXvm2v5AT
UkfcKg5hcSaCsUoi1Iys78fBb213C3UrUhT4WjQ5knQRQu2PoqlYTamAuLcpPCfa8q+xUeacBGKl
ILYL+o3K4i1jKieTCqS564UEw1VGb2n1Uea8QPZPloE5BIqS1BYzebM5Ah8CZC2d7hd+5l9AWY9l
vYZLu37V0TeNfCHEr58BXzFkKvmXUF2ZO7Tto8bdSszh0/TTIe59bs3qFz5AgknRHsdMbhUaHgMT
tsrvNow97iZvLhphOlD7x6UeYR+vo+dfMRMxJS6ItBBOeCoFIqZ6iDVJY4m+kOCUpAb2G8xUCUg8
UFxI4Lc0lhCwCI7/GeKDJ9IA78KjhvvJPQEdILjtr75yHj3ttdBT+wxydteWL62vCZTjUWL0RTGQ
zDg4p4YVbvk8CHcW5yPkjSFZres5EAU60BRvGZr7B2J9LXYcoP/1wFBH8/+A8if7jy3S95m94HaW
yR7ieCR+WHMvFigwBRc5t/GJ8U/LesVsxjUwi++l8owNU9Vkoi95OtRRXbKmtdErUTdQOkBxg/P3
BcxhhFsd0lEExdFlmNblEBFWKQWLv6SpVxizfrKw6erzSrRwwq5x+GNLOgBJnERwDbelpnfWzw/v
3F/9J/ZxNo/GmMu6bvmNZZzxw4cYZnZ6IRyb9vOlJkgDi9C1oeqXXY7gEfi+k3tbvKCSpWu+vKa1
6LKk/v/ld4Th34KxI7pEmFJj/nJv30PWDcd+cUZ6oMlqh3/M7DxgdlKaZjOwWtnLi6W8nuF/MyF3
NF475lWACNRrqSjdlbmYD5Agb/BsoHdGCsvwEdtjpi7+CGyC3GypF1s/Lrrx0ae9a/uAipXa6d1i
sK7JSTQdZk8pwHXVvS0dG/LHM5ZdtYDHj+VFu87vlNsXsiyFO5LMD7f7RtghAnmhkiBTmbFIGKfd
eo9A6mIqtgYrbyFZa5fHC4DWsgsk6KB4aLteoH33o7L37kZy3uHqsMLKWHmQm/v+DLoMAsXMlfE3
bN4q8b2S2eaKU09dWu2SgVUPHBOBNdcDWaC1rv3CwT1lVf1aabWdiw3njqjTQ7pkqZjBhyLd6fzC
f7d/H7ED3KuHYAvO4e4/XkxJnoEzQtwPZ9Q9j3trWOnQ5ykiwiO89YibMg7th2xYXwhzPueMlzfw
omafeyy/lINwUUJWEYf8waICGvlna9wGpNl71Pq9c63K2KHcxb43E6W7Rc51L8pUcVeP/IYr2Aa8
/0um+jgECxbYKwsbfJHpoUoTldLGs6LXnEe13VwSJAFjgDqVS3iwPsacLIJQR+koSuC8UwcuJ5OF
PU/a7X8RpZ4SN9jUHDH1F1ZRyjRCiZbZRgsXrRdqt1q3KdkWPWK6KRtGqJyzDQxt/LEZEesFs4Ee
mA32iXBjGd+QPOWoMFOEav+SIv7UOPKKb5QKLxH+qP6vwLhSHiCSfT0DnWI6wvCx92lxpmFuwDlC
XmP1gr2d2U89bdgGg8R1miId8syP5dILFZGShGWVIbq/cnyh8zMhIk9anTAPXKfwvRzrW76tgrGB
os3bufV5XCfCfCueu8trYoK5GB3h3PpKKUOyGb/+27l89ALuvRUeAUOEuQ7Uhyrij9/YRcMwREHt
GVA/7kmPbh9saLxgDyLBPHUB4qmagVGv8eNLbv1GCGkohkMgBbXJHhR8VY7PsYpp8KwSiz+jk8GJ
USmKY4EPn2nPpJBZjQg6pi43zKw7YBuCQRP6N7cumWPQcVcOSHv0Gh/PMhkKpzWGWN7b0DXvq6+d
Ugu/a6eQisU8xoFB0Y/f0TR9r3GQNwOdJSZG2DLRd+g2kTc7DXNASEI724A9cSrklY5t59oNwPt/
h3OELPgmswEhAG+Ir19PKlnAn1f+AOE8P2CL5uPvLYzuduQ7otP/GXpz8A1y5ra3+V4Q00BvqKmJ
mudmoVsUGUuHI5b9xW5WseHkRn1PEkiInfxxQvbDHOMebAzIexrcy2yAxdWm4RZ9Gxypwia2W0ty
E4nRFa1mF7sXWf5fy7hFCiQuCg0vgTcYGiIUWeZS55kUtGMQQ3lY/bJIZWIiGePWO/BEC5QTfpjv
B+OaJAMQm0rnPtYf98grEdaOfWw/8HjRow1vF1C9TSFpLgg8JDhRUK6aiSa7H7eR1kQVHNJhJRSE
j7ukzaXyg4bkf0dIoo0jrK2g9ON6mQs6SbUDZ2tT1/WfvlQp6jGTg3n/ZyUHFcJnSsof3+lTWGYl
C8frEYqE/N08pr3kNBldBtdn3+EgBwDnHpOOZqSUexkekY7u3rEW/T73oLkls886b9m31aJwBhc7
HkJS8sYgMw+eIXPX+z/o2Uo8QcbTJN+9EnKzwt7dgUx37bwNw0n60NIDRG5OHozKVdhzbCUKIXdw
GG75WV9n9+EgJ/FX1aouEPSmYu/AwZFl7JASmG9eaODzWYKxvBOCUnWm9Fqz806c8LHyBhlPYg5i
yqb4syOU51pW93kU/jpSeaBxMogXGxEcKvdH6DtiRpMvUMjD5ExigArGSOH8bm6VsjT0mA4Qh7pf
Mjud2KbVEifn/7DJKeVEb4D1g+yT7C6diOlI4CE4PdbOSov44Z6P4O+YDKdnRcuU7cgFPuPz6nGg
9kOz5hEQCKawWwwy9so2x/pUga005JDWBGfMVmYDpM7G2lm4tYILwuA9BseW8nKW084W5KYcQCrJ
hngdSYqb8/E9f3O0bTACCVXKkceCuKV7f+529Zz/9X+gl3jKM5FkaslAW1j+jmgP7F5aifbY/isL
OqUXqfBTlI0eAAS09tlE8JQ372FYVowTb7gXGniC8Obu/TnZFzSc5hpxesLKIUAS30n5ZATLiGGP
huVQfDLyWYVrkxeIWT4utM45MDprMZTofkPO65rDaf9qfBO4GggpQ1igTING6g2ESYLzfP8NaI6k
t4c/9ulbYBKtlQ/iEYCwixvuMIvj8gNIrGThY/8oLfMtMK9a6Wz3b3S6SPeekecBF6XjcNR009VQ
S1Ro9dMCbFRp44Rnc0uSoKJZrbumQaGjjFEXNJOAQ0UhIi2Ihdte/v+spVPa01yXLKbwXhBd1buA
6syfNMjvR23Wg8G/32XVYPU9tCpiHVqhtwEAHydsPRgXv2xh+Y7/000pEIGhI0AeGLDLt9v756N8
Ra48QzzHzLzFqm/dB13aGyWeUBmrV+YJHzRswYsqpPZ2N9OtOifRVd66VaYEieRf1/IE4n/RTZas
qye1GLUDaAlZDeomYSrmc3lYDocxcdOv1TylebffpNrdkWjfjVoO+1SWWzN4sq6Dle6Hjk6Dq40n
kYRtgLIKrfZrAhd1hLqr3UeL5GFERr5ivwB3Oybqa4uyMYmpOvDnsKBZ/vgaWQBmkN/O56380VxY
HYpAdMEH2jQmB/D4ce+YqBut4R/Zwo5pDK5FRJNoJZazByFVEqQPHdHfXfTguid4bh+2t2cRpKvd
JMQEPZBFC/+OMuCKmGx5CUmMgIaTIAeE9qdlCOHf/Q/kPMoBLFgVXrv4H1HHxpi6+dKB95Sntlcb
R7nEgc7Xch+p83rXRDK4BPbctFrxAB/9p3gWvhbUQT00P2ZdTtXBRPQ2FvHKkVf1O9wVVb6D9pov
5GlDtnYoaVwWDp7hl+4VrnOGiOaZ1o3DDBey0vshkLVwxkOPvg+HF52W1Zvq4tg5z/OL5lNKWTRR
ZFCgOoyRY4rK/FJFB22vwwxRyPfl1CBQs46x+1bdITzyC2V6FzsjMAsqw/xixj2lCKRU9dmhqE5+
mfynT1lEylkynampKCfEVu/OSjSC2D6je/GR89ayW2fPrAJ41DS1VYU2VMmVoQyXTxNi2TnbSc0m
O8OeL3dxKquEyaPmM1sj/mjQ2ZC1iE1C2WoG4yidFK+CrhcFLXw3YGf0K3lvzaj/gu9FlzdHKruM
AzOROsOi1uLFTJDmsLR+1QjYLaA9IE/3pzvyppnYpoOT6YW2h+qDjdFsm7dCqQ+bfQpG941ZcGQP
lk9I/HHm4phKolmUIv/jU5f6vl3gj0KudpPJXBWrEUjTw9wBqpG4k8yca6v/btLyjqeG0glYmcQl
dceTfSzNXRieSEgLiEuDZQm5zatSCOuhh9b6HqAGz8MqDSvQxMbN9btTq7G1yhF2I+13BIaJwN7F
Mcic6JG8uaDOHecYg/gJkHwP3OM9CPGXlbPb2sxaGZm+glr9noqEEhxEvJw7NqePKWFGrL9rYISs
2pwwhUeO/4uSnke8hQggIUEaX3+G+e6Md2+AEf49ljnYX9GWwmmAy2muwd5tYUQOft1TiOa2F//a
tjLHBPPN0tQ0P3bymTYE4LLzgWQhmyyeRn4ZoQZVTwvGmi14clqA56kTcerDDvNFTT/PkReyc//O
RBmjfOc4sc1thxnY+XsxlenSrv/cZl+7asiFP/B+PaLvskbPj6ZC4qa1Bn7YEnpXMI1RbS0DFL0C
bLeiJ+xq5seLM0LhWgTIkjox1oIKGPzDgr3fdLvqvVV34JYfuHtilsAexoR2IHhwhFdZEmtyd1sL
yNvRCTGtYFxBVTrZEJTLbXcZrccIDVwW/6vXZJsLNFAux9OnCICRcQmHQtsiwFHoYcgW5aDH3kYE
Mw6/c2nG6r+jSgBKdNbCycxQxAUVU9oyBsE4B14MFLVtngujfHhd8VubyrLFGNKuuf+t6LQqwLRh
jtUU17V6HVT3/cOUDVrvop6eU3Sc+tR/nn6UtlhPH7MMi5BbhpIhnE6CYWWyy6K2jOhS9Qb+9nBO
PvVQYRkL98/FlY3P8wppctKfIpbohysvD8ZbvWaiO4RVsmm2tn2uYL+3tHXhG5CJUTe3VeLt0//t
fTSJRnLoo1/49UEDSyqFAHc0GRwMVuNZFoQ7kaqx5qRoxEQTg4vymuvHQq2rWucMg2Juan0O6G3O
rT72T5Y2KBu13Xn0zeOoD0FXpNWhNGZBI67wE4ZCvJDgNmw1co0YnjOmxkvZYqlr/t3oMerNbaqJ
B7bTMElTZeH9Hc+nJa5gAcWVvmRiOSAzk9LB5uhUVvXX1BnkynAn5vyaNxpbEVAPBjyJafx+UsIc
Nrd7vhVwZ9adjQJMomGyEs4SsXdWYvFe3MsyY9vmv/ZN5CXFxlgR4Gr0NYKalzG9ikp80adNLy8f
f/1GlNrhBFYnwGa8T65Nzk/WA2+nrTIUUlSTCIaLleR6Jw+cEQM1A7Y8AvfR7pwj4IKESLOq8Kgp
ywLFtvVZpg+CytZWQn3smCAa8Wfyhi+HyT/KKtgzOuhlswFjQi2iiBNwl9sx+aHXCWT4fZsfBWON
BOjEdwY9EdERJcThw7wP5x+wC9p24XgxQVp1dDgv+jN0tFHOVGbmBfzpxR8NBb7EV8yRZEnDq6NC
3PCbxKGSEs5ygfF6ECw0zXIgE/sI0fdyRUHW8+c/bzwXg57suo6Yj5gtzTjlEEmGkticPEsnERkR
7+i+WWW8EVAoGaxwr7Xd0l8xoeV1DU2Dt9ihgCw0uWq0Si/n189vVylb7VDQFXvOZovSVL2peEja
rbHJbBGIS1JTBaG6X5IzyOPtXxD3PU22oHxrcZ2eV6GYuJZM7E/1woPlT+alPqVgCaUuq8Kg+J0y
/gvOMh65WUbKU8ABwfIO8cl7MAi+LyLiOjiJMSpW47NSubeHUS2zyjhoEABbPNeTuj3vdT44d6sr
YBz3Md34JLqaFmzRK6EHOf6j94hTC73TloNzn1chUMHgmBtgkydVOtETDCjbPHPxmbHiAFyiBU1v
NGAW8i/OalfwvAcK83M0TzEx00RWJ9MD6X+18ETMWSOG6RwaMpeiIqxRpgFsUchPFCucZRky/Iqe
CFIwvOmN+4/7gnkth+eQ3B+MNgPYaRunnDjFJt3PFLof2vSAcAD1JERGtp3KZvsGK2pj7J0ZB3hA
C8HIyWzIbtlW9EkhQ712vvwBusOIWgAcbC87qO/FvT3xGKLiXjbwOiBJfVKbbEeVcaQHnXw4z6On
ZDFdYBZ6Uy+mLM3e3sz7aIEYA9S+h2f7R2JJHpYOX+/3iTM4P9ZJ8DiKXvhT6wQpxkOJxq0vj826
tUZ7wdOcoCwWueHDLx52pghfiGrlb048WK1IyWb3E0UqRwAAbovs8f39h4dZg9t4VY57zevgZI2l
H58qggH/RdWpSj3zTPJW4OWSUoyGPCA6qHZJsxIFhqUCgufTJ4KFVW/HCetW+lxohG1JmdhiQc0I
oHa7v4FH3Q1bOcdg34PGz9sPDqzzjZ8sN1s+SyT0OMyuybwaV/8eMoRUp6zjRiJKrtQ4PPuRmkrO
MqaIf2nQHwqR156NQndED59y06V0nIqIKbKmg3PRTmr9fIKCPgD8Uv+iIZOu6EzE7UTR96rJ9t/R
Rz8IwwvXav9wEW3mpCKwKScvVQmEmuCM9OuPeX7ei5MBL6k+Vymxp4x7PijfEV5hIoUH0J2PaVAl
11cgtLvjG5xqNQI7Z0jUdlTadjNobKBx8/2COKtpnAipQBzQiLYz8eZ9/f/X6nGbaYWYIPYuXFZq
OojcrS1GfKS5b0uSUZHWDIgL1ZV6H93IghKyVTAhbrTgrdkkBvTcTlrAC3mDdR8ITPl7nH9wTuwC
hIfUls51zjK9PJxAqJLqBfSU4rABhqd+xhH3C8pmEiN+/m35BPjzHth9FI/fRzShhyzL6kMJ0bAM
4s2jcko/dwD25JMW4RpeOLj5MGieUO2NCYsQvelcG/3umRTZlQqFFDzob4BUIC5Bu136LQb/8hD+
Wu9d3JaRzpJRGG4coY4nFX6DZwhej/wj+hUAJmMKo7k6G1QuyfBK672TzSaTA4/m8n3z8qwKOmx/
/G0cQv5Hwia6z26ODGCCuqp+wn0o0AhvdQtQkyQflMb4MsMChKrXGIMTFMgRMn/LHIczhjbNGXGh
1qhYVYsCNxyq4LcOl0MAWa9ixINo/ocufAZUBeZTagBHqNfGXtWDArLmIA82152+xuk+mBn+bKfy
cYq1N6gUEoPnAXOiOUnlJrNCNq6qw6Z3ZAR8fRQMPjDU2DoE7Qd59XXGXFYWIPsBM4kv9w12Rhnm
3kXMyyy/BCD3Ppfwc2TNcTB7tXJZfvwNTbgk4xvcbYshpfxeXRLoQ0btmFhx7zqJgk7LUXfkFoI4
D/N3Xq+wb+78lRVihkyR2rjmmLAEisQftyweUBPFNyInM+/J6j6tPhfYy9E1eTwGJGGcYAfO+Cnk
sW6lGZ607xpwBBn/9UC29B8rPa4SUUSf4vKkTZFPPljZzWVCWMFdetbMnJ6QwUGYsoWiPyv5e5Tp
V5/cl08ZusXgIuyu70DAVCHTGNsiHk+iMN6YA9cwMVv9hbriD7v9eAisKb/9LqEh5V9s87jIwZEk
uBl0ajYJbHMwv6rf1ng5DAHubVTTcWGIP0mBHhtRhVLRs4xsxPbKW8U7cHmXaVOBR/K44+84M01K
USvM2jyaTyeQJ0pSFCqgkUaplBTjnoIi6ymlGGgX0to0Joa5h5qxZUsPIznNNyw4u/TOs89YeWdG
lKrxTMEvRkX0/ANme+wWyzJMuvcskht5vwDvCdZkWRYc/LLA1qQbCO+wDW/dUUdIgDFIPtbovi2b
fdd5HKGcFhGPA0z5RN5O/lMZGxRxMfPkpG0h2qoZVv+lhV4CDfnh1PBO0nCW47hrfWqeHAssUfXQ
a9gHq6pLdMkeTvstjgDspj5XIO6DmWQLpjpXQeRkQBkDEk61rg//br7ox33W7Iyn9jS0f+iJSoNt
wrBzu1SRAlM66lGuWHebL6s9wwPiQj5PJmREWU+NHDckLcJ83byKe0ZPhWjMlqvejCREfRVcGUqY
LhmlWRZhONo1ry08orcAnDhw0AYWsL46rkcYUOddY030WiBVZRzlfUCG1yW0oJ8c7nd18NbR0KJ/
B5699xSH4ZDTVSUj0cEN9ABUkwqimkUDAJpBHFqvjXw2tsCgJlpW6o8g7ky1EZ4HC3F5Wd+lhK72
dk92L7zVgLa/zowI5jqqx5TvytAEyLDfGZ+EbRTEFOHjhuhccQWAb+FNONIZTeX9xJU0ikKwpb1I
n2fVZ7TvgU1SEfv52hHpYmR8g5njZ9B+qlBmFcFBKqMR0f1dZSY7h4xClusBUcnt2PhhG0ymQxgu
ggIyreVHl+zaY3XbC2hoWIo/Lm25nqH4ddcPhn+7pKI7f5FiKfeSWgGzojiLKQRoKvYyEfzoMT4V
E2RCH6FaXkmxPNt2LyI66wXbsUVeqZDd8lFomnyaD0QZ4fu8MvZypO1by3IpiVa/RTVuMsU8z+pw
B/U3Htpse52hjR/Cw3x0WLUEaf2QvTt9O7lx32v8RlKjDYPO8lLzljQ0VrJTiia9wnxiXWNm/S+m
10MW/GLBVCWT9n3etWZks7v/xcsWz8diZPmP1B7fNbNbZpUUNk23xbOn2v6lfs+m1/+8NP9WQDnt
PI793cjrpDkkjzi90lro1J2Y1O0Uq18eFt+Gg2OQCf956Kll20QRYLd+mYcGCaeH9xXNH0YdHpIn
ta4lfrgMX7ECeVWdnQr1pYgE/5ZNJcyiG3qHuuGKu7licwSGJInhOiXfZ7cGD2oVW/FbgecdZOkR
Z4rcMbQAH7blupRpWeO0CKA/0rA1BBHvZzX5r2Z2kfOjElhmp8UCe6mogl7iLQj+2aqk2supH7t0
I2keH1fEn564IbXadRXchisOwyAiX91dqTV0Cu/7wDHPtFeWeF4ToI79rzNihSppv2rW3HV4t6sV
UIKAUXbpZBsp6D1Lml+QbnIod9x55uevlFSS1ln3iFmAaKDav3kSELBut2y9SqXLD5A7Kpprd9v9
L57UFV66kaUolcXVjn7w/cTgoOjAEeBw7MMm2Lgnm8J2sOC66DaX54qRFx7JiSxvcrj7ekCGgUpx
W5PKYWlfU2xrK4hQ2CVmKBFVvZ+3wHL1cwfofnEzXbnQH7IgaX1DvUTMR+Cki/OQ6LkWx4gK1lkY
Qn8n1OMD2LSC1S6q4yVXRtGGltS6ZBGOxu377ryGQPX3xL1/PnboMb7ZrCMu47OW1PeFaKCE9UEu
sG8SdTixbtyqDfcWaT9mRxvdGMtqoO4l4S23HyL8639uDqwXXYO8/UB0KXD0Cqc0H5VkVrjlx3h/
hpX4Amz2EDRnnj7+Bgq97lX2Cwj2Sf/lFb48M23bkOgQCuzCwyqlvROawn+y0qQ5Iqwp6YlSD5kB
bbalPeqhP4mrb2wSRJ4UbWNXoCRbfY1ggcTOze5du5EFCq5DrPJAGnNj/DJwrRS8dy3Dj3IqiZWZ
IvROJpi5sJp0bMnAXtXHL9VqIlBpV1vDY9ao1CocJnPjwzQt0EZeKiUwbdxUUzy5bFCJNCd4AyZR
KAiZyDD8sCJgxPtfKYXPnoUZhoXSccjIsF5YTUrzP6HDl11emOZEHI7XeHomYp0ErbERj27dpueS
+QZlwibOsYVTRwt+jqjWOQlfItc3DboWq4iQn2XvxKJkt93Le92aZKb7RXpPPrchqm47IRTSl1ib
wOACV8fJGMceQzl2zKVgpTZH9W3+rPeUDIo+qeky5MLPpdbL+hhQ9cRRubOtMmCfj829VJFOhbJH
kyvzT4UEG0+uDTU+LEGevu9ZKRgX4nEULmG6DckY6ed0Yq+w4M5wxkZVIrJhbUftGNNKL3fkV0lQ
NDQHm+YliOIQ42MHBlx8Obq7yjn6dG3KvJsjoQW7rYsyD2YTg+OfYlh/xC+EDeMG1kzKYztXQxn0
e6MF20xOGgyILmUHkU0aPLgvyy9hVMX95SmFVpJ9Jf0l4HN8bcWiyNcnVNa9d5QEmJBCAP9hTTHl
KvhY83Dz/rOPej38LovaYNyUNEWkZ3rdX41PW2BSgH6zLWQMWJoOxcWOZqxZPN1l/E/cHr7Wqjyq
pHZ9BOz0pA1RMQ4Cj9DHUNaFBB3VsijO1Gk4TJNIs1i4WYlIPZsXPskgMbrDPjCu/J0//B6mhk5C
dTlbFatgvhCv5EeWq+ZXhNAiOAaPqI6XFwsl624z7XJCqTZTa6ipDW76TB+qnZKuxbTA8xPfFElk
6Wf7z6QJ8lT9lkKp6QFcwfBgjzoFZYRyT6EUZV97hpIfL3a3WuiWhPBRAogjG2l8R9ghhkc15iSS
8b1LjzqiSLl4kbIpwJEehBHIcmsqLlMN1EkXrs5jiRE9PPPlnJTO/TFsxaAOq6dDdajgEOpZunwQ
jhONPZOTELmqu6oHicPYgfZVp6zA5FvaFO8fw9Rfjz4M6Q83J7ZKMTfdLMr+DpMKXAlwmom4KU4I
VwPB+eCMwivkyrIs1nVrba/aFfk74fwZP3aZs3Y6pn+6kfUVBmCrCxuIGShy6LJQG5BoZPHeVUT1
00eYuOw01nR2CEMxhclNrwqhwG4YBfUjuzibyZX7FyoM+Uz5b78pdt1lWu6N5CqpFLuqvMjl8FHC
u3FaQ96hdupMdebjzE3OfvM5PeNPci1P9J6BXZ87Q1MBFu1TZviRDMK2MMInbt0wu8pyhm6y6WHo
N/XNyPejIBiTqxWg2fLek8IZNtpsvSwAnYWWpg4JJ4++8OsA1AX+Xk1D5/Ua31irTt2X9DoJGNFl
2/jRvE1oJrFruExhCQTtpKwmscbSLZHxoG4SFmkQUDOXabZGzFuf7eL1GzRuXmOMUWfkBVddLatr
EOa/mmlhWYyO2AJnORsfdpHMSWJNuVzlA4GXg2piKu+HUOz/0kiTY7iwD9l8Y6xmr+RB5ZTTxYeI
c7jT+tl81td2FpZm/QuW/TOJbtpSlp70dnwPtM6DkRAC/WRxuKWWzXLoyygu3H7XU8DOtMS2l/cx
alzDWw1pLqJzqBq2UDh4x+PhBtx5DUa86WdWFnWxw/VZCKvYm4CFjmDVFDtw+xz6IEJ+gp30Jedk
T/lUY/MOha5I67WZtHHYHN3t5DFT+ScMAC1kN8rQ097QBla0aqPNxA6ah3mlF4Oe+irpmwTbdc0t
3v9/e5m4+j25s2xF86/yKawip0rT9X9nzOBu5bJ+w6v6hiF/TfxWhEs7Io4mIlgBOBgE6OKJQ4F8
JkEWaDoZavjwL+ShTh5X2hRW4oQ5xHLwk/51unGa+u1P53QrxabfnNUDmA6gchORs/XHsVQfLLz5
uiWPv6tcxDNssdIWVwPwzwSUdc6oPtW29JOMsFFyOIJyyBt/Fuxy/W/iirVz/GJLnGASPWVfxeLm
YEbMbeAIhR3jcuzIa9ERvq9SGvGd5E87VTClQFbGqBZCwbXS+mhP+5tLtpJpIcpdwEHZRdyhFj4r
kJUOeOJW7gqQUlNTWtnc844LHTc1qszImR2ZeOGWPoFKxCexQvj4++9sPt6WBMpZsyw2p8iNBzSR
2F77tUxmqAPRmScTmBQ+28C2TYpr9MaIN18uWMRxZYo/lJ7E4zJhYgM542ZAo4EeIhSzhWZ4zQJx
LQkb7AhTfFV9aMltv1fzctN/0vZpMXgDCE6pHFU2CGLyfIEogNCpsBxVus/930b7i06rnFajVldu
SfTVWjkai3OhoUPEsKd0PFJJ0RkBgVGaPRcCh7Lq9TJLMk5AXKzEEZEucl67/tWY37suhhiFeOIw
pYGzCpS1DvYja5f0eZ/DbAkqR+qY+ccIXIgzZ/HRwWzvMaNYNWS1rYYtEUkiqmtRjd+jMDq0ZCxr
chghmBD+srFSCR65lCLax7M1PzRPmfrjgx7KhUv1gRcLAth2+Sq9bKmJYnE74QEyjxEYWuCVA+tD
s+C9B3wWNa1OIUlbmJA/nG/W1q+lqKoPKsbh3r0xHTrfWlbqNyk+SVaKW55SSyMYTb3bY3Sf6Wvl
RZRHLHlm/uMWYLT8jVlMsUqpuYl1ov4Xb4efM/DoA35hRHH/GsOWbfN71kMF06TeO0jK7xKrYMIF
lLRVcxH3OLn3tZqhV9b12Fowhs0wk6AjqkQsjXVxqWDZZ+FTmCDWb8f2KJvDB4DxfeaJgbGIeFf7
WsI9xCvd4d92plHmfooaAyMI3f8XapSfSNWkjTOztL/puLJZ1O44JOMui3dLxt0XdSWcuhTYlpq1
IElJ1N6yWUenMFtqm0HbP92NkclZTNaIH/9Cv/yibY/MAko+5sYWB/ZPo1jecikeyO/flfoGpjIw
p0rOQSpGBawiFn6qHRNhxOSKM4YtTTnLb7g3q442V+0EZylJ9eo5u46iHdelnXnjETRzaum/4/3k
urAsDnDTVJ5h5taPBqLc91S/T6uyXHc2sp+8Gy39QUDIkvtOP7Lf8q6Q8PZyY8kNtl6UD/AEztOE
xlY6p1EMB1kpp847rWREOKwXCs47rb+qf5E67GK5ELdoN5iWHWc+Iet3LqwI7CQ032LfFWjLV3bJ
ftSMM263y35yPALiTQlnjwUPmBVluWOPUWKC7pk04vjasX6L5A8oPyRw/i0LU/nlpX4mntDEdKEI
lUIpCuM4LNjom+dO5c8/A93hYjzL9xkji0u/YIpByQ7tPGCDRkCYR3j+1TinUnZ6d/+2YvAnQWAY
f7B1k2KvUgmH2AIPzxwQBkoCaC156pMee4FqVHVz+XhYN7CbGLNOXbE0U7lgIcskWo8gcx3lFDpl
WxP6f0NEz2CkDZKsPKHgOk12xepcxhvIdJ9I8kRxkaTC1ktZwHRTJTCFOtfDJIm2Qsce2eVyTZGa
0XczpM7n4LVVvtOMcihRB2TMby8D3DeRVVY3T/20pTdVj4ub+3XpcrzfGySopwNCWW0DiWOH9Vy6
h/j40ntQYumw7ozA7dKo6eXMdx24MU6V6RrgFPuZH+YQKEqxcTm+Z9ucE45pm6lJqgXPbU1lbPEa
nmuu+DjF+EBCxysoY7fu7ZM0iUAfPOKGfLByQ/0Sg40a/h7KGSJrYArhy7P9crQIsqSW7bOArNge
LB5TKu7+GzNTbsI+L0dVtRKTnPbUjm7atgNeXjZV0dL5sHfS52GJIiC5EnQ2Foi/SnOs5CK5jd+j
FOv38BR/zI4U0RVNGDgCqR3fvBMlsk3x4tRYODoLDYeH3DWLTwvvVl4t10ctrxbehId5R4O4VO6x
OHtCNdOfxzFzJkJ2qJ9w3zsazmmdv+LsGYgQfd7IJbK0Ue88Urt5wm1x9bNdW6N80DJLL0acPV11
E+0+qu4UiEnRMxXV8mrdcojSqaDAVeGvLjeek8Q93AXYzBtlTnIT8jenrxxQjAXELQvEypFKeYDZ
c44+hM3xVXIyttgERIHABm/a8MA09ux30UTXX/c5yTpqr3Wub9U3VCUmNlSqOKcPUdv4nT/i3rMa
2vax4xERvu41Dh30HJGCd9S9STq2i7jBIcqQf7BAU94SIlSZ36kslb0eVdRdK5OGp/YCJXb3N/+f
hOvdSQoHqu20Gu9Nj5qnu8qatR6vy/dgtuitBeuj20w6A9FqowLMDjBZNZBas1gyHNeDWB36WRK0
skjqLjC04DBbuPpGz3NnsZdvtpMIn3VDSj7H4gO645nmuvTZVBtQQPmxPQrQZZjHuLMtsTqmzrOT
OO2unv9Z4dA6Cj2bMafCGui2dz92tugD3yOEEUEPG24Y1hcTbBuloSOmQ4f+9L5dyWTHNMc/D85r
ma+JX24cdUTlHYLh/tesvUfyTrGuKW2POtHNmugbgJHAR6+NouJtoqFLiTWridZyAm6q3aYlWDVZ
z5m1akvGUwjWb/Og+XqBxUYs8tshgV2GCzBpTNA5yprw0Qjz/yJRmCn2hUcCzjg86tyiq3MvXzCw
9MazdSyX329RcDiqvno0KSQo5vGsCjYoeZNB8PG+VI8IrsYBxDQhHSHKQfSZoHRB+T1P60TlsNRo
da5Oka3PKVsgpQUt97xEjvaH8xeOK+jr4VjaZoMitMwC6r8Vu7TfrunkaCyUf1GbMuQibGmF6Zih
nwKvahRPf5hYneMWUORgisZkVoVukbtDz8DrHVKzdn5UGMfRr4+H4/rvM7f47dM6y+aEvrF8Ro5u
PgXyL0p8JoCUt5ttp57KaEtyDZcJQLKB+2Ouwm3P6v2GO07zBEUy+Cx4xLn1P91tdcncRLhlSyKA
GdGycCKGy2yQh8V5LbL/5G5rjE+qhcVPERilXiY5LBVxti0rPx0VxMBn0uzEiHxf0/cUcXJn4vfR
k6KCSYHk2glu71hJyO4ZBxn5UboV9jibvPuDa7cNa4HSNYtfoNDk8Kd4J31tYOm/80Wa1FbzB3cC
BVVA4fZFeCP9I/id6iH/YGDOmThXTloontQikmW9wNYoEBCEUUnyzESVKfI8wnYK12VKV5nwz3hi
Ux10ESOVv3JIIiGPwL0jVxKk0JHEy0frwMcMoT5rLQO+RXrcg30c1cVTtm3D8ZURCg2nZ6HUcDlm
TphmbhfR8337OUUR5DdhNsjTItIyWfgRKhlWVULU1mNHqN1XSy8YuUM7ib5BfETYSYbd+GK69Aqk
qpQZI+prmT97PYeu3o3SrL3KegAKF+ZHn4rpXex2ey2PHztuE6KKy1vVngd9Zewtee/WBiyW5GEZ
GKNYeFbqjMAEDZsxdBhUiPQoPF+SNFZQ104meGHYK40gbImlp3Ae42FVPJk++JWlHve8s0WiOWa9
BK4zCv9KcjSIO0r1r8/JCs5dqPmpFdvdLYbP47YvnZpe0aONy3vwQpPP9lRG+s+t88GB4YZItAWF
G08IJbDJ+Jj4dfWBwu56LX6V9BgSr1RL3Sf4I2DzLilcpn9zFeKSUNj4Pi4Du59hFxXq8M8wn5HM
Y0dfkS6MeZVp+/5Z9aLYpBJepxyLEnaIG4Q3KBtFscxDfvAh8aPynfe1jMphExTWm/X2r3Un/K2i
e8NgtnARvaemA2HyuXwjsEvFcGcsAcr7li6Z0b0TTgL32OU0r+5O73V2Ls+0Hjxi3FtJ2F1Hala/
urqFgXnS2jpjvBstx3GW8Li6E1L1inEjlJ+YtRXQPh6H3G6UeTRnNK/CNl9j7W5L3g9jmOnIq3pO
VIIjMzKvlSr75VSOCHXLlaZRDVb4YX+8uyepoZOrHVWII318PTRdozt4brgMhsQ0c329lHK8zU2w
YG/lapHosleM6PxWoaClXcUvit7jjAPwgPOThoj8HBXYeXJ8f0ApHpHwskeiHKzBq077wwa3GIRi
I6p+OA7fCC1obyfGE5uG6IMnj/lWLWj93kNZWWCs4sLPrH8yPMSXGDT45snY00rl4GEUlNswnl0A
gjRkxkCyWt7Oy7b4lw6Vq6L3TjJhnNEyonwRnYqHuN1+39Zmk3y4L9UggYZt88MA/7ECLv2leGnU
RX1ldBOzj0gaO+YX3AzwCZwJ99rcXxROf+LdpgwjZe37cTv1x0ptJAGu5BI0mvvhpJ0DLeonufyC
3kvc3CVMQl/524nSEhxCF5JFCyqCry5Vk+7CG9z2hGL5oH3xf0Y1yURZ1G6DEQiyobpvNW8huNBm
quZviI0nC6LZxdxt0yzyQJ0wV+MVtltFQ6INZ3jvOinQrJWrpw2yEXgUobpkyQX+lWMnAPBVasbS
jOoN9KrJ2PmWU59EXdE0oykGwxtFF+n0UGFZW8bWqKnMnYn22J0+Lw6FzF1RpIPISdbCIDWaeOTj
cHsGvIl1gt/f/4aV2BXZpI6AbubjqZtSfFarQU+lzQOyNQRl+jFjuLa3lankYCAxhdJnO7ZAOqOB
Twy0EFfmsKMu3nG9ZtGSoucv3KBYwvyHK/LRZFjUxJJsbx+TzkIy8y2+TeqMgepXlNYr+Z9WWv0H
mSMxQH0obuqL6AOFC7apKj14/mryVzAYQzp4l/bZypOMSjjWQgPapTZkEa1061vrDHnGO4JWIBet
q5z1TNI1wNoy0uQk93dABfHrAzYi+5v286xb9sdSZ9Xj/FlGRFZcxdhJME9Qi1xsF5dEfUOy4DkS
qraF2jAEVyPD94DFlbJTpsSGAdeX0WbWJYKXAvnAXrEF52TN/VKXLbFp5FrYqp1IC0os4WK125AB
Wgs/AHcz6rhuo1BAC279oFtVMHsEyg4E0xeJLEopMCNm9t56vJ68b8HfsZMCcqMEmXh4BX4WzLuQ
LEJA+z197+pOVvIvJmvs/0frs+k8loLbuwWkiVrI+webRmPuTqVFJzoti51SJ5dgWyS+XOj1d4z+
6AapP7G6wPOy4ETVjgquyY9ZHXVKIVtIelLfA7DHWOo8i42vU75VkhqLWywBNkrDjxBmi0WQsXf4
zOBWdiaEzN8BoS4UKcqIowlvUDOmyOyCJAWtNCbNCRwYVaLp6T7kPI4nfNLNj+42YiZgMkGJwBqT
pbCbUTRpQB2cynnK4GPpv4Q1VeCRaMgehNM6ZbE6MEF9nM2zQ7eC8AupJGzJKAnS876bkI5U41XA
AUA+C2wb0OYF/DZNsYFyBetDUv0JlmjANcwBbJ+uRecI1RUbxBWUt7Y+cLti+aDRbzfogV/Gw8OG
yNgFbDbKIHfaC/MYnrI/W52jnbFKBjr1X2eWXZc5fka3OVXKtwBRDX494oqzqADoj3QA7Ypeek9j
RteSyTPn/GiiI4WZPja9AkddYavzNpE2Gyv1C/+FaYbOR8RTbi05DO/5/gnI+xigSBdDxJ25irBG
iAjonxvCpXXG11RrRT55MbQEJpnVlAsCw0z++kQ7XxgYlpp+PbhKNQ7Jgqh0yhgREZ9ojoP2SoZK
OnWuTHGs/o+cCb+DZLGpHHAaRcMWW11DChODWAazoEVuhu0Ek223Dqcv5iIP7hMfnj5JcgIgVebm
J1zMT7yI2PL0cRzZxO3pPfzN5yRcorWqJ1UcYVYZlVAV8pyvXHlhtRFxqTtpBM3S2iXoPOayaJXJ
UWme9w40XxE1iX9FcmBEiT/KlugtZgC8WkYIk/TyXsTC1R9PiLjtu3tbVESsnTpGkTKg57sL5YX+
kAEaypSzjXZAsT1A3nra8tLtZjCRI7VRxSS+6sxEJS60o6nX/eUrkdt+lQSblm6/DMndMEDISPI5
5Jk0AzNfQHmyQQ9riNkU77VxR76HO4K42CLX7H14KH/6/LzXZTcz9rc6QQnuArgfxUJ+5uMU22ME
jdtB5MZsyMva+zd34JyBjD0Sx+guaWAJo94wkgOTbOxG5piePn6F6XDzwaBUXWuTeeoJA0c4OCKx
rKql6FMGAJbgbWrcBG10fT35cdoI6BJfc/I/9A40UNrOaw6BCNDSs2iZw2EOS0UVq5ezMsOmlaDa
oVTQDuqgvtgSus9pUi/gdNEGnKfK/iYE8yJtkX/kyXWZygphZlhWpfMl6hSm+5V7VqIv+yZ+X2PV
I/X+SRKOR3GVNXNik3KRTd8hFj8agrfjazhr/0J8CawfgF2H81nEiWVSu9KQkVDbGjwxTtfOFO3t
UZ6OOA5u5uL8mDkSd95MzlYD+tWPZZlTcxytOk3T5gpwtGfNAtUdVvHqmdOpMBcE9jkitncHpICG
Jdu9u9VnuipPGpp1AwFTrZMteh4EZfCsVi5uN2xAi0iYq3pVt8s8ZPpKJ2GNYvHyL9DCihHgeYso
v7+auh/vs8EVOzCzCDDjEwQ9Qfcf4NFa4hKhg17bRyXx+R1bnItPFu06tpIN5sUBQJYKb8NeiBMB
3XuKypct42pICSJgv5aFyN1KgNB20Uw5aHZnQaGEx9cW6g8xVxsIV1zQxqc9skS/fzE3h8YomP57
EO9tQFJ6C+XjANbNA+WcaBec5uyiyaSLJgk/Wd6vqB5sojBGWQ7IKYLTaLQaW51OdvbXqrV1KwbQ
Xfs+iIVJVyHUVZjzKpTnfUInIRhb9mB4c8W4CkQlVEbkrqvDRT42HHpLUgsYMg0un6KZJuARRKOe
1Ek3l7F3YtHLkffa3pQ1o24MOFMm36PN8xwTvQozQ2jsN6l3O1Q0bq7gDZavh3m1BPkOPMi9yn2F
EIdNQh7E1j/PXhpEFZI07x0eMVwC8DXa80AWFxl6NhuyVhcTIO4MRP/RHfhQWpWkR8/k6yBqZ8t+
CgDNRJtckZBuzcqwNgJRYnImb2ehqzis2UgwMbw2QosqanvoTopUGbpaoMSeRwNlkacY4UsRHT1f
Ak1HlraPp/mk7AW3UeHvV+nsB+vtFO5pDf3u5NcbVVsnYo32BP5EG3fE1kHnhSV7qABNf9zDp1or
cnVfpr8gRWq1AAVM85jsLbuW1TWaSDqTFFZdvNXDb8bc0czUjGSpi8zc5gFy1POJxAsyKjNXVJ6q
06X+20a/Hi0ypIU/4v2JfFM8cBfyxFN4B7wsXOXZofm7raLG4TgS8UkfM9J6GlyQTjmDTE2ru89k
kZsdGBWG6jjBy6BrmUEEOYYp9IhUbxdxwYEUeiiSGF8LVBcAp9sRD+HhQSbWcgCCpcSvozkRWqED
5ZjzWaUhQC1Wfp9Du9kJp6cFmC/4qzIF0Y68rntdKK4DVk1TAWxtdFDXdLFlQxjd/9jYcUY2f39F
q/PZs+Gb89KM0TcLy0bs0oW585l6bo1zTqcIHv2/Vgfp0Tc+a6yQby7R5J4oL0j4zhWUUUl2NvDr
uG/2gyDElvy66Z52lmUEASB8X4883+iCeD/JFIz4v4ZmOrUd3R3gLsFA8++g4YULcm6xco657yqr
7ZuuLYFxJ6OtxKdJxe8ormVIe8n2kwMoMyMEDXsIehijjQaNCsrPZiCzo+IbxFIzn2nUjNShfkYP
zMWWpyrT3BH+YI1hGIRu/nEEvEbZi60P+LJVA37WYeNzcFebHaxxTEvISpXJuyiRRxy4oeV+6cmj
61WDDXMfYH4WvjeQPnrAyxLD/OOE5+HBPpN/tiuyFOV/dsyCRG2oAgVLG0yKVc/XCviKovCF9czD
jZngC9fthYrTEwaRPyiqPTQdUMXWEY9gL5y08Zoi1SC52tSj1DRdlxiDyN/AQX/8YNtNp0DeIiRt
Kk5d+GjZnbYX0QsJgF3xsFpBZH/MdbDGGls4uloprQa47uPpFddVxuT25JjpqpLMCYJYgnuyM8h6
8TpAQari/+RT+p8FWwRdfML1HVjWoa2vQvXjfmApokOP3K8jNxDqcwe47CJ2jiKLCbOapU+F+ct5
/Lr4dIMBf2+HSQqGmrT+Z2zMNxRO7Kv7nSR5q3AIdAOGVx8qOFpwKpitFLCIV3Mt4oDfCR+qtwAL
w+TQPjld9HZ5H8XNKKbUqQBrSZ3oZQfgVYAmIYaUCYx7KqbtyktdL/XW1Lf1F7HSUkRJ2Ca5Cdv5
kdlzhgqQdKjQPYPODIe6BYdOSEmepPAipeffcpyd5vMkSu25JVgbvT9eYIzK+oPUS9q9Ue2jJLj+
k6juiNytpIQGnSXBTZXJgWM+o0G+ML3o/QN0vmA3tcxdxKkm+XJF2M6W1dk5823moxS5XR7Lnryb
vw6NRqgXgBQvh6qQGJ61KyV50/rfPy6MTfZtHOp5s8G0nbH9jY8YvuSoDYSmZ3HcB455q7h7MX46
45VtbQY/zQdNpfkzpTKvEXZiadeXShbx+u6Tkc2QQZH6BmQWfoSb+8MBPV770n/XLlxFYXFHuZrc
Q2aIz6QGS49g5U/jXjpx0tFKSTqyXGtJ4oPtwep01vb9Qazg1Fy0W7TE1NI424OEfUKepVrdJ0hP
8GLgrne/+X4HTXq41CS2DLLnKsboPGxfSA6vxUFyHAjcrLB1Yr602itbOG15Ncz74M5mnk43Rj+i
LQVmlDU7rZbUuQXqYED0Cz0gWNQ/oweLRI7yijDn8uAW4OjAWSNWgnxn3hx/pooSQSsPblk+2dar
udECaaNTSC3ywzQsamOPD4VRX5ODy/EOSbqH0HQ2Tx29BmsE14RTxpqjaGp17uyRoCT7RUW7bsr4
VYzNVvIxx9A4aLiEn1dAi6XX3Mnw4mqlnI6slNBn0HrVIYrm90t4Zs2CBsJXuiZcCURb5LpqZETb
rjNZ5eA42DIuaKZ25FezzcAdtsvPQt4H/0dDLwgXN6PRXaIWLZF+h6k/sn5p6MJ9Kq1VDe4F5AOD
qLgyeiEGswGWMv4rHbnXTW5CMzaHXDfrU9EuUyE+y6oPb7gTy+W0oaQduC7Xubdy2SLcUP9cLorI
McmcWDxV5NoH8VrnXWFJGucDcKLV2JQf/NZNJKD4gI4vaGhrQnb02TDsCocZPYR5xQXYMgb0H2wk
dbptXI1Rz4gXmAEgEH1MSqolJ4eI4fzlcUK9velOxYRDCjg3mVb+H38YtjYhnFDsVgmN3VSyesA5
cBVrF/gcY6dg0ExmuRQrgue3AeIsN3GZjDgynrtAgUkzkD8m4VdJcJwf0mpm6vAa6S4T2cD+xAXj
XH2AJOWU7p08Bfmvlf+vuHRD8yRspDoRgXdbCRoqO4f4qZbtukIKZPp7/xB7AEfKqNDZCKem4gS2
gXOdA+mo76pcrI621fJVg2Emy1cLBlWLrpVd8G/18+/lo//nNS6dTPoJ7jVtACMeLxYpECIkzk9y
/ejBuZTENTSBWwLQTv5iVhMdkS7Dvn/3ieni6hQbhMoZnXeVxXjoc8dWROO9XVQlGxNme/ceieWp
0aSrjm4idJPzcFIJLflD4J729NNvSDFGRp4kBvAa1dEY24VM1hrfp3m7fwqA8R6ef9fZcU8kHl1T
LS/VE3noMcX9yaC+uL2R/4ogWtRTcFwM9QF5B0np7DuAF2/09AB6p1bNwHMmDKffbjCM2EH/9yvq
EDnsdx6wwqmg1qOKJ59vjP3Y+RhT7rf7NYZ3EHhjVBkhvBqYSacbMuNTnqJ9NB4183KkeDYTV5Zw
7X+tzJoEPN7ndrDrk3Omgou3ZIBsp2LxJAC/Nomy7PeekvQNSV5q3sen68+dCCOUJ9rdcjOfdGvF
HD1pnK+C3UhfizkRmdOB+NM2srARB8atLm+0gtg43AOMo0j0GHVIWxMo+0qgkkPRUchAvlsEzX5h
5ODF4zLH5ILeUTKx3pNi7DLIzd0zvZkzxRhGCbXufzI9eomYvAb31eIiMcjtq4BaEadK+K71urvz
+ywuIXbVELiAS/Tk7fw6Io5od2CROObqGs9E9oSItefCQkQqWTgDdW6Lv1y+zDD1KD570dJkKd7M
cQ5H3TbeJmrVorKtL2LI2bYUlMMotXjWdNlWyVOoTdPzPef/7mZxs8o/NWu2r6DWWOKpv20SOZk2
PJNd7lgMooY/BQptrM0a9kDKGX57vgROLw+zEhRipUaWEoxqNCAIvM/N6soIHTHsG++xYipc5AaV
YyKnlXRJOJXQO+YKkAFkFEeCZlFBXIzlHcZJljeoY5qixo/p0Z+HbYoQCKakhXsuT407VEqB/8J9
kQZyM6vFYexh/pKCLggKrFp8gDZKQOHw0xUxLr6NpxF/GIz5jil3Mlq4lxkVOXzhMFVPmrA+v2yW
kxC/qS+qx07gwgS78jMAgJe8Zk2jYXiZhep854avbrIgdNRAPSRBNUfmsxyUKcwKpSFXmthJVzlG
YRKVeDgS5Xyuki1n8WmhIP9PB928pm7LCwPvJnp8hkkzeqOGk98AbqbmMqdlzTc7ia1KrCC4EXKg
x8ZapcKPlAJfmEOS64SLpFDY0jJfu64fXwpT1owKKZYJtSzgyxzARJOa8zRAMPRbnXAHHwq4Pkh4
IGTfAVi2wvv/roz6DUv8xI6p+PLNy4EdZU+6F0MXhQtQzP8dUpW2XZIvAyDDo+Gfxn+e9NJZWGj3
5K0d+KlVpuq/fNNyyWCKJAHx8GWnMi5QQn1iyLrXAfpGfGnpc8D6EvTevjGsa9t5PabI0qHCP/Y5
xnPqii3XxtAnAUq7GOTOCGBytAW59W6AAe6BX3uPZlBbjDrUHESLbkosMUax1jh6jdYtKPAIBPjV
Oe1fphQfmvWaGFr6QMRDcbaxiCs6OJLbHd/upfELY0tC+KGh69dSwH2DKOe6vac0//T5ac8vFMhI
nVvw3+JpaxVbZOtQmmxAM6E8RBPY5nsXNRxKYi2npDOQGALE1ajK9Z6yInZatPIECB+nto6t9rFc
OWFLJ+69fbmlAd4IEvfoFm/codN058MYorhu71qYtuNes1yZGd59/I6o7s+oTc1e2T5eTTikGxAT
vGHkfoheKqqVGynTuy8ZMs3ImbFMU1MXuBkl534UCnjdPLiSJZnPkbwVomBa1Ytsl9Ec9L9wMN9/
UKmjIKvRrfehWws/4nGROQyocNb/KiDM/EprrqctMV+sSRIJTkTNhhEcflVW2JovsnjSS/BXcaPT
gMr/E5BK2vUYzVCzyEZXDLkykBr4ydmBbBO/HtvVGXfn9ZhZhy5uodotiMfscEdddPMO5HQE8koC
q7NVJU2HlMewTA4XwAdGxob0oKSUq5NLigpASZtDLUwDkE5T8h9hxF2HPGltVt5HSrqkVzSRIWx/
iIf4M+9X6M9begurpue5BzlN2cuOsK1yj1A4cYH0JGCqDB5/s+5zc1uYd/QlH6b48HvlZS5Tc9ql
vZtYMBoWflzR2JFVeoM4YsLlbw5zbqST46G2r7yqpCu7eA8/zyOemN+SAxSBcHljiR1iNv31lLLo
VTMpEYLvdCqWFIJTbQRcK07sSsp2x/Ws7bsz62nbWtIM2XigtSl6K7JwoYEKtS5zcoYNCBEzEgdd
dgn8OzvPWdHFsQFTqxx6vCVhczTsdqq1lhmGfih5czEIKDs5XWozge+wvad1ssuVQ7RN8vQeEKpy
lYci7cPMT1zAZfeEucUn6gJRTf+/pszWvoWi+vG/7F2DwdZA8OKFWpAyYWoBoBgNTGC+A8isKsA4
5aHplxAIweeAzczPfyGUOcIt6Cb6TcvqSV3RzsxH2JGeW36iYDL00XrKV3r9nTbxJiD9fEMrgBzr
mtz/JyZ9nrFZZ9XrehD53/ix62H8xc71wfJoL5fTInprhe0eShQMVjgBsYCHs3jSTRDszG1wDppL
3ryksbPGo9fDwf1tKGgmX45zUSUzp16S8ipaafHi453SU5f3d82LvEtN/Oc5vP9VcruShAhhuxjq
5P3CGZkAf507hxTQeiU8CoXcH6Y2FZ9KW/CgIrrisD00teZNC8G28lHG+jVGOlKI6hoYaI4L2y9k
bIOMp1OB2Qv92yuXQxOPepE5gpeGtI3QNVDa19hDKvGCKzrG9aws+q1hnR2ftRsSS/26mi7FSmrx
xW4oV7qxUz91xUHckmcceg7tdKP2jH0xVQf1snkGGgrdisSM/r9Y8Wq4j/1sWh22ZSPCUNvfusDf
xNAAcPEQA95iavczeIzAy2vBh7GO6kYPipmn7perf4dAb/1XuUvFtjp4DUlCl16UY9vm1PmBJrYs
OXa8mBbTuwx/KFvIOT8lcOWjnvGlspbcrQK+z0wPxXwBen0dTN9maUi+YFLBWHkotzDRxanC6hk3
R+bbDfHWdK+e5H2rLerz021DzkFRFye/pWGl5Y5gAAlBbO4xMPrOVhQws4Mo41A3OvNjTtOJY+j0
wvPygKK1+j4c3PtKEjN0RYrNhCaPCEXiAwXD+3vojHO2f3eVEFPbBRv5a/pwoBTsnp7wCNVw/leE
6upL7NgFDpTXUYG73eAMxsu1x7LJ9VaBrPSU3jZhm0+f7KDV4v5ONh9M3gxEL+3/m4olIPRMLgZ5
dTS+1J6VJiiVfXX7766pe9YTvE6LYX9t+1phww+DfQCklFyIOiJ2Ggip6j01XjUmv6SbdI+tETch
HmaW/wLryuI+UeyH0eA8QgQWAi7W+TiSSpqn/tenp7tFvT1/tIAqcSCPK347OjaykosSNg7FHJtL
sbCyXOIkeSbrZGGmHlZ6xe35itQnntZWMPeatXRMnEeBAAESvg3HsCSmbjrX4siFVg1l/U5XK+J7
mMNxuLo1AwGvDz9nQUT5mSE+moVd3/hhlErRewHAMIjjDrWp88JLSuNTLyMe5QNY5xdarf2RpUo2
ovxKV7UxRUIF/yJ+QIKhol50Kkh2PIiZFWQV2RW32ijV1GyQMOFLBzgzlGfsS3zShsSPI/N3Z/A9
oxGw6enWGGzttLKOYkimpeL8b/GaWVdGJcXa5DVb71FIoI6sIreS3NoaxPMqI+RH237eaQgb09GT
sMNZSyBCvmFuvWSwlLUKqaJfdv5W+EhpSfxvPddUaZaVOCF8gGq/flxxIFzJyFMBxU0viOc5ZXkR
7qpFeIfhB52niJ4VyEcTC/93EXKl4vMr8jZYrmvV6yCWODq4So6I8k0U8GVvAZ+QAOshoblS8L96
4UU5k/0bnDSW+d/7yhwf6F/MnEPTdNDdkZg+f7oGKHc4QtRQpjSMgVBLjZu6pkNh7e2ljGo94bvo
cX4B6PuWGswEuotZo7qyPvR7QLNYDkDvKXLZzb8MRssysyFzOIHYQAHkS2YGEJ6lft4Yfy7heGaC
q76RDFU9QZ6nb4aws/CaTErXv+Ka8bPVqfi8YxzCDXB84hjhtACx9U+K2Tlj9EES8Q2yq5b2KfBo
AflAZP+x4EXvYl2BVQ5SM9Wbf5oSTcy0UpcBHBDbRXfdJ9VfogaMIjEgmAJCwO9CdkbIwD90nIFw
X30Ql6YepYNkpCvBf7x7ngspK2ZKWNCsNZoFnDfaGO10sdWeac4P/tLxMD3o67mmczHgV+u2uKIS
b5wjk8MAMaOVcXkRZEGo6RlJ3f+TrQ4l6dG+0yN+K53SiND4PwRFGcX8wq9DXW8uviKe1OH7HE7S
jGDyuaVFWDLaLgRiM+BtazlCFvjedeNv4tOmSYxhG7IHEngUgbE6HnZ0dGSoY9wMAugKI/oU15+8
STuAVhgLcQ662SzXf8riziJb9/bug0SD5bOBgTpFy1Mf8krSye08VJy6KaHyyxiZtMR00XFSpfHv
w1WGWFjoHPzr9YvlQ+C6SBGE+IWU/+PcChlW9Kw8OgUwgThwDpMWwKz0B5nhK26nW5ZfoFB0I83h
6JSGZS+ZuLKy2/+RdATKZu+0e3++psXDp2IsQhqUQ8NP/ynlUb6uxyl7/2k/SPlhygw0RJUTolOh
YU20j/z0pbe+GnAu3AbPKpf4nRfOrai53/Tevn8vSEZwqkODzbHw+ODxNxAzZb4SSpvAnAIFB+Ba
tfGYZGb9k1LkLlJE8it5pvMVJKrqqde6mZwFCKUSeKSDOXDDuthKR1u7Q5yxV3nFXm91mvSUh6b7
9FtQgnItYpD72XLVlY2LCLO/NUhbBOkQ4UoU4QjVmKv8+yMLQHOD+KOhpngroJKXQ0ofe8pXSjtn
hhWv1HJ3rzCBNa+l2wRSUBhYTL8XW+BliEKfBmECe6cCnfBJr8LBIRTrb0tRbAuIPAX+wE78PbII
sBj7mPm+JTyoqDs3+oU+9L7JsEWtteda0JCyN49R7xAlTdYLexQcKZTtUhtmDbtlO6WD1Qq7GUyV
iOMkRIaei5i3KCD/WIijg1SSJ3syrCq5MzSx5QTEcPkcjbJaLZ1faSFMDIkR6+JQgF8/X9RpC3+G
SxO883g8oFEQfO3yS4XrQ9jfntFVG7y/6gzTwU/1yVyQ0r7ThiP89zXrKpTS2Qpbq5shBnD1g4iu
w4TRXBNSH0JVlAy6tdk/ElsgbdHXgTl3ZZPRMj3GjTMdoUtOw4+DIKFuwuqAXtUXwaDjB1sFvEvM
dviobdvEDoPV6U6PDiVZKtnZ3O9yXH34SliH/6iQV6PnEG5HQzfZVzXL9BkKymxXlvVOMAsdNxBi
4T1G1XVcJmdpG6ihSPNqMGswMBkMvzzqRSPDEKY+0l0Wq68maVvz4ul5IsnPE/UeQzLPrsEIacPw
I/cgBvd8/R/qqGqankzqCSEkD9hDlLLWQBjfzCA/mvi5FzRUbC/ovmDeCuUWKCXMfuTDPmRNicQ5
jN2yfq2tsLStp1RB2uRjvz4PrtYfH1N6oQ69Bh2eU6kBNkMZUWOQ2WfP3NXPr76v+4Za39moeDTR
lJq7o/ppi44aH/tsNN4eV+98KJbXMVUuOzykq0+u5enZtBmuHtLQga6aUVq+3KXC4FgYsKperlu2
kda6+6tTPInTUgI4bTrc/XGw6xh4UOwKkChExHD7lwDJFYNGdulKTICRovxP1TYQYs6Fu335rzPP
rgSDf/Mon4GLfHmN3jJ2Plo+a53BnT7bPAA2x9hb46LJqC9W5x2asw70Wog/wRFTqoHC5dEt9z59
j0ewsmAEXfwF6ewBPFsI4Mx1+jrOCCOpHRS73IWXcXy8rW6rsWfOj11b63Zlu+WSHlQfIK3WN+F3
4qpE8NZClC4f7hHL1GgYtTw2G3PqYUtsPdbm5CJf/kGJuGi7+W8Xirn7ZbOj9LiZIOw/OAmohEU+
PIBpiimzkrQ0lUOwICYkuhVcv0lIrzyvqc2XC4SgHAzqwSfgUXEFBLxBfn8a4BvtVrl3KltW3yNH
leXpBDUT86jexdSFBu6ls5QFsaT9+bn3oPrPl4DCFV9h1AEdT74/ePyanNDj0u4YMJVTbcilLuZZ
GFetN+W2MttJhzSxTRyq5nh1LgwoVUb5r70supqB06NSjWEILHRYpJIe1ZElzN2DqvishOLCRrzI
fmx7DXT4KvbjHLRVOX42L0oP3BOBcitRk0OKHsCN/ZE4JB1sFCsn1BBvqqmKZCHKO54+HJuHifOX
XtcKn131FzMUfTTslsVJduOby4D5Q4hnlOOgXsXYaR8W4NDiEIsanKg7DoEdyDGXTHjmLEJjsYD8
DhNeUf/KuQD0SLTBsz8rRBGcPJ+CZv8a8lOMkCtcPSb4mNf83nzB4atuGsxK7wVOeYZTIN4/o85w
arIksG7BsXX2fv8bjvz78eSmKgL+oUPH+424G6ww50yKOQsUdhanTbSsRhRnmywvbwWOaTYgtnGM
/THMQRrscbjLrJ0on4E+R2lFaNEE0QxfpgNeKHu6FY9CLGcMCuRLHqHgGX79WvU1oNu/kQjl7fGG
9aQQnDGK+6btdn6TtaNnlRPjrhFyh7KQaV/V8YOaIJHvpthOOEdbuTAK42Jgas7LIIrlk1L8In2X
TSQ7E5sdoYc9AM2urdTRk+AYM9vLXu7QPjvfZhxJgMKzsSFd1c9e6BzrEZTLLbhMmjru5NWWb0LN
EPYLfQjGcLbhfYcexN/7e+9M9qYHXA6thEiyq3wb/rdUNy9PZrYbA4LwwiYAlzPAPyYP9vh/TC58
4lgv0myQf6K1TKRfpVZOp5vRjUSLtJ4MkSxIQVozLIvVdIgoOyXXyZLD7SbanD8KTlmu5q0Ye9Iz
0JBhpM4q93PJxn3LOA/EoWZ9UDS+/HiuhUkL33c4quFgkSkFZYz7/LD17pxhO3oxMgRRQvENhf0H
eDldk8BTSEfegYvP1cl2yxGO+XmbXTyjzZCc7ZJiXQ8N8RV/EhQTO/Fqg6WqRazE0ELrd7aOA5mK
zduLVZ4jQJBAicCVxQ4+N06Udw0MoauGyv31VtJSFJM6Zw+Sklfx/GuhT144ADCMRuuplEGIJctx
Z/AOFZ0ziP+8u+tBO/cCqoNn/WT908+QtL7k82e3RQFsMDJBWK9bc8GPxgaTkgRIPj69rI0rCHeC
GIjFGpnzTjG2fQNQxS8lPw9I6oLFP22Athg+SHPwMNHeHYP7kfzDLga6ve96qWNxBZnVgzrNOR75
FKw3dmqxDF/4QaFYaO41QAJa0oFIkKBaJ5JYiKRnLRXygWDX8TyxTUwwxH76MQ9HGiQ1qUu+OPsN
yAO5+ar/xUkgjdn+Chkdh8e79mw7338TGisFXN5LP1pFTJ3uNrIQR+fWZLTSVropjL8aKn3n8kmO
yhISzCUXcBoTpjRo0mQXoiRrzkyZJUObbdnYf3Q4MhIHtL8r+Zlxw9fomyDJGc5VgAL+zC/z6a2z
VYKgbiKSsV+66HJ++wdHV41uOL5G3GWXP+TPY1RJxwqHiEifFcNvMzos4mia7tN1JmHV/uzCNBzb
nLsY/IZlQA7/zvvZX+Q0TBQD3MucEyycKOTvvQ912+gYDYZyj0u0m1pXfXLNo7d22R16Vyxny1r7
5EKPD7+TxON1OCMTGU3C0p+WRz40vYq1UEBvpA9Mh8OUB92QBQC0K3q32GyGHDBCRwAI4MlIKUDp
3WiW9Oqvm5lxVixDkKr7A53OkZmzndKHF6s+cWwvC8brAISEn+VDe+5fdCd3iLUf+vGefaGhNPu+
CTs7dQ+o3AvHo3e5FDGTHaFtNzY12qEWTlDfY5LiNwq3ESYrzLDrf6PLRB9C+TEgDAJ5h+3ST0pM
qRxiFY8nLIV2jS/FlGBKz3lPx9Iyi2QSFG1LCvZNC2UxkUtzwC5wp0mwi9tzl+XPwZO8RzIw8J9z
1jgdle1ZV95057TgRL+EXV5iOD4bGTLOFUALsRnEjI1SmmcyNpL5Nead2iFl6DF4hyvfsp3vx83L
gqvfaf1Rt+73rO6dac4hnqJhs6FlX7PWG3ucev9yCferlGxmqybmekdLNUTQJKpJTxz45HJthflM
+D+2BLIt+5iBpDqQUQT+uweS8IYkoM5y6B7wmVwbrOp1VahVKA9UrB3XoOMJxVcF9aELE0k5RaAp
SDiWGc0mwKZWoXzAX/aor8z9ebUAtxB2dt6hFEu6Xx4xIba0k2FfYHgAvUwG3RGjVk9wGP9uetsX
T3itqS4qNALBE6vCevTiYT1PxxfSTqRrw+zbI8XztX0wKuZHW1cgeQHrrxU+bVEqC1c791RNk6/S
ScFaUUCXg2kUNL4xE+WkoyBLbxOjDM3xq5ZYTa5KqEmZf7WiqNXoHTzrhD7OyHZDnDsh3SQGDt6R
6fzx8vL4+TTqzVN6LrELg/LU8FJ7GVd3ZRRlRReqJg2HffgnTvudl+VDxrjgchvCPswHypc+Nm0W
PXpdmVJG99OQu6UWFEShlmZGSfYJELTnZjklDxqj/pYqVRUquTHJgEbHtNFI6ThA0QZ0uhr7iUkY
k2UJZ9TKrQ01Q2Ce3OYka43HQ1/uFPAdpQNffG450zB13NO/GS530dplBNXT0ZTkugoYEr2Lt/60
ESEAuSUaO+G+tRRV9WS7JMoRya1sNgJl5TkseP2Nsixt3MEJCu3FoEJPB5raQHRy6Y9EKlAzrMw3
bqXiwtXHOMK10/mHgGmvFEPzd6loBancBEkJj/V7XORmftl0nRYOobrsKeCkb0TGf6pKb3PguHw4
WYiH4vH2zc6r2OxHnjIY+/evRLohsawt/VqH2K4vVfrZl+CpNLxHN+mybSSCxEOIUhZgeVQ4DYKV
W1MIa7tEOKKxFdzKmDl8Ciw5vT4Hn6EPdGLHbvhNEVfCuCtkcZ742AzqtKqcoXm6fcWM0UoL9AdT
7JQI2yMlsUC5YyIrEMedzip9BiXNrV2MtuNDY4wRZXSPeR27mQrOk+FhRygEnStlhmqAq+dBZu2E
OdHPCzIiRcL8hyAvpsQYgKxb8XFwgg3SdvC6x3Dmc0utuDTm76HSN7nTclmriN1MPoY0f6qS5xj2
vAKbYYe+N5UwmHHd/s6Dlz79IhDCEf9aAj7cMRS/D0tnWijPX3PcqKsKX+8TY2TTSBTWhwKXzd+u
xZVtOfK+VFlpr34785HOs/4RBZZOeDxUxeygakQG7ufX/tM3enOs1LmPCtGHfff9YgjPhxtjAvW4
SYN7aiVWJ6CbM0dj7ui24d2rWylFwZx52YNxVOQxEfNyi7JWGnvh94CV83uI8m3ypoyZW58q9c7d
QpUvE7P7atVVbVV/Zq5G5AcxeLl9w6Fvgt0gzHT3dsLk0LMeuj8epSy3xskzR6FdW2fCMfi7oww1
ttQS5ZEPyYylS5hSGBg4KMKr8gSryfq+V7FwNHKKu2UZJchT0D6emhHxs87RRbn/hQ48QnOyn187
Gfums4BNtpKF+lHfDLWd2a7D/R4mzVxAWWG2B2NKJe5mtlYpd/5mKMcgLxO9yiJq8ucS4ZRiFaIC
jEkyt8DtHYHcL+wZ+UQriCEBj64vcsFt82BpAovniycUB7f7LxukNi4l8tz/GvFSU36ty1+HYkSZ
0ZyHRIAaXuZjBjJ+ZY24ZMpTQnQl8MW3bElINFyy61/scfgvGLNPEV0+80MtB/Jo3I3FAmkZzNuB
k6+muUr84vqZIjvQeJUIq3bchudXui5dTaY5/Y77fQoHOqkSBBStuNU7vcfh6VDEUEBqE4F3LX+a
1ltFwW3LjZQHeBH3KunvQJnlzcx7V2xwjfdX/ISvKxXCA5Wqwo1CbUd4SCjyfQWN3aXi7amit3Qu
l5nDlazwTX2CVprH1xpdnjUzvp9Xaeuu2c0kzpyYoaKDR0G/Nr+KMNAh3mvea9alUYztHQSRvrqI
iN9Zt0zGZiaAJLjK+oDeJuWiLHv91hxcnApQ5kRoOycQf6gkdGYgVG9FRhym2gYAUIGcnqtTvbbo
+1lBlfYajFklXrigN5EtShswhuIv6nUd/Hx+kzmBax3KvqvMtAYQc1s/H+aYBFH7OAEuY5so0gLO
EiNdsk0M2P0QN9EcFltFgXNf3efDrBUaXj7zunE04A0tB22tDJbl7FWdNbweIMAzDsx9l396Wa4B
ax1DE+OiSSSVt7Q9C9dm2a7YLNY1Ldnlz5fVQukx7cfO6GKTRsU2skzMDL/YAuiqoWOtfYgltAnv
8EqUktaErYXh83WZmGha8WWdrutd9qadyTx98IAHpqFC/r0hx48cb6npM58LxBO7CMEE4J1OkHy2
Mbhi3ugsabXKByz6uJDh952w+rgxHPSF6hs4yFq/pRLuMyx+5gJ4YHfQQRzobOWTzQR7ycfNrawL
5b1Uy5kqIyudqRxJDtBbLPkncOV8sN3rXGwpvnbVifYEb14hRHvVMbGWodSBJlSVgC+aeFm6ibZv
PdouNECUCMUU7Ra5fZCponCdGxw+VEQt5IVpcdYnnyhtDmJM78hg3EYIIm1gZVPggAoMdtGeRDcz
1RciUqD/YfTSVCoS8f3dp9ibgBd8H9C8Ye77IxYhNwIwiUV+xcM6RQoppd9dTEEPOutlNIbAqXvM
BkEHk7iic8JoM/vhV4Kft2c3nl+innC0kflymN8ExpkEjxjTJ5ZS10nA35xmaOqW4MKzabVFhFIn
DlhT8/7d/dI4WuL7t9XPLPpfoB+tqYXzCjs5bNBgxF8WYBQKu2SEKzT8IeX/W/+J+SN2xB6gs90X
z/nSbsNoI6IscUNNiC1pgpPsm0Bf9F6eybh78v1QRsSTYxt5Ug+uMKOFU5X31T5N9j+pD2kfVsvf
1MmWLehQitF7QbDKhHA78zRsCcR6cMAT7oDx3nsKE4KZpMw7JiWhclb0oErn5mYD1pJyOqEV9h24
qmiwnh9Kgve9Cfaj/U83vm5jOdNeZ8QxKclJxwvFsTr7Ug3l522gu4joqh7OK6MxptlWgDWgYxd1
S7ClPCYVoVzTtEq+ehDY1X7ZjQ37E51YljF9PDPipFwkmGIy79vXe6jcnJtBMGqiMnlYAZcVQO9V
Mne8iWz4k2atoEGTJXil3OQlxJxQVUr9p3Qd7VjGar0dhyuNVcTlGMSh33sHwl+ko7RHiclZNGjD
+Nh3ZlUMzKlJafDVP0eyzKN4hdIYaMsPjhajC0nV8Jj3Vbwy4vdcOWMr6OFlM6u7Ky0J3zr7ZRIx
gf4/1ZCEWlj8FJWhShXyfsEQQonATGSbFLzI84Y+ukAViRtvxttAir5D1A0PL7SvqwP09nmnyQMe
jtj6HfcQDMWfAyThpJr2ojDQfRj2Tv9dzafPT/R8FFL8hTWVnVPxejlbQJRatreffwEUjMInH70e
YIlo18UnrbqKKvBLs5upu5NKzCO2nX8ljMkAOaJuK/ggvBsb/R7Z1OGJ1/7pvus6k+XsoT4+KiLq
GVYudSiiC7IlAH7ZsVaXFJs/kcwsaQXpc0jJ43vz6N82TNAyjBrOTzg0mTgERw5xMI4KwgMFPVGT
Iv6zU+eQsqVWYtIXb1jgzDU6CQqXsNvJljiyOMJLjhgJafxyfZBAqVda+XZOyOl4EM5rWXz/28h+
L0hG7w8lOZFwJnc4iQcd5F23BVgMmEw3Qe5oIH+C8N60pHYLmvfklaQ0zpq4ktFPZr/sG3W4Hodd
TLIcuBhjzW/UfyRR1CaJI4rv3++W5qI3rCDTc3xrQmplLa1alcDp3s9ImkfYJI8XfITM4NzpB3E3
GP7FqKKfhInI26mVj8crFABZd87ijime0mQoOVkb1lxmwckKPuOeG0omBI1coaekNeOp08SYTUIH
L97UXtIUk+7kjnLAP9Ic92VrsgHjlG3l+t+pR/iCd3NzYpmqplQcTca/sxe0ww36ogZ4iDdi7p0l
faI3ahzjMSYkCplItiTYSCS0qb2EGO8ECR98vsKelHgRi8dyghm2ilIEJhYI7vPKgBaU5Uhox20t
y3skIH4a2dCkdTwM0grmaRokcsHUMkacDD6oKwXNg7S+lkut7ft72mUYAJPqhU4TdH3rYeDfna67
0pg8DN6X4YPLYAlliXh2X/+UM0ViA0fu5hTgc8HYWctR0w7kbb4JxJ8Y2LU5m7+OwledaODVI16u
janU4nbWBgYFSqihwymSrYz3yT+C5JyrgUAoUQWGCvxN4cyVX75lKiE5+17W1G1/OM3qlkJo9fOz
G41SFSXePRfjuBowNBh5quMFnyr2uP88Et8WQCxbwa7Mw5MvJJ+Ee/WfA+2Q7DDU9zpG9RPUOPq+
D1DMansxnmpEsFvz+e7MSXOsYY3prOwhnTi+I1NqZ7Ra52N/XEE/IsMa4XbbVtaNcnxyFsME6TGZ
c6ooYldGzsVQz5I8EA0zX5VvBYqc2pmTckh1+G4uU9EJ8Kd477hBXEspCrp16nk/mdTz3S7uLTnw
S6hrTQhbnPddgludZg+Pgq7v0uNfkizGbnSdGUwhLUZ/+m1304g1cKluTkwYAjzGIWFH9GHpviOE
S2DVCmWfMli3iFwBt28t0mi1voMMKlGkTpv4JoKcF5V5tcGpD8knaxkRuftSN+z6MsJr0iNFBEB4
rFBweylPXlYRbrA1v0X4hPhr0w0wvPrT7Qw3tvX8jOVMUMpaQpez6tPTWrGJSbHtqTZ1Xpp9fafS
TSplJjxwZJJxylxeBBzVka73ykwwB18DI3RMLMDf5SRpEbQ/3j5+COXAg14fo4b5t65FQNSwVjRU
IGBz3qchDbJLgxlpkJDsbItGf/CJiP0ctOk9X9P/XfQS64ukg9jDJ7Ed6kyXFHGdYEMOkHSRTja4
ufORcwWRZ7BtMflwZEnquZ15NJQ0O9IWUkevNTzdGCue4o430/+9IYJxHygE1zsv9EFb79eNFtzP
AMwFARhcvplI051sxNF5nakQ7j1RBldEAwihpB4HrBOutVA0sbZQfU1f444Sb2248XuWAShx+U1N
vOho84l+NrdiDhb1To05860Q8eCV/4JbFqmbfwUoAmaWETvvWCoNKjYoV4MXrTnsN3lS39K9Ny3z
hTEmLhqPgp+qmTCeq1w0YDVA9ga5XwJSudMlTO6atgrJH6bkkzedtrMM8E9yemK1S2v+NpnD21Nu
Y0aah/DZS0hWGk1ynXJbadyUCcalIImivg7PG8Na0DnEU7XKMTpvj+CWSp4Ukbpt3vfDB9qTLW4a
GPrfJu2xdbou/PxMN56RKzV5IU3wLMpQRmhd+AJUrNUi1GceCnc7SNd/h03veCMovOj+9jr913R0
JH54LMrzAEiqnnlNhRm0vaG2X3fTfwGmabu+VgbRfzbrLjm22n4tZ/2mMpevA7TwQb35xXxOtRuF
x/5xsHp5pzkNSBGNZHShGiKwVQZYlrQncVmVkObSaGtAR8vFt8C0Zz+mq0ifg08wGq0tCwz2ep4S
63HOv+eXqm+hA+qyJF+hhGINii2cE9tYIJClmfqYrCMIzRDHg+P+djKV1zxc5pL5gyxes+r6qgmB
xTI1cQSaErJMuHG1pWs4oho0tWkRLNUcL3TVZ8ygzog7WykFamvq7I3+ShnPECfIm7DV5kJSF55O
RgT/4UNGcAvU7suMPxsN9u+hYSayZIc8MT/Y/WiFFaMbs57LOjk2py3rQqjOL0VPaMnDb5Qktnz7
6HYAGhYQMNrDjNjRdND+NqVdvOaKfctLXdsthFmCqTv6sf8X1W25oX6ZN+1hPx1dBeMFURtvo82S
JId99qthKWcimyBArHMDS5gWcpRgnHsf+opuFQEz5jHvrnKSqlmCFE1tkogZyv3bpd6VqOl1ysxe
ZC7ctWUXdZFkI+C0esmGG8UKFZ3F9lQq/K6Vo2l2bqBkhU3zKe31X2SSYOnxezN0wW8CgQ2vQfEg
MMs4tnWmREg33cx2IZVrBVqLol6oPMSMUsburotNIj4TBafRZ56ckyXAzkP0TDpIcRclyNPeetJQ
XIo8e1Qecft6eAqib6mXyWhlHIulBRJWnl7hFCYCW3sxOR4PYGUzmXrG9IxvPqu/95bPPfCSyXLl
SYC+UIT9P/OlP/i4F34XEkd91U1b6C8OxugKHYyh+MUJKY5vBvDWwUpbBsgMaeF3J93GuiZjVDsq
03tqEj5NMoZtNFJqFziABxUaGpBqMcu2hm4nFl4WH9CzI8LADuQingz4DltkzB6fDTbuw+BnZ3+f
8gI9Be9BgHFlWKyE7S2blE5y64R+2pjbEDfxZmk4XDMHYref044svHjFfrXxngHKp2NqtuPBbkqg
iEEZD3uTTpgOafni5QgYQNTa0Ahxfc5d7Uvrguaxiickn2zP+FTQWrR64u1gH/arK/vhbvRDE7P8
tX1TVFSJFhytCcGIa6w6v1rLy0pyGd7ncgaLYHGhdaMjeiZHzgHNcbUgMM9IIjWZPAtW7zuo2dPd
00n45zNCNQPX6mtNTwJoqZ4PMMV0lGyyPcViBGHU2a81+kITSRM2Z2Z+MF6A+zPojv2q6T3jopGB
HijxvZHE6/sdPVvy9yQyBLCUOrwGKi9wQeRX74j/38UCm31BNUIR/outDYvZeUdWXzoRL2PhfJjr
WkaKFZw3/os3aNIGaZlf3qdtJlvnF/4FqWNhxGy+hBH2e+NW0J8ktokaoUjECWy31DYAGkKCJvu8
JG5P8i927WMI5mxxjsshq7/bKn0XfqU14f4JoF+fB+/Ff3weV55n7UJYsW6SCWso4b+fi5TNdElP
mPREg9otCXdkPIRIsiiIJAmep5Qkoyejd5bbV5uzZFpHGbmg0wBIzJ9uSel7PttkF/ZDs9GK6kfs
ocSp9w7nOQJolx8zpjhgWmfuENhCTRavRDwqlqX1IUR85SKrk+4g1zc6lKbB6nL+2NK0bnK0PP81
Cx5Py7SCmHM8Vt83NyO46kQmU7zCt1b672i1BlDspp7wXC7a1nMdXehuhVLwaW0kfqRBRfu/m1c1
c3VjaGK4o4Yss8t+2imTdyIlXlYlP0vN29dGqsWCJ8hjBJQEZ59ewC/oJHTD2jEQG8XjY5NErDTO
VzBNIKoquTePq93uzXDROstVDuecxz9WGUw+Iho2DsMJ4cwPODEPAtvWn0h8Pea0xiT2i8FNox2j
oVa+PIrGLRXyYTOQRNMJiaxL7XtLE2MlzELZRUkmquFj6xXzyv3v46KIfixdHJC/Rpcl+aDaddFJ
JV99mVgqY8/lQnxZLEpIFCEU/eXWjKW2JazvhrdKcmnzHe9a6vnNtgyoLeTxLznoOk1S43vbXZIl
cDzlUu4qQLyhvUXcov9RSb+zodn7xnlwceK+zqX0Y3ClqKgfZTHfzHHYWqp0fIU/5BPFT0/MVsOy
mOZpmwoe0hl+jBeJ2jFpu7+PTXTjv1beJENzvrLSHr4scioViLmJAK+nx7rxzoJEDSk6EZgYKku6
QJE874n5IjK0zMz0nfmag7m/T03OweAAPuKQudMDfIgx2opfqWbcvEtOhLlNBYD/UBDwWWrdt1OU
pyvB5tY44LlD3ymdYehujPrtTz7npjjgXWVzAg9+fSUN7XIGc9b6lnCRBk+xFw9j7kE5JBxtE8eA
mOuISC9vle+oiaNQkuzIa6V4jyVy4wsyI6KBsF3UGT1YDHgEDaOMTiDL+upNWo/pinoyuJgZEkjJ
4nbWXIld+0pA7qJO9KaHhPw3XPdZOZM/VWH18PO82obTQXHE+wU43a2TVLl2U0Qx24r6SludjPu+
Vu2qrQXFlpVTbj0xU8R5trDKR4g4tQVP22V8XWwI6VYJEOj8Ef9EFjmRfS9REX0QHSGm7i4HWCIj
P3P+nQ3gADYO3NdGVX54e4LI4M5SAoNsH8Yt3s7p2uYBxwof8UUhEc1zCxpFmR11OL66i2LYmpho
ba3OyKixtogPR+gJpxhl7Ul/qprNfNjhgy32XCP2hXdv8XBL+0aGB/U5S4dbF1pshMyOeB9B4yzG
mvY52F/Q8m/mjhyhERyodBdMeP3ZOkCQuMRWvuVTh2z+2MJtWK64qGW5a0VojGXA9T3m6SjERkXq
3tld2aYCp6jU49a2naHF1boiDMOCpYL/QohslpAOe1+rKkJPUUe7yAxWOQF6ccAJQzCNmhR0xB+K
ZXj7C7HS0LGccgvIVi/Bguyw2fYBcZhuJso8g+Jm7ciK/UeSNpYrhU+vzvfzHZ3LFIPPKZrjdIvA
vDuawXXQsScQS05n5RVfpZu+CDms0ejjntmlPu+gFvPzCFvPQ0m3W/Z0Gi1zs+Dmg76j10PRiE47
Nk9mqyAE8al/s6hQIHfG86adS6f2rOPfDHzXIsFZ8HM2hLKoT+YGXWSQe3CyJlZ/1qi0Wj57YjW8
kTuuWsSXMvXUxZaqf3xW/IYylaePjNo7veiy3D9O2mhbV03cVnIf4Ox6msc4sKs+67Ey/eTpFgsY
IrKJsAK4QrruDBN0wVZqrcMW1kalt3nbzwacNowkmPKbXEO1cls8qBzPrHZHgptvZBhV+pPr3EyF
rDmj4y/7GA+6XqLAvCilH7LmCuK86UZy0UIGilcX91LNaKWBF2G0gP2MFNoKGYNtVJtOYpK+R73T
ANIoIrX5UuKVztvC3E7hn8g8bxeFqY0KG4GOxF+rerUBFl7bijOfw3ngdbbvl0/9V9umvZJuaCKL
5wblgRg3N9H7BPSPcvlnYmbrbKtvCaoVx2Wi/TeNHLduu4BrJGTUkHKiz4C3rzhxIiIypaMB4RDD
WiKDl9ZUxj6v5RxvpmwGydeNSmPAO6LcQlkgwzilxfuPy1V4jQDpWqbdlfvQYODpoeQcWHq4YjTm
avVziRjBpuvGQDDl5BwTEn7wFx6S9pO6aT4PHPZCCQPikL7OPHmCEbrp/S3mA+T5WeBsszWjpPMP
DpzvE9UVvWL5egxXFTrWx62rtqrh1YCgd1mEgQXUUGpgM/+G2Cx4PiVzhG2UZh8QMebHdLbAJxVx
4YqWnRBvE5nAGR+8ogKUDg/nEDxxRQjQ12XbTVA1nRZFYfJywa4S9YtY9g0Ti9fCPLdEPfuvnQNF
jq+X+Wph73PZRNIVWTQ3ONskNrQ1zLXpt6yWWffottod1B7KMpfX9deBFUR31OyKNWvk45RoZ2Kr
zCvPiXCAZv/x25xnBJnZq9l/rF7+UuVhOmwSa5+S9Y+ENXE5HD/LRlA3W/xlUllfl8MZ6Adiq9X4
3t9QKQdld9CEe7HWPwG3e5miNwyFB+ATK5x5U7S92F9IVYKhKh/M5qIpbRQnvez8UF6dwr5eEiVq
3KkW4b1x+wSf/6XBGLuRrFZWwxbaogd4GUIVPs5BTLnIJZn6qNCFMheDe3w1TNtkfk6SDuZIm488
7ZoCHkU+tHGF8UlIRf3UzgCctYlCPkjVtXt8V++0w0FrFmqlPh76zgpOa6a9SKuMja3W9KPPMy2B
zV0naV5OhAWTfgNLif7bT0h7Na5tuwslw5cESSU5xSgF8A2+OUOKoDuBAcdhiibXQqQOBohJbNjO
W5aj7DiGeZkoAHozdA4scusTjpPmhTrBy+OuUsU2rFPxGiLslEZrhugzpH9GhpgVnpEAzfAp6R/l
DYwLMC49I9SCfsChsw1XkTRgTQ0OTHpjjl7fhgwlAg9d1coRoFMtio6oQQ5m2po4oJwwwUEZylLF
ICw24V/J9Xyx4P1GOvkUl/tRIDMaOUxHlL+TgGaNw2YXJTe138fma4ZUZgtIPAPpRw69y5RgYokM
ySi3XwOxX3YHt1rtFFN436raI4pIBFmKoLJ+soe5z52fTQKq4rSVECND2WjQJ0sGnBOPU4mPN3/+
bV0rxdoh6CxvqE7jmjO2VWCkaHNEKs/EVNLdrtC+pwLMS0eVUmBahmhrHOPiNKAxHmZRdjWCY5H6
FoY9MKC0IRVfTHh3I0oZevEPS9ecnd1EDfaGAqUR3jp93EKDEGe6eiUPrrgAH1AXabeijn1zYMPY
wXliza+20hTH6Sul3FPMTKuGgCmjkcKobbH49TUxyvts6exzqWIaPlA9yUiHxezSAMKE+W5xczdz
qYG0xYi21QtMpyYo+WQQvDA9rAKmSXEDi3XKNjU0XXz8+dn4mu8G7WJ1wCFBWALtwKW9rCBrwvGO
DAQo85hyGtOMqicMm7AsROOk6QKgj4OI+lflJxrslxiMhVrzJFZt55q3qeDGMSe3lFsH793L20Yk
a+WLkvnJUwbMqRIOv4ho8n/g7ZoCe1pSZKHiRhVpoiGQ/NKs6VOrCqK8Bicz+vr1SlztVNeeTvQq
eLk9wpRS5FR/xVHgzvw1SMK5wTO+zZLAGOrLNswfgxliGuhALRGU5Amz//qdyi6N2ofT9LrHj7SM
t4g6SfeRH/+EPyoW9O9WMAag9U+HcpQ9MuCcvwcXcE+6azT9OOyFzwETFn+Lh13F4HUfU/c3Sdoq
JFQ+FzqybRBx/q44TWlsUHmVTJjb1DJcxI49FYLFef1tldA+0MHjhwJg4W1HTckSBKtTNULiv+bd
iORRNO1W1FIRTyh9QeLQZI0JpRaEt0IMyiZeoGbHfH8hLh6bTzyd4uVk40nl5b3bJS8NylKjRS9y
lcxgQM58riKy+gluGui2LMWW9onM6tzkBtOp7LiN672QKnONk6D6yGs3xysY5ZSfph/BS0GdRFUj
yFXMCOCIsf7AOWWJOkXm4nr5e6HTKbC3hpeRTTXyhLFO1bCQZMdSFNiAC2fDMdUwIEPPb0qAf2m1
rXH3GA9E9gBXkJnk/KUdMNrNMq3mlDKh2LYjTtNH8QABBVSrU/3Zif1t0gvoRevQ41NMWKOHQ3ES
hKJSfNlYoPiQ9Wyzp/l4OcuIjxgvgEI4VqXrEL4XE3rPvHgK0W8ETgf363YXpILJ75wTcWeh/v2o
ZUngkVdtFVUBzZ1X9LUX+3LzoysVfTs1XeIrkeoXLfyUeO5+fODWmlJh3eOFJTFEtLyedJhyXPjR
FNXVoMzGVA1cXU9J8pL3BpXGa4MGttnG78qM86QalR6XK7VUUe2AWGDCHkEoEk4ol2LCH1JkNT7C
Wyt5ScKYYYqYWaqtvVOjNH0gaYMUwr9qrYrJGDGTZEc+Ug/Ugm9vCYiF37DkmiHhtvobO2QalIEk
rwxd7viqOjDbd9PdLrNbH/WcLOsROjjOriMmhY3S5Whq1iO1nO2KBwoM8Ua1sN2JJcl/Ybgb1K+K
Ihc9XGMl+FExNUPaYmF7xfhLdTCcUADJJs3HdwHB0ATj0A8QokFhthuY1vLtngOEerzSqexFMxca
3lxZgbH3sOTIPWxalelb5MM8xsS5HZWklECaFZeOQ7K2tc4ztIF/f6zxn79xeHLcMcG/l7CHPEah
skbCKGcTHRBYoiVKCT/HYBmYrmQthq9tocCcCwALBwxvDPDJvxogVqtaxqAqlEGTXTooLRBE/E8G
uT+mWknT6FEpMOF/pprXZhg36IdMR2AQT8LQYBXU5xEgZgISMl4PtDaPdPbG4vpfbMsSyjutlbJ4
S8Dd+qDG5XbNBELv6qDnJvAcUGRJB84sh8IGakk7rm2Nl8rA3kXAzZ7Td5UqZv+JscHsGPMWLo61
b3B1DkbEja0SqfQFNWOYlbZGyaCDmuS9zL3TkOag1UF81vMemsKknT24azfDyBQhR3/ReBoPZUsC
E+hyn1OEKLmACkgtPV2V3WaB2gFxS3eY8TUMnSfyFLstwun8gzB0089vNJ/cheV5hmxYP9EwXzW2
36CB9B3hrGv16bD/3Pt0Jvx2OgPUb6C5MsaJNIfGMfdPkpsRFyDIj2j26jkIOTp+ABxgHtDKEV1U
Fw0aA/J5yz8Co1UX71RjXfLWDTbrucu0+ZtOT2OXTaiMdOxwHfXqXRtTpWeunSRAjE6KKe5rtfQU
8BnHtrbqYfbEnlth9AH+QQl+N2+Uu+AV/WzHV1pqDq0H8XAzDvIBiDorLOl5XanVQcVctTW6Ol6b
50grhPs4Mbi7ePo2aLzHyWmkKk4LeRlE3kJB8yyrpp6kZmXaZwkCmpBh6eoeS1XcrkIX0tSjt59h
/eg1ieyvEMtKwDuqvU9MmjJ7FrMA10wvVsfvfIrcO8daV2aBbFUIn3n0jAH4lJXuWUi9LSeLgDRB
xxGw6x8nDw8pyd/Rc3boqv3/GCALA2pXJHR+aAxHPUg/2SPl9VI8vEr5JqPLu3CmffsCJczz+PAT
SCusHMjTED+bWtPjxnUmRU3SYGBYCpz7/fqzLR4+22EXsfPFlcKt9xOxZtc7eVsRjKqtvtx51GWe
7oPT6lD2MnTMpbhsMxS0U0auut5z7m60bc7PE6N1pSWYEQ7MDucTcKHfv2NPn+1sFoDFXXUkB40S
7aCYwJZFSR9LjjK7lxn9TmD1rTreEOmJZBKSAmH+RgXcPeebRNg5bCSdo7a7LeQLmoCAxexHiWK0
th7DoIzISA8lIUICApWEvSMfHYgQNJV+3ylfh/4v9HOxPxG1JG6M/f0kTKXjBDnnX6zq3Gjy9iuM
Te4FHKMuqiWgQ54v4rpbnKitMhF5tRFcZk/g6EAEN3UIEi285McmGDNjiSV+FgQiKkxrGQs3EDr2
5zfdkQM0tY3GYXWPfOdulDI47MEWAlIocNpRfKeiiNdSjJSf1t/BktwupdZJ47ONDA/5xdUrfTJd
9Av9BT6svuQlQnfc67WKtBaDNFp3bU6ExXhQbqIvFm7CxRjTs9FLVnfIuyz/lmyOUIWpvXpjbpIm
YCeD0pr6fQVgplvsNfqSfP/LI2a33DH5JADTsAkIv6YeJ/MU2bw9RW9Fhoml3g2cZ9C20xDkFOzv
wAAAHlNbahYPv9P6BMxO6UTNKNvykJ+8i4xAp8eDpfH6Q6dwqS9p23rpNWx2MSL5ekktKFWHaGny
Ru93vTmzwptK4JR9IruxE/D0PuLOtfE3f25lzqv0piY28/EQv0GPT1x/1pe+y5YFFzk2vrgGgeim
V9ZxcLQxNEzxKKNl5l3xVCCBJqkYO6gPVdv0AbPaxSUn08nB/Rjf2TD9pnWAtROyu0zAnNo6dm/l
qM98uVA6GLnleD7s0d0id0tAZNUKgxd5tMbYIMcw2oCFzKowfsdukQb0CC6D7Fb7TIx79Vztq3lo
tqbL2zoJ/oxwGWfTWhaBMgO024jcY2/+4ndxgZLlX5dH7eDfHgu00PgxVx63Mdtm6XnXVWoepBBh
609rB46uxdzU35D9e7peGnKXQH1av9uxASExpunuIcsoCO/NwVNvQivQOorSRNgQ1KFAdnXd52Yd
EQeKCqYKUWTdwa5Rzl+gnZRuesm/SVyTPrUKcuvLI7iudGd56TFZjKhr30QfD2Pc5RerXsdIGLyV
vji0wAV09imuMcF25o63LQ3bhzUK4crZ4TOxloj3jknG73wmtrsHfnuQRfHaVyxGYvYTbFEiveSf
+/AWzi34qVdJO8cJ/Hw2kCRHqKLybKnMe3njsT1Pxh/uqoH/fjTt7/wxHy7SPtxlpem3tjPANaGT
hozauLIOddA+p6XJqxiVcrmjKoiOTdlR1jABWlFOlvMNvQK4XjLQnl5391FMVYT8jhm/7Yy63MAe
zlCYdyjCToAJBHKnsWDWQdgUAJwnh/FdnKbyHld9kx54aHDfrWS5A4xX6Dfgae08082UptTXCXL9
+cFJ9SMGeMxUaAh5TcdLNxRSjKREEr7KgHkqrLMnNFT0hLnGKf0cz1v4riYm+S3v7PNeJu9tCMYT
k5qVU4kQVNnTDgsx2zyu+Wfw5Zadbkrz5TYhKFAs7MNxCFT6X9j+sfBoEtIpNgchY+Owrl2l1XrG
FgC5ujAGolrySN/SMAsx74E79tC7Jie1/10hyLh3gr7m5oZCZGx6T0oHTNnxOu6s1JNyquHonz2Z
seDH4yCHCT60SsJQBXDISYJgkA5yateiMRjn7OVXmrOt+QfZgXEQdet/jurJMOSr2MQcsifBWRhr
eDB1c++1jpVRGnoGOm5hvG/cKn5zqILTZwBmHodSLsoK0AYrEobk/r2PoCfrpiAIIzULoDTv5zWn
d/q356HesV5bTJOPLmwK0aSjhI6GH/JMlVYN6BRko/I17n3xiS8tBwOUg53CKqQW3+2m7Yo2H3cP
CpBIJoxmkJGT07fSSge7ZKPGpBqrfw1QccSxrm0WuEODm3bGPpcP0h1eLCFqQIng0rYC1EUxLROW
QaKFmE4hyLU6Adp27gq9HHIGggsieYmjxQlCVEu4f3oFhcXoKE0hLxfhBscnx9/g6Cb1RwaHPsYb
+fbprkKdRvj+7wF4Wpbz+3dkqm71hf+tSbnrdQDvfe+emXVAB7FlSoxWRwGtBfyzbitELHcEzmrk
bwV2yKiiHmdc+mvIHvX5b1pLzW5q/QsYdOf6B0KGSguLUWaExDGYFIko5GsijYx6cINDxvPJL+dx
LKDhghGVP+GStId5gxYPINVr5a30ak8MQHKOpcwPyV2DwI77cnamGu2exOb7eGLzfXxryog20D1z
eYYtaT6VHikfwhsbfxLbZNo/eC1WmKFIX0/tLdUhvb2UTjNHAEk0HBjWZDKGmjp3Kbxr5QKbPTO1
VebGFeQN10XGujNZ87HYhKX6Kl5oEkOvSPErNCeXjQ03MxZBL1frdLTavqWysQsj/6FnWPfiB8An
EIRkTY8ZcnQj7zoaIy1LECv7E2sWujK5FNLS8iwP3VEv9xdWmeiz14BPqF8NsOUWZk53DFqarKUa
3Ef5VTSuVoqbmqz0EXjDuLi09aLApOehPaorRkaXV9WEmDpmcZUEnjTT+j6aTbJNRiniZOsi/Twf
nMKuCVnUYuLOuKFnJPLmzgD9kUWfhKRSkRd5NZCSQoG17a26KvKPHWbkKiKZxcMZpVPFwImNXXbr
wutVTpg4Z7cwMf04DV8NqaYtd6sMZe+yscre4wt+dOIEgvHBeUXJxrzV3/gyu/0Id+XWxGyQTd3A
y6Le55vMLxMY5/yXC729a3Cv60UR8awCDdJ1ub0H8PurDWtHl7EVAsTLHGUTerKTiUT+aM0sTuFy
gGEo2rAAKclMwcSrFt27ITzcf7Q3L7PDIPuHzzHFhaeYsvnYbiVirdUUcK6aXrkvqt7U2zmD1NFK
LT4cnRIWZX1oFPrOrhCFjWOXyplpA4Vrceec/3SCyu/IfFDClrCsfI8TRt85Y7hC6Aq79LOUGkUi
d1HO2d1dhO/DEbWFHsJtHvXoUiBbFDKMszhN3yarEcti9O/zwJPzaguJON343Qp+weroZEdxFUzg
VZrn5QQ2SkE8fqz1hnl05T+CPJtumKqDn86MicsaGBcGzBBf461NMlguzJ4NqwiKBaH/rsrZLbey
Uesix8tZOohWcIJNU4tq06ABRG7MsAjigZF3yXhaWTh8CMriRG8nYpp3oMuIgWQq6U2To6LmLTKE
RAhVsqQRuFVBz+4O8QK0B7E8Fh078r/VFWwFJcLIcCSEFxx+J323lgtz6irMtgZT3GLgrGqXcyz6
H+jWXzC7G0XJt8Xz9medmKm9hi00DiRRGZggu68iJa7ppXHL0Gdz//IQBi81MPsKT63fdiDaGsNT
6hEOLAxHeC0qnMB8W9XAYXYhx2h/ieL2Ed6yHPuSLmb7UsvH4QlrHO8pe/OCtwID+O6JXuFDRJiy
khsTsg3tKeZTlt3ovC//6QsYe+b7sya3ODtxz0uZCijkeBQhkv78WS3IUhJatzZrVgSIXOjtB/j7
nvhO6OUdP7FJ9B2ZEMJclsu+JzUCT8bogf8KZqb7kSmFWswrm/5f6b8lwOkP6SRcn7dPvUkmduZl
RNdtrXVx6NiPGBRgux4dQrvsUiBC46/MSC63xTufTmoEuh4Drda3qCtY4hrBJJh88QVz1CPcSDN3
JzxRoFl845n5gdbqG3QMDLBaUZncU6qNRaxl7LI2R9c3I+Tti4jbcJdOOT6hOn0tVsXg29q50Dhh
cQPGs2en44FOhcDLMX5lRcwNn9pxD8bw0Rg+Wt2Zp6QdNKfE76ewUgKqM0nR83YQ5D2bOu3d+ygS
HUn61m91y/iRU2EbymFgkv9f7GA/V5PUiqf+smL/vy1LpxpHA/j904pEJsHSt4tfFogdJ7Z+kyHK
DyXmMWL45xPrcBrEVOf+Ft17ByZrhG0t5pS47GuT70og3YP8cTmiUi7hAjSBZb4g4iA2nLoUXtph
SjXWS0EmsuSrQOyi/zc8XejcddDcGR7D+LHZRS0rDVL4ILCjGKCJ0IKCjRmZEarz1O612froEFkN
jKi56C8vj1Z19sK/HH5AihR/ued8T7EoUxPeflHU2orTvU8krsZaxgBDalDul5RMJrAzdMlmiWfC
Xj1Izc+DOsJOh1HjEsK0RzyOsM5Gymg8K0h0HPAHbiijAUojf2PHSXj18cJQf3iCckDHJLuZr0gB
ke64f+J1gsln4U+V7zd6WrUjp4v8oy9TMhGm5918sWHXEny1zGeWSlIqr4nT+Bl6Pqb0EjYXvIlV
hftcluPcX2PZD/O8BBRQAGCqMCvys5667D6l+4vth7Qw4qN6yRsabzWFCB+/b7Y3C+CvrQNU5jx8
pukzK/wuCvvqg2HBw0dR+Da1w11/cL+TfSuxiZAPwWFMe8FaBmreoP9ODbISWr6tS9hCEilK4XGU
zmmPUeJdNVx8aSHO7iPCSX5UFAh1LVU1rHfoIGb3CtG3B3VB8dsCz1YK1dVXsEQ8tfNF1dsp6al9
EQ0bDfr+LrE0Orsd8330XBVEz3pC4ocmNAS4DC/fhPAEdeA2ZDVp+yZrZxzC6lq7dNMnI/uCat6O
xfGYi9QeZTev+Vx2OtsbppTinF3jlPKLKvrcT9HIzSCVBhNOD9EoA7YvCjiU38I3vigwzjcUz+ST
dPghufmQjzVVPgSoaKXHCn3JWvcB1v7zWsOCnTcsqGjVcwkoI2d4SuXpfCl0Tqk6ucBDaaabT7di
fWfoCllReZlum8bt7XoejVOB/NSvtEqCAQjJMPdIBdOdf//d4/vmfN6cgRTYGaaKfqzHumCMyOOf
D2iFuVEk2Mg4anzftdW/CezG7hjY5LydwjX0fhCxVSNh8dpCOTO5ZsUFwL5niUThffKysxNczULN
iLT77Yrfb5yP5OaVgoFaL4qOwrkXIPvsICEZnOT6d6zKmpMhn47POq1jBfELaj+7gI+/HwVsZ+Ox
xbOEY4YKKhyt7MMJ/vJw0SzdMlfrKclEvCTLQFzjXm9Bkxf93OWZotkUmEot8VIf7i2jPEBZ76Ly
sMH+L9XFy1/u9IZOXy12bPIvlNbTfEmDvIjBGLnP2B9GcTQIFy3hcAWZMvioiqpXD7COcuokkNLF
17Lye2JgDABzoootD+9iJQnI6dJMMR9z749hbcJM2Y0YVCP2oadusBPaXhHTrSyfIwa33zZ6by8f
Oz/mUnQ9+/nz4IQjof0a9YEG23nPPLGAU8Lk4dAOJ0E/alPxxXWTr1R16q/D22iph9ss4sD6PMkw
b4kgIPQioGbS2+ldZvD4f/EZKIK+cFrlQoA3uUVGABHxCd4hvyDAVbmXy0ZYitZi5aR3t1ncYuKl
SlLTltqMxMMAuC6u2131Zoz6xeJChxIlahqr4rdgIW4Ci9HY0+y6kCI0svLF8ioYUfGUm4A+fuh+
Vyh6T3z6JG4hlFi/w84xHz65T16enyXm0idJ4wOxEcvEcIyC07vcLb7dXvzH+HXEoVfrfp1i6q/S
rBedOQpxXUPPpHqPq0PgEBlqIl85ZdAMiagbdBxPg+WMkXUyvwOE2yVtZYLyaSvwij5cRbvjWQZU
S5snTw8BVaIwBVKhZyUHcO5U3AoIg560QqYXwncwR1B2dIjGvUwxf+kJLI3VdXKIMYsQA6Fli8RN
QxRQfJaWPWpAvRTU2M/gwLaHPAOGkvWXTw6YvPQOp4VM/RivRllUOLAKSN9Mlhs+5PEoKj2rOX1O
xaTL03RFkQ3ZJ0XLhDK+CdQiXXiGMT7TG6DLKz1wdHbg50leVrZruE6N7Yh4l/s/j0QGi7YL9q8v
ejWTU97nLX7QYz4gkeFSvjkwl4PYRNo5WMoP/H892bJH4LL4V8EoKP7fAgksnWmZsxxx+cANjBuD
J+lNOBFoLqzDfXWE3xgFST0vCyv2BI/IsxwhFIGyJTo+X1Ku3aJh56URL/QgFLUItyC7mvDjbbNJ
ILrgPShkOipJC6LlTK5WTBW+odqgVnSGa60VmiwNRybqMEn3vqa5+8aNO+3k+zRDoIwuPmrG1JKr
g/yxeCuW8s8XrwZIU2xNUIDSZJUVqjlkbRBpF3hUR3L0hEwwcGm506kJztKIrzfK9BhPBAKEZlU9
W0odhpM4bEA/RPW12w/F9EHjLt/928QBooqCWjeYjuuP8A9VQEGO/iCflsHVtK8a4WAdopQmjixu
oD2+K2Mr85WxU8NAnG4sTwWX2dLacNpi06ZgOY1VnSvoCwiTPdjzc42ODKkqltM5foy/PHefFnYO
q6qxkQfhe0jsYnMR55ZaqanEMNMUpbanTQG6IYHstsjoWHlFJK9W1ca8PgqfMMoyukt8nBMcincL
aECeGhSriMbqLjADDbnqOVs5DLha+hxrAXTPh4Z1ktfgI1BNibdV2FQX11duCCH1BvBKNfbrCcY9
r4qyLVZoXnyyKBZqTMi+9499k/oXIn/m2jklO1F09YgNft0H5ksDBczTIwzQiW8vLn5sVnIbKF6n
AFY2kk7T71Ruz0yg9CJcROGjxBA8stoiyW9vGVMh+zvLPfbddvC0VLS+gIgWbiDH1WS67G+KuTG9
de8VIoMEYSx3405d/fsuNEbFA6rxKfls59rMLwTilL2CM44ihmk79DB4EANzBka9Pf5v+DsdqWmz
/bS6q5QZvet5mpgvrbD4xQMeQV1QoNkgJIHcGPkGauknUl6XPLB780glxpw4iRTWXIAmirwIA7zF
sbEUnAN0fdQU7l2Su3rAatuh+rXu+mvILOmlO8d4Dmq22DLn/rVwi+hiG6oUr+2AwnnFulWUiMb4
mB0Ro8PTA73uVlBAYJLH/NJIcmXpngDS8IIC1rYO8/BTayUeWLhAB7Z+VoKu8O98i8PlkGDhaRSt
8894XwMLxl3nj+ynW7PzT4+FNqNEZVgSIlmsrX5dEKRnrMIZuMcdyvLVF+xukbg83g5+FtNrlWMT
3mM6L22DjvI/z6aspVtKu+Do3wU3TWYvayuMAKxzlAih9oZn3/h6ZFNib8sPby1MX6mPLVjLHBTE
9bskWvLYHTEzoOj1FugD9bNZF0S3CXK1fzINSGd3eXyiUopFtpIsa5i+INAS9SVxXTw+JsVxrvAO
izKm8Cf+zs3N12wfv30e38slGrF0PJtHpe+u/paUJIWDjC+ni/A7EkilifYWtZfdZBObiQwKht97
T4LIT86Dz57PSisq98ziq9DHxsdakw4HPUwrGlAtvZ6QeNtICoxQ30zkJ5WNR5hKnB5jrBb1R8uP
/fwMezWp1sYeycBUw5iEivg+W8TIf4AwmdW9j/rgPyd9rHq2jH8t3BWtY4aXw78YVoF2Dczzu5Xr
nrQt/f010K/p1HElMe2E8/FEL//GvyHp69tnlPlloLRp+j4mGv0HH0KLFG2ztvWJgKSywPACBmQE
xC2zEGkX2aenEEAnsa09JSTkiEwEcextMzAzFQ0qsTo3ZN6h+Hy4kHESgX7zRI1Wjji8FEv7dhGz
WQCNYqupATMilcIDD3SEUzB8gpvVtS9lBhphqSedMEVuWtnh34JQYMMV/ZHURyM2ZOYrNq7p5MCy
EtUN0KzrkLHtfLkxEDz4n+L9vtRKtl0LWfNipJ6qF7iF2hlB/aZhdyKbyBE+6nRZI7VoI8NIMfLM
3fOvFxfx9aX4DIlaiUyzf2npj0iWOzDD3tox+8HVTyiE/iBnifaHoBTZRv3X+vOCR3/Yo36uz2df
nejYW5I1xkvkEDM7RkBGCy5ZiBphAs2XG3nL3DN0IHckCvLOAHBvAEWz/Hr6Texk1HVmcJkUPLjY
8bBuOIXN/tXV3wslEFRxAw5mhLqo2BBmrOqnNNpIpoGUEa+xiw1R7bmgAMPCdYSXGbmx5Hx5TG1K
WlWwsC4ags+6ixy+6VEmBgAeccVu79TKgRGVSzeX+X8foH5V0IEQqWnOZkjgoSzwK6NVcZBiwcTS
NtiNTZXjmeGLJVfF/dU0NS7Kve8xTt/BDMqbd3+kvlgRSQEsZBITKrs9YuS7aWXF29uCbsjMmcPL
6cL1ffVr7bbhlByNktEVaU2ShQ07RJYH+35QI2uOeYR/JE/2jXqbw3eMLhTToYQjr/aNPr5PB9Z1
T8xz568IF/mnptSEDm3EsYcOTJamcJ9bsugNYcEpcy+KPdbz3FOct+egCRuZ96qbE1of7eSf6qx9
bB79ALGUAJh/oDqzno2fNJ/Bz00VErhshegst+HAVhe0BEvC0LWyzfKdLoCHhyhGvFQOYqbe0j2F
Fd8p6CjZ2265dXOEYsohtnIOCB68p1GLEHS1p+5b28awdcmzRwD53695O3BLtK0bMDb+AC/7hxeK
LHR++CmwtrednCYx030dZAEXIhKnV/vesvCKVcStT8NoZ2HdtOly5wn5GjErlhj2pEm7WXC1RQjN
O2gDa3Nz3wLZPnvAtrMenIEizZSKyz0njrkg5z/LvQy+x8ccXlBqkWdVN0eHhuFRpjXbNJrorIlg
lOuHWx/06Y8oezBqF6dY07fZIxypMARxc5rjID/XfBJbL0ZMsirojpdWgLT6luXVSsFNxdtUdi2N
KKEYxwBIjIye8FqJ0iCfdYNQiH0wkLHfV+NQkHZC0YP8chHRJPwA0zgR1S1TsxidAhL144cOeYyI
a9ix8llG1jsYcIIIupufzGxD0EGA1s0p6+EDtnJwa1MqIxRcYsDoB4xx5IjmJ50Cb/XSWcLYn4Mh
6IYM8fGO5i4ll6SzMLwKfSCpfQ+5cvLdrz+xpWNdlfODVQyBhe7NHoXIde2M+S9iscAwBNoOii0G
FsVgY3l+n8QM4mf3LMHADqOExZMQ6C5y7PTsyOa9Cfv5JGCloavLdYEfwsRFyrWGV9rszf0FR+TH
DEim5YaLRtBX/q+9hZniuqvWRbsqJ/mLtCjxGDLDqmLNao5m6+aMkh2mqzPNsP/kbuWm12/GB2wx
WcXDN6TlCMWagDCtKIp8mmrvuDBKzCRT6RYjDzrFiDdZWnU4ztTsFAqBVmYWHHFzKN4G2cjS3953
ztxDT76przVXrxaXULsZbFYEGb2/0jECgE8NnIWNeWyFjSdIm+5syYvbCho9DGtaqS6tJMNHb5lz
qJo67q92P3mbsm9OvNB+nC4jrvc7mx9zfmh8q95g4HS2Vroyj/6ho3XbXzvlRh4yzZ2YFRjv0RgC
INkd3aa8yS6qIahvBpmDJFr/DtVAbG5KRuZUSaE1VpXJUFqCt/r25lzabo9eQTFf0WJhu++YtTHc
P4XOqU8n0Krmt6yxq/vKQohOaVQfP1ZwphiSzHu7JWN9BWCjO33HKRxGnp8t+fFmjLiThAfOU0xb
jjBp+RcT0JKo8jyoAZsXE/oGWRsaH5v0ZoHdMCDH6TtBwyhHI+S4U49xL+vb1MKivubEea3SKDiu
d6XjQomCHMw7Fh6rJTYWlzuVUYhojqD64cw7/gAsKkfvIY0PImPaPZpvJioJe577c5bzStjCCxFM
KRHjNy2oqfi2MAB9fLaQiuZXmAuomjuodWYb4OpeRPqBrpcQY6WoZFyV297iVZO3U6lSUYCiVTI+
5qSPM16e/FcQVPsudEtID8LkXbigiV0h/xb+c1snOCO3lVceK3tT9OQy7YMwrf+s77/AvUs17zXO
14rbt3XAoLteGa9wcwkYTLNdX++6bLvbFR9/5nq5KmzM9pWGlq/QBWX0ilmCo8dmCL7Sv+X3XGh5
r81KppIaF/HpZfhjnzARHMUlSMF6BCTvh2H5W9zmiyPAxJfEJaE8zbTfVrwGYXFbfyl3FQ5hrsDD
mAYJ7ayubgXUG2EUEqq636ZrB/zoreY2q9u7dRsNaVc7iJ6lEEFJBpvgkLXeqAA7xJ6sCg2KiefJ
b4LVROmpeJU5jQPkrQQLF7RLUtJsrUqQrV06pExVBc928x5LS45AT5rfuSSvGEXTDaHYBw3V1cum
BVmNS+87APPgb5YiUOaNdFF8oUl+rV0Nnxv1PRH5MDiOpxW5bfbFmGWrGVljVpX2WUoC3yMq/w/Y
1+msFUQUDSUSY582lkveW40G+65L9SY2KwPgVEQ9WegOJXXXBt21tqiX4aL5u6l1o8VJN16wI2ic
+qtwwaBY3a3eoB9bIUDXRPfs5TELchyPxVJIbk8Z2KNnVvrksL33OHbcaiUwAs1YC4gfzqaktREJ
MDqrLf3oVbWcM5mZohpVB/owvzfrQj/sczE8ArHM10U4loOs6rfljRMlb+O/21sex7/p0ynbmmVd
ya5SL52+kbmLBELNHh7ESRtETRudTbmfNOCON1y4FBMmPvYFfv6SndqLmGPGVMHGDGn/cMlUpmn4
Zcb4roWlTK4cUPvE8r3DYR12L+7IFJSyFe98YUNmGQX4b27UWQ87F3bQ/c1m1JlvmbWrme6DBdPJ
R12F8rfvmTnLLtQp7urcJ+eKtgyaVnM8TVv3xg6mK3mxq6lwYNVSd/54JSYTr+438ZVTOCS5m4Yv
XpHxgBUqr26yd4NnhjwrNfnwwcPnlkQxONxqDJrIUSzM7xUcFamYUG8m/B4mtMcXsBdUm3DFNMMi
Zqq4H2YvmriMPnpTg3tQvKzstHLf+q5s0FqOl0Lf7jhP2g3rKGZB1YC6dmbcuujgpvUwOijYRumD
b//1GIQeB6Chd+LNs8q3SS8ZiGIH9XCYB+bFegYBbI56YiSBz1UFDhM0SXqhZNj1+O9xOW1o/CZQ
FjspSozld4d7O/08WUfkjcoH9+aREd1eRyK0ZyuMrIZWGPDUraw8zNhY+JleEqwnvfdktBSaIXJ0
AbE44/iKcQxlqph2d0r8LVIL5cOCqT9IakJyJ9GGAq3bcrGQzXfPI39NMzVxynRzRglQFSkq2wru
tCVBbMesTkRWgaLqN/veX9Uqr7DyufasRiji8b3qirna5TOXjy3dsEmNO1ffK/dOWbUYgqRg8q/+
ebbZXONmSh6h2VRWNW0uJwVgY6ueQ7lm9hxIaeaevABnr9uLNyw6C3MnAzoFPNfbiX37DymK6g4U
vUfFgkKH+6MZ/b40unX9O6XKMs6NzIGOrkqHrblEdkfpihcsWR4CiaNdpK8lu/oyoo2xlFVmIqL1
3DDFjFN9qzOnma+DHSF3b8Sihs4NRpRTnIKXTMQa0jyq1tF+PJTSaK7ZSCgw+tQ88GIj3bTroIkP
da60Wfpaa4l6Ceq9fLyrD9qU3RXZEzRy9bSARQ8BkTN5s6csvzbcPAqH5GEQ5W49vXto2ImmzI3h
XSM0bDWMl3+b7kI+4DpQ8dF/NFk4b58Itkc6YHr4GbSTVA2NTiTvAECpmhfDnVk4rFZprQZFsQIs
9BBKshkZ2hN7Rb6i/3L6u/JmafTpDwPljICOLAqK61eBa5txzbJP3mYcl38fiD2u/uPhqvERpw0a
byGYxdAmj5OssQ745wOJyXhxxST0OXLz8H5T6s9RrTBlYs3BRPtynvvpdIBibwg7sPK0tUxEsZcP
jfx+4TqlC9F3XcqyIP3k9oAai6EbOgOnsDXzapbibyK3rzIyvBmkba1mhAP8Ps/2capNRcg9rRgw
QWofhLA76fmGY00KWVei0N+jL7T4r/K35Rmru8FHoqpYd8kWnQTTonqTRh/jNL6zyfIW1bkK3JXY
jp/UW0osBk9CQQunerlPIKt2LTKH45UAi7UcHSlyZw8qrR84sEUhySlqshVZrBCv9atDC8z0AS+k
Ufr2I9W69PSUE3O732szlHiTUuvwszR5gsvNqBVjIwOKxoakELMJPqoGo1gx3zcY99B8z+Iysu86
feIvtqPQjAZmtBPrIkL8B+RKEfJOUqbJyb8LVkLfYBl7tO2ZIZYvRfhMBI39cGZ+XmuTxgkLVbPG
hutSQZeiG4GMAc/nYHroB6WLkoPwPLLGBMPRWuKX6VDPuCCPyNCC7V1w7vMQS3YMqXYk+so+oECN
Zv27s8qKAurD7bK/19zTeD/O3o8bHN4kTsas5k83Y1i4RfMljqtCj5c8IsOIlvmD9H3WnofGEA/R
1HQt6CsKRstlW/lwBhgSXPGZX4cb5Uc6Mz345SpyAHefdqnnhz5VWJFH9TKKY+j/WQ///i0vhSCm
JkEvE1OBeIAAPpRE/4+CBpl3j1T/+pgLqvuiDGcizJbcBe/GL5lMKVsAGqxbyj5061CoE8WenhVo
9CB2mx8FDkEZXu69A/fqS7dqwcm+zqNX4pHwowlG23XBowNL4E7jXxuoyMz3sjP8HiSKW3lDETBv
ZvrE5gzhPdktM3kfWeV4zf3vVPb/nvdBBpKplKQqkcdPaVGe7qanYy5CZhurfKCcw0St7gGtTZGm
zB4NL1WB9UWfIl0FjwR8xH9T5OiHsZ8OZfjB2YOwS9ErmR/nV8ZIzrltQCXkG58PSCaP4CsG582h
/SD8NL58kxpR4FYE0IO5zfQ3dDtNGMzx4y1ylXex3yeiXolxAvff27O+Y9JC+NIsswcI7Jcbk1eU
b+owrlEdwiRAQCPiyQ8Jg4INyZPa0EpOiU6jKNx2VYjqZAy/KZoAtsUgtJVQVpElh6BKzpn0zR8Z
xanuii7aXVvSAgvFaHR7fCavUwGbUU/RffP+ncmMJMjE6CXxAYJwsYRySqDKdww6e/+OPUbqGVBf
7CNi5J9xYFtWXKEKmCBvaPngHreY6YsewjMshw+BeVkKG0AsVYjsoz+7/ODtGMZVWTkOvsP6lhKU
3eGcjhx24K3TqW24H3HlIkH5asy/0GhGWOq/DjdgCScs0csTcxBGt2+F2ToCsj97dTdvlKKMzopD
YvIhbaH7ASqtdT4WrP2O5bBSLoEY4JRODaK7NmxhUdExIuGl3uNOssgR0CQFVQDHX4OZMFYYZNM8
c6GpShN1yMJNCCGHxX13C36cA8W6e4BsHJmM17Y9243x43tdDMEXXp5+hAiJNavcIYLaYjONZrwF
KQtUvhGJoT3EvUlYyT9zVMgS8ZmcYAVK0ry4QL9rgTWtLY3wxQgiv1zNSoUN08TFzDpBJjCBTPqP
dafwr+t0XHPFROSZHnFhN130iN0XLg9+5oRMcQRGnAw5iI/4Mw36pxgz7aDSy+t9n4MG13CIOQQV
B4dHGNJO3CzR63SrnFUzJEucwHF38NxtwEklTUH9nAdIRpgr5Hw384ohztZ9rJCRlx0iNsIKzybi
vI8aU4IMAEGUgXwtWB6hIcjtaR+H1ucAoydS745SrluWHNU5ONiSz/6EZPkEgCClmHnu/QKER/u/
mjVxnEitYph20fM3hLhheszW8zxy9HuVx2eHJFjTaeN8dDV8NskuaXviTBHao/ZyZuqJHDVqm79I
uJqRfoUYAu1gCwNs5uW5wRC5Rrhom6gOxGqMFAa2V9HNl7s+dqEaY9nNN/WHjGRMfXnEb8C2K6Pq
+ai6m+nL6mSE6WUwXr7Z7bKQYheey89hY2y1rz5HV/dRkyvlm6fr5KHiORIMf6NM/aP1p7n25HSD
AQBnBr3Wr4nIemrI/rXX3WUlNWioepcYKzi/EVJKWCcrW6vW8GRARNU4yb7ODTnb9x3C+HBK66QY
6sU2iytn5J8gEmu1JTu4XijiUgsQl45zuStQNzV9DTS0ICh7GmYvPDXAkBvglwftAp/8bGjwbf5w
g1Y1fq+jOxkUxmHMB/G2SiS5mWCVwguEEwkLn/WeFOsBXxdas+DGe61ZEuliAQeuc3sXq0LvWEnp
iAKMWu8HFVJE2E8sVKqAIrg8GWzktSoDMMvgIbH37UKEckMJiqCgRsa7Ko8uyZRHtNRNzujt7WTV
43BEJJRMkba6lobBGG3jLGn/DnF0137gXItAM6T1jpcOv7zuWVVjbTTOVkUk/u7hyrkqXDCIMMm6
FuyMFTShhSHKAoN/XbhDmCFT03ct49YX5LsUNx1HRec8xwc7u1U+xOlQii4BOwZOVxRA4z1Dfqei
At1KRk/9csVI3Assk6Y4pAHTGinhPIqa/xofTt6ohHBYfLjECOcIjUQSSLqPMlCA2aUj9VOMf7bz
CxUg9AWfVv5s4FyB2nneGvMZdDFcl3B/ENFwl0jJ50AjprPY86b7ItPVPvOJN6YOurozGu8EasP7
PnjAbr7vceBw2ADCVJRx3WTzUn7Hobyg+/H3ySZpTJrTZlt3IlBDnNAVZ1HCWh3QKP4wnZLgrEoi
VE/+jINz687kOiQ+QnwHezE7NfHblWSTzDW//BwSbwQC053/C6q7KLaPFvRCM1fAOwyPbqeK4boq
eT9kt+arE/j6bLVIqNuzxMnKrNcMKyVANhrya/3+rKWCTPz2K5RbZn5Wl11O4B5SjaXHtcIze6PA
fLsFJwhQr8Up37Bsek+bXMBvE152ANt6ZZ2rtd632Z0Kcziggho/b0dpYO3spWblrlzSHU3eBfnz
8+RiK+WtzU8QvY5EzRXsdR00qUB8tJwB3QcXRA8q7Pt/DnAuRn+HzUZm150KLTymraYlbvDRdA8L
JcOD3Q+MK15EZdowxQB68rJ+bppyvDpjm2157zHbtAPtPBU8tgR9A9EzIGyjNPHv4gsil+TfwGfL
yr5eL1+CZIbFEZOtW2v/7EfEJD4vyAKtZkB8+jcBoE2ad6pOG4Iw8bFZMec06CAGl2cJ1qN5lFPT
blAEN9iUhiJ0Lp3DsCny8BFcnH7qtahpNqgCbGyFxA0Vonp547j+MtCnMQoK6Hl9LWUmT7EHcE4R
zLe1zkmnp0aGwsq/VFxULOxEc5wwCAQHzA/YRxO4kg84PzPpJcgkNvoREJQcR1Av2Gt6cyicxCRU
s/ym8NzuewCC290KV12nS0QDfur7cYFwXOV6nQjVbc6bXFS98W+LmRodbn0k42Aa3uWE9AByyHMD
kNU0LTBa2L07DnmVivtrbuxdqRRqD2/1WctCyta1AltoyW3dColOxhY/qtvMjq504CyGNEVmjQwx
JRjh07hvubcFNAJ87yRfRWxjM9bMyFJx2aBkhrKKnkxLT9WBaozpN4RtTIJiSAr3xZBoQtAXEcoM
hhN/bdNt9f8Mokkb2RhUrfxORgyigZbEZoRUEMGGm/xxut1rsINx/OMXsBIG3lvo0EY4pMG1lXhY
g+bQ7wEJf2vI94Wo6iHpJLcSZfVaq3qomPLGNj96QXi+So+Os33k/1EVOa9J52FLKbd0frr7L/10
ZExCBeR1fYeYztqFv6kKDPNGkPRwygMg16DMdoEdaffQDiQXYtxy8SSFlUxf3oWYQrXQPJRXSVk4
8fSjaEa60GgN+tW2p5TAZB3om63Vy8fDkvJMQNj6DEQEzEA+v/egDhSj8TrqpN2ATTZew0dDGXGD
L+R0TXee/PpVb6N97coE3irRd3o9J2qAem2ewEtjUcUppSXQsasF0V6gRftRy41dnH0VjYMNhCqe
EdZ82n3ddRbJR+VE1D56qmd8zWuIoUkgLBOx0R8Qjx/vTJNCMr9XmUq9j6pMZt7b0+9rZVLdnMhx
71mGNXVYnYDfgHUcI3bZza8xIzl6Zdu9+0CbEBOB9WITVKTvsf68kIWuuVMNQQD4Mh0HaC9IAcQ5
8qNPCqmhI3sZcIzB6N3epQ1HeUxqkz0GzE/ohNJ6apzQaVYvKrpw0Rt/1a1l66+9ZfnnYRhaKgsJ
mGi1Q1trLjs/w0JYUeEhokhl6lqjjbyev63MAdWKuTGfK0piXiIxPjoMQM1QgMaNwwvhbC4PMYaf
rr6Ozf+ZmHjNGmlYZ1FzGr3yK54RMWXGu34MUWbcH+eFeyC5vMlOEX92fJhLQANaIQb8HxT4Azcz
QHQiTPj3r9pd0Y0kPUZPBmzIyFyWctu9Ffi8C768TySbY0zsfJNdAYt56aFGDAVXC58P84GdJt62
W/+3XTpIINHy20NJAJe1Q/gjPya+rOFDJRsg+QZTR6uKg0Hi0wSsMcOCLo97B66smUvZiA9JST/a
RCG8x/kgtXOyKyE3IzxmvXozobGExETkUU6Ya550XPYpe5W6EuYaKfpeCCTN8nT7jHPfVUEH6m82
aeHtSozgOXB+R9HB4HiTMIKFOAMEkXwmi24X+k0wj4p+hT4EiA/0E5hR0GEfxjhF9FHnMx8HNIQf
fVGI480E1YP12WKfUyCioep5me/7k6jyjw2Q5V82affrU0nxbl1Z9OA6ZJ5J6YgVIWD8Hl4qCxsb
SnPMk+2usysr7fE59bUPZoMb4f0BmGhai3vLloDCZEksUu5WCj/RqLsVcnmCVJGEIsuYd547C+HX
+a7o4+jAF9OWRlsZzeR6KLrOn0sZgkWJtfIO/RJNRHXpU1Tz/vEEL+H96XecVLGR9GHkCXd+cnE+
+7pbe5k/t2oGFJz4C3Sz+EZktcr5F2L7PIJvvDs1xjEdejz9lCK6qTzdOSoflEn4MKa786tIATYU
TUbrKy3kuekxYVlYl1ImyCJOEnV6K42mNP0K3ctTc4hlLmjf+VlZ0uAAuytTWw8JApA31M6h1EnN
/j74Xs4RsM/NtfBKX5DCwJ6Y6J1sva7Dp6oLxua3/soFtSoKGCLGeYrIiKDltSBCVMbCFZr5W7KO
r1SFPxO1psfOHER/hm6NniJf5Ll8lTVJXIXKPIrsvaZbol3G7G2CsiHO/rwgycOKeHSjozt9S9bs
3/453AwTYTjP19msz6IselLLXjZ82c8gwnEgIbaEuZME/R9eLuXz1NoQfOlRr52o4UONfrpMSv74
GuUdbvxa0kH9fjmbnD0P8zjCz4VheByiqf2MWBcoUphRXeqK/pyF7xsgSh8RotzhuQkBsUtKazGu
25URvwHBtasRY/31bxSFmOz5JmOzC3GhMiWmpuOn0MO2ALjrKNPfHKnhwTY3TSI/Ae70WAZ7Sisa
H77wnGwmpBhxTklwVohjaDDRbY3HK05YDw+cqbdi3mpY8rBt6szc0ZbaCcPhOdiGUOcgABi/bLHt
Q00RGanNHcqWnPuZhEzNTSCfMeFTRi1uwafSgh0CB5/bVWLfoSI7nKSVRSfAsZLuf0XdvtgQyGmv
3yS/7IZm3DAoFv5D+kXGPtkLmNDWO3f1JDQn2FbSNvBHN99icqMlOrVoPItUvAW54nfVgaYg2Gsd
kOK4AYphw+MF0HxyrqUdoPDzRaviTPEalYwt0aH9ECUNPkWgZahjwMe4dDcyqstOJ3T55E85U0Gs
mc2wz6MYnf7RyCjj2t4gMrbufCoeUgo9taL1T1rEarSPzclL/05i+z1rcr6BqJZCf0O9+ydKAoe9
lSHGPQ//Ac1FA3K3/i1XF5J0cQjZNbtN6nwVJ3oHuLL5n7anqeS/iEThbhFllnUBT2D2F7T3RsTw
N4yJSWctZNuAmoHjz6AuKwiO7GpQgdM1cr+pix+P06Ujm/fOmEgzwFLPyZjhC/ddWqv3V9++WQW/
2WDrpAV/G6Y/gBlhzmh4LjpJGK9WGOKba4kA7KsxysS7xwQMnM1szxdxQ1U9EnJhy6ErAzQRFlRx
xKBCl5j/hCnhVg77BCfgy6Ypyvpz0Ddqn8oEL6PW+LdMKoRxDd55xrOMmMscZFJqIMuy8rSJXAU/
MvuXhoCA45yBqvZJ4rqzol0qxTHVNGHuzdahCJEQwdQvstcKgfp98siuYh6YsrhRxhCmAFjtW9Kv
v+Znlcg+YJPW46Hq1lNJVv7UVsOFcLlH/y6KwTD+oUQA3HoFexpS1M0n0T4Uaw3rvio3XESM38OI
sW3Tn49d7RV+/W0ArLw7j/1CuvKD0S5BGB3XjUA/kqx4OYJezldJzZ68fXN497QthCoeNmr7b/pE
3yyRsgXiiVCeR+HsPjDqLN4fteuU5wFnWPXv5v42qVMwkZUI6jl1qF9vQAQLwM8O+bmbVrWBU5on
/6uaTO3bsyfsOp8wvctieLr8ZSRfUEHmxKl05iSN6M2z3NdlMBYWdZwS++kz4/h39Shrh8AdEn6k
LItXqTSVWlBCwvp/HLVjyR4M8lNX3yvRCzx9Jn4xDIYO8eHkWmZx1ejl9+S/lBWFSQLt4EAZOeHP
ZOXMI3Wlr1w202kYQNOv08t3+Gyh/YY9xz2Szytnkt3+Bw+39PnkRgB1mhv5kZBlLPEQQ8l9gPuD
7S+FUq/HkCODUmUO1TNvB3HhsfprYyrruSOl1CTgc6vAe0iYQC/1PmCQwmqGEictJO/QuzeS8sQW
/WeQ9j08ndaf20UO1rmDFzWIvL5sMRstr7t3FhBzJrNuNbQD9XlrvbdA657fmpiZ/L8iBXozv6gK
GGXe76+lY1LeYDgrnUxaE6Q+z5XVN62taZGkhDrivVHWfQk90EC7Du2QFUamLD7Kk8aOfz4atm3W
2U+X475ltx80LhZs5HP0M0s/hgjqO4hMoAnPkBxfRmHGWdp4lOirT69VDgR30TWrQ7bhTSl3uZ14
1qsWv0NIYyT8AxQdcGBT7mXjOX7pOlO7hlBx8U/8Z4ByHONQ6LCeodkP37tI9mKMA7wUtQpAK+39
ybPCxc/gUcS/OZs5gPCVHLGleG11iEcdr2uJlgwBOxcz84cDzOYNWBmOzwWFB4xLfiWb7FsJCWXU
kDZ/If9vz48owCxO4ZAR1LVzJrjVU3OXjZZzG5WOfXvdcuTt1rMQyadj3p1pzWn4+PGZ1mR46a2Q
b+KOcLPwFnrHf7tl4DAjVamr+ByZcjCdT8RhHwUrzv7Vbrt45cwxFPR2k0yZtzIh4AkqBYJUq+m4
/FlrRUAMg2H2MbbRwvkhg29clvyHHyqI0R4kHnYnAFdbfP8bAcl4SPnwZobBP2zuAIqn4axMQoJ9
mXExD0jA/LLOdXg6FiYiNCdrVEdgl331PXXbFSw/6xmxoyQZxk00fSyl4Zo9E3KUecEBqGWt7/od
CGYkoB1Ga/onID55X7JW6862/HxUovnZcnZFvEhc9Qkj1S9hrMFNYJExOIQlS7dN98mXaeyi/pTz
EZdk9WqJEcuVezv+Y1aKlMnuX6UbgpmMN67hYF4U2LrBJD7Phe3nmLaLlmr+sD3Y4MU4gWTbJFTb
dUKQTT/g0DHFBJGxZ/AWM3GPCb0+sLa/ofbtlCQNmPFFAlDE2WI+Zz72N2YC3LKSy4OXlfNszKHF
3PHAGy2w1Az6MzPbWalFhkMgUv/RuYl/ChiniRm+h/A/BqU04JGl2eG8sL3vkhFqFvPSti6ELToo
QFbLbdescr25F9MkDU2EiKn5yN8UoeAm6Ucqm8dJ7q57w0H1+n+FY6wVzLVdHB/ZK+icRLZKnDP0
8LeRqNoMcLEPn62EuMgY9SB5SBBg7wZV1qknLcnuffECqc2fv8k6Ur1b9X+aXPXkWVU5BI7cSrm6
DIKvTlorsxMx/oTva3NinHjPE2aO5t2B6ntGoYkQLgIoxYXFJiiK9Bcjb7AM4IYju4TA2zXYihYE
8gnJas3Hq2Oz9E/qC991i0gvKmJ3Uz6soNV84Lokh8JA9iTbEjJb+43Zr2iig7k4YtNLqwL0OEyL
7abEsyUrVXTBmn9AZ9lY4EvdAnC+FMmLS2OgWEVi8FG/7grJFbaq2mtZhRm0n0khOGqdUVVJShil
wSIz0YJ2oYJHBHjrHtFxNYVT2wHzgbqcbAb5OZAshIZ/mErRukBmc8P4jfCeKKYgJf+qDT200JkZ
sxpAh/tXKEFufcwSsftDxUe+qTZxhwnLP4mwDnGkiwghBG8LBYF7+KWwxNQEzqD3gJN1l6m1kzlY
eGPpjh3wBUtYvc7xSiqUEjwymOyVA//hkaRtqkwGpa/x+DtYVe7dqJnOLNBTyxFneWbL3PSQDnVh
Y3qrSRMH0IAXKvyi+mQ9pOp5fY0witUsW9QYfWLOjOFO3gFrDgZe5tiSSFuYtEvG3+N+P7bjDPXF
0qqkSaEEe46EKG1CgP9VsQgxW4kg77QVJIBjhx2O/MMiv1k4m3gclHee+BUXMoOVVe6DKqxNOncr
n/IsXPVnFKAXosLLYAgBUHSKrKTfaPMbYoNsMCuzLH7NIe3AdS3QjWvKiiZJz1E28K475S03pQHD
7LaQJeyH3YQkqAL+lhe8zcDgtdnLde60qtz4t3j/QQLLfWQMPZHf/SWNiPMS+IAbZ3nKALkI/VdJ
G6ptjlrAOJpUBUql/OA/hgu3XF+KzlNRRYtDrHzm20PJbGoTNDo5d1DnGFg0RlkU7jDkuYhb4f1t
gpU66EdAJmdGfWoAoBPATne61PAETyPhg0S505Cz+8dCjZkoESK4iAPqVEkOd1aF8k1GUDoBE4Q0
PyEwdeHv//+lcjWiujLqVTKgBzD3zD81dV/f3VpYY02lWUwJg47a4+bePtucy/uS/PIvveLqawSl
g1YExjWUvVhBnFjkmekS9smFFZOrjSBluEhneC/oYsx99jdRSAxJmu7Dq8Qa3rX7DaNVaDdGYNXZ
hWtn57Q+bf/M074noa9mYExOmyMBZPeiiFk3MU+NbDajTx9VtjnXJ1lG0DfdQO7xrHZI1ny/JyK0
7UhxmzYzpvPhaqX4NGZN5Oft97GLE8UASNLVCO93fSDreQ4DaobilwlOtccUG266Q3wlHLRvKk0F
YFQbFWfJqRGXbSLeYHLs2WwWXglgIi07esGZIhn6SXYltHC2elnWvOC9kgr9oIDSgkQkGpLUiuqd
tYxqxx9gY6bR3O9o/UWa0M+pBb073VXlY9Zuk7qFLDICS9IF2td5ByqL0WC1ND2GqDGso4z0i8M9
ySPCUJOkswq5SIcf572/DApyaJ8jlmhqwfApJFPDh+9ehdXmKqEqlze+6SoRlM/3PDHLufA+NURD
3o0bx/+KR1iQtZIttEiWYrwP0DtqAP3B1z3tHzjsDkqaikK98w+bL1dd4cNa9g6N/lhb9t+drxG/
OmwVfZ3ioZSC/QkJROrULQKCnQYH6ZG2nuUI2G4wjcMRMImPpbp1qcALOB/qVstBKt4hgRH0AyL3
lRyooKdBIV+n5i9VJifh/yUv0BovwZ9ucRcywkuP4wYKsCVxgIJ7A484r/pvqccaV5y+T2kwjWLw
AcLzTpkZYx5DqNSmRC9L1Yobl+E28QhWXbOQZ7+KvqK4BedYRlodMSC+0wR/IhDh8kWUFmdFO4zI
lPXsf1RoIzOxnsL8A0ncwD/UB83clDl+dyPMX2U3ndn060tk4arRQPwu+av8xclJ2AOtjTL57nsk
9q8Rn7O0zImjuZnf0r8Q2+rZEEjGiHF3ByI2DN/qAEiYekGl3chGi7fckB5W7i/a9aEWNLVsHL+B
8Fx9BGm3w2mRH0nxrAI0HGWovxfqenf/XAGr3JaUH6MX8CZ5tkz2r8NtUM0Thrg/09alhVjwpFm9
6ZTzQCwOk/9yqyliMqha2czSzTCgWwKCchptuWaRNdqfCUAQ+6n13Mh76PdYursTAoROYqYyNuA6
DVvoG2GMAyh0W4JQmOULMWx7kbeoW6LIp5HmUEvAKPDWXSuQ31r+fsQPVKjd9ZMl/ivBAjE+gm/x
Xd5c4cvBedDrx52wiqr174eN0NM+CkYlmEyF5rzDmGxQQtinnV10FoVd6j820syxFGEg97EmDDg2
jZNeBPSxckptZ+bkXxeyApMDZxg7Y66TkzwiJkfXs/gu+yWAhlCRpznKZGTDUcqm1TYuL0aKCjaN
u4oYyJ/upjMWxUX3GaTFdlq58O8eT4vfsAeS688WmBbtoMzZjtCwPk1bkCXUott9+pi45RU0a7XW
DIG50uccH7YuuGes2brCOD9vUEGiFGsigN+hGDgffU0LorS4UqfBmkC+0+THbXzMIjbbnTlUBPEs
eptozpEPZBVu8e1/M9YaSQ0WmNm4rRu/i94qWptf0w8obLWBBnVfhUy40yIqP8bAaXerRAcNXOAm
JR4PyFCQyPEEYfSA3RKsBpbTDb1vcEwgycMPai1dlIc7qcP4oisTOymPd0p5LpQjV0J1Z2zttUD+
qTmBrYRQOevGSiVKf1CgGnqILVApM1Jplxkk7WGskh/ql4KBdDSJn3vGVVPyP4KPpG8FsMY5kobr
9ULVR1lKaa8kN1xIhPg7F2t+qkUV2zeDuG911OAgkvAUEzB8iLqkc7TfNGwA7STuot688asEKUGL
xoP787wtgf2/og+pN+JmjIQRI3Ut7oFElxbohTYffmUyFursO7GwEbGFfKNyDcx1n4Xa4eSU0xUW
x1FBRg2ydyv0WHQyhYCHHhO5V6AWkNwpmx9DTHgqArmtYxgJt7U1OtLnn/hMm0y4+H+fd5BSgJcs
NH8hz/1oSUhI7vdynaplTFPKsj09Fd/iI6G/QB+4w1We/305D/4lJeG/eUlL91O7kS6XLZsPFDoD
y3ztQh3mJC1bNdhXfEHT8F0jnBwVO85VoFERBSLf+1JHbWT2Gd92rx2/7FsBNVXNHQS3T+OT+W3h
uq/uLqukjZxAv6u9FL91OF0GrdNSRPc6v1qV3nGjmmPeBa3N018TuElsmltef+V/SCcO85TGJRnI
NPQMNkKLpwYXGhaSmz298AMn9kM2jcdFYRhOx01+anWgIA9skAfgy6hfGC655/3VluLWspeovk46
IGj7PL25RkrNgpfB3coBhEqgCM2tyzhTYRzXYQLdjIwj9dIhynQbvJAS/aSemZ3XjhGqgLURVEQ3
guEM5O4UZ5zgs2re1W6/ywV2nyHpSf1aanZyDy9t0PkjtcWfbNYSeFiraSJXFsiUj2/h0jVFcILf
S9dzUCDUiyog+cCwIxLGyBE4FpZAu7JwtWNk2HvuI+otqkFRcauV6cE9fLKtQKuGgU0kozRjgL/b
t/l0RKh7m/nRgGnQNatF0hvYFuIq6rZ41JgmhFntVJUDbwgnIk/X+IHX5zP6O++2r39bLyGE/bxe
IdMVg0zhMBNMsMVZantE4p2UNFMUSoTqEitGOQsw2rXjNrsTN10O3752P8tKXp/fCb8sD8OWpZ/R
+mj0YLPQgRCH78dOzYFtFRcWIQvHgIk3ucH3/i3CBpxUMw+6SY12m70UP9ssZuj73j6wzrXlQIrd
mmb5lIoaAcRQii9VsL757LzpNdEkXAat6tITRYm2Qtc1gqiZicIn6Mwo1HIVd5xGFmm0SmJqv4pv
M40bbqHhZr5bqIt9srbcvKs2x1E594nz/0o+RW4aePzCosqY8DVm68nvwHqnDq94gekGwDeBTbfe
rIwxxq+ayR5+3If8/J7rohzXI8zux176679PlkQ+ZE/+ytTItCb3zSXRF30y53puHRHGl8etLU3H
bUAvyeFLxoG4zXq9XbLVXxzmUBy9Z7OgycU6FE3/8tgFTg8sCwSNDOWOCeMUtnpdxeYqG2+Wevrd
C3EnBKU7MvN3ZIATlgXFr/aEzWvTKQc3QistI+x8Il6/NJ0oJzgYAxQJja5wInFGqMvSpRoVZopN
/t4jfN2iI2xg0VdOvZ2KJL8AGlEn/GaeI/pyyLx3wujN8TZeRIk3YZEmj4iIXtvQ1qxD4jy/txx4
mL8b+ilJAU02nZdyg7Lily82CfpQrpQZ2CTJqEpd9RsFJR0iLxrN2FJbXiJk/lnJovVoS6Fyo8VC
D07e6DyKPZD5e8pA07wpaLZzBYgjZRD2Qeff432BPURvIeNU8VOsnGNuuuU09APPtix12HNQJE/J
wYpLrmDom71OX7OHIgAWOCbSl+P/FOqYkuinGRaQaTmnO3F6ukimeqqZFdgSQM5qLOITYr9BYlr6
UmPMfYgCEmJenprpWm/qdTTKLjYoCj/oLLuwda1QRWp/j/Oq4RPlCt+3cJ/vIPi8ZuZtSVXcYlMp
etD3G+/6fwXfuBaK1/0gZKchCbOwXUPG0VZYp3DgN8KnenEBPkm2MmZ0UHuq294G6iJK/gp96F9U
Yz4c8a2CqNEP+GZVv+Y2wlqxIPr5saAH4xYHYv7vGIDtPLx4u9vBkxeGZLpxqfVE5j4hwrLVbOWq
Dl0C9APyLxIi9LiPrIww2BluHySXgFzeSOcDY3rh9icFSVDgk9AaNRA9i9iKppA+fXOgtJncf2IV
eyMSYil3W8emTTHvwk2W3jwbeBU0Y2ztTWUWiVB5uG9P6iIyzY1yTVvNMF7qHvEglaydzbAcdUfs
o+9LOcC4RvIBEiVH4chtIiSJ5cpdVUGUo22Du7eMi6ZiBU2qffSFMWlrSEZo/9oY1fs0uh4fHpCQ
5JNocDMaYLoOH5zTN1JJO/0eBlb2NZJ6T6WgfsA9mQCrQVhqrHck4C8mKlFglNuQH0GyMqC+pzJB
5aHMyUb3wQ3PbM0qUtvZjq1cTqdH7v48/x/y0zVKAXhvZTqM8D3xXDvPja1jni61IW2UcRwld+ug
m454UgwGEEinudpJb/YPi1FKISwSr2c/t9kRmav6vFYWpvNtTr/RR/Kxfro1YP+firr0K8phtLCA
eT7K1z2EQKrhd7a1MKhz2xYx2g8iP8C0X6UluQ617dcRtYK0fC99XTQPL/BBumyN5fTufuQLcwtr
DsCSdR8qI2hqS6eECSW/oAKYBMj3ZWIHZ/5HhF5c4cFlMHSNmoM5/e3f+QpersGwdaxPslcxAmXF
wbdvgj7mNww69VQGBjZwIvtm9pMLW7YdPBCicpJMrds/81koiCY/ePwg/F+KHq0w0HsOgcIXkZgJ
JGIjYL/wjG24YYcAaK0BNVIouDpZs05e1gpRGmZ0JruwrMhhdbJdwnA4ci0k8uxe0QPEkT3Xq/BP
sE13Y8Qj7/NL55uP/L/IULQYz+X47oCihRUEbHdTOi3OxTaNvejmrhX3A39Hb5oWj3ZV7uvxsoVJ
2vjroNq75CxOhQ5CKUfo8a/OOvbjn4apKS/E4LI8drT6a3LOggFBc2/yigbK4BuX+jG5ff2bQzog
yTfoqR/OrpImmEvRfkHWeVqmmsR6/SO/ZV3nNSvOzCLYM0DitVMwgqwKEO6iXec/iGMUI50ADHx3
qlfx0vyN62NzAfxJYVP/aSwsLK7duGsqYB9yYOr7hmoyLTq6gfya9B4VkaiMNFYzyo5KVvC1T7ns
u18VfPBE70LxxoOAQb2sqCZYCDqjcUOuuC+6GjN5O3LHW0SdVpU77WOp8y1NQkvoYGWKP5pX6rVa
5H16P13AT4ZtT6LSO8Wvrr8G1zMmy1tcIR3tUXVRrcAOuRiXItOg1lGgWpnfbhwuljzTR4d03NAJ
65OyyiOYAS6+T59eJBagPVwAG21gt3HHKfgTstp18D5V9c+vFJjRVFVTYgkC70MJSfpKwergVvSa
PDQ9EF2YTBXk7ErXFAqXo5E/+9sWuglIxwoqGqaVyV7mqTZbgOCM9aLw31ZKCFVzn8m5/yDfZbEq
gnKFFOIfNfRzVBVb3EtNTqlDxZbKq8FqQaIzW0lJm9L8/EfvkWowBImxHqtXzZOA+bZfyvQYArVu
WD7Gfz+rII2KuE4kKbbxc9eGZH7H8+H/CsxwNsU08xubUESabkCmcgtFgP1cfqC9O+PGtyWZh+gn
3Ur3FsQYo9fT2HVzTXA+Q5lMXAuagXJ3mcD2c2phD7mv/BL7GFuFTTUG5QUHNxs/Df9O2NGONQWo
7GvxVad/BcJFRFvK1fBFubOJHdCC2BnH6GMIepemxclFgdOM4RQzdn6o+YmOSjrBnCBq2SMmTRJe
Iri/rIkLXZIJ7rcxotoLtIp0TaDH3821TuUC/qSY4+5Z4ij9jiU7/snBJUKJ46pw1ThzdqQqoltW
2+NcmH9+yQBAe5/vUakO9hlS5if3XSicgyA6s2vjgGBLf29ueyweRF/VEDiLALbV2xC33867Flea
s0BAcswA82Lo4ouqfoFACGGvULl1W7+JhpyKLNCV93Fq41HxUlOCpnF2+O/rGNmc+mvg+qs9Ypli
ciiGyKf0/FsuGN0J43vrUPxi/4GEnkBUj3fFWAZDxT3jmaP9EyHoMNTWRCEr8xBu4Fw4XK9Wp16v
z7aWDEjAYld/ziBhnpPgEv82zk64GaAJZHlazvjLLZfrZNi8KgMvsLEsVTya6KRvtKUUr5+e8jmM
to+Mm0LK+wx6kvgnfZTrO/PlvKyYeRqks4XIPfnDdNv/5KcaPOysqx91dRj+yLzslBzpILZQW+3F
ZejoHrk/IP9Lj7+lJJqOsaob0a2exCFEg1l7/3Xx1NO0uIdCpDJMxieevPc8K2kpZwh0JjQ9Y6V/
hHztHi4FImOGOVV3gsWU+L3xZDotDzcsZiLLth8qN0dlwAhFoyxV1rlc2F55E/bKjQwXsDTHAlbC
nj2to2QgAE/N9OQ3wf3vuyf6+l1HV/5qXXQuHUtTqUYp4WCG60T33TsvEaImTyrUU/a1MspyMSut
ntr0UgOgkym0nju6pSSNQL6x3gCo/8oTufDtOHHMk50Q78zyFda9RgHjT4RT7rTLaJWv8X7lO++/
z93/9mceLu+t36mamrlUrcoWXuwrMcF/q2HVabR8kG0t+RkdaOVNWPKCFqtTIRchUnxgpAGsG0On
31p6qB5uPAkAS9eZi0YWC2T/7hM+7OHwCKNh5oGSjAwG5uS1NJFKjmY86B0fkuCM/m/0hQBkZnQT
YtGkrAASDjTYcQYztR+9naNn1whb2oQU4U99uCmvS7K5O90//9EM8Rp8eCskBaKC+V1s9BWtfbl4
xzNbrJjcDl/gUVoDMK8AjHj5pawVgeA85HAMIEH3DBE1nKY2WJrHNnd8xlFabx/jdzvbW9p+Rgbe
bdMNjElFwBMINuQwM/1ANv5hccPjJrMC/tuuXjq/cnxTgvSFZi1MW6GvfxSUX3Wx7KB6Gop24jnI
DKN6PtZGFvXB+dEM9kBOyiz/MQvoTtfEzyHbFozpX5Nun2xtqgc+mIyOzYweMtiHYOMIgekPF2UO
CFdOOxKX4BaW8u+qw6LhkLKeKfqaMSJtKdgSMWbMd++Ijl7jevKoxsg5ThlbVkoLF7qn7z1rLcBd
PEQ9eaw6evrgrDoLZ2Da9X3soYvBV6eQ8P8MiVNnUBdzZ17fSaHOnDMtBcIUvE7ASttdfH2ilDKk
XgDoOYU/me9lITC37J9kcEaEinDlEBQ7Wt++0KNT1YKNCyH+9+cmBuFDF2VOU++isemzSzpghc9n
heMVvP42t/yaGlgz1pvcgdnC9p0NEm65QwgGVbr+1kDSFwMrPiv5+YGQut+HU50CxsYEYMCs+6mh
GWswN24N3j3fNmB95K3uH4P0n12ea2IyxpgHLxzJU+5cCXbJFBzwG9SGLqTRyhKp/7GovwtGYqC5
MzUYKpeN/oGh01vB/7Lsq17QKi3Z48NMpjUcCweQ5136xeGK9b5RnXJQg2qwhIf+CGPbMHV4Rxfk
PNtTQLwLvUp8E5K2+kiq9l3ctQi5BCRwtjlJKTBPsA3zhGUpG3k5XNyrdTWp1VoHBPJfopj+w07J
k++sTDE7G9PTgOLjyDqbPcwU61JytvAsUAiEVQHvXt4wge45R2WMKuGEFWpk5OYlvkWzvpAdLCgS
hNlnd03IK0iiCcmMuSHF6WFExVAWfPCDdCpVHFmM4XKbn9ALr7dkQQ3sjFfCrbPlGePgooPf3Lrh
vbwcTrv3ziOgDZ83K9dQCBLFdc91wNAoPW+sObuv0udqQTzuzlPc7qR6EumvKhAKeM5/r69l/Q7B
SPN9aXvxokyEBur6AhsxWuTeMVLCyyheiOFhZiBudLZwjCZ45rlDxjV/GDconMsmf0417csCtI7a
aV7AJo9FIjk3v5X+fFbF513cD8WMlWzb2P+rwWF1Juiy1Z8wUfYzeY8CGzyUbn9KV6nRvcxSVQGc
2CtlimfTNsBnBuPboYsdEjXXrllV4dEjjX8VfZR/IQ8CsEoOKD5FhkzQgXBqK9edmi/kAH5fHQ4B
JwHONi5wnCyzN7a1Hd4IsmbZZeT0kAB4jsvNMdUchbNaE1D+dxoNMKwMPefNMl69CRoE0BaLO2OL
P+YnpRUwZ1ga7ZNTw7PCREp+VFLRTRUocq0F2J7TOtX2uabCemo46kKRjUUAmKFtXB3u8Wi74AQD
imReRcTSbzTP22nPtebRKmqIpp7rNWU6cszYTiZf+dcbvACu4yS99Le61PTEXejA2ooWqnP1PzvA
ceV9mNVkNc8pcHEV09hH5AMJaweaN4pSXi4GX/rtLZwkMN9lAZLAR2NGWjqD71IX0PLYLMq9cbrO
GH55nWpVToeyhUGlFj7Z/6Bvvq4Phv2I0AHLV51RCIwhi1T7M6OPdJm5JBEnRSofYQvkKPXv5j6X
o2oyuCA45P1MBIYKl+7KmrUcPTKqDYt8tleFJ3wDCAbFehGG8gBs5+Avn9sB4pvQePzfaF3DtH1w
XzPjsKoP3CfRJCMXpWgPI0bBJXtXaGUj71tpmnL72VabJ/TUbytp6CwXbr91LIhTcPZctja8Sq8E
QKAhUsapyUgV3n35HnFwQsFir+wmLF9McKR837c7lcrCvUsuF8UMcqdSpUD0ifm6Jv0gHBRJfS9e
6zbxbPjLpyFB62I5m0q12Xx3gtmi4PJwzJ0XOKScfr3Cn9EwdJvxluwFmFyvqojQXYjG6jm+89hj
Y+vxhcLK1RUXilpAjaq5eeUs8yA6bNTZpOUxhLPdr08BKSi6OtmhTxIUYhznQY1WNVt7d/9Ya9UZ
7516Op9YdTitgWr+cEXs7gvPB/idtMPL3e43ExRjiJo2MeLIRAd80XQ3/Z+bK8mii16pYydtdRoc
YFE6WvwpS3g3JvfrwpywBOdhKNilaKW8lASIWTe8Ic9o8cXCnjgOBs+p7nrNluist7OdrqFl+unu
RjNE5Bcbhb+drnW1MiA8c8D5nohU4RE6EtxK7c80LqniodHQ1u7eiR7UQV0dDWYyAaA430tXCwKL
kXc/O+goTdC46unJ5ye55EA43XtQesP5iC18H1jd2b6La4BHxyCtl9CUtflAQslo7pYSK8u44Jd0
kUpsPWJSWY9He3I/cEh3n36X8mmUaLF9E8ixd2TBvZM0WCHXo5hCpdRFpBJkRBJ52BOa+NmpvQ3A
ZN+WOzgOV89lxJkwBgb+t7Li6gENYh+kVz8oiXSk0WmU34UGg1bLK/dXQuUzpmKG8f1KA7+K6Z67
nrEZUILK+KHRmBQvgYU8ShibvZVNY4rtzp7OnhNh+S3tP0g8S9YirSH6QRtlCXc1feivbJYw8SOu
2E+vItmO/mLKBF3cvgM4wxZj2hRPBk9/IvGuEIKVkvayVLgoWN+iHyLyLjQAhm+vmw5/1wCWe4Ji
0KOQeHawCD66XjBVE2IEQ5ajyyz2mhdr1i06ID5FFgETYtNIaR2n76SGBF3o6yRMo1gYihe2OQkx
2fR9Lj9LDjl9hBCsy2wlbVNGHtpvQduiUw5cx5vZZTmcPqa+FVJvqJhw9bGB/Gz8TXMDFTNEN/9a
a5NQ0OC4P7N8gGENudai5sg+HBpB7hFNIdOekn0pGyyFIdVS+20WPEqTAHiX2PfH7aJ2oMR5xAri
HiOROSSK+CxvMoYP8zCAYzwjBrV5pNOj/x5k23sjAsrn7MgJAqH8DlItRml8gTAloUk5zt+qxVsX
A0ypcFFKk51G8jYIAwnFhgUxDEoEkF98NzrIU9mW4uU6pdms2xbW2AEr5PexmcrguM4CWyFc0AMD
pVZ+Cmiwq5DeuxtSOpN6pvz6Ra9t6gatUp9CjZjRLgHSramvzdUvXS45c/4m8q8xyC4NNcQ21WrJ
5mZDo3WI4kxteSsY5qxECxFLFZvxSqgMm6146gJqQsK3zE0OOtn2ZbAKc669n50COb0c6FEi2D28
MoYM+BA7ASINl/7SZKpzWMpVWt9YljildwJnt0mcFdYTtyWvOwSWPIr0RwQXJ8GmNt6567vn4Brq
ZILKWkEYui8htql6l450bjrruo6ZgyOl55iqLRiPk2rBVNBdPuc9DX3dnkkUmwrq+5NX7RwyzzoK
+316GEj2gJHTM4ciyQcA2M3tttRopH6r9dHCsBRjjwDAbXAtMS8B+80PAH8amn6LHR7kTmxruBfx
5FZSU/wQ8iYEQ0I0KQJoaKHJrsr6gQuQVjxpaIyhTh/Uw43IigZjlWWkmbERbEhOx7bx2IJq2aoy
UxDWAek1Pz1oQ7ZKqpG4Nz4YjR3+XPoScoqKwxLDngbn8yYotliQ8i+bEupajYu8O2/9l0nBOjYE
ZpYBO5w9qpXvt4YJBdVknNiL6mYqHvceqiOKb+hpo390eYah0Id6c6vJyuLchltiZIFMAKJ+FdVh
SC/kwQHcT9WV+VVq+ZBbH8HLa0YeHZgVm8M2ZjNhDDb2m4G7/bCh8bkqo79gKzd8ZCbIrSWFHMzI
W047JTpqxv7qY/kzjlZQijQvWb4+RF7GjDARHx39w1WzKy1EVYjhQRj97ykfTex6gbZ/5KxgucJk
VxLJaob5sb1z+py0ilukqV6yijb28V8WqiNF0fU1qPEzkYdlxXGsHwwJE42EGbejkMOrk+iJXVbq
W+5QwC74e8J0oglAhjQdtJR7nMOxX0a2csBlERCT0uYsw8lls49FtGgp+uOXula9+5YlHKSJLyQF
4eLpWD8hKSqio6Coo9ly3Od3uKO0HlUIhmg7kAC1SOfRdnGV6A+9SzSa3Z34YyOTZl7HUPB4oWeD
9t7lrKmlvDoE41qRGDQIHTOsjW5NxuU9XzjdLn5c9I6rCaYJZ7e2u/44bpe0faSHo+yn+uj5ZO9y
pf+motvG9+D4MyRfC0d5iV63TYxUhpLNrouwskqNANidTufhQ3B/sUQkUH3klnDXiFUaGPekrid4
UIztZrIabi0/3qg/LDqbuHxIbysJyT9Ql3+aTi5mRNH9nmb3C/ixphT1wvyTHAGx5zQQX/xVK5jD
JKsqai1AjWb4ZUSR2cAZxV4o0eUBtqoOeTSbc3wQf0ndHuBXZiCE43a6vWF/w6/tbTzrR0VATThF
7ICLxmlXlemF8UQe3up1eSB+xTHNK78aSrU81hxd3BVmyg/xCjeOyNkt/RPPQ0SsO+KAxsQ4LeDC
iuZ4rsjXhipK9UcVSZIiyf6Y3begzNVFviboXTu+gamnmpl4/MJelOE0R0cyw22d3Nk5U+ZogSZ8
9XWPJFRvU/Oq5SX2gjhnFOwaNl9eYoKlfbgmuEzOomUjI/XDi2J0x78uYc+0DA+2kmAghuz39r3k
8OIndpO5TeyqTViQrISqQMQsTl62D+3AdDO7fcO8PDDAx2je/2r0G7QVrU4s0z93FG3tJO4c7vgK
4gVcDUxX2SkuMpG4m+v4jjWPGRsX1xBlVFzicdFRhZTq14rw0S/CrILdmNcoGfVVoqeS+VPWfTwy
KbAMykHcgUoO41vlZhTOYNvWQCw8SiJormQoZLerJ/8vgbed2NcqEUXiwFqTYhyJJ3JMX6qVGlKw
tUWuFJ3vyPeKaqgIsK8DJ00vA/I0AM0IP8IUZfNeM4m+A7hnUbmix8ARO6CdztdiKhpEyI/VCiDk
nKL+3jbzabawmz9RBno1DzTLaY+n39TQrSNP9nCAjLuujZBezO4saAZgPopEAJQo49WHwg2+E5Cf
16ZpIqxGlRSLVRPEv2T5+pn/YD9t3v6ZWsm4wTqzS6IzA7cM/GGrhfQgVcOb0ISrugXdiberqujn
dnuhulV9yf/QSE1VW6IrRquF+hPQYsxTOAicT98foTtB3xyACEFN7VQPio5v4c6d4zdoivqOKIV7
oQ/HA82nn9L3mDk1fkNfPrMjnwxanfRdxREOhaNQxAZPoSXXmG2c+DMFTbf3ZABqGJARM+Y7OG4T
GDVBRsQiwU9wA3z7DjxMrJqDz9fc/4+waTFLxPIoqvT7tkmwkVW/ZEZiRCamuwHlywGHCo9C4IfD
Wi9OIfXv+5I7OSRFEYkHjwTwnHptOG0aREkPw2MtmnWat37k3lFqZSeavybntwERcAII0pwdJYPw
d0u/mJM77Lr/6F0GsTmvfbw2YDdRKVuraD4GXNHGCsisO0dSdoU5j5hYx9oj2qsouvQAUcAq+8K5
qxEXC2yB+38kBQ5OQMtMaV66xKBaBOfyw+717rYXZxsHpVFMm5Y3OZ7rQIXohJj5cf+YKnQ1ME05
qMm+Y44CF7ucgsRcj3lnvtFGDrSPfA3PWO9N0BzCpKHP1iIuY1SgxE6kHITgr0B0TWCQ5Qm9Xav+
kAlNcAdq0359e6bVzpwm+/a7RhCQZCr87faUu199XlbpyVW+7i2Yl0Rztxpbi/rF/MoQ2VdkRqbi
FDG2tY6TFrn0BrmyS1z8ASrrYEtiKbCiyl3LKlJdx9M/1SJ4TMHecZ/3KWWewJoX9qdaNsV9q2Uy
Z9hypKWGDdtcmyyhPFcmKsanJm4Kubr5q0f5wL7Q+L6OSCw9oJWQnbSHLwHKRz6yF1drKZsRGBgV
+duuPYzII7uuOgxabUPPYp9XOLfbio6baGu2UpHl60sl91wR+m+NeUt//u7qvw5fj6cyVwREaqzt
clBvajMXInpgrAe5GrtDXWe2UieMJzqD7Q1RyPCidf+ehAUMxF9/cE28GfD2E8cVX5m3lm/u/hKF
NL2mrugZJmTgD/pNwgrZQ/RQ8IulKr8VvpZhF/LiKROsDQAr/2gfdzoJixbDh2ji4aZDd3nyj0xT
hWYdpx0hi/d/nQo8p0HJMwm+NJupmiIGn5tz6MZxeSxxsq7KURmsB3r6PiX96QlIjZdu2jqFLfA5
2WmBEc8dppD6Pr9dgBi1rkhC5uWJ83uSZEClEIEeeTRAtDy3Eg55yaQeqRsWNUBnwsVX4B1gPYDs
ini4Xm6rJj2svjlYa1ztiXkM7l4z00ffLjEmLDPtJ8NVaUW4GAfeySKdDolTTSaKIMknDJjTSGPX
0ARA/GY9iB2zTW4mvfTpWk9f/yqWu9SG/33Hp16LrPn2MeKUc+sVpKidWfX7rLmxVaaLfu5ba4e3
kXij4qExrTyV0znq8/jVs6mvJWGpNMRwTrEgcJ5mUp9IhzxGYW4Ti+Q8WF/uyHy4+xgkd8U+4iEh
pFI1WvV+KGL+0zPgGGzSDFcuvhkqTlomC/sJyLzg87PTxsZjS7U+UJeBC2P0XtS0pbbndEv7yrmw
FLth/nMfMVBEsxra1dmQFYS3oASxcJ+S+WhcABGII6pdB+vcLaZbBeT+sG8hA7nzVsibKt7A37mP
6Ya/IOt8kN9YIO95GWQZz0n2m2GVEJDMz9ByQuoQdWmyyjh6P0f5RKpGkrgr+kUTFpDSBxke1jEN
Ik6CTKC4TLgdD7oOyHIuUKIgdv+S8A8UDLJSdrv3RXbkCzxg0pV4yKICBwRAg+10XSBekFzGHeTZ
IA6m879WZQ/ti5x3XPEhxqF2ySf3iUYhJpzlynqOPxSfNVomnbq9Dfz0nYcobdm2o/LVcq64iBkG
BrbzECGemeoLChIKmd1RuuZzcF7MWlivpepUQPzMl2LtqMeEGgVBhOpzqCpD/vFhvuQLRYzjtpU1
BqmblQ7ryzTYDaztOtqoev+rgGpxK6XK5MLHAnWhK1gh/h57OyyVVerU30Rj6dXKCq0yIzE0gkJN
GQIwVgnc8ucau9VajwQLTlhk9D6fW10v1qOrUssdn6ozJFVzRBGnUEtv8ze4Y2cCWniiHjjHLwmf
mcG5qtKowDm9xgPLKMgJBKxAppjEOdEXBuZsnuE49XMasy6Da6Kohiif4bbFEvjzSkfrcdu23fDf
DDctnJrjbz+aCeNVfT0+vuxFfPSgYXW2iUiQnmWUyec/L7PGM0GnpFqtpQs7ebskY0GjpHi42R/j
AXk/hN49LWXdrpPA6tJPvxjlgtTPxwx8yeG8jckOPOJcAOcgfqH6Box+VGwdmqN7mDlZ3IFkNPpT
zm8ff121wn0ywAU3EI5AUMDJAM+84FuXFolOD92hWuaXCiu9XKo0EzIhIy8J0nhwtCwRvCH2HmvI
fRnc7ddv8LptBH4f8eTXvSmD5tUzkQioWJmEVOabz31cXpnikXGHy5J5mErsawwiOyXCdk9Qgz2a
iaUftEeCV87wnEbWxaiPiIvnAtqYPGC7BkDyAF0Yg9lhk/+p1oVVrSp1vEGzcANb3/OOtl6LmyHd
KLprp7gQw6hcl7NKXbNBmXgb7/rXUu6mTRIlrF9fZcr4DXIHaFNl7ioOhB2zzWcmQe4MgsN2b+OY
zvLLKzUCpuGzk6Gc9Z0l/WBCtblyFPVo7JwKW2GFzndYCTsvNfAh8DOv4Cd8WHEN8iT+vLZn2ZzA
92/w3lYbwhhEytjyfMBgyrwXn8ghPl2E9KkRwnHN4p9ILVE9VokvCnEb6e9AgM0XaoUve7Ck+Uf8
nYVoHYTWTNiasJqnQDIZ8uwFVg40wSMKcPtLwGt1mugaEvdMJaTEEjG/Fpriqj9G3kpnr8/Bgcu8
F7uhEcGSrY1NfONH5zfG1edZkKy093etjsPRK4WFy10Vu0T874IZcHYxGRinDjtIrcJWEyNjrU3B
OLQsNIPztFMoxaf0LSS5weUYdPlRJ0TDtb/HR+U2lGupjhUwj+OTFlZkbi5l2WvkO1knxhM2D9ld
K00jUHqHiivb9+UhfcwM/Kjsw8kE1hgdOduP95zkJOdKBnsp2XpP7J/tPHTS4pf/zn8461KRgiec
PoGI7gsSW9Ar2NOp1OfTFKkp45HMHkzHyzm/Yb/ZD9vBk24kN4eYQAalCqJax3f8RnYd1SGVz5fO
YbvDqpViJwk4Y9/DlO5W43SpqZxiWXA2sU9UlJDkxEdofx65b4M8+hviAI2ckfEB/xS3wuWh6ihS
3aYgYOXItf0gdwUm0OjW5SwEBPqR3P3f8unecOLj5omuYlKmXCFXrT1gMP7XwNLLQT+WnwOKrWYd
aLV8VN4OdTauB4BwS8ZZg9lotZ0E/NNARLjaYJX7hgfrztpYUzjdQtI/fSQlOd8Zb2RyZdwfKMvC
7crUlGzTC2jEXyzijzbuMc1Uq5eQ7LKCn5l8pXwfq36ixDzBeYNjXDrMRS+6J377XkHYMLlzD+Wx
Qy4KELHjdXF5LldGLrZ4AFr6OBsprDG5r+aE0jyM2xUnkg9xaSnmlgz8xRZ8GvXyh/6qEErsdbpI
WSXawY2d3U1GONoYdPYp6xFOTxqexDiQeYy+liPK0e1ZPUXjsuMvPtI6dq/kKRLKUx8Pf/RZcUpJ
lavhzNzrc95baYjUrLDCsyIGQH6LgVPXPrk46NumO9SqqRq8W99zJVkFGFajSNGKqiscg43VCmAN
QeUg87dlDxhpod2BLoTpLx7h39XbGSYu+NcRd+3pOTTAgiYH1NUw0eBwCSSwNTqw0gWIvb4SFy4b
0snwtSjjYQ72Mtsp6wNsMa4yh10rDfLxGYQI9XTEkCcsGw8K4ulG+YbPjnVSJ68HQ7MA1OiVS9KQ
8TnQdQMHvOPXGRwPvzQJ4FRBXMsxgrHYa+3zrNk1jLtxGdSADBBXYL22PpQoh0Ky6c5AO8KNvAOF
EsLBJkvfM6Gi+nIII3YwKZtnxwW4RLrTLPMK3LJMlMES6FuebBjyQfB8fRkBUN2xjED8HRUkMagP
Ieln0fOQpZkmOlooLMjgimsdw+huaqqjAvk9Q4DHqDJ75VZ8ltc/jfHmYAd4/NSC+zGERs8LtufQ
965naphK2zWvnUXVlDnP+untkcvzGgSl8hJ+y5qu5OpMEnFzNfkhkRT1GzR/NP6JYQ0KNOXS7wg3
Y3xisFZEiTGahk9LCesaaKqvWvCrz+2jvA5CGnUq/jsDAZbRKDzPjmcvjoFznSWvXcezJvC9UGpf
ToZ0pMhPwyqZHmircYmu0RoNMw1fnLZZeQQF7Gn8vyGeLylqhsSa5XgXkEX3vkFTgiZud2IXtpXS
jTYROgGNDm1FfFNvUZo/pj9t+wl4sfP7yQBsNShCaWNwrVzC/zmErhKTYszzOwLLspp65EdACJLS
pwiZmnC4x6kcCndcsP9Qa0H9zDuft6PtORwX00+JUUBv1eUSvQWBf9IswEWdCZgnPbcgbxZUgwTx
8+Ul6zx5GfyhuuJqiT5i0QwIK/qsP3gaN/mZbPZxBsy9mSsBVj+9iPRlMEI9yzlvbgQJKa7JtqIu
plwnJTmUsIoyl4RElcfl7ptwf7EQenc6vhnUM9ogx4XbEZNEUyAZCG51NFMGbpKkJkVU7mgrFLmz
9Y7/1ct8HFTAVHxJ7j9klg7zrwa8rM1qCUZoZmSV5CV9kay/2le8hLqJvGxBIaPbQFu4uR1v4k33
QOVyzOvJqqkgy7vYaaxcRQ9SO6TGVY+NKqLdXFa8RbnAIml6RtsjXTCRTrtQCstloBgAFl6Llmco
tHklsJQDj+l+n8FULSym1XA/Gp2Rnh9JlixDVLO6dqxsbdSN6t1onpMrab/+pNUqDFJbVpMhgr5f
rsinvX8DniazfiEPuyhaC3U9rJobFyReLCcbHF/LtiZVpPRLr2pNstGyrH/VRxCTzO63NzMyZk0z
vxSnmd0do08EIC5etKkpRxkmgaqxvfXO04GRq/OfbUUEbBMQO5/1kmON8q4msH2lXJuqOSGzDKZ2
twNl3MtQUhLzcp8CM09ZuSbD8AXtt+IFoJZ9/kSOKWYojPxH9jSJLd1JcypeW1yelYzeOSQ4gmss
MMoX4HyKdA9Q190/pRRH3xZqXn+MEMzb7S+fjy96pomQRZZ6gc5n2Kw8YHJvD4xq+Go8Wu50GlzV
OB09twz0pV1bJsc3ptZwx1NYOfIyU6VMTXTE+iNjh3NCuPlCtnWaIoZqzmeeTDbiLWxfD7Pt0x2E
q5S4TZ7ZXP0vkllk51wzquZNlFwctbTJX3Frm8YDk9onHcFVxeF1nagHOVFH3HNDqt+QNBMpMkcj
Cjrlf+LFcMbKQmC6H5nc8niGh4vFgs+G/834ZvXJ49eTpHuAHqA34q55YuCxgcj+Y+AjfAq95J+5
XEOvxelSFEq6xWeJbVfIDD8cyzR2iffpt7a6rKd27UZ8dO/GthqAW9m2g0kxlAxCPOfMfFJo+tfQ
fVn9ytVXrk0mDoMlhZ8RY6KEJhkxWR3qAPPPDmvFLHO2cwQsgwHouGxzb/TMN4XTiif/sqYEAYtV
Jx1jkXP9BQZhFHcx9aH8uyhtvZAxqvYFlruBkpeWOpd66LpaDg8dGpWJAjsDUYLY1oKMuZ41Pf+f
DOnWaT4MqxE9liExMVjGFa1xy2Zu+4FD3QGo8wLSkQ68Y2kDkOnyA1VKfjhRjhuoaUlvlhOYOoAR
ShLGZ/2wxYkomb3CPsSoOnXehZHOgqL5b7jFvdz3liivEZHBBjmIwhTAJ5f6l/BfVnU/1cfeEk7T
0PS3iwKiSwhwYam0D7+HYDTK4KLvNjtxlubsm9j89oAvt3DzN73DKgV5L2wB7f7vKB/CwzL1GzLU
PuduvdOY5j3Qo1rVwoujoBIz13ZIYw226zc4YCimjSRts6vrxzxI+xrZ+tvgMJl/mHwTesLDVg0m
OP36dqHTM2udH7wjpjRaRbPVVYLl9EE8d4mC/0kdb0OKxKU2rwwkXcYC34FlBCFY8/eh/t+X5xzn
FlQXeToTUEYUUYvtOinOvYlAYkQhhIJ+INDcYGQkdF7omjnFcMiqX6eiRWzkhC/MwS+0g5g+NTWP
30RD8CRbTdstF3XEQ0I3a8lzmlNLffuo/GLbkKDiHmwTnJq5GJyX8eNgFqaQDj4BoVbe0yO0HMlL
9kZW1NLCpnKvGYHbHCUo2wxn0AMRtkcTicx+b2V4cIcMg4Y/G+Yko4GyF9Lm1dzjh2JpMa/bC2lX
9iMuv+ZqStMYMl01ciA78cSjaDz0Lb8/M90dGEX8RCiY0zTu83CpsDtZ8tLICvOAwa7qAS4YP6gT
/UjJe+Vi/HlVzd2oK98mqSK0q63nNF7MUIM1Y0whqCziTRp8wQDGjf3NwLnjji2W6kwjsBv8ofUn
c1RvQZRCQ5O21upx1pUSruQQRZtvvfnfh5JJ9qY8kbUtcOsTcZSe8ojPJIjketPk9jG2ToKIEOfN
zORBTvhXFRnWNxRE1gZYxcwtWXPFpQUhHruQLIalCjh9ZAVvN00l4nPM0nPU7PLCQQebYO7p5inT
tpXtA68HV7zgB7kcfyTOzAuytkSeNKGfL98lay7cTC/48Uk+lUx2WWRTHaUK3ukUrichyfry/AEg
hBc0E+Yo4uI8loqdHExNQ14Un4ZbKJSG5lNQfw52igDMVv/zGId8A4HmTYQC7n7l7WrhAzzdRGMI
uP9//ALxXy4/tvwOmMZr5LOAZFehghbElKnV4TJeh3lyX88BE6gfbumabkyh1t1P7CXzgAkwOAyy
NllrJVZH1woUOBdnzK1fScpMVlXgslG+adlMxICQ4mddP7pf7D8Aw9qgYkNMwojsb8vhNLhPDGkU
w7reC/Z3yZUTa+Fr+WUGf79jCXwdp9T9OsCq7JePY0F5bUrC8w51ykqkp5Gj7ybGxAmnnx5P4lc0
QPpvxcuqRiyyII/kts6zHIrjMe96oauqXZWk7+jdnJK/cYRiVQSyjQni0YH2KunhrFo9KOiScg5Z
bE8Pyh5aJYSJIA3DnZXkHn8toe7JPZ/ZSQwjDj8O26QxvYg74xlMW4IXzcuS6qVP9Ax3RYLLnQ2X
v+NSDXeLWRimovMpbNeljabo1lR3CCoEWEhkWx1bPXVNtCJK8wBX37Zs8GvxDjEm3pYet5Alu2vT
rUA7wnJIgx/ikawOT1+kSbJ/zFlXSmiwhSWVWRfSxGk3+pBEk4JOWEyOpY/sSJYbKPanaCMnXIeE
IytPOQDsWOrmdVng51KId121kD2nT54as0oKIhn0d6rT+K54WCqTTQCljzMkFAm4KRxWi0QbTBfT
iF/HekP+OyuiHVAEmOcNy2oXOcw54b32wUSAMtUfo32nJV7hex73j3kEoGbHAWRlEr0TNN4K7cvB
KQiiEcYJ/cS3KfndQn+K+lT+6YUxyIkU1fkaWeLG2FdmQE3x2ej4+w6oE8+l7QkYn0ZwIDeg9Y87
tZKFVxxzUQgwawVVCp71Ywkxd/DDV2kab8VOTGm2hl052JUokZBglJZ/+7m/9dpbzgHK4fGGNtbh
k1PsMKRYK0m7Hykx7EqagA8eQd1kk/4oGMxVtICSlYBdEazpofG+qQUazEuJjFp+bk0svORB0f+1
Vfl89CjQ1VvnSwHfO8InXcBpfEAxeFtW9C1q1dlgcSwjLYoCV9IZV06NBGrWeRw5tX/XEHm5AmeX
AdRwLh7e0NTLAXWVIje5VVE/+nzN8dn/lfMRYETc8fj667lbva8dhEwC73aDdamjgLivDAbAgdlL
zg8e36IF3nllrQuOjMHkUVss8vFxuICs8z//FrOxZlGa9jb4RdR5GtqH4fgdB4LY45xrRYmalm2e
vHes+W0/6QS8jbpNyKQTGeAn5Fe8+a2XZ2cvgl5oBBAfRoiFBiONlpChFfPcgFtzP0dKJP2itMl0
jpcqrElnmBbFB2IzFbpvoSh+9aIw++ZEusWNS3FO5x53Eg3oa2JNP80/01TexkeRodg3ckjTB+mU
XzorKQSuX8ywFn43rkGQKcCM9x0chePiRh2hqxwx4YyqlCCKE4IG5T8xfWjxOEBO7xMWYHdeIpKl
MzxhkecdHwNAl4LnDClh/nxqRUiMDEzNrRVvzls5gDZH8mni5teV9doZ4MBxTKFPi3NFmreE7aSq
eLKk7APeA/WjMVEy40t5WJAW+L3/Vx4/wDHNTtLEDxAzYHE2IkY9fPx22Z8L8LQvfh5/usQ9XxOZ
pDcztJAUdApDUInKu2MHI1XeRcsSB0zNfU0KuHDaKG+BeINpncbfFEjB+Fo8SnhZ2rc2xvwQR3fR
l9yBL5QUFgaCLsJXIQozz2ewOUyzWzIw1022IQ1HosGbm+BQSgkZGBIAF0e8GzgETT7bYvC9ZNKx
Pg/R2MYizVvcmg5jV+bBmeNVevijSaNqHljD+0Xlc3SL1qyZerGIPtQJaWFcsJGHaaEiUFM4vR4/
/Xd+7/dfKHLbzUQPzGWA/SGbzuxE9ayTCFzKwKIJbJhkAOCMQEMtJL1b4o+ow0Y7nS0fvXjuyAhl
eeB9OKtx8M7oqvuk0bYFoRebvkuCKsu5gmdZxy9tgCYsximSQRjBAF7pidBfKXigjeM5Fr3rtiSl
OH7f/r5gHDZ86XXSE0S+bvdIM3pu0G64QstlWX0VEHn44b0UgYVGMp4HtX3oWePw66sZdozp08dp
BPmVzvQ4/qepFMAAKRhOop42EH8XNgy8mX3aMybxGgEZ6Kk8l11ono1epClqPq/jm5+aOH+V0EAP
zstTtDD5R2JXrbPdw+G7Z6LkfdSmUNct1TbhhTGhz9QbgwFQRI6J6Zcnyl/xp7HmBtDRj+iW+kup
A5J1yqgppvh5A3LsAUpFhFA5rJaabla5330P6Fv1QVmm/iOS6g8AllqxuLjp1JtGDH8PcywaXD6T
plGABIiyzy1ynO0EubxoJX+NwzJZ7JWlAWTqWdcPwuwsY4LhS1W5fGug4W+q4SkxR7gmzLgUCmOw
OpqvgFhL7xIcoGpakHUpR4q6CIPg1sNlb08hvaWG4+A05Qe+lgcoos6DR6uEaVVbDfwZfpQ2DYmQ
u9n7FTE/gqQss9LI0uzP+wRocSB2vQrEZZjsVRSU0lpbOwsLlB3WNbXA3Fw8AH+p8O96fuY52Ze8
ShL+n0Q5RznAwZSklcQBOJfgQ5IrXblKk3jR/fZHcgoyGXba7bLiuxCKjXXX7UVBDmIiWZWeByTX
vBFwEr7gzlJqS7PC54Lp56QUxD8Oq5nU1pcOrepmX7s/1lYaID14exgpJBrxxuXQywfyGi8Ar73g
0X7XhPT7SHXaop0Khmcr3RqaX78pGQhzpPxmoJk31Vt0dcI3M/MXD2kzxxfzJ+ZzQMebuyarz7+J
mtOe105MxCbtgqJM0jFCm8tqXIYmGu5MBOicK/YzObcLs+KYAEXqVMStsQLaHGh5oW5C3UxQTVvJ
F9HOYIRi1XKqcEewbn+8LplsgE6lTho9t8AlEXuWCt86UXEgitumkdMYtZSO9fyxwSSS3EGYwNzJ
64xqqATQyCskS/iRcrK3Plh19dqlvSR+GdMwiKMspIYeT3jgSpjuH+3Qi7my+nMrZsxpLdu9YghY
nCN4T+Pjl2Ouc7D1Elu2kFN5Xd47qARj+tis5GucNZCIJehFko9ZOLFefi6oxGicYl3jvhrrFNCe
vLXfEJGeZd3/iDn8DXeALOT9exPUm0rtPSx/a/yz+RRsVgxun44pejwt0l12JgeXULxEyCSG1Njg
xdU8oQanUb9YrgUIjfi+EYoaPtb03u4eZEOjLsW/FzYrIirMLR8tMiRQeVCi3YH7X5FDb2hj1SU3
8jhGiKJilwSz2/VCpfEsyexg03WN/yFryl0CyHEvRXX7sMFdh1eSgMqEI0rUroBQAcbtTWtn/zhV
35QlihkUw+RWyezOGGQdjZcLpV7FEdlKzStrwzngqIoe/9v7IxafXNRhgPHTDHE6Gr3ZUU71j7zO
mhmDkPRjaeezqU2RvuEdbPZo9difYP0EQcKhCaS7PTE83HfIf1SVzRf2WZ911CWZCSUTMPv0cviC
ZUD2Y1QxD+zJwHnHDMGFRveQEitv6LuUFE1BYpEGj/IFLdElXSqjEQT1M/kWnyNT8umzI5Zy+tGM
us3O8Q3vJ2Usb1ZIMc4xrffZa9WFw5wetC4qiXy2rn2yG5QH9cfNCmFegk6JF+KwC7HsPYWy/s+l
Pfcu3x/hnqqWsAmbJyxgK0EprtzcsmFdyeun67PU9JPgKs2T1wVWI8O5/pcpsl6+2LFA9/D9tQSN
wMtAKX1WBKcMtQJi+J6/2qsBXOt7OKbNEBXapnPMUHMzMg4nJ/Fk/aP/aHWH9Sdwjbr9BfGPhzK+
6MwvFMSgR1M2GWlAP8YXdqSjRXJDUxiv9tla/9kdjz7JfuinJtyYY7pl+N8I2xyPxuMUSkdA/EXT
krPkHTLpPR9Fbd/mIAfzKZn11jD3KsCHd9ftaZEU5x8r3vGG9nZrmqzQ/Vv7GCDoW7kv/CCmXIgM
9fIEi17k1wcTh1x7EPpSxqZw+9lk2t7dv9IoPbddEeNPj7eWNlSj7dWjkpU4avVufVEjiPHxHJBh
FijCKUgrwnpAujIM5vfGSYFLCq/TqmsYrvppTBicBtDkGjBdpBH2A2zeQCzXlnWYb3oOAQRte+Uo
nUv+ccciMklJmQ/M/kXeiQkjuj9OPWhMERLHW7N8m1iu9oKSXqFjwU1pDswROUHKVekn+42oKDKZ
8EsX+yk5PGnhPOOLyUtM/G81INgv/1jTrtPbtECl25JrylgM94HxpIfWN+CYsPTIuXgIyNDYOc9a
v+saum1DnTAgM52p86pSxH+IA4D15nFYJTtgJ47uAu65hE53OiLGyxhgOK53aM+3QDkLYqBk/TLA
jw8fCiEUrGIStYls/8tVq+4BypE9lI6OgWR6KNflPur9s/RG+uLrjFcDadOcVls8yrmlgV1RsHbH
cO3nbjpEQf/IdIM75+nqdFLORKiytrI9YqE3txOSbIKz/IpI4BbNEEDILJtafY63ZY69z8KBedKH
x2GX3Uq20dCp3GaWWAxK2ndcjXrdNzPWuykxZ/BUyaxuA2G2xuaX4LHb/fOSplycotCXWhty3QDr
z0pmYmwh1dKJOs7uwDxqmQVdEKUtVGqGkmfZq8xLcRjWdelzjUuVofDATAtb0nZu8IHOzqeO1EfH
W66W0Ugv7QGrfd/HfIi8P5zjGu2R519ZIl/jGx9oYpkxmr4sDTrrFaSU7CqkefyycfE+ert9htB5
goMmUmY6WW8FfoFZwkjGJWE1M+gGHHg7+y003VBgpUbSsTFbY84BREIrARe+M2wPrr3YdIM0UZL8
1Jq30EW+ih+2hApdz43flXhGkoAG8lJitMxVoulXEk6JnwdCJ+0ME1FqQVNXW/Z49simmullJSFr
S6TCjh3HQcg6s7ZmE9GoiJJlV0h0Okddbj/Y8KYujHmsHU5MguQJ2p9MHTR/+hCFVSWaccj1nKMR
GtAG8lfovO/bsAjKpzZRQ4NwLCpb2OPfbaFMFJlLQB6B6QUG5yTRmJFcuZfI0gTbPyGMhPaG5vjE
VzDSLHzmyrqCoA4YmonbJRnkykQTmdCN2+b7LB7PGNX/wAyzzQYsv2Szc5VdOFkGGS8h4RwpMWTX
lZlcUN+PrTV66sIB+/fVE3PJF6yz+atEenRbGp1+GDqZCDMFuMlHgxxx9vkJtapUfFy0eSwcyzSg
9YrRCIzfeE66lMc3qRvd7RgX5GUnd3VoaXhULnlLZ2DZ53+P1+PAMoGZKT+R0SksNjLF+Sjd55lV
pqArsSkCMJSMSMmkQV7QUn1O2v/ChvHyOkeX7KAOb2niUIvstZn2TP7JCXfD9pBCdhMW+5t/rK1g
Iqct7ezJ9YB8yMQIsllv1qlgERnuyS+1Bcvx6VdCOzZWVSH5xe/HQScH44R9nyULt1fmPn1SgWPR
0sgSGiFdEMyFa2trLR6ob/PH9ptp1nPaD11qmdYGljBFsPZuFD+7/Pf54OWFGx0iEqWTAbi9+Pyd
lvSDpFIqv3C40UJybhYEo1HSWjCC7GlU02YKmzvDHxzUgNmrWP62Yxs0sQbCQf1QPbC7sfMtplk5
WeCcX6BJhu4z0uSRM0dED2iSaqMYrLWn8cRfg8SVIKYN1jMXsQ06Aj2JmIaJLPfuW2WpDBZY80PX
4weTMpiFCGvMIEDEob42ivDEoAdJawi2vUP+1M6MCwKcGybKNLOO+P4/9MOmaQCesGfkpEqvrmg2
rVQJNPRYTbFp+HHlN99XDwk+OcD1QJc0vLaUGothNVZKQHVDD/ebcJGe55bHy/S/pT5LtFI8BinO
CBLfokzEo1I00hUgaf+SLqtwzMC5lW42iPSSNS7nfzzgfMOXrfsFEzILd/wEy0y8HsPIHChTa1wQ
mNHYFK26RyHSxLi8kMc2k/SkTf1wyYNkDgG7J53uTKGFwyVAyLo6p77/Q8EJawAqYp5TwtG8grlZ
KMlTiZoQRLrCVRbtSlrdWrRxJssISXa6LkryLXehM7UlBIpb7z1tm9tgceFonCcSO4MRdZeZxh4R
cxZPDRDzZ4sLRFMgFfvLHaK04lnlnStxltdeUg8fg/inaqQ/bnfhhX1bERsMJJqj71MkwPQ10pHl
ETfryYzY+VkkUnKT8WcQ8Kank3HWUpLLN/xKy/NKujvEsTAiCg1KjSgpGjMmOwTGaEIVJsn2Jmol
2mgy+AlG5pCAFPi0TRZ4VXKXG9jAarzuDreoSyS8Rf1lzNoI8OctNKvrdCaTKZplMNC7AJ78mKYh
wx1zmCZDxQrYIvJcKUwVFVWCkXVLKyB6kb18tsEgEqNllkTc0eb4I6ZPzgZocleySy9pEYI4u9hP
GBZwzVm4isXtbISv78b0VIJZw0q22CXcWn3xM5ZaapS/NPNIWJ5SHmN8rXrdvg3H6wwwZ80mRKFZ
QTSBOgfmmTXcFOUsbmZ0bPdB7JT7cD/AhbB/B7aDfLKgdl+VV7fCjC+IIC1HXJCfm8kzI1Crq92X
VEcK1krdvm4lZU3kdyLr3VA1tZpQWGxNMznlnPhVX4bZohkcdOVeLKfq/9HNIf/54CZgDec4aGRO
3S5XHSqb1UfMzJNVTEuUIvUCx7pWiHYXbC6YFnNJPdtnNwGHsQ7Pweyc4tqtbLRe3stICo3PfKDJ
R0OAkYC9TndXXkEcvnXFwuSKIq/lb99E/+2YBNUNOd+1zrfUV5qGzegXW3xtvXbcbtQyOMEs2E9B
vKMs9Xl1ci2fhP+A6ZHj8HQWFk/q8bzJRZOGOqtkxSqJSqvfh/uzK+z9yEgQ9pz4/cUU9lzwWymv
UZEqP/5tL3ETNPDVVOVun8neWSpT6w5HloOgQpul2Fj/eUnZ6dEwqjlmL4v7Y7ndf+BG5WY3au2Y
ttW8cLIl0bKHM3//fpZ/nL7xe6jaZIQxZ82N+JX3AB0Kp5XTebpKCaZm6mrzfnYrXTx1m/oJnJ53
N/lIZ0s99Of+OLvdPBZDDyODFyK9aPPtXKVeNo9cLPVzyoeJwxVCsrfXqkVU+HPgfdM5al0UbBad
2nHNA9ANfZtr8SETSQ9UJWS4xGTNMaU+uTpfoetUsFDz8YDI/OHnP9fs5/ATQbsTKQe2JHwe+dq+
bzuEYt9LcsC/qQzXmX+YTB1+rNJIJgDxKTRZYixYcLe59n6FhnStOXYJLgBiqMIco6q7isq6d1Yt
bbVVCWiuhxs6NShjXDpKOpZa0YijgDme6c3kbB7dan47xSDayL0tscFZ/2u2Vb0TTaNCfTht8MY6
UAdj5JuTI/wWA/LhoYJwqwPa2Rpw/S0xxREDqynnHxKt2isy7S9DpJ4WApTvuaWLKuiN6J0pAagT
+Os5uzlwgv46SgCVQ9NhbbFbMMQHsArzwKjZn3S9cb2W3oYf+F0OJ+N+CTeElIoFQ3ZCW8V6IVfK
vh8fpPj978qXtKk7pkQ9DB2VirJeGI2joDtdx1qdOzS6BYZPROcvZFqGuU9MaIXQoUhLsh1/0m3N
mjdvuBjPJ+sG9uGKorkg8v94BsnWfYcA2xxPRObIvHPWuin1eGa5xs9VWo/XXKimboC/VnTpKhHo
hr2r4VXZw7jymZa0KXEJK4bmoUvMz+qmrPZpzzBYsb7bakuZvByZCuhLNV2y9qVRaLwWRziKVnEC
h0llA2y0tBCsek0y0RiQ3HqOqRBZM+r0rr65KaWwh+ZgpIN0epAnABGDiAwkbzruKE7knhdx+XCA
UVHXAzKbCiWwuT1jhRPeGdrfbCzeorB7jWqy4FPpBHXbvg0GyrNIAggzhOwBRwqq+33cOl5TXJwv
0qXMUEEefY+a0SFB46KeRyCAYbtvyHvI4zMPYBFj3cwIXuJAP9zIDAw4mAgNNXJAd/tagW+Ysg4t
H9oApn7aByKQjKeCkBBiMNuHj/PxhW1VC+Bfudd3511zHRinwkRKNDjgj8OwL4zv8EeriKk/X47l
N7gLGKlCpwnb7Nh53UbMW6yd0yNN/HI3iG7LMlo3lelmsGROlcSbu1xABMxQqKcL/96tH75QPobP
ELR9ksccVvvRoignL3wOJ0rjnPG+YrG9g01sVoSfXwfv9M6gqcvfl9Bhes8pAhA0np/usPsMzRu9
TAgAfH72XzEauwvEKF5KB5p38Y5oB9qvumU2rW/bT9Xb6cqpMXAhE7tubr7wtqfPUnOH7xLYPbCB
h8LcxIAkYKS/qKhGcxWTxNNJQ+n+DZaqEil0HjPjIvjfjlqZHcHL08Dlk3kCXurdXv/IQFcD+ceK
fJqx3fUzEKrw46ojoekcbGXZq5d002pxtsafaWrWGXJTH0sJanm1oB0RenFbpf1WU2YC3Y3Uyvg9
QLY9BthEPeLY+hmCYiYQzhAJI4Hob9vbl/ewa+bh88u0H31YHgjgEjV7KfTpUsnu5N7tTFs2k/xS
u+IxwlWCPEve2wZ60sL5MjLIb3caW9mZLHVOok1ZqJI1RmS2WPK5++66uEV8szCikhAvUcJXgt6k
nk10xI2+Xjrj+5YvBXpN39wakUfERKKKf2TKpR1Ifsg8pyKBI9cBeMCSg/0X5lRvsTuS3ajcBm3i
uEAyo98u5k2cz/YiZtGwdB2jtf5XuljRNNsWXTJfo2DUDPMuyBSC3qeURySR3xZAe2kwD0kZdKVp
OzYdDnUUAPcMcxmIOqG8XKEAguKPihftxMlhogyvEc1AqncA0JYu9V2CGMbO7HPDTDr4hFdVwScW
oNALS6WlkolWHQdaqu0UsY9zFAZAlTtnfPmZ01dYnEFtjyfu8xnNkII0NuYu86OYtrno0aCwriOX
or88DckYt8mwf7EFEdhKrxKdEDqPiKh8p1DfqT7bGYyc48knBXGQubqGk8jApiaZvzaVUdzwM0qm
0Q+JwuyqPcAM793rmHSAje4J4lFEpxIGmFW7ed4mD+j1JyQ3bJVQLfrlv5o1moiJk/l9c7YWuEIn
r9DUG/0drEJbfKs9IBxkXBd/R2y2ZMvbEKeKBlV9+lzyYnST0Kr17YXwLZvEw3BiE5C9lrmHrKYH
ye+w7gFvaPIjKUpv8gVMvClGb0fbkOpHGBc29mmtYlXnUm3+3aBDa7ZdbZ4Ocn4miRXIUoJkOt0G
0AfJi9G//JI+ClcZ/T8JkvWk9PEFBKmvwQFkI3FAeG2T4cQ1OtXyyEtQYpvUfFxLPYnzAD8TPFlk
3SatK9GTqXJJcxNA3w4FKFtOoKCEstmyi2rxr3yGJTbgq6On+qB9QW6nEEw6gUbJ4jpsCvLFwKNr
C7BmBw4eeRUOKpt4cp4g6YpDmMyg6ngGLRgxTzo094X/OgncRDPSxjDDG4UnGQw1S1q1zhd6BjOv
0jbN0qDtO1fv9aIj8T0Hb/JAfYfSEK1hUyJDQO4W90JlB1mTjxg2Z36K0aFU8FPXdvYWNSNUIL+H
487neWQcaSHx1EkhOMj4trOW9tRU/PoA0bqPh7SGa0q0ZYUxi/OATRKLoTGsCHYo9tAcKewmYcL4
kUvAVtVVfgfJ6mUe06lOyD6GcinQQ2ek/Y/c0KJ2rwWYoRs3w2p3nHfEXA+YatuQ0reteAA8/CFD
+3YSKfTim3F9tgHHdNkTd8qRrA1rCHEfaZqm4vNEaITYAT0vmAXGt9Pnwj18RC0acplRZyo0z6lR
CEtEQP2ygCRZ0hr/vw5gzrDeVHI8XZi2LVtED7U1U/v42BO9A5VsOTzMQriZdVh5bJt30ob1Gr+Z
tuyc3lsT9DdzMuOCYbzsSU2ObMggAzVP53lRRxOntATOxGCPs7SAkfRsvCqothBu7jxQYDKv/2CH
2p2DJL9hRkJgQQ4rdroV4eHULO785yK8Dli6Awg1AHr7bK2I9gZ7OYhJ35D5LeWv0b8gFQEiBdS+
71uIegJjoI0QTTukdPH8PLEk7icv4N5JKez4qLVgwUFtthQ2WysKKkju0x875b+QNrU8j7nlWa+v
H9m3lssyS5lbPlPPJnDTPrXewdRvkRTNeAo/AKNXk4IBH3JXVFJg+j5ylxX548QsDJx10JcelsdR
SOrMmV/UwwsUEz2mexg1xZSlyga8kx8q5S3PdSuYn0w0zYzYaNM4rL9Q0dSTVq7w63pW/etu+n1e
t6TegdWCrFKXo/bB0kM+utGkIhdSNO/fn7az3ot25TlFBuvVth/BbIPNt+0kwHC1oTL/LPzgzV/N
40Udh8XWkuaCFzmFpAH0SwMlPwgee0DGW6Pl0d5mfnRx74BCyZf7MgeZLyhJYu5b4pzbA1ncztUe
ezfrq/Vl4MKnPeM2g7dQfMKp5ahtA6ifNIKHSZkjOOa4pbCwi0dkeWDnbUlZI+SdkLqfS9VOblf/
hwlmSbf8CRPRH9/Gdzc7sBsrOesbJzJ2vSavsw0AyBvzFMBxCarmfqPIo45hfqtrtJzVBAJOITgE
ihRnd57/ecmPy8DqFI3q9bu7i9anyCI2gKurjucLTagOIZmCti+G4d9hWFaBxmtQq9OSNlTfdCHG
bGTGCmEGCDAN5pRToow3+ZYAaTeP90KtKnFfqghcs1r8hLuE+SEog4pR84RkHDtD1d42cnUIowwR
IENdr2KFv3DBmSN0MOJosC9xFlp1JF0h6aSrlYYX+71jkswdc75yxWV6gLOSjWoxbcTkrwipyQ9Y
ltDFubyophjJ/f3EfYL6/UU0E31ks8c3rysn7dJkQIykptgK4R8EzGJ2j5e7DVX1tZlkrZPi9ASn
Ry3YFv3eZ+kcC6LW/5PnGRdpmdT/wMs25C9M5PK3FKXDgMUobQrrbxt4cUAhr2C+xKz/EY7ENXEF
2/xZec4oA1CzMj4btVQ57DecNP49R4crTXM6YovzYzoajzGvxdOw3A5cPoyOTNfM1lFX8EgbUq2B
pJPiMPBBwkUpD9mfJLa7iHbaenh3IQUq2084lltLc25IaI7V63r9Z4giUJK0vErVeUhrt4zenXoa
2N7cKj70C9PFGWq3jWB7N69SnxW0S6IcDeRyr7646rpstp4S+Zd7PP9ePLuc0dz71c07cOq/Sel4
aubQOSxsossRhC7rJl8Jz63zBTc+Sfk4IDDciR6MlfA80g98l/fCAzNvc2+6hW9fWZ8vTuCHkwf8
4eTLLZnCTQ/xsR6bW3tWz62NVICWmdCAp2nj16FA+LHfZx5g81HR0nou0c/XxT/sGe5HO+27JVxN
23PLuv0G0aaQnkehVCk6BGuf89dcXfTEM7JNZkavO3fpq+RDhuanFHsu4mv5u/Jk9KMLXlHRrO6q
KfQ1zDSFrdD7pXgaIN1k2G7dNWMsn4dZjeaLMqId2o8ltleNt+hMPU0TUUAvGgCpPVDknk8gDIrn
v3nTA+K9GXftoEIhsB9bWYCjwX1URj84+zwvakrFegf1l+7li1ifjiErBKq7x1WAmOWDdiwQFlcU
wxExxU0ZN4S1mPtqyJtxpmZb0KONVcL0fw5w8dKGHg9gHAUrtIwu7NR9wFxzIpZWCMNc4C4pvwUa
Z6zOnzP3TVvEnmv5WSiFXRTdr1ZCeDg9QX5uTiMfPCPDb+4/H+YuDHN5oGulmqNTzxJzEyr978WC
Qybephqnt57T1J56ulY6BH3QUF3eLfUHI/A8UB3ZztV+wZC/eR6AnVgXeVv5yS5VNRDv01amYEvq
zw5GCAicfTAw9gmkHC5LoXA3CH/Sq1DxmEjOOYKKSM3qHvy7ji0j4c1GQJ2c5JrJLSSZRZQtrdFi
vTnVrTiXIh1wbYH03adlQuscRXFDFHusMkcI1xM7QTnLA6w1MHSPLT1BeI7BlA+fQzmljmjTe+Ef
Zn09eBD9tE4kZkkbXmoCa4wZiYASW8NYxn57xK4AIfj9OaTH50RTV5GiWHT4TXKSrEEcBqYxRmjO
zAMLH9CIOr5tAdfCRGRDZSnoDpZfYxx+CEGzVnIIFtYtCSavkP55vDQqFtaqcsdoTg0055usWwwG
JFBByHCKHR5CXvslSrK1I58u/fd74POTTnRAGIlXSzmEwEYjdbfUJKubjHaFG1f+kkbK+9gZSr/a
OihaT9sQVaC/sHr9PT2/LJL3jwl5S2FBxowFdrAd4r4SkRmPDUUKQPs2xVKQerPnBVO3mopz2Ttg
qBBHEYvPKqzbrsQIGvYXs301jVoUJcKVXkYSj5ox/JhrSxK+Rz9IeOJBlhhRBBMYt3WXgfS/pjMm
sZ6PZvQwEoCMRn06dIBIkJ/97mX5mrRl7zltKZ8pm8ALzBJZyAA02U40OBuBrRDRlZD31xdi/LZ6
CuFPNA6T8ZD442koBSerB6c2M76Cwi82QrXSLXdB/Lh9JBSTNIianvomN+A9KgXwidtl5Oi+7u+0
TkFju7GbbRw6K8UjMt/pdZL0O2GRzxw4Pco7l0ECaf5/vpLt9xwHopeWxQsgAntfhR9CbeYJEooW
mSePVuIAnSWeTkBQ6PyljixRR1GXFl4KlLOB8e8dJkQm0j+ZU27WGA+dRSKwsCB83NO0lPlvgcLP
ldwca44aDOK7ozx1gd13kyXjE+SsCjafIXJ+JW5aCz8HPbiakqM103DmUSkXmCiEc3xTyiDPywlh
J9uZ6qXvRDOUYksGgphfJFX2jzqDC4z+mwQcR5KxY8r+o8aFGJyCYAlRL5KiT0yWcEtslGNtoQ8T
BDQKocQZ+DBe20YcSPOLZBXtjbcTM9Khvslf7AS5TKI8wJe33flGEbN1RUBVGqu4Gs4mXr5dObvz
xWAu6gC54dBFI43TGPMqodkkXWWwYe+ebWcqPgJkED6I9XV+/4pE8ZXI/dDOsW2Dy3PFdLFKau9p
1s2ecWsKarf8BIh2YCsWN1rF5zgbB05nOFe8WElGewKBlKYjdDwfZ63KTcbKjcYYQwGNd6NZf8e4
siaElSgNCGoZY/+Gh9x2WYAxpVMmDUxN9vWeSes0ol9qw21i71AHHxsvAnyz4dGhn4lAryR6DFD2
sORgV7evdTYvgOvLuFVJlG0ft6ZaFuYbUmeR1d72bGOE7nt66SKR3tL9ik66N6ifG8CDoDFMUEGf
8Md4SV2H6p21tLa/KzYl3JnNQNPeL9kwm97ilVkho5+vDtVaFd1jGkGpoov6z5URQkldjdq2Zk/C
U1+8Ih7CnBVee34o7cNTO74GG1cBcvJ4UeAZeOtIRkFzmkhTozHzeQ3U1d9Vh/Xs/sxiQeD3JZ03
6HAtYj/MzqPmJUAWXzpP7nmKwBZsNfYQWlXPnYInDWf+RHfifH/+TB8MSnGJSkI8uOAjhkMgfVlt
doA46TR1tZN/sn5kQz0HiVuPsKIbrNkI/JM+EhU/kkZ6ge5t9emzKH0x8WIjzjN6fmy2f676bCpn
5sr927PdhceqJBmFABqh4sOk5a0wOxXkTnS11rqDE34BZzdOIpmuKLx6RKCUehKHZhsfpqjkf/F+
og5H+ePgsq92say5K8e868Jt7sO20MuLufg2Co+YbCLxgrHdOVlKyzmYW3EIrSaKuBsidRY7IWOO
boE0Gv7f9dWJe7nRvnH5QyVQ213gQhiObJf1KsmXpvmtJpIzoCG94dIbJysRH1hUjanZpPEJ2rPu
GZTO2n9JuNvzpEIL+hHJveGCYCE+6WVyEA9EN4dokGPtewHf8Bhm3yoehsT0cL35yogf0cDJVTqL
ID381gYbBSAesJKr1gJlZ9+TZTlBLC22ZZ3HvrKW5GpTB0X3dPw1rxUV3gOKpb4f3I5BcgOFnO0d
vERuyGKQe2JoVC9AmSDyR8yGg6m/ToSsftinxRXg1JVTfBMqsu5KFSWhrNzpkDQc2+HjS7EFRBsv
8QetYNxpO3MD2b1SgGsRvtHdof1waCv+XLZPrHJsEctXiZCBnYSNOwOAngGUf+lOMHX2YJx0h9Oa
Pk+f+7FmZwEhMbZ7PlYvz65iQGfvlkm5d97oHC1YZqZOJAp5VxPI1mlRDbyAFWwBkgOtTDyWILf4
IUILa4Y1hPjp67oAsPkkCgNpAoVK1EUntQ7E4wAr5aRHoI3rlwDhLYMZe/alQ2UEWQRrpLLlCJgI
ygM+HojowtnSj+gZ7Iir15sU8upU796/Tfr0fnpWeUIAf6RfMJmF65bWEB54A6FYfH9STdkU1zH5
iTayGhjOpzXC09xpOkb8369Z6jAeoCXS5zfm8VJOGVDTYq+eeLeMnwmsuj7wLkpyjhYcTGlHiPHb
N20AG9Ini2e0rzne9UR3g0isyFb0pP0YNQwjGGXWfsihuQDhNPRnEUY0Pa6SqWM+hL9CJwN9lkYw
v9lu+epuira76uIADGHDQCXhRbHC8jauRpDzoLymIF25XdIEtnee6pa0UD1hFahLnbwxDOwprwpz
12Pnou66PT8UCtQ4pXPrDmZwHL5ExTpUlqGsVnY2kJi9cxhD0zl7ucOzev1j+fKHCi2/EYPhW4dS
05fcXvC1VnOCXurl90tLLNqx0w/XBuQZ+5FFgP8Y/W0Er8C5JPm6grDRSsx9IHo78hLaJSlexr33
nQhEYA5Qra6VGjKAbh20sKZLDa27BKNfcOh7/X/S89fSuFhSydoc46nAVnwV8ppSQe5/OwgR4vY2
hJUY4PR2ZROigtnj79EyA5/FWtVmdRaYX63lLvaIX/BUVhC+C6LnWKhIbW9tOCCvBhogEEvE8biR
dulgKn6I7Go+wmJkyOKvZZPmy299E+h4D/ymhpy/7rfCH2xAmqUKbSPzDP/LgFBP3zRYj1hVP7jH
c2zbFeWBNVIOmcjkJmZEO5EVIwSq5Fbmhrh0LLu0KXnkv7/qCGNUHdVe8eoUfJoXI8JdWJNNQrMH
mlHq2CuZBMgsSVW9Me2+eHwASH2TwFO9QIYGgsr+Zc/4JCEQxXp1BWXa+REgZb4h0qFFNZGSSKVU
JTEduN9RP6MLb3tAeH+smosF5B19Dg1VvYz8zDVwJjk/iMw4cTTWOx29H/3xH4DMiJwpA4EtWoN/
i6t8f2IGVgtKPwhJb2/BwoTEurS7pKyvfoz4iM9+vD/vecFeL/TCDhbvA1VbvoiFL7qmqGIS9lcm
BaQXkfuo9w4InAtRKYWMx6KOaEA7yjSTyheT/+Pji3Wi8bOAjuw9OU6c4Rj518/lrUXJa9aCtTHn
oXwCfJHB6zJGIGfM5wpy3W8ZELFTgtPmuIzg653lMc3mouCeYgp/3k3moRom8Kf9b6HXpYU0IgJx
sSecFTomSkUkdpeefqOVIPBa8rsfoF/GMWiWH5NulOChTLl7E1YJEpM3RD+y0C9EiJaY4x3UzGuC
Kes7NmoNAEiO/hKaR+kZ8LG+Ce+1XlOhWmygpwG/0ES/qtRDjt810r6hVR/1HXNsM+o60d3CxjDJ
ygp/trHJonHlZ7oeG8ulG8vcc7YqFQissz3mlXgBeNH7WYqA+PW1QPwM4HDSXTN/2w0OvDpaplyW
mGCOG/IocM1OceXcF2zXYA6PtnBQ/Bf1WvLkYmIUxzQPxQ9wypLxpk1d2jHqqNofBOhDFYTA3m3c
Lj4xcgZVmvAD22WSeMDCrV0n1f1bb0asX6UDuh//NNQHQ+krBnR9H9kucqQr6/E0OJzvHgVtzg1S
++Zqz3EGClGU4PkwbBUaubZemvGueIfFtClT0O6xhpm/JEKe0q5z+YjfkPWgN+4Qv0XdpKCuWhp5
eiE9ZwJEQ7w9kt2ahKCzAlarUwA+wjyf54ElD/aIqMjXQDqqHBoQ/eG+AmCxQ6jWPpw4UFFuHpgV
inbuzBCAFtgw59meOKGi+zmPMgGn87Cr31Pb9LZ9WTVyTyuAvaPqPphihQ4bk4nT6zOUPhoIDBn+
SL09KLIJK/8uiIoVyXXyWSYa0lIFhysSdrtbiozIQgeq8a8ta2oIXrUpJThUIYzDsspwikpUcHJp
2YCYmNCmsgY2dX2hJ3Z02G+Ou/Rw8LarP5bfGuUvitu88atR5IeSdoHbJwVEctfqlJ6OkZTMmh+v
qQHb5mE2lrLk+ilxpC71UxTzfr9oBxAl5AJJjOXV2PX6pQ0gyG/JqLeN2/Owct+Q8KKFqohYOgI/
5w57rqQr3tlJyc3zTu5VG9qbXC2uqPQX9/VpN54Ch2IRi0v+xiIO4VZa1PeNurn4C2ivPW2M6GNv
LJ3OD18znhah4Gr/cCE+YhsbbjP4Jxj6tdLg/mf0ehy6fA4T2zSO8/naU3cXYG9vfb16G0LDTrL7
8lxSep85yuI5Ak5er0GZF8FuEEYR/T02BOfeffH2+LElL4N/2b5EN8gBQ830YXuDd3N4cg3I7iGK
wNBP6I5D3kc6OIj8PIdmQIflyuAcp0cylmHkEr9ZWpSTI8nUS5SxFxAnkIffofZV6oyIDGnsIyWk
VfMzvPreD2W4DJ9I4asvriwRjkRFwMX2efBgiiUwHIjAIcN5lYW6ZXi5r9d/nWum2GiTJ2qVBzbS
FS5t4ygS3fXA3EUh49KswHUjc5hMFLD2nXzGSHF+lQYhvoRcECeo+zc9opd51EoJlh3GlmmiVw+V
+MNTsVEIXXR/B+uaPNqvEVEpFAxDB8+24ax0urs2uYWdfgxRE40a7e/n/aokVh+FapnTqzYo76FH
47Zh9yf13G0M2GvxDrbxbbPOw8LRSjDYXoioXwUdjLTAbuJDKkw+tuOBsp7h6Ha2sRRQWk2ayahw
GDFsCytWww1NswRHpS+vng/R38M/DQEJkAuGzu0SXtwPoqtb+U7wshClALcsT7nT/30+rcCCXpUb
zDZTfd3dFVdnyHn8vyDVAeVicy8RMS1LorIB6UdKZYdQw952GPWlYOviCfNrHhgcQcHyDqD/kQSR
mdb7XLcFDVXZAqNF80OWBE/d7hXX4kQcugmu1+0nICCVx3a1u7WUkP6/UcbZMyeJmyzmO/HBFJn/
qwS8GbuVk3BRJLnEupOFzZIXeFshX8tx4UgIWgmEa52vBdojJAdfwrkGAYr5Nr0d/b0QeiwdK+Zi
eWWWW+oO3VL2jlifv819eN6nYbv71N6+T8tXrHbv2kNoZa3s4hCaXfWiAQBAO0M8cFVgOQRHfJLF
c22WBb9CqSCfAzz3YOYH3xvIifFsdtzYqwgGKUMq1V67fQkEbzlhJiAgF8AwECkGujwDNLyAIjhP
8sIETS9r3CfoljILrYSnf0Nts/5c+5u53goMlp2m9lEklchaFa2sKdDvwksIJqYYDu/XSEUeBziP
7jTraMVRn+IVLzxpyJcZ5YJCVt/Wx5JYKOXaz2CWAhAiG3t4vF+nmPKn14xnBvMb5Ngn51bSrhcT
kuhlsj/qLrmsf8A3jPXN9K0br8m14aZkdNoUodgkU3Z5mNDVEOVuLh6y6kg5a9xexN8Yu5YuVqQC
CTZZN/8QDVoDCwkB8yhrFytP2s8/PHLIjQ8qw4xT6/+GwNhjNzUYBteU5iF33vm3dV+JSVB5K/C7
496Mrd28OUefpxx7YR4UrjhhSmrbbpkhCH5h2ShXWv62uVdL+9r/MjWAptvnLhYXW/OGqDlX6xmz
E8khaSBCDKjWoF2ghmTXJsHPw8mzTbhK5mAM51EIOHNsDlcKp7A4zNohX3I56XXbELN6egyVlCaS
y8fen1U52qiz6vDfM8IU+o7zKXts/20jJ+ey3iYQ511O6jTAK/FMT8wVd+u7TG1wq20Kz1ecHXEj
yh0E7RJz+guQc1q1FEyAePkPhyWaHNfS5jQfDrewfjfsnq2wDtzP1jBXWyyOovnphhgV2K5HJwTn
1Kn1ZariPF/MGhrSXvIjQKGf6icXvb57Get3NtrlymxdrU6TpIYC8fJlgIGzhZKjAvqnkYJ9AOqM
3EoCYbNgJmsE0ZIKXkz5AwnsxqfwMa4gR1g8T+kdvJgroOqNa3dQDvBOSo4561q6mNJL9ILn0dFa
lgLwEaGoBWuBeUuMoJDx8WzjQW79mKPLb+Ql/F5hPC8nUWvsdNWUrcKDKCgU99Q1B1jWvl7+e/PB
jt/SW+TGzuV6g411XKatF7ti5rxgh9OSNinaU0MRz1iQsnOMIOAhKZWTJpHdxEqd+lpxScFQl5DO
QI2MlGnbTCLQgcEqmUIZmMmwqEf0JB8hDBdcSyb8Z1cKjeRob4tq0PpZpugCX85yOA8sI0bv9TrM
JETXN34Kc95izIGDxD2sNcVmUFXgoREPJIvJziHvm6+KtifgrsE0ISEZXAzFdOQTMff7KeaY0lEA
+pXhDInptGRZCN3M1tgmDCiHLuSiB2b6h/00WfBeYWpHw8BujzToQL+we7KSloHVex2eIJVRVd+v
7dVnV+yJ48mPcBOIujDatUkwgO38XN4eXxCoJoAbWMszmwmdrcHwW58/xj6VFzCLlamI+NhP/MFr
6rql/qB/IErK63yv4RigrNCj6hy5WJmDCUc2HzuFEDLC+dJPCgx1jMESjGPGjpq6z1l4hHNZd5b7
mFawlMrWhnqL0K0Rh8E+zl7NpxHMqFTzA+jBABLyzseNoT2I8Qi0CLn1rVf8RQQch4+KwPfKQl3r
HGLV7FCUkhIAo0t57BsGKxuDh/jLefrM30EKEcSGrKMJmP0ujIukd3gOZlO/jADZhLB1ExZTsUyv
wiaDnIY4rjpL/FQzr8BoLUImB4KAB6xFSuqMK1skEuKWBsU9qL6pLKseVKW/g+tB/kbzmUZ0N8as
VWXrE16A0sz/yHnzKCcm9lX4FF2x61GF3mL0Pb83b6U19huPJm/9WMd4aZr5Ad7JmfKDFEuKPRnN
OpUTPN0gwz6Yl/XwTCbkwlx7msG9mN/f6UXBfjyqTDsX4/zIHDsftshlmxaJMNV2X2v2nmoPg9/v
/KIx7NQjgXn7n9CeEtVSRlDVz2QLkQdjv00yAo9v+ZoeuUkmHnXx3jveL6rs3Ann9E2+WBVRDmmI
9cq1lnSrY3qdKbN+tesKtmAxmNPN7S5uISzy0FZodxwbdw7+dbHngGwulJTcJepgjMZ40bQW3rTp
Tt5M+U9zDNPCOdClHGF6cfydBwu6yCnG4IFSVGVp0viHme/zt1HD2fOyK/pb+/2bJ7wc0xOeeyon
nuJGvKIGH+qvM7tpv6gBEuZYxIrIU1Un3BWWGKxMnolGCSiHizxpVGnA0vsBFPO1JrPm0fw0EiCo
xeef2flAv3T21zdyZ8T411t2DN9SaugleRafW3wbbdk9P54LTVntliKjbKNYldrL5Zc5V5IM2Buo
QaqKT6ErKpErb0wqJa0BBgRXJuU7kjPYjC9BO4ZodN9xVYuhZuhc+AtVAjhzN3XH1xHkcyVGmOnt
k7O071isbif9kEXUm7iDxMCU/udr78uGOOG/o37c8vP8m/hKmJhv/I5n4vN2aSxcqSf5xmuJYj9i
CsEZxDQa9aFU2g8O0Hw8mByU0oVpd9dyEzNXD4FTMqPoyqCC6yO4FaOPEy+wApEnfIw+JjWGOYI9
WVdbMpkx9cTtwKzePQbOQM63QNqPGEHlI4oBnyvM2TECYjbD5o+iH89mkrPo8pcfPbFReNaikTda
VIBmjjWs62F1TqowgFSWSOS4PMoHSka4jH4r59cdCKC9qr32EQUSsfwx4NY4z8UPiCHtpm1m02q3
mOAk+xTwjsiTgZwNI3yfQRaWfAPtPhyMCCNC1ofA6F2xPCVG4ziAz+6VUd+KJPs6K4ZsswGA7mkj
1S9fLwgsZqoLHAjr3ohVjR8Q7+K00rQM2iME12tWbHgm2qPrk1Cqeiu9Zu8zA5Reaby0GgebYP9+
TkxYoysrdo4K4mGYG3RwBEbjNFtZEiv55rhCi16G6Kjwpk2Lni6xA1YHZ6zAZCsHUw+ZIvEoFJzg
+RH/oVBwzaVVKDKmf4RpktlLo74bhDhM96pZRl54kuoz8hkAbOw9FsWf/ztcLVtKDdz4nMAiK+LV
iiF5ubRv4kVeGlHhuY8bSHL02Evp0C2Q7S/4PG5YdC6tAJjJgGacgvl5113obMdiQKdtrY2pH/xA
iL83DKUypFQKz2zUS2Hv7M3dgfcUdMw/EH+vjgblgM3KpeGuwZPnwO/Z0cWQJugjwmgXMTZc9UOE
G/9Soem6oc1bk8lBrDmZhk3FEvs2KeQ/iwPx21lJV2rD7tNnQHRv6k2VSSeCaPO9YpgRG0aJsvNh
ttLxyWN49PJCYHyaeQrD5Z78qbZIzpslrH1p84EVSxzB3elqenSz7V/6eo4Qq4hZRdG/JwDC5sjN
XlxellvCGbhWOTfAOcPH83K4iDtDOtNQVLQFaFFG4W6mmNOylFEurEDosAxMx4Lvd/vv0E245Sqo
Td50Sn+/OX4ZfGpa9+b0nrpy8pir17BxgUoKQUpwcUgUZAfsTK7gWiB32ZsmltRRSqhlrCXjj3UU
dXuMAERGS36sQDADy23th+YTKAHx2fSc8puQ5Cv/kuui6QeEeYbqRtt+JSEWaHBw0aH14IcyiBKb
JO0XFhDRLwM1K2tr0+1s+z4011ESIvTAJjqUgezS6pLOcc/7EOiA3trRmm53z2qYltUjIBD/P1Jf
wMnhtdKh448dQnvKtiieWwaHvBB1BzjVTTqQntufGB/mO5dmw8nBWa6xP/dVYi82/FjJc4ntvFqV
qUgwbkd/342PvNaB6OItUdhJsZHQCHmbWqR/jpJv5P9XqHWmTd5+R6IEqYwV8/KkIJ7W7efLMLmg
Mekq4PEL7pFfoW5fZGxggti5U3GH1dvgwsWKDzP3qKDGzfEsWLZd9d+IL+gTVFdkIGYHbddtkoQ4
qsvMiAH5S164CqaWnzyZ1Y06LyF2Gi3z8/f1wJr+oRfK8eA1biN1Ft+ksROscuJPCAkv9dSljv50
FrpDxd+CuSXyv1P+hLIhyQOaV7FU7txZF79YXYSD8o+t4N3yE6nNTS5oHeBP+yHQk/KPo/TPrvcS
dFewJs26qE1LUcI5lwiwNx42ISRoMZ2tzdvSx5Cuyq2tCqrWGOmV0vka/I0rI1IWp4BzH4S12mMW
vm2oh1mHCeJnlxRPj/Z7TsECA4jTQmNq9NBXXrm143swGoeYwT366rYetrrtcyW/5wpZE5lXYdvP
sGS7QJky0hVsJzBP/WtFgTbnM4zWYwspCUMeCI2j/esBPGOiR2tCnQ1Me5ZtK5hQiwL6I6IpQrS6
xUzTz51HIq/d18UaTt54vuo1lihQs+C79+HDKUYFSSOYZ/SVqsH0PFDkV/wzongdWkl7HZd8ehus
w5UMXFa2qaoI/rxc0J2F/5uIgtg0o1NoWjfd5DzHoZIZkkqKgOXk9UHZT6NamXP23VauKFwXTwTj
KdBOiHmj5+Di81AaRkvcBv70LVVCL3M5vMvvuIV7gIYb6Mvscp0sb5efiu4lbCuIXCJKPVB8RTxT
t5WtBcZpHuxMZdcg6K9GiwqzBpjGJelU0Mkf75x14wGIdqmeQIlUhu0l9+ioNUwjObQmeQrAo4A5
eC3ljrrxakSr0XsE3VoYbJWZ6mx8VhhDUYx3yxkloAw88PNdXJefWk03eemEbCHYvVmRt8OJEQeR
a/PL/9wnVbXEI6q9eIyisHzJZBUkTfqL5XCD+XRQE+DX4vkUfO6sovBvC5qE7wSZG19eJ9PVvL4o
T5QrPchM3lkpmnBnFyPwGtQDgW8XZsSKYcBFc1a1Ogux2yIndvV+lYT9HlZNl6ttbLT+b5Ew3Z26
90VtJOxFoAscfAP8sVAKTU3UbhBXiGokj9lAzNt7YFHmu4huuz1PxP8sKZFq4+QKui4wuHUpcuMq
I5zx808KGUJS0ItZrnENdvFnYzPObmr9TEFQe+sOAN++3Ubj9r7V5Gz6AZxnbnSARkFdYxwK0m99
QdOOP+bqw2lh1MnjmwrtT6gaOKJBwAS7LMX49NgFf0kFlePyt1lTfwVNVCwdrat1x4ngvaM/BP2a
JvBLs/69Z5VoT6Njsq5q+OFRxuaZVNEo96RUwaltxGmtST2CvH2WyXNlHauN2dAka/cOQVdxiwHC
I5m9hKW33gpdEYFexLX5pwThLhtljl8Uv3/7E4yhjrXegtdp7q5KXZjxeitJiJmyAIpqud6ZqCnD
N0drnsMINS+zv+91C1kZiAQpgv5qMlTjBe4MKbiGLRemYt1vYAFdzyEe8STqqdt6Bl2NQgtQZjS3
Yk86EyH17mCrDnOfV/ye+nShyZCZhvTu9ZIGVplsfSuA2vmzdRh+f/9DSk9P52xmcTDe15ViZWU8
FtQt48PXupjGeUbj79P/xXKPjuVoti4p9wxkXElj89U6N7NPTQX36BkSPeS4aRK4UjkaXE6iX0w1
C3u9y3mKVUsg5mKic0XURlib/X+p53arV/NpAjGr7AwkBOxzRkASgP3ER+UBekKGaTT1WownuC4n
aM5Zg49oA+ZyzScUTJcGIHr+rRREBc7aoa3+watiAp9Qi2R0vmp4Mhla390w/TulZ/wKARjRz1VD
xLC2zsBoyPANlzBldi5+M/fMK4I1eU39qWgrNTug68NsliGgBM72pmEMY1jAR2eA75T8JtxQiYVB
n/vq1lKvWJ42HKrpJYakx/64+3RzEP/QIBgu4Rv1aMGv7m8rqN6CGCmV9LsNelmPOu/1sIJw6FNw
hENquq3PjiSVm9rFRZzSyeKJovGM4uint/kckr1Yc5SRxUIZUa9cHqDQTDvNiuCre+imWLRuh+85
vRIcID7Er8uTyH1nc/wIlhHUYpYHFzmos8VDMnz3acAHYu3m6Q2sUTjrvgeuG2iL9GhjvVun0ekO
SHSnY9OjIkp93U+6f6OwNMPgx2CxH2ok8KY0A5TzjYDOP2NomRcjM8Ovzi7640A8K31/KiKoUTzA
5f4ri8v+QALtXy0txkpYLtmVJiBKtKfs7fPkIsxyIjzGrYF03fsizUmTdAhf9pkfx9HqgQfNyXe2
XE3tLXxAvlxUUJnV6Rx+yGeLIfN2FV6H92RJOFyAGDgjiGhZkTC5Ug5eOTE5JtK64KLIoDuTGiKS
xwp3ffyD0bDezlMc2vQ0/HvCnNqiGzcioKXgmk2IOLKoVIuq82vzef3taxKbNJ93F3GNoNgzMAyk
Et2Q2UN+hNpNfEXzScITcPZcy0jOHS5J7tH3m0iXNgPGt34QsgZuuePAgLJX0pF5FxicSCLl5Wxx
2m74+Vsees59v8USlwppCDcR86fG5tOgRsd79zEcyY1KhVprGLEXK9xzk0iorZWrU29odkY03qQK
GHvgL9wO5VhNH65ELgeEKXBNGu3xBK9F4sOfFLl4K089y2gmiNKsABqfO1Ml+NNdcOfOg/pSniqg
c+Cg0JShDuFBZYfnpfD8n2FT1SbOGo0+pQAZYflk51/TlG9HVYbFil+JRIKF2j6GlQ8EoLnFi98S
mvPoZYuxGs7mKTaOxLpC3uyz6k2T573ZC5gJV2SRHiAq1HxkLJ83IYVlAnoNPZkUuL7jXtnAbyso
mfoXN57MyHDAdHLTopWE/NYZpCYyew4k5quL2/c80smszabap0U28dLxUrx2djHofi9P7TjfQb6F
Zelt61XlvYGwbd1QhMq/vp9tmunHKeYVLkjiEFgpY5p5PSc8YukPDsRmET+MTpkrATA/prAMPgO8
yXh/5AwF5pCue1UHuo0vUEx2wiBxU+7xHeC01TOMUTWp5WFOVGfmkyFXEOBzVBfSebLPwDiyqvne
zF0IHus6u1Qc/tRYJ0c/uydvmywsRW8TcgTOagALif4bmTilk/TF7gk/q/Gh4DkUJqGQK9teLj5I
GbX9dCVyoXXlcZvge8vftgUT9X6XALi54i0i2HjGPQ80BuGjWiJQMtPbDbTzpqrxmKKHtsVDa0Qu
0eDk5X78hHnRzRImqurh8xdz1g2r1uQuLi4JcYr77nz5yopWBfYmyN0RF50vM3OFwRW046qMOKL3
BZ0gmvuq6qklVmhGr0L0VHeUkAOx4WPvEn0X+nHBHcj7KN3fv+UwaKFE3qBTFtSwy41vIiNTZBlo
h0R65ir16wNl/pqqpOYxrO0CEMT2VYC+yOp4FObn74kFRZgbcKtC9oFSfm4G2NJ77s1+swXm3/WJ
43A2Gm3RkIHoTI15jCt7JHEZHNaENhTocEbuEGYloVniYBEJYjX9uUBTk5K03DpLh2TtJ6/vpVWM
iY6nKvOlQPq94Luhj2q4ATZ8cLPoeOjtCK7sPaYzUeA3exDGz5yTEajI2OztlZHyj8lygvktCEtz
QAmc+/gsDSxbxTFzB9/trqs/BY3z430x0Pigrj4mFGfZTqXnoXvhijcsuzKUuknHjnIRe0mPEvt1
0O6PVBv+p1hgiWXT/kEdWYBLQuez47jR9Ub9VbPopleSfGhp6ZJscA1iYat4/uOieGG6LuV2PjLc
dx8eNH+VgsI6pu+90Qyv+L/dMqSd7sA0SPk+ifD65EO1Jrz8ONU+Sw9usJ+Bw0ZLvmu3DhWGzXxu
q2r6TpVZ2IEXBxevcmD/lTB7RRS6Z0FmqkB4YybL+mhBZ9XIBtxMRqJ42gVmNQyqhWbNUem78HcI
EXiRBZOg6tJvnZdEpfbCok2mwaknCOWWvbumehqSV3f0Y+5oeeEOPyBcczc+6dmU1iyWpEDEX5LO
uqgBppT2CDAOXXUesxpKHsIiL6gBK7a0jMha3V/wjcTn905kWh03CAWclYNcmAcTax0mScY6qIkN
xWlda3kuLgsPPlUx0QMXMeC2DtgLqx6u1FGA+C9xWIXp2ZuYEr50gwcjfSNZUk7OFKHAdlYp7P1Z
FtzBZwERp28B5WZlcOPs5+uSQ4oXukYzLPLU3LGhWIpx4rh/1XKGe+9MJ9xybiYEV0k1THVk/cA5
Spp1mF++C0jB+a34L3MOeLJvSeqQqlgFIshUSSQ2XBAOyIUEx9vm966SdLpDr2lN4e3Nckmc+yKo
AzEQzJUEP4G7ZXDGcTEJgozB2MDlZe8Gcw9wl4tnvWSMbh/nXZtUqSktnjkGbB4EpHv1ZHJEsaqD
8KBVwoIfZdcp+51JBMtUBtjx/KGyKPk2CdR6njptca6GWwarc6j9KUlOkn+8z7pN8++BFLyZO7bp
35TiHT7LKWk8CFNCZtiqdOExkZtR2uP/GrZ53aC2GT9+YlCjUeSEvaCezL5/8xVzhECzo3oqzUUT
UgK8P2XXhhAug3POTK3RL07Iv/B2V3nAXCOKQ5lZq9dCGXdYnlodMhCj8JToZ/BSqhBXG2FlOyzS
qMTVvDItchzvYz0dHtWnT57x48mqJDajjC+zsSDnAyv6nCDpna0bXiRhVPP7P62nMH/TzMPXJKrY
E1vuWXu1RIC1TbParUAuMbDOQCJDD6EQeEb1bPjktr9E2TUyEUn1oRUQbdJzDCypO0EvP6otTELi
vvysCp9K5XDQb29TXdQd+2CSvvF/7Ye2xjN1R6w321Fk7aHzO11B4AlN++OpdGYRDWZ9GyrfVBaY
NjtIKHSk9K8WFeIJEQRI40U9/GcUgplCBYwlZ+zWOILooh54zMaJSQOrAiQx7lLcVaPbqhhlC0St
tK/v5Z4sNc46HDaiZrFefaVX06VyPtGR7xYkGqRGxPr+QjPBbPr4kO+Oi8exzSSU6U3sYZxspBQL
NQP2+q2U8323LrNZxvPDd2XNhIr1pL4bIDXE6kA30yYPOe/ifaYkkkvWoDFDU1ZUYIw3KVE42e03
W7pfa0smG19deP3tmx3EQMnB2+4T4uVcCoR6rpXWachYO4vz88WFtPguc4stUAYlAqvFndSXU/71
jbImR0JUifZv8WsMFSahQ3InObQr10rNZFEWzRRi2C8CuwEKLm5aZyK0JTqwuPM0lNrsNzN5YTuP
KPI3TPmw284Zzgv711/u44hkWK01DKQ/8hAwps7bIpaE6jqqGtdMSCoVrX2zCacmZpQv0JuqMlle
YugaNZPzCWqDkZeCVZ1puemMQOflQj0eJ2uqdcIDJg3z/aKfO95A3DemB/ILTemQv8nbaCkUNEt4
ui8GXVQvGuBm9Y6oPiC41MbCD6HH6b/4U150A/Ve4vUK/s45fs5PEXY7nNu3hb1QfS/LxK2foAro
75A4a/1KzmUo+eRJpfBYYDlfHpnXYhl6jNzF6MMaYbHSJ1TcHsdAGPzTAUG10xgJSKTc0S+Ug0Sf
ZnbBnk7+WDa9qK1pam0Lzgu8G7RJujKDf8a8b6FaJEECd41GpYfqJH3jnDnqNNu4UScoWLJ1yX91
hcz4hv14/W2aI4CP8Jr8fxkbocCrzSDcFb1IYnwGiyVtSeQ6FrO991at4PSaUOpshyd99M6HL8We
uMIkirtCasPLMUJ2BBxp3zoDfd6VsD0GvXZ9t+LE6OQok2a5OS5s4md7yzv4laFfuTLGKZSLFLKH
PcRxtXD/BkTwGpkDPZiZkFhSub/kFOPHs2q6jjNwIurfoN5g2tMQZnmeicCQHmnINiHXQycHYIPI
c+AJIdcsV0m74Ld6XsYANu0Pvpwv+7nZzZSoHBmlzZkEcJjw25lbMdTC2mc4vbeiSE0W07+4kcNg
T5oDUx8RzIsDzKLBYFVrNOtaZ1wzc2+AiHzkpoMAc8vCFd5h8ZphHsors9lCFlMorJcW/ebRATXi
m44n5u/uelxEx6A8bAI6yfqr24U5Nh8oREEBeFiuMVTlwdHR41QLQ1yHztW/ie7FyuXAgYE8t7BZ
5EGJgP0hilvTCb6TEtBBlYpGSOYs6uYPu+4p44/QoEKpW73vZM+bMCxx2/fYtWFn9oDpY1nIz9D+
Bv+ZKZGb4S4EU3L6pPLOR+IiLY/Q8oouXP6kjdSU5C+0JEy3ra+EmGYZoobbTUG81x+eWCKvA5En
Y0zfbCbMZg4lPmX2/z2TmQ6Nr0VuI5edJQgJtZAlSXyFZXdmhLITt4y1eYET98R61sckmEQ8udAx
iAeJoW8c7TZxoIHB+RuInWXS3xwrnLLIaiYe3JZop9tvpg0NxbYgw0rTykUZe0wof8UMcG0cVkL+
EnPPRQifAoQonatZC2uaGCDRKPU5VJUgvsXL00dsKv/pEP/8vU7e+vS0lJwbEqZ67gcv5E6qQBzN
gfyTbr4Y2dUo3jn2ciB9kZM7/DPsVW3jgw6SxBNvsp3sgwE9+9K8bBhE/reIq0zMvXP3D14DMguC
E5JNFryJxcVx3y/uEVbc0WfUCCFTMjE2C6wEPrmK76KW6Xl5lrs9pi7jqvu1ps/ym7ikx9Am2UfW
DIoEzheJ/ELW99me/av7s8ZpqJ/kjW1O8s8ZCzr9C7aSn6zn6/8kTIJ50UZxZ+E1PKbSI97aR/Jz
87luj36bKhTZ5WeHTibXovAj5W2WR7sA19VGHftUTIIfCuVAMrCxpfaBjE/uW4oQL/OM6tQ7daV+
cLuOCfeW/knDsypRFU0PxfpD2t2PJqZNbSiLAO1O9KEQyV+pvhSWZt4WGtPuK99pm+dI1fdAedxx
DWwZUhmHwaN+93doy09jD2FHeezPgwqEfA29rvTbvNOaS+UCGy6osRbqAstj0vlwbCTjzFKjQlvU
sLReR3dQU0VD2PYAfrHR5uwj39OJFIKgarvisH6ZuYmtWE+FaQGBhDUq1qSOm2J6DjJ7WEZ99KiI
kxQJt+IHOISmIQNXuSNMP75ruAuJIkfPIaFACfILi89vlR48sf4ogyOuDn806zd0NhOFcJED+ugs
n9daYZcH0e9IN4+zKJj2eFHGvTdVTZRVVRI1AB1gnx1Zf0uMyP+qdH08eTa8XvwF3wLipS25wSc1
QTvlJPl+RISvS3apgZTQFgZGrLcEdJBnQYa0gttxyvVRqZhrjFFiKHr20JI3GjunRb9lb3io8qUb
YmDGpOPGdVRLI6PI2sPaYSquGeHqIgLtFrkUg+I///AzhqrgHQKYPxeCWh4TsI4+yBpO40e+hw7i
wL0iX6I0R4HT6S3wRN8sU3wXMQdFRGNQwXI0f1A8fh3dV4eYp2qE8F/3IELcBLgFa5eUi7VrE+x/
YOWzQA3DIzQl5nO5qfprat5sOG0W6ylf7APycfEJurpgXJTVCcxieeo550qhZDxB4Fc7JwfTX0kC
ffe/z3OfxhSbSIBTT0XIMgfoT94GdCPYUovHkyqdHZIp1XBb+XIjNEojRGcksnDmpS9cf8r6qqyd
4BYPx8Yhg3jOKOn3CyABXduXc+zYgG18cxbeI5Q2eLDoSCtGSO2JGot5f/IGL/C/61vlysBFuGsY
wQqn2039lv2ExfhK0hngmuAMSvwJwkddQKwOxAGQqzTGAn6AEIMYaOgcgeHVCxB3MDx8cTIc+HGS
u/rFjvAzKdOOUsIHVMWXR9VOv1fxR+u7BLKrGHNhANdq7Z+rnNmpgFYKXPbjn4YYS5e2RCtSk6iW
DQHEIQZf0DcPFEUbJwS4YwXxB+r5NwgvFKch7f2SDSEttvN6QjJeLgqMXCCcMrourdwHTtXEAo1c
p9VcGIP+uHfGfme2Wwu+s3fs06qFrQoYzAAcL/JeleLT2MHD3bZuy6BUHIQg3Zvrj/sZChuYVaiN
0lBeI7bkzQiT5B1Oq7RduMaBuyIwWYTdZgbJ5rbntLcGYcp6dEfyQHe0E3ZnFLBHz+e7wvXUI4uc
jqD+0h9yhYCb4U/kKaiGf2E07c6IMRJrN4UcrXu39XDPR1FqCI5aClTZR8Y16bEssWLclarEZCmm
8f7J29UiUliUZfnZvUVTri+PZJ2RY+kZPgMp/axQcaseMLDP6XNPj9Q9ho3Q7ZM9EErGbTmIoVzt
GP/lPUW7aZAOVyt1SYaOne8T2HT+rWZKHTHQNfvUDzOtfB7+y/TYnImpm334iZlj2sy1VKhcQt9X
SWYGeRb0FZpl8bMo3q3vpw0+/Kb7wiLEPqygYg9sSZqWr0CN3hplyoBYKqxuyAKVybDMvoksR1eK
ChYC5PP7Wn2hNV5659KzeQOl8rkPq0wvYpgoR3OL5z3AnX7Iqx4O0LNtqjK1h4BsnxK6OZuhrorK
5oP2d2SH9IjJJQWWAAITy+rhAM3SFuHgC2Uor3Bymir7nR81QbqJfYjeHJY52iNQYGNdByZ9d6B8
upKNmdE6rcNxCRpdhI2WlsSlptgtV8c6+ngcw6dGEcYrMb+31ljvR+DzyxgS8S9mWX4ns9hKOUHm
nJuJpbMpoiqOmckYM23qWenrN4mer/chJwREknsceoEStH7CwbzRQE3XlQXXjM6FwuNcVNdC0YK6
LCE5w+MWcmUqPiZpDD6zZA3ojdN+XR2LYkc6kir7C5vrGSe4KdlTUOJfgy57jAd5v/wiG8mX4PM1
ZaC14FfCxvKwx2HzQHDyG7anmlIE+6n+GsC1xJZxducMzpFJ2yQGu8WZMJr8q2DdIkc4tb8DXfAH
qaTGfIAKI0d6l2ljcZO+89P+QBsHwXK5hEtBvmO87grK9QW9VuzhcLh7CLUt0i07XwvoEwfqjRMi
1M5U0yEvPFUuhQPKyrv2Wy0dDQBfB+/v8K+dx1F8sX+wU+9u9BRYPFcKjHvtBs6kvQSKXRKdUMAt
VB7yhA0KD4uCm5pl5k/Vzy8pBafzJOWgi7oz/YXaxRV1QiWtNMzPnMxUrD78KNThfc0299wLAlFR
D0n2GLpdxtqg6cQNBZIsKawyeDXKcLktKHCIsuYL6U4kF0KVpWfiF5YV48Q+HwD3TSHWiRnBGnMC
HYhn3AVTzMAL0Esj9EJrD+BrcBdszQvdbvgyl9ogTJARG31vRK6EXUEkSGvR9LaX9QLID1BvLZTv
NH/2zFysqP7J6KxXzNEf5aRBSFQ5otDDRHuCax4OGAKhgk06AfdbUcYyWHH9CSHy4NEUU1sTBeJj
KA9qycRhfJMxBUMDycsuUblyfOL8glylFSLQQPH5coN+GPxVrxX56ZEbF26U40Im7+n6ZzvozZu6
UtLhM2EvfodePSiveo+R60ICrY1RQeAf2SW9T9Efmp1zLm13Vs3LRPievdK+mHeQA9F5zyTAQDEp
nEwOgm6336ll1gdbJatiL7d7LA9DUiMzc+fsavfG+GZLzU/+/7AT3BsXhAtXdz5vo6XH7sSzGI9l
CARe1QXInGJZiY1YuuwO00UcUBQwKYYgdNaAflDfK+cYydTa3ICjKLxkZ0U7obd5U0aYW3DCBHMl
loNBkZ+SgA9s92feTLM5NQVwTm5tPteQM/ewAB5Qo66loWiuNirvcbg3KWtXlsZTRx5G0Dxk6ITM
o1oL1qgS9caj5G/3zD5YsAEj9iyDf/SOm57DvdTe3/TKjswpYJOxXWBJsW1bGxLxsz/QeueVuZX3
vu5GSMvfW3lRo9s4S4XuLjYjfea6HXZ1MFFuxO/zaAYpd9zF6K7w0GNv8vTPyHbMAPeqjBC1a47w
eYxLG7D/ybblfNKkI89NS63nrVr010pN4N3CKizk8QeLQzLTXy7/HI7GXWUAABL2XT3O7SAZL6im
qBY76oWEFmw3uZxNTWT/iL6GVycUCzbyGucqSE4Q3Mv2iUgvF1pvCxQ48zPVwlfUF+9hTYBGcLr+
VcgIEw/8+rlyqnKNrcygTwMphtXf7zI+dYuu5+XmjbbMeEr5Q8IF/6694PBFdcHHDrdX+oWMfXjz
EjFEPqw+z34NGFzWCO5MdYMI99Wq6eQB2So9RqOylRir75ptJsoW6Yg7bOIyzfw89zeIPBSiAIem
eQ0AubEsttryFJiOfacMP4X8oJ1R+SXSgyQdPqHisdEh4PUMsAUdaLzOECXWScZ92CcPJODkUCks
wDz6P9r4+pWI1DMBgiTHGfcwM5xfOm/5WT1Pn9qaAozoiErUhSVB/l7w9fe9xeSI0KnjsbVmrBtu
URMxJ4jQBRqyqxpq54J7fyqSupDCASerYNQHfLaQjORwIHdVUEQi90sMNBTCIlBPrcQ+saUAQgmP
GIcJjlJHVs2UuRdhr7ESxoL62P7tdnLgU+/kvUnq4Dadpby6/gWn7+LEYmTgzW1rZCOvdaCl4VeF
UmkNV7q4DJSSU/+F+7S2FgdhfCZ+foOm4Xqd7TMO2oL3ZHehPrmzlUrCF839qovK4oLA71OOJ0cH
/izVuZrjpypZeR3U3Q2U433e6bPdU2RLkeuqwHeMnCwaJqEjvnhXTy4/2Qf6hNbl33X9C4l9ENFp
xBm6LNIHLProy7CB+IEL3jXqD91uHp3eVVXtaqGo9kSGGK2rGA5/YQrPvDVLvPW7m3r6p93WM/3v
AyMO3FVpzLyTWiSFHXnicPute8XGTBo1hz5iBODyl32ciYAAuyNXWUrYKi1CvzxLNbKNBTFHwsG8
LbpUUqtJkTR4Rw4yEkLLZODLpuj1kZH1Q6LdqVf3vVMjyZiutNMyEQRxuTqPu0udYswFtDsrw4HK
W6ZRAkKJjG5volPaWGiyWDuBQzc6O1sEFSxjMg2aqKeplf7CRwn0FsNRDxT0Z9Upn2EShbw737Rq
nKUs26+jmIhO9hkF7fih8ynn8hvkcw0i0+rU8/XoyCJrUzT2rMlOBaCJi6uvp4+5kDq1ofc+831B
pRnyqJdJeCqhEGBIQLCofo1Caq5dj2rtiVe8ty68EcQBXDDjvzD2tcWPlAPaitOQgeYd7zHrc91k
K6pWg13iHziBcwfimwtTod383l0ICwF3/0yQ0UF1HwQwxkt+gFl6eA74McfUmpIqD4qrl85A9rvb
fwkIcZCjdYBiAUlur2A8kauRXBv2nw5MoIH4xtYT2kbR/QMF5C854i6jeq5Sp14W8xarDU1plQoD
jYED5EWXgcCDH++tQECxeH+RiiPB08bfcgydJusSC2oPYsWrhLDQKfQBLMeACJnGwNxr8UVqru7G
9SBRU6HDSJ72K0JbqV/6xp3cyKsveud8ph9x/RkxXjFIk4LrCIHLxkUGCy8tbkuDKZrCSJLFmWbR
c26mEuu4V5BZADD0Kg2Z7avGNoECqqNBgAast+UalY6oQo5N/0mYbxYmKTHV5osdAPbAtwXoj2V/
kmstdaJpnKmGyzsb5j5guMjwVqHnV7foIb06ifKjtYE+Az9Oy9edGnM1seGmwCozPZqrXyZwB7hc
yzt22S01zXIIhOuQPHASokvtAHY+TUBPIgRp/hNObH6XtVXfIh15KNscP6WbN8q8jgbiLK3PFDkQ
MM6vRRjGxfQtZ74LKf5fRsWEb/lVaI3q7WU8kGZ/cUMH1BvcjNBP4JTPU/o3jJmMrLjgH7HocUuP
gLVsoOcCzOA15YzhWzjjfQOOT76P9xzS0C+CZliRnA9soncwxBmhF3oBxkuQUQPFkcz+b1+c6H/E
nr/8OLceCiQWv3M9LvH3RzejY6Pqh3WCdfaJaqlr5Ud9Ed/cUWTTlhwTnV11AHh+Z4CInFH0PxTa
V5R3arv/oxOPOyb0e4nzlDA+rdusHbn/gs2bajcdBNd6ROaajG0b2s25stxosFv6Qfm+PLWMeO7Z
AE1ajhg3O9bz56IzkxjR5UEbL/sDutHa9ju/lXBS+Ddj5iRj8nN0vIydnQN0aruADZ8g3qZjLa7W
fdiX+yviwqihHkmVToHRKW5EVOZPPdbAFqMIa7q7NiijmTLWjnE3apBYP57qdy9PoSfmXI+HGius
YfUDuoQLXRkvh7MlOj9j+rcJjcGg0WL2UhM+SeiHCZQAK+GEEFKdPEB8fc0h3wBKMWI9j9tq9Uhn
Q9lFFHVrVwFP9U6TLFD4fa+mUXmBeZknDdQcaWrD2k2ammnKtDHGhEppq7oelgn7YgZasotnVyvL
ghOxHm+0im7B2/HE1hy+UmUeY/sEz7UjTSbgTNEQhKzn5TuNFp7DNX1i9QhGPrRH/oTZkpwLLMQR
m5RuuMOW+t30f2KForT5fc+KtHCyqeYwb5HGQsU3wuwPygiThiASShT0D2u/D43CxaYEr1g1LBMK
WXn1ndpZA5vOqFZs1/GIHfLNXH+cZNuK8IJFKBRCzZTS/9DlyqsKGjQeriodFU6Pt/Ia5m/O2ZJx
+iEytmihMQ8Zs6NaNEyYcLjW3DBmoHElS17uGxaGbcjdCqcjWXH2zdSF2IqNHkbQwyCfszRDlDZu
mLzKFVjcHSbATI77GSCXFpv/PTcn1y+UBivjF6gpvE4jVcyr+s53C4TMU3u6yJ6M7d37J+oEbdxE
GqP2fJ+bbBELkwHn8z6rBKTWSw2GVYfWfjPlvseieYi0KD8aQa73sMLEbdVcNdktuTQCixdH55vk
d9HDtzFcETBIO1rx7L1TTwE14tTGyVw0KksHlElngdvuY6GPhOaWAYc06w1ttjTiwXrvMr0AZc+V
dSXqpR7CFhALM5LT+I3+O0zEHBMtWQv0IbSYoO4DLOzy2Ax4pLqHo8t4n78DQJ6Cc77mErpSSKt1
0+RgBjAd/R/2AXMZu0lTZVsq2fe8aHprGA/Y7ND7BemTTifYorf4QiC598zS08+TF2qD0CvlOzJ0
lWU5y+XhmkUmJdeqHmiKL7yeKGZ4qMdPNfMUeHRNtbOOTFMzyrZBJVtRnVDyE/JHI/MQwzLBuw3B
Ah19B4CZiUJi3V6F0OaC7TddTBnKRAEiVLDsdvXX0h+hNL++sDSqVYMH+78zVPuWhh4FzM9yAvCu
wq6o4JyO0WnErER4r+BsFxG6NOcxu+K1EeEDrgtHoOQODwNuvpIDJ55Oo+Sa+LI1u9EZdypHl/SH
r8wucbWUnEA6h1x937P0cTu/KespfxT0eE67GWAeAUDGJdEr4sbEqxUoTgqoIaVIypPEZ5kubCJ9
OLf5fwaPV/ISyj/VRL7a5+GXirKKEgrkOxGRp5BODtQh7uPChzQoEYzfrDEkUvxMMYJgTfXvm8h6
4q1nDl8AK2Ix4m0vdOFLqaqc1Bw0aFa0LqIpOcdTOEDNje+togbeWI7vX5id1uZUXmimtXiNv5/p
gs7CY4gYfPUbb7LU3EcObcnQlwXNjm+Fxz5U8bjl31ki5iAp+h3d0gm37NZ/eDHqoUSzjCES+CUh
tfX7DXg4mrX7OSek6FaxIr8ON98Zrcd6UmnVdg2EVgkoBldF7qkoveRtbG++H4MIj6R+YT5vFoGN
5ZHb4PsvQ+6j5vYdCSrg0MX6yzeDQbodk07Uuh1XQhmfi8uzXDitrtgdLRTfGMJhVdAM1G4vH4h3
tY3jXH18JO1IAy13uG/lL3f+x1PKpQq/KgL7QtDanDaInwCY88auuiC/TcRFHd/QQNu0T39Ag3CY
kOiGZgT8LTiyzOg8nysZDWkqE3JWqIVBLtHNgOuDAVcAkroLHFDzl54xpxi3GkZ8orsHUTj2ai/0
IZ/cFuermFjD0TIHflFNJZS2qpJtU719gDFgQVYSCYp9jVoafAN03zfaAgGyd7VjA0xBLxhAA+zW
PAkQB688KILepP+ixuF1qpQndJEGWmuizaEPNR9Km0PD6iUDxMc7wa+nE9Sm1dYwv1f08PKskolt
PIyHs9X0HnWJBc0p94f9mzLnRdQtY8RPBPMazKmKB3WFy4Xe7wpyUK94HNMR30whHOP9s1Uhy5A2
B2hj7JMK1+ZV1hVn41VHHKD1ANXbq3OWt03ikK9GGnElnV5u3pwbX5LnYU+4foQj7vrBC/zm4fAQ
hjyc7b0xa8Tm0R6kYbQe1x6p32P1XH7xN8zZQcgBIbasyETmzj6z3JO38WhXPbYggfeehhEvf27v
u9Jue5H5pjKLC4JgfcmvOQhFRjC5HEyCihwTbD1G/mq5E/tjVW+0EnuOhkh5gYxVTdylDKRd2xxY
TUFIL0A35pWixA5LMXsP83xFsj80ZDkdArkc8oDKXOyNZUduIE2bK3kF/Rt5DooJLpp8KW+N8/Yp
yHpWASu488ZLEwD2QEEdlCfVO554euuBQ3JX1nJgG5Vvhm1PHwS88s1VNeoprST0DMkL9FsCxlXP
8/+U7/tpE9DITSl8OrdYCQzc0cjHxqblFNfF7IpEbF+mriQYKVFOJrq0GQA18HbLAb2kKdam6t1X
WDq35/qgbzeo8iq+NovV/bhczqcdJ6TtsCWYZP/RrzNQan+y9CJINjBnqoClVo2Fd/Eo+gJ+Fw4s
3U2LHdJY/DGypEgNhESe/xOiS5hhsqMhoxBVjk3FN+ex+tVkNUbbxuFYdB0W5IZiWvMpeLrbACBY
hDu0ywEI31SpyrCeMdOD2J18DpjcLI7tfK1XVbKdh53ZCMMvqvrzxNF2RevVmyOAIUfZdg76ecIf
JiIoq0RDrxQANFaq8ACzWe4C7PLQJdCFXIHm+c4CL6NjSxv/537XrSgqe0B8QUyPYJ8c5cYk8aIP
QQ0/ZqkSvh1KJrOdl6nTbxfrT8F4hVogtb9RY12h43ZSI2Jr5E37YfjvKtV9UHmj9z6tUpUP7z8R
0GcJQvby/DAyPjz1J4kYOBPNlX8DiRTXUfc+G7/YcmhBoH+SSaHXZXdlEdbGng0V40znrZSCCenZ
Zlz5eSuS/4lj1/ANIOuVuA+zFbJgH9l6STLbxur8YI7lqkdu5eTCr7jitRcfVv9nyQRmm/7M462I
GVJFfJldy/3Iu8CZbjWcleueH7QWSjJONJgqM51Snny7mXnYvT6YgSX2ZVv68RumXtEsCcpGaEL1
vidvc6wA7Y+sIqAoL4Dy1XiY4yliqvVbBCcPOyMp14zzPdVQqDFDVdj4R6Lp1fSnrhttsQ/cRS96
t9a4TTfxI4d1EGONliN9EzfXKT17I6AYIuMwbakMpRhly5mWYINvtE5tT7SQq6FcsgFzlWR10F+n
c4I+u4JNr0fR/Pow6DfGN+EwkPdZeC3he9MW5NHVWaBbNQtQ7uZ1XDRMuQ0azNKwPwpma4gUGinL
WP+Cpc2GNGXTv55VVcqVtxUS7Ap8z/WzjLP4KlaEnsv0M9eaeXriuMzv1WvrtnM+2lWShnwSobFQ
SIstIohm4uLD9bftcivsDrShmOaxSPe2QjQLxMFiyQ7zmExO9HQNKvYc1LtR4I4o7o7pXgk/BIog
jZhLS/DGyyvlRA5LZYe7OmLTZi8bSJBOnxlA3Yn3VqWcmkBDaNnJ9TvIlo1xlLGr5s+UfcBrHlsg
o7P9/Vi5M8ccxnT8qVM/w5cXlBAcwE4pIb5ETg8MUjWQry6xIV/FjfhYxuTmk0sXIJA0LqU6hDgO
dNNGlUOAK9V17D5t5s7Jn6Y9spF1y3Md+t5SMXNuJVq/f75krOkB3aQbg7ZTK3Y3RHNGyMx0fPup
4t8tftqXf8PdX33N0aS4xDYUyUr+2z7tgphdLKJyjuvDQgAz1RMk80CaRQuKv9LQjwpQWFCyyAE+
lao1qmIyJkOhuas9UOYF3FKuBz7z0f9BCvYbnyWdkHHGJDnP64y/DBgTDcBokvjTfHaDYb+gGUyi
1K6KYUf24Ho6jmqo3pEG7CZVW4OmDoS7XSJPrIJyDyWe6uUMMlXvsJspZ9o8C3hxo/wmc07/flM0
hFg/nyTvDlgCwKHZc0lj+GHzGoV9aDHak4vk7H08eYT/zkROKAhjmQw+VoDSd27CaE+n7XI8L3jA
GkFUPETf5KsHXgpblatXt9H7nWvDqSRQb+kxIcnCQvu+nSDlKgvxJFkcR4U926kkAj9o4l0ygAde
T6+VyJQxH4CFhm+JEhRxFedS1VU6ByAWulQPhekmQhB1tsAXjImANXFYFpvm4aDyLjhpAM0CNpRO
RlKk8SAVwn3PbIEiNC33DINvf7kHXAEqGzLgsPMnZpfG4bSnManSzDT5msqsHFoatw6dImXdz4MM
prN5JS+QFBAaGhxjwHeBoTs03PkK/DWmMiTkXW/EofEWBb37/SjQ61whTuBa4szniM7nawqQVewh
xxgtv59XMCdR6WshrEog1fnvG1DRxPJw5QqjJDvls7X+2mPiH5GC3OZUS85luAYiXKcPg0zm9mcW
DdHa4IOAJD7Rrmq3DPCO2ud68q6fh/S5vYlEYFfMgNEWZyfVVTlOkw1Dv7Ou8J4zodG0R7AfvXaS
uhqAAD57pDS0Fy67AbhwjibTQgvMaUY4YfL1UqYP/sk70O/g65q8A6Mppgon7YIfbxKMKzNjsOw5
9N0gRbxgHJC8v/a+/ruScPcJ37C+8OX7HzsbNpFHcghAiiAEP9qfKI+QCebEIYAO8wX5JUHFE5o/
SUOpagQG6T4UhJt56m+haLFP8m3IQxRCjnmw7uexgrII9dLsGOATGvy5d3h56SbaaC/cLMWe1hsI
7HL8EkyOcocyUeD1jV756vzIN+FobuSCx3EcVPhY3Zc/uQM2PNwqACNVZOquRo+gZfaRc7AvleSb
xA3j/XdUSQNuIyAnFmYDN29aAtwrr6LW5NUHID7HA/OX6vxgUCSzpD60hlLf5Nosa5epxHG1+na/
E7G6vTkAn8AhtjG9VA4j3jdNg8Bf859t3LGyY7MiWc7r1swkWp5y0KdWHi/aY32ssT0yU1HoO544
q6qzM7z2+i6wMWB1BEa/HRq/QXjRLxklgYpQ1L0TphimOCmud+Q3ZQsUcnjruNpMCTMaXvzKbpyd
gyfKibMotzTZb5rC9e31VjbZOP7KZdC6zAnTxXeT9+JH5gtFB7K4JAxJjRn9AhR9AtQWh2QklaIC
f72RVOHWiXPr7tyT78TY6otunlnnVT3ulQ0lGU8sBrUafl/NMS0VgqEqcKjHekTkBNickqLBP6rL
0VXDconw81SCNRlDid8s1dcZ0NxqfaHgZzgX+2+yG2UYSKSJJt6l6BPJale1VZJgWIxQS4IP20r9
Bg9KD3RzWsiVhJ2NdQxVe/ifRpQHkD4XQKPl4tK7aIhG+NptiTZmcBz7A7f+n6kSlViEyBewlkmY
Wrp3hZpMwzP5MBpUHcEkKqXHF17DHLx9kyTJqbgX6HmPGK32M0agEbmV0yz+//GOMchq8yqLNbqL
1fyyxTODbOTnZDdzTOVVSre3cy3cnYP4/Sc09RpsSwphvw/y2uygRMTLjq/+Y+LIhKkuKpxmvi1E
zAxD28AQ90BP2LdpsHA4FQa45oasNx4eL1Pb8+LbP8RXf3kZmKks6LZAQuea+E7SP2pAQ7mrJVD/
YR3Q0ln0+rKsStMCOnoByfnEGlAhgx1lFCilCQZBDEgU+znYV+obSQ0fyvO0Un3VGn/Jc1boDLrq
6jkM7NbVbTqqOQ3uGBwFJb3j1t1Davd+mpbuZt0wTMxZwXA4DnLPZgTCZjdW8U9ErnX9A14aS2HT
QzgIpM2cBwFzUszGxHhvmmWHX1Mnh9E/2MSYwpx7f8ed2TCM4XA0shNZVnFWcPWvAi3eITgblIh5
vd91eZ7/regHrAwbTwYhB7alkcVx/FbPR82FVWznAj4XEdkpsEVtXeBIQV2PQQ2iN0ONYdz2LkL2
LuvK8fwcA7OcxfIx75+lcyQyg7zO86c5DwJuOjNUx+uQ8FlELXFx7fopZU0rgka+tucNQUO8G+vU
wxBqTetwW0qjNZsAWZkioDMK+UZKVs7BYXrfJaeX+MiNBe/1S8iGnlKWTdqvwmzrasgPD75OPifs
aM1nn7O3deuWlLDP9KbC9aGFXxsIvsseRBeNg4ALAt/0qmcN06L6dOUq9Jai/wqBHpSZ1F3r+tUV
+7/3RcCqK0wyoTGEYIqCRh8GI+2ZEKpRkH/fdtfdbPVzU/JCQJtchZ4gN/gUhYaKBMfM4Ybn7jFu
VeyIfee6JXqsCbO6haVdqMahTfnX69pbG/kJGlz178JutK0V6EsCghUDVuRUgH14s5L+yO5JKPkn
90eB309gtpLuvnr03WgDPKDeeZXDUxkoOO3O9mcwT5R9VLW8/WhoO7cPQmj9C4JuQef/2+4nIa/0
ffKg1DYj7XgysWqAY57WrmXY0kI5SU61hvgefgC5qBpD+ErjWCongynKbAy72z9tuxco+1yvRF1l
VWW1rZ0zdy/zRKTKzySYFU/OGy53nQDKn77pUd79guPzsd4WMk71z+oWT0HxAdoh1QEMF9rzLgLp
//QEE21R1sqSuV/WYenl7LGsrFEP+Dl17nljeCUqPY+mTZLjFCGgMPfjpOlYqrQGkLTS0T5IdxHO
emnBqXr+RtwNsTwmFwmKX1iSLvf6RhnDRxqrPpqvFUsSuK55cTLeT7TVEjCaZUNg6JlZwAB+cDky
WJlMPjM+ErSWRCROiaiadKhHT4fZuVRCfg/V1owQ7ebsH94/MuG51wIW9Dvy3KfV+XWOT1AEmgvb
IcHuR0OvikJ2K+BEqGjY3vUJWC8B9HHUte0bBvSpbaeMfFklVOXSRCa8TFLekeImZWdLyFROjy1X
dKXyDSzer1DtKC47d0MEgfAu5uqjJYYQrOcEY1rDt6uyBKvueWV8jvZ4gu1v73GkCs40kQKf6Vgy
8aPB2UkOAZKJMKgcQm8643gixUcpfz89NeAfyc+p6tIkuvC9Kx2PPIEKI2J1syS8BQ0UAKjYVMoY
NQ2E0fSyyU1qiHDidQp1Cc+RN+Vns8O2hdTtmyYXby2bKSNmEEMQm0mxpyRMdRsHkBxHSTUzqnbk
207dIZ0KkPF6g66UN4B+NKJiht6XHcdkRts8zchIzdy33Ovyk2BI/QQhBxLAX7O+x91FMdQCzERK
p1zxEmV+XEBEare74nndBiznyfAdcYBnLDX//BI41b9s+EDyhxDvdPf2D2FFTOMcHzOOPWxOeSTz
AZTBTKKor2ZdAipDRpVstFmU/nWXRHufj+WjIvtayEz5YCKLSn0NfqSybZGJ2Aw+qYxvT4paRj8k
TxPTWsr6nDKFphug1NlFjwt3BiqJjHHZa6Nrdxar1tw7NgunKzIJ5i7BsBFQojqVKiSoiw2gh7ty
KzoTsePmWrA1vHkwMysx1To8Ky7pKEVilMDPXOxRSfLotP4Nw3gHxj+ryGtwv0j6g1XExmkt24li
HQripFWlscgx+euQhnNKL6Tj8M4fFwrDKzJ9xw0rUwlmi3+k2exrB3JuQmcXkFhMrZcyfXjL7HJp
Vmkfn1aboiFxa/+OaAkLywMLxKT3CB5bFADTFgbCZGfU9PhfP4KXiAE4p2SU1MQpf5RRRHB1IuYn
R2aFNMwkdTJgBlTe82NrnGuy10Wadg/1MiBIqSyzdTC7UduPygow8Ehc6yMdLKrZxyeYVf4UV/6F
ke8dgmRkbOtT2AM704pMbcJ2P/6AJCv8uuaghdyPRthgThDCDCEEpd3eR0cu5n0BIdiFuIoaQAIv
icBpMhLTcSy8vD2UJCTLVQK99FJATdRla7hcpprMrkloiP0ARMZkmdoRoqrPQg8kZqHGIAKdTXTr
wlp3i9JbP5Uk4khuf2IiOIo5OTIor0Oj1g9BiF4mv4DeTfGWrE3W/jxWK9ttjwFJzMjHkdTAJ3Nu
9iRBgUxLnz72UPFfMnYXQYgilZDNMg1uZcG06JaZeQ39DQTvXGPrSRkOj5oo4nts4gn8SE2b+Gcf
nM+ZZGFaBv4Tmh2ndiFuH5lfGivhZXUp9gLxgkikD+rfKLTL4JFcUCJCVTqFKbC26wiYKPAWiQNY
05wBjHE279rWAGwxPedTMzm33UkTY7LerSu9/5Ekq2afQ9ubwOMuQu6HIBg23e132oBXRD1Tzxzx
ItkjncFibugrZjHEHnHluQujyxucyyKqnmzS7+Gw6i17WeHLQoRbrhHYj6GjBAK9L59mD4KWbBJj
3bfvDUlwNaMSAvAUIVZKoc+SCRhwITaEzaD1GgV5uGdO+fOTbPu8g/vNKX8lPqhxb51pFVc5tS55
gLzqMUcGvoOKWLEeFYKlA7a//X1HqZ2t9NOEcWzljilPfDTnSycUZZ+lvEUk3mCBu76k1bbdRi0v
hRdQH4znx4s8ym4oAfch9s/jhMts+6FC4+saYLPOzDWpFNYnlAJhisZ2Ew0nUFJQWYV3s5B+9kE3
77zVDHy61HvhDCwtePhqNkbxMlTNA9W5s2S9YOUuUTwNVPbRfarRpkV9Y3M2RBDgeyietV1SFD9z
T/u/w6s1Xq+RcE5d8Gjjst4W/Jd+5PfnhIAClIkwm5zWjRxz5o1e4eTp4YYX10GZB+/eFAwyP+SZ
yoSJQh6auw27BimmxCUMHcQIRkyi+SafM7mxmzwxuCEADKtqAQPxQ7dAe9wDM9abkkQzGsCwyhYP
Vv1iCkJaoecs/wPuDZYIOVM9u8PecRUi5Xi2EPp/TC/AxCxOxC/4nkC3qr80a9X41YucGPjJ2tC0
fneiEGheM0cczIIOQ+EyMrw9hrw/Lm9hmO519mhk5Iu+KXzIS1igFm17xOfToZJdgwlVRdN5dRtv
V2HrbfEEydq+6E2YZkhEWrs5tbPvz/VfcjvzP2OsgIdTljyeGHYqSFcjzhg+0Xpi/QaLjLunU4Ls
7w3xrH69MT882QH6xiTZDLHAMWJ4PimwAWUhFYSi96fBcjllwYitlwbqwkSqIyLyYUbmVN32iTpg
3UmYFBbb1tGzp26MzGywO/uojpCX+XSgoi/kF7xUDBCmD+awpZ5r4xmnspj3ikiCTfwZC3+84JxN
KhqCyDZVMDiuJRvFgbAtx9oSaq5E2AQxcJourHYazd+Hh+ilmE7yqPW/yD1UVpqsFu0hVBHsPJy5
L2A0SivVntjp7vEqg2l7/BSzWIfoqhuBp5W598sHdmRefTSpIdgEtqT1uZcTMe8l9LFJGlsXXwIF
IB6RVmP+65Fho5FvcfLqTnvYg5zF614tAVtKUB7Dz+wbV9bxDeQsmGn4mR6jLCJjg0S4wHY59LD6
xrBKEM9ZhNVb0sFSZ7LiygdLmi1olTrIn0nWM1n62wP7OjGjMqVpHTxtgfBgS7/9McLSqvWoZLkm
mqqpwXMKR75UJWZODe+UhVm3O9kQ3+q07pgjw+KYBZjZuhgazKsGOI4VkdNE9Kr16jtZVzfLtDi1
LCaSsAmBtvQ9mf66gOWKjkmysYfep0a95+kMfb1mJqq3iS8ZUypOuYta+9WXjLGaxSfAwr/uhakL
3JWvHQSRKndQdeIBD300J1qmS1EbrT+325gHu5mf3k+S1GhYn1x0RMgum210Ekc+PzgEOtP7CPld
41SbNsm44XNjFrsLlbOKKoDnvVnb0NS9p9augc42dxWrsjirmDrKvMKoYCvbvIuMPZPVgthkzm7e
RiMY8dbzSYw2s6QmvLF3pgapC7Aj9ze3Kk+2IHCwzxc1s/BZBOQ9MRn9CPKdpI3PFdLdxq52ydnB
6KLj1owT0YGrZB7d1VfJ/GN08JEoYCXl6+6RB6tkYvzw4wXjuMMPb4YmX31a1Ev6uCm1yWa8cFzi
DLbx7EGi4FBMSGVWO3plNJaz7ZWB4ypbaQIXhKPbIssKzpvabHZD/lMfKlZWWGNr3e/3G3dMg/+b
/Enc+iEeMVnIzHWsq6O4nUDymvUI25+zEqUXsPyjv40BHaHTir5lqDDdrP5Y5PB8IQ2x1PimFQ30
32solfjCB/4/eoIitYV2anwVXo5Hp8OIPA+1MQmMSLdxDmFBoBJuoFvBy9xUXhkwy5Esu+FR2jUB
1f9/HOwNUDPjZ57JoVnT2qSVLoUaVmbvBb0gtn4YNkYJ1wYg/gocQfb5GvR8AnB1BrNa3RuEy+Ou
GWVoXifvaULTZrLRiIm9hndblcynWS5oE3d3e04glmeoB0FFhALTbzeEN4BCstQniugb080fn748
pqjOACjWeErH+G1ybCBqImhI2EWVrGR9IcXZRBmkv+fnUhsQ1+scPhqQgrM3Z7Cxq5yxpFO5yiIT
6UK99aglHMsMlBA87SCFswQ+5zeYM+Ik1wczahsV6ZwY/2VXI6bhy9MPpUJakwTou53fkJkKZVZr
RDVNxMwBk31MpwOtIR2YTrCVUJMhTNScD/pkOL3eWN4W148NFRNdTWGWlKgNIpvDuKMZmg1nUMt2
lKVyr2oP1J+K2l/BW0srgxX/Frp9Iq4I1gwcm78iRQJ+LBJrF7oDOYAGp8tigWAJ+odUVP1+ppqO
CZQEXVnzG/l7xmc2x75F1uIy3OD1gxld6O/PeXIiJP0YgZ+UsDOI2YjD170+Wgn3/GwILZS+XQ6g
U54TQSQ=
`protect end_protected

